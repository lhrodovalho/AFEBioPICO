magic
tech sky130A
timestamp 1637857729
<< metal2 >>
rect 5520 16595 7320 16600
rect 5520 16565 5525 16595
rect 5555 16565 5685 16595
rect 5715 16565 5845 16595
rect 5875 16565 6005 16595
rect 6035 16565 6165 16595
rect 6195 16565 6325 16595
rect 6355 16565 6485 16595
rect 6515 16565 6645 16595
rect 6675 16565 6805 16595
rect 6835 16565 6965 16595
rect 6995 16565 7125 16595
rect 7155 16565 7285 16595
rect 7315 16565 7320 16595
rect 5520 16560 7320 16565
rect 7360 16595 7720 16600
rect 7360 16565 7365 16595
rect 7395 16565 7525 16595
rect 7555 16565 7685 16595
rect 7715 16565 7720 16595
rect 7360 16560 7720 16565
rect 5520 16515 7320 16520
rect 5520 16485 5525 16515
rect 5555 16485 5685 16515
rect 5715 16485 5845 16515
rect 5875 16485 6005 16515
rect 6035 16485 6165 16515
rect 6195 16485 6325 16515
rect 6355 16485 6485 16515
rect 6515 16485 6645 16515
rect 6675 16485 6805 16515
rect 6835 16485 6965 16515
rect 6995 16485 7125 16515
rect 7155 16485 7285 16515
rect 7315 16485 7320 16515
rect 5520 16480 7320 16485
rect 7360 16515 7720 16520
rect 7360 16485 7365 16515
rect 7395 16485 7525 16515
rect 7555 16485 7685 16515
rect 7715 16485 7720 16515
rect 7360 16480 7720 16485
rect 5520 16435 7320 16440
rect 5520 16405 5525 16435
rect 5555 16405 5685 16435
rect 5715 16405 5845 16435
rect 5875 16405 6005 16435
rect 6035 16405 6165 16435
rect 6195 16405 6325 16435
rect 6355 16405 6485 16435
rect 6515 16405 6645 16435
rect 6675 16405 6805 16435
rect 6835 16405 6965 16435
rect 6995 16405 7125 16435
rect 7155 16405 7285 16435
rect 7315 16405 7320 16435
rect 5520 16400 7320 16405
rect 7360 16435 7720 16440
rect 7360 16405 7365 16435
rect 7395 16405 7525 16435
rect 7555 16405 7685 16435
rect 7715 16405 7720 16435
rect 7360 16400 7720 16405
rect 5520 16355 7320 16360
rect 5520 16325 5525 16355
rect 5555 16325 5685 16355
rect 5715 16325 5845 16355
rect 5875 16325 6005 16355
rect 6035 16325 6165 16355
rect 6195 16325 6325 16355
rect 6355 16325 6485 16355
rect 6515 16325 6645 16355
rect 6675 16325 6805 16355
rect 6835 16325 6965 16355
rect 6995 16325 7125 16355
rect 7155 16325 7285 16355
rect 7315 16325 7320 16355
rect 5520 16320 7320 16325
rect 7360 16355 7720 16360
rect 7360 16325 7365 16355
rect 7395 16325 7525 16355
rect 7555 16325 7685 16355
rect 7715 16325 7720 16355
rect 7360 16320 7720 16325
rect 5520 16275 7320 16280
rect 5520 16245 5525 16275
rect 5555 16245 5685 16275
rect 5715 16245 5845 16275
rect 5875 16245 6005 16275
rect 6035 16245 6165 16275
rect 6195 16245 6325 16275
rect 6355 16245 6485 16275
rect 6515 16245 6645 16275
rect 6675 16245 6805 16275
rect 6835 16245 6965 16275
rect 6995 16245 7125 16275
rect 7155 16245 7285 16275
rect 7315 16245 7320 16275
rect 5520 16240 7320 16245
rect 7360 16275 7720 16280
rect 7360 16245 7365 16275
rect 7395 16245 7525 16275
rect 7555 16245 7685 16275
rect 7715 16245 7720 16275
rect 7360 16240 7720 16245
rect 5520 16195 7320 16200
rect 5520 16165 5525 16195
rect 5555 16165 5685 16195
rect 5715 16165 5845 16195
rect 5875 16165 6005 16195
rect 6035 16165 6165 16195
rect 6195 16165 6325 16195
rect 6355 16165 6485 16195
rect 6515 16165 6645 16195
rect 6675 16165 6805 16195
rect 6835 16165 6965 16195
rect 6995 16165 7125 16195
rect 7155 16165 7285 16195
rect 7315 16165 7320 16195
rect 5520 16160 7320 16165
rect 7360 16195 7720 16200
rect 7360 16165 7365 16195
rect 7395 16165 7525 16195
rect 7555 16165 7685 16195
rect 7715 16165 7720 16195
rect 7360 16160 7720 16165
rect 5520 16115 7320 16120
rect 5520 16085 5525 16115
rect 5555 16085 5685 16115
rect 5715 16085 5845 16115
rect 5875 16085 6005 16115
rect 6035 16085 6165 16115
rect 6195 16085 6325 16115
rect 6355 16085 6485 16115
rect 6515 16085 6645 16115
rect 6675 16085 6805 16115
rect 6835 16085 6965 16115
rect 6995 16085 7125 16115
rect 7155 16085 7285 16115
rect 7315 16085 7320 16115
rect 5520 16080 7320 16085
rect 7360 16115 7720 16120
rect 7360 16085 7365 16115
rect 7395 16085 7525 16115
rect 7555 16085 7685 16115
rect 7715 16085 7720 16115
rect 7360 16080 7720 16085
rect 5520 16035 7320 16040
rect 5520 16005 5525 16035
rect 5555 16005 5685 16035
rect 5715 16005 5845 16035
rect 5875 16005 6005 16035
rect 6035 16005 6165 16035
rect 6195 16005 6325 16035
rect 6355 16005 6485 16035
rect 6515 16005 6645 16035
rect 6675 16005 6805 16035
rect 6835 16005 6965 16035
rect 6995 16005 7125 16035
rect 7155 16005 7285 16035
rect 7315 16005 7320 16035
rect 5520 16000 7320 16005
rect 7360 16035 7720 16040
rect 7360 16005 7365 16035
rect 7395 16005 7525 16035
rect 7555 16005 7685 16035
rect 7715 16005 7720 16035
rect 7360 16000 7720 16005
rect 5520 15955 7320 15960
rect 5520 15925 5525 15955
rect 5555 15925 5685 15955
rect 5715 15925 5845 15955
rect 5875 15925 6005 15955
rect 6035 15925 6165 15955
rect 6195 15925 6325 15955
rect 6355 15925 6485 15955
rect 6515 15925 6645 15955
rect 6675 15925 6805 15955
rect 6835 15925 6965 15955
rect 6995 15925 7125 15955
rect 7155 15925 7285 15955
rect 7315 15925 7320 15955
rect 5520 15920 7320 15925
rect 7360 15955 7720 15960
rect 7360 15925 7365 15955
rect 7395 15925 7525 15955
rect 7555 15925 7685 15955
rect 7715 15925 7720 15955
rect 7360 15920 7720 15925
rect 5520 15875 7720 15880
rect 5520 15845 7365 15875
rect 7395 15845 7525 15875
rect 7555 15845 7685 15875
rect 7715 15845 7720 15875
rect 5520 15840 7720 15845
rect 5480 15795 7640 15800
rect 5480 15765 7605 15795
rect 7635 15765 7640 15795
rect 5480 15760 7640 15765
rect 5480 15715 7720 15720
rect 5480 15685 7365 15715
rect 7395 15685 7525 15715
rect 7555 15685 7685 15715
rect 7715 15685 7720 15715
rect 5480 15680 7720 15685
rect 5480 15635 7480 15640
rect 5480 15605 7445 15635
rect 7475 15605 7480 15635
rect 5480 15600 7480 15605
rect 5520 15555 7720 15560
rect 5520 15525 7365 15555
rect 7395 15525 7525 15555
rect 7555 15525 7685 15555
rect 7715 15525 7720 15555
rect 5520 15520 7720 15525
rect 5520 15435 7320 15440
rect 5520 15405 5525 15435
rect 5555 15405 5685 15435
rect 5715 15405 5845 15435
rect 5875 15405 6005 15435
rect 6035 15405 6165 15435
rect 6195 15405 6325 15435
rect 6355 15405 6485 15435
rect 6515 15405 6645 15435
rect 6675 15405 6805 15435
rect 6835 15405 6965 15435
rect 6995 15405 7125 15435
rect 7155 15405 7285 15435
rect 7315 15405 7320 15435
rect 5520 15400 7320 15405
rect 7360 15435 7720 15440
rect 7360 15405 7365 15435
rect 7395 15405 7525 15435
rect 7555 15405 7685 15435
rect 7715 15405 7720 15435
rect 7360 15400 7720 15405
rect 5520 15355 7320 15360
rect 5520 15325 5525 15355
rect 5555 15325 5685 15355
rect 5715 15325 5845 15355
rect 5875 15325 6005 15355
rect 6035 15325 6165 15355
rect 6195 15325 6325 15355
rect 6355 15325 6485 15355
rect 6515 15325 6645 15355
rect 6675 15325 6805 15355
rect 6835 15325 6965 15355
rect 6995 15325 7125 15355
rect 7155 15325 7285 15355
rect 7315 15325 7320 15355
rect 5520 15320 7320 15325
rect 7360 15355 7720 15360
rect 7360 15325 7365 15355
rect 7395 15325 7525 15355
rect 7555 15325 7685 15355
rect 7715 15325 7720 15355
rect 7360 15320 7720 15325
rect 5520 15275 7320 15280
rect 5520 15245 5525 15275
rect 5555 15245 5685 15275
rect 5715 15245 5845 15275
rect 5875 15245 6005 15275
rect 6035 15245 6165 15275
rect 6195 15245 6325 15275
rect 6355 15245 6485 15275
rect 6515 15245 6645 15275
rect 6675 15245 6805 15275
rect 6835 15245 6965 15275
rect 6995 15245 7125 15275
rect 7155 15245 7285 15275
rect 7315 15245 7320 15275
rect 5520 15240 7320 15245
rect 7360 15275 7720 15280
rect 7360 15245 7365 15275
rect 7395 15245 7525 15275
rect 7555 15245 7685 15275
rect 7715 15245 7720 15275
rect 7360 15240 7720 15245
rect 5520 15195 7320 15200
rect 5520 15165 5525 15195
rect 5555 15165 5685 15195
rect 5715 15165 5845 15195
rect 5875 15165 6005 15195
rect 6035 15165 6165 15195
rect 6195 15165 6325 15195
rect 6355 15165 6485 15195
rect 6515 15165 6645 15195
rect 6675 15165 6805 15195
rect 6835 15165 6965 15195
rect 6995 15165 7125 15195
rect 7155 15165 7285 15195
rect 7315 15165 7320 15195
rect 5520 15160 7320 15165
rect 7360 15195 7720 15200
rect 7360 15165 7365 15195
rect 7395 15165 7525 15195
rect 7555 15165 7685 15195
rect 7715 15165 7720 15195
rect 7360 15160 7720 15165
rect 5520 15115 7320 15120
rect 5520 15085 5525 15115
rect 5555 15085 5685 15115
rect 5715 15085 5845 15115
rect 5875 15085 6005 15115
rect 6035 15085 6165 15115
rect 6195 15085 6325 15115
rect 6355 15085 6485 15115
rect 6515 15085 6645 15115
rect 6675 15085 6805 15115
rect 6835 15085 6965 15115
rect 6995 15085 7125 15115
rect 7155 15085 7285 15115
rect 7315 15085 7320 15115
rect 5520 15080 7320 15085
rect 7360 15115 7720 15120
rect 7360 15085 7365 15115
rect 7395 15085 7525 15115
rect 7555 15085 7685 15115
rect 7715 15085 7720 15115
rect 7360 15080 7720 15085
rect 5480 15035 6120 15040
rect 5480 15005 6085 15035
rect 6115 15005 6120 15035
rect 5480 15000 6120 15005
rect 6160 15035 7320 15040
rect 6160 15005 6165 15035
rect 6195 15005 6325 15035
rect 6355 15005 6485 15035
rect 6515 15005 6645 15035
rect 6675 15005 6805 15035
rect 6835 15005 6965 15035
rect 6995 15005 7125 15035
rect 7155 15005 7285 15035
rect 7315 15005 7320 15035
rect 6160 15000 7320 15005
rect 7360 15035 7720 15040
rect 7360 15005 7365 15035
rect 7395 15005 7525 15035
rect 7555 15005 7685 15035
rect 7715 15005 7720 15035
rect 7360 15000 7720 15005
rect 5520 14955 7320 14960
rect 5520 14925 5525 14955
rect 5555 14925 5685 14955
rect 5715 14925 5845 14955
rect 5875 14925 6005 14955
rect 6035 14925 6165 14955
rect 6195 14925 6325 14955
rect 6355 14925 6485 14955
rect 6515 14925 6645 14955
rect 6675 14925 6805 14955
rect 6835 14925 6965 14955
rect 6995 14925 7125 14955
rect 7155 14925 7285 14955
rect 7315 14925 7320 14955
rect 5520 14920 7320 14925
rect 7360 14955 7720 14960
rect 7360 14925 7365 14955
rect 7395 14925 7525 14955
rect 7555 14925 7685 14955
rect 7715 14925 7720 14955
rect 7360 14920 7720 14925
rect 5520 14875 7320 14880
rect 5520 14845 5525 14875
rect 5555 14845 5685 14875
rect 5715 14845 5845 14875
rect 5875 14845 6005 14875
rect 6035 14845 6165 14875
rect 6195 14845 6325 14875
rect 6355 14845 6485 14875
rect 6515 14845 6645 14875
rect 6675 14845 6805 14875
rect 6835 14845 6965 14875
rect 6995 14845 7125 14875
rect 7155 14845 7285 14875
rect 7315 14845 7320 14875
rect 5520 14840 7320 14845
rect 7360 14875 7720 14880
rect 7360 14845 7365 14875
rect 7395 14845 7525 14875
rect 7555 14845 7685 14875
rect 7715 14845 7720 14875
rect 7360 14840 7720 14845
rect 5520 14795 7320 14800
rect 5520 14765 5525 14795
rect 5555 14765 5685 14795
rect 5715 14765 5845 14795
rect 5875 14765 6005 14795
rect 6035 14765 6165 14795
rect 6195 14765 6325 14795
rect 6355 14765 6485 14795
rect 6515 14765 6645 14795
rect 6675 14765 6805 14795
rect 6835 14765 6965 14795
rect 6995 14765 7125 14795
rect 7155 14765 7285 14795
rect 7315 14765 7320 14795
rect 5520 14760 7320 14765
rect 7360 14795 7720 14800
rect 7360 14765 7365 14795
rect 7395 14765 7525 14795
rect 7555 14765 7685 14795
rect 7715 14765 7720 14795
rect 7360 14760 7720 14765
rect 5520 14715 7320 14720
rect 5520 14685 5525 14715
rect 5555 14685 5685 14715
rect 5715 14685 5845 14715
rect 5875 14685 6005 14715
rect 6035 14685 6165 14715
rect 6195 14685 6325 14715
rect 6355 14685 6485 14715
rect 6515 14685 6645 14715
rect 6675 14685 6805 14715
rect 6835 14685 6965 14715
rect 6995 14685 7125 14715
rect 7155 14685 7285 14715
rect 7315 14685 7320 14715
rect 5520 14680 7320 14685
rect 7360 14715 7720 14720
rect 7360 14685 7365 14715
rect 7395 14685 7525 14715
rect 7555 14685 7685 14715
rect 7715 14685 7720 14715
rect 7360 14680 7720 14685
rect 5480 14635 5960 14640
rect 5480 14605 5925 14635
rect 5955 14605 5960 14635
rect 5480 14600 5960 14605
rect 6000 14635 7320 14640
rect 6000 14605 6005 14635
rect 6035 14605 6165 14635
rect 6195 14605 6325 14635
rect 6355 14605 6485 14635
rect 6515 14605 6645 14635
rect 6675 14605 6805 14635
rect 6835 14605 6965 14635
rect 6995 14605 7125 14635
rect 7155 14605 7285 14635
rect 7315 14605 7320 14635
rect 6000 14600 7320 14605
rect 7360 14635 7720 14640
rect 7360 14605 7365 14635
rect 7395 14605 7525 14635
rect 7555 14605 7685 14635
rect 7715 14605 7720 14635
rect 7360 14600 7720 14605
rect 5520 14555 7320 14560
rect 5520 14525 5525 14555
rect 5555 14525 5685 14555
rect 5715 14525 5845 14555
rect 5875 14525 6005 14555
rect 6035 14525 6165 14555
rect 6195 14525 6325 14555
rect 6355 14525 6485 14555
rect 6515 14525 6645 14555
rect 6675 14525 6805 14555
rect 6835 14525 6965 14555
rect 6995 14525 7125 14555
rect 7155 14525 7285 14555
rect 7315 14525 7320 14555
rect 5520 14520 7320 14525
rect 7360 14555 7720 14560
rect 7360 14525 7365 14555
rect 7395 14525 7525 14555
rect 7555 14525 7685 14555
rect 7715 14525 7720 14555
rect 7360 14520 7720 14525
rect 5520 14475 7320 14480
rect 5520 14445 5525 14475
rect 5555 14445 5685 14475
rect 5715 14445 5845 14475
rect 5875 14445 6005 14475
rect 6035 14445 6165 14475
rect 6195 14445 6325 14475
rect 6355 14445 6485 14475
rect 6515 14445 6645 14475
rect 6675 14445 6805 14475
rect 6835 14445 6965 14475
rect 6995 14445 7125 14475
rect 7155 14445 7285 14475
rect 7315 14445 7320 14475
rect 5520 14440 7320 14445
rect 7360 14475 7720 14480
rect 7360 14445 7365 14475
rect 7395 14445 7525 14475
rect 7555 14445 7685 14475
rect 7715 14445 7720 14475
rect 7360 14440 7720 14445
rect 5520 14395 7320 14400
rect 5520 14365 6965 14395
rect 6995 14365 7125 14395
rect 7155 14365 7285 14395
rect 7315 14365 7320 14395
rect 5520 14360 7320 14365
rect 7360 14395 7720 14400
rect 7360 14365 7365 14395
rect 7395 14365 7525 14395
rect 7555 14365 7685 14395
rect 7715 14365 7720 14395
rect 7360 14360 7720 14365
rect 5480 14315 7240 14320
rect 5480 14285 7205 14315
rect 7235 14285 7240 14315
rect 5480 14280 7240 14285
rect 7360 14315 7720 14320
rect 7360 14285 7365 14315
rect 7395 14285 7525 14315
rect 7555 14285 7685 14315
rect 7715 14285 7720 14315
rect 7360 14280 7720 14285
rect 5480 14235 7320 14240
rect 5480 14205 6965 14235
rect 6995 14205 7125 14235
rect 7155 14205 7285 14235
rect 7315 14205 7320 14235
rect 5480 14200 7320 14205
rect 7360 14235 7720 14240
rect 7360 14205 7365 14235
rect 7395 14205 7525 14235
rect 7555 14205 7685 14235
rect 7715 14205 7720 14235
rect 7360 14200 7720 14205
rect 5480 14155 7080 14160
rect 5480 14125 7045 14155
rect 7075 14125 7080 14155
rect 5480 14120 7080 14125
rect 7360 14155 7720 14160
rect 7360 14125 7365 14155
rect 7395 14125 7525 14155
rect 7555 14125 7685 14155
rect 7715 14125 7720 14155
rect 7360 14120 7720 14125
rect 5520 14075 7320 14080
rect 5520 14045 6965 14075
rect 6995 14045 7125 14075
rect 7155 14045 7285 14075
rect 7315 14045 7320 14075
rect 5520 14040 7320 14045
rect 7360 14075 7720 14080
rect 7360 14045 7365 14075
rect 7395 14045 7525 14075
rect 7555 14045 7685 14075
rect 7715 14045 7720 14075
rect 7360 14040 7720 14045
rect 5520 13995 7320 14000
rect 5520 13965 5525 13995
rect 5555 13965 5685 13995
rect 5715 13965 5845 13995
rect 5875 13965 6005 13995
rect 6035 13965 6165 13995
rect 6195 13965 6325 13995
rect 6355 13965 6485 13995
rect 6515 13965 6645 13995
rect 6675 13965 6805 13995
rect 6835 13965 6965 13995
rect 6995 13965 7125 13995
rect 7155 13965 7285 13995
rect 7315 13965 7320 13995
rect 5520 13960 7320 13965
rect 7360 13995 7720 14000
rect 7360 13965 7365 13995
rect 7395 13965 7525 13995
rect 7555 13965 7685 13995
rect 7715 13965 7720 13995
rect 7360 13960 7720 13965
rect 5480 13915 5800 13920
rect 5480 13885 5765 13915
rect 5795 13885 5800 13915
rect 5480 13880 5800 13885
rect 5840 13875 7320 13880
rect 5840 13845 5845 13875
rect 5875 13845 6005 13875
rect 6035 13845 6165 13875
rect 6195 13845 6325 13875
rect 6355 13845 6485 13875
rect 6515 13845 6645 13875
rect 6675 13845 6805 13875
rect 6835 13845 6965 13875
rect 6995 13845 7125 13875
rect 7155 13845 7285 13875
rect 7315 13845 7320 13875
rect 5840 13840 7320 13845
rect 7360 13875 7720 13880
rect 7360 13845 7365 13875
rect 7395 13845 7525 13875
rect 7555 13845 7685 13875
rect 7715 13845 7720 13875
rect 7360 13840 7720 13845
rect 5520 13795 7320 13800
rect 5520 13765 5525 13795
rect 5555 13765 5685 13795
rect 5715 13765 5845 13795
rect 5875 13765 6005 13795
rect 6035 13765 6165 13795
rect 6195 13765 6325 13795
rect 6355 13765 6485 13795
rect 6515 13765 6645 13795
rect 6675 13765 6805 13795
rect 6835 13765 6965 13795
rect 6995 13765 7125 13795
rect 7155 13765 7285 13795
rect 7315 13765 7320 13795
rect 5520 13760 7320 13765
rect 7360 13795 7720 13800
rect 7360 13765 7365 13795
rect 7395 13765 7525 13795
rect 7555 13765 7685 13795
rect 7715 13765 7720 13795
rect 7360 13760 7720 13765
rect 5520 13715 7320 13720
rect 5520 13685 5525 13715
rect 5555 13685 5685 13715
rect 5715 13685 5845 13715
rect 5875 13685 6005 13715
rect 6035 13685 6165 13715
rect 6195 13685 6325 13715
rect 6355 13685 6485 13715
rect 6515 13685 6645 13715
rect 6675 13685 6805 13715
rect 6835 13685 6965 13715
rect 6995 13685 7125 13715
rect 7155 13685 7285 13715
rect 7315 13685 7320 13715
rect 5520 13680 7320 13685
rect 7360 13715 7720 13720
rect 7360 13685 7365 13715
rect 7395 13685 7525 13715
rect 7555 13685 7685 13715
rect 7715 13685 7720 13715
rect 7360 13680 7720 13685
rect 5520 13635 7320 13640
rect 5520 13605 5525 13635
rect 5555 13605 5685 13635
rect 5715 13605 5845 13635
rect 5875 13605 6005 13635
rect 6035 13605 6165 13635
rect 6195 13605 6325 13635
rect 6355 13605 6485 13635
rect 6515 13605 6645 13635
rect 6675 13605 6805 13635
rect 6835 13605 6965 13635
rect 6995 13605 7125 13635
rect 7155 13605 7285 13635
rect 7315 13605 7320 13635
rect 5520 13600 7320 13605
rect 7360 13635 7720 13640
rect 7360 13605 7365 13635
rect 7395 13605 7525 13635
rect 7555 13605 7685 13635
rect 7715 13605 7720 13635
rect 7360 13600 7720 13605
rect 5480 13555 6120 13560
rect 5480 13525 6085 13555
rect 6115 13525 6120 13555
rect 5480 13520 6120 13525
rect 6160 13555 7320 13560
rect 6160 13525 6165 13555
rect 6195 13525 6325 13555
rect 6355 13525 6485 13555
rect 6515 13525 6645 13555
rect 6675 13525 6805 13555
rect 6835 13525 6965 13555
rect 6995 13525 7125 13555
rect 7155 13525 7285 13555
rect 7315 13525 7320 13555
rect 6160 13520 7320 13525
rect 7360 13555 7720 13560
rect 7360 13525 7365 13555
rect 7395 13525 7525 13555
rect 7555 13525 7685 13555
rect 7715 13525 7720 13555
rect 7360 13520 7720 13525
rect 5520 13475 7320 13480
rect 5520 13445 5525 13475
rect 5555 13445 5685 13475
rect 5715 13445 5845 13475
rect 5875 13445 6005 13475
rect 6035 13445 6165 13475
rect 6195 13445 6325 13475
rect 6355 13445 6485 13475
rect 6515 13445 6645 13475
rect 6675 13445 6805 13475
rect 6835 13445 6965 13475
rect 6995 13445 7125 13475
rect 7155 13445 7285 13475
rect 7315 13445 7320 13475
rect 5520 13440 7320 13445
rect 7360 13475 7720 13480
rect 7360 13445 7365 13475
rect 7395 13445 7525 13475
rect 7555 13445 7685 13475
rect 7715 13445 7720 13475
rect 7360 13440 7720 13445
rect 5520 13395 7320 13400
rect 5520 13365 5525 13395
rect 5555 13365 5685 13395
rect 5715 13365 5845 13395
rect 5875 13365 6005 13395
rect 6035 13365 6165 13395
rect 6195 13365 6325 13395
rect 6355 13365 6485 13395
rect 6515 13365 6645 13395
rect 6675 13365 6805 13395
rect 6835 13365 6965 13395
rect 6995 13365 7125 13395
rect 7155 13365 7285 13395
rect 7315 13365 7320 13395
rect 5520 13360 7320 13365
rect 7360 13395 7720 13400
rect 7360 13365 7365 13395
rect 7395 13365 7525 13395
rect 7555 13365 7685 13395
rect 7715 13365 7720 13395
rect 7360 13360 7720 13365
rect 5520 13315 7320 13320
rect 5520 13285 5525 13315
rect 5555 13285 5685 13315
rect 5715 13285 5845 13315
rect 5875 13285 6005 13315
rect 6035 13285 6165 13315
rect 6195 13285 6325 13315
rect 6355 13285 6485 13315
rect 6515 13285 6645 13315
rect 6675 13285 6805 13315
rect 6835 13285 6965 13315
rect 6995 13285 7125 13315
rect 7155 13285 7285 13315
rect 7315 13285 7320 13315
rect 5520 13280 7320 13285
rect 7360 13315 7720 13320
rect 7360 13285 7365 13315
rect 7395 13285 7525 13315
rect 7555 13285 7685 13315
rect 7715 13285 7720 13315
rect 7360 13280 7720 13285
rect 5520 13235 7320 13240
rect 5520 13205 5525 13235
rect 5555 13205 5685 13235
rect 5715 13205 5845 13235
rect 5875 13205 6005 13235
rect 6035 13205 6165 13235
rect 6195 13205 6325 13235
rect 6355 13205 6485 13235
rect 6515 13205 6645 13235
rect 6675 13205 6805 13235
rect 6835 13205 6965 13235
rect 6995 13205 7125 13235
rect 7155 13205 7285 13235
rect 7315 13205 7320 13235
rect 5520 13200 7320 13205
rect 7360 13235 7720 13240
rect 7360 13205 7365 13235
rect 7395 13205 7525 13235
rect 7555 13205 7685 13235
rect 7715 13205 7720 13235
rect 7360 13200 7720 13205
rect 5480 13155 5960 13160
rect 5480 13125 5925 13155
rect 5955 13125 5960 13155
rect 5480 13120 5960 13125
rect 6000 13155 7320 13160
rect 6000 13125 6005 13155
rect 6035 13125 6165 13155
rect 6195 13125 6325 13155
rect 6355 13125 6485 13155
rect 6515 13125 6645 13155
rect 6675 13125 6805 13155
rect 6835 13125 6965 13155
rect 6995 13125 7125 13155
rect 7155 13125 7285 13155
rect 7315 13125 7320 13155
rect 6000 13120 7320 13125
rect 7360 13155 7720 13160
rect 7360 13125 7365 13155
rect 7395 13125 7525 13155
rect 7555 13125 7685 13155
rect 7715 13125 7720 13155
rect 7360 13120 7720 13125
rect 5520 13075 7320 13080
rect 5520 13045 5525 13075
rect 5555 13045 5685 13075
rect 5715 13045 5845 13075
rect 5875 13045 6005 13075
rect 6035 13045 6165 13075
rect 6195 13045 6325 13075
rect 6355 13045 6485 13075
rect 6515 13045 6645 13075
rect 6675 13045 6805 13075
rect 6835 13045 6965 13075
rect 6995 13045 7125 13075
rect 7155 13045 7285 13075
rect 7315 13045 7320 13075
rect 5520 13040 7320 13045
rect 7360 13075 7720 13080
rect 7360 13045 7365 13075
rect 7395 13045 7525 13075
rect 7555 13045 7685 13075
rect 7715 13045 7720 13075
rect 7360 13040 7720 13045
rect 5520 12995 7320 13000
rect 5520 12965 5525 12995
rect 5555 12965 5685 12995
rect 5715 12965 5845 12995
rect 5875 12965 6005 12995
rect 6035 12965 6165 12995
rect 6195 12965 6325 12995
rect 6355 12965 6485 12995
rect 6515 12965 6645 12995
rect 6675 12965 6805 12995
rect 6835 12965 6965 12995
rect 6995 12965 7125 12995
rect 7155 12965 7285 12995
rect 7315 12965 7320 12995
rect 5520 12960 7320 12965
rect 7360 12995 7720 13000
rect 7360 12965 7365 12995
rect 7395 12965 7525 12995
rect 7555 12965 7685 12995
rect 7715 12965 7720 12995
rect 7360 12960 7720 12965
rect 5520 12915 7720 12920
rect 5520 12885 7365 12915
rect 7395 12885 7525 12915
rect 7555 12885 7685 12915
rect 7715 12885 7720 12915
rect 5520 12880 7720 12885
rect 5480 12835 7640 12840
rect 5480 12805 7605 12835
rect 7635 12805 7640 12835
rect 5480 12800 7640 12805
rect 5480 12755 7720 12760
rect 5480 12725 7365 12755
rect 7395 12725 7525 12755
rect 7555 12725 7685 12755
rect 7715 12725 7720 12755
rect 5480 12720 7720 12725
rect 5480 12675 7480 12680
rect 5480 12645 7445 12675
rect 7475 12645 7480 12675
rect 5480 12640 7480 12645
rect 5520 12595 7720 12600
rect 5520 12565 7365 12595
rect 7395 12565 7525 12595
rect 7555 12565 7685 12595
rect 7715 12565 7720 12595
rect 5520 12560 7720 12565
rect 5520 12515 7320 12520
rect 5520 12485 5525 12515
rect 5555 12485 5685 12515
rect 5715 12485 5845 12515
rect 5875 12485 6005 12515
rect 6035 12485 6165 12515
rect 6195 12485 6325 12515
rect 6355 12485 6485 12515
rect 6515 12485 6645 12515
rect 6675 12485 6805 12515
rect 6835 12485 6965 12515
rect 6995 12485 7125 12515
rect 7155 12485 7285 12515
rect 7315 12485 7320 12515
rect 5520 12480 7320 12485
rect 7360 12475 7720 12480
rect 7360 12445 7365 12475
rect 7395 12445 7525 12475
rect 7555 12445 7685 12475
rect 7715 12445 7720 12475
rect 7360 12440 7720 12445
rect 5480 12435 5800 12440
rect 5480 12405 5765 12435
rect 5795 12405 5800 12435
rect 5480 12400 5800 12405
rect 5840 12435 7320 12440
rect 5840 12405 5845 12435
rect 5875 12405 6005 12435
rect 6035 12405 6165 12435
rect 6195 12405 6325 12435
rect 6355 12405 6485 12435
rect 6515 12405 6645 12435
rect 6675 12405 6805 12435
rect 6835 12405 6965 12435
rect 6995 12405 7125 12435
rect 7155 12405 7285 12435
rect 7315 12405 7320 12435
rect 5840 12400 7320 12405
rect 7360 12395 7720 12400
rect 7360 12365 7365 12395
rect 7395 12365 7525 12395
rect 7555 12365 7685 12395
rect 7715 12365 7720 12395
rect 7360 12360 7720 12365
rect 5520 12315 7320 12320
rect 5520 12285 5525 12315
rect 5555 12285 5685 12315
rect 5715 12285 5845 12315
rect 5875 12285 6005 12315
rect 6035 12285 6165 12315
rect 6195 12285 6325 12315
rect 6355 12285 6485 12315
rect 6515 12285 6645 12315
rect 6675 12285 6805 12315
rect 6835 12285 6965 12315
rect 6995 12285 7125 12315
rect 7155 12285 7285 12315
rect 7315 12285 7320 12315
rect 5520 12280 7320 12285
rect 7360 12315 7720 12320
rect 7360 12285 7365 12315
rect 7395 12285 7525 12315
rect 7555 12285 7685 12315
rect 7715 12285 7720 12315
rect 7360 12280 7720 12285
rect 5520 12235 7320 12240
rect 5520 12205 5525 12235
rect 5555 12205 5685 12235
rect 5715 12205 5845 12235
rect 5875 12205 6005 12235
rect 6035 12205 6165 12235
rect 6195 12205 6325 12235
rect 6355 12205 6485 12235
rect 6515 12205 6645 12235
rect 6675 12205 6805 12235
rect 6835 12205 6965 12235
rect 6995 12205 7125 12235
rect 7155 12205 7285 12235
rect 7315 12205 7320 12235
rect 5520 12200 7320 12205
rect 7360 12235 7720 12240
rect 7360 12205 7365 12235
rect 7395 12205 7525 12235
rect 7555 12205 7685 12235
rect 7715 12205 7720 12235
rect 7360 12200 7720 12205
rect 5520 12155 7320 12160
rect 5520 12125 5525 12155
rect 5555 12125 5685 12155
rect 5715 12125 5845 12155
rect 5875 12125 6005 12155
rect 6035 12125 6165 12155
rect 6195 12125 6325 12155
rect 6355 12125 6485 12155
rect 6515 12125 6645 12155
rect 6675 12125 6805 12155
rect 6835 12125 6965 12155
rect 6995 12125 7125 12155
rect 7155 12125 7285 12155
rect 7315 12125 7320 12155
rect 5520 12120 7320 12125
rect 7360 12155 7720 12160
rect 7360 12125 7365 12155
rect 7395 12125 7525 12155
rect 7555 12125 7685 12155
rect 7715 12125 7720 12155
rect 7360 12120 7720 12125
rect 5520 12075 7320 12080
rect 5520 12045 5525 12075
rect 5555 12045 5685 12075
rect 5715 12045 5845 12075
rect 5875 12045 6005 12075
rect 6035 12045 6165 12075
rect 6195 12045 6325 12075
rect 6355 12045 6485 12075
rect 6515 12045 6645 12075
rect 6675 12045 6805 12075
rect 6835 12045 6965 12075
rect 6995 12045 7125 12075
rect 7155 12045 7285 12075
rect 7315 12045 7320 12075
rect 5520 12040 7320 12045
rect 7360 12075 7720 12080
rect 7360 12045 7365 12075
rect 7395 12045 7525 12075
rect 7555 12045 7685 12075
rect 7715 12045 7720 12075
rect 7360 12040 7720 12045
rect 5520 11995 7320 12000
rect 5520 11965 5525 11995
rect 5555 11965 5685 11995
rect 5715 11965 5845 11995
rect 5875 11965 6005 11995
rect 6035 11965 6165 11995
rect 6195 11965 6325 11995
rect 6355 11965 6485 11995
rect 6515 11965 6645 11995
rect 6675 11965 6805 11995
rect 6835 11965 6965 11995
rect 6995 11965 7125 11995
rect 7155 11965 7285 11995
rect 7315 11965 7320 11995
rect 5520 11960 7320 11965
rect 7360 11995 7720 12000
rect 7360 11965 7365 11995
rect 7395 11965 7525 11995
rect 7555 11965 7685 11995
rect 7715 11965 7720 11995
rect 7360 11960 7720 11965
rect 5520 11915 7320 11920
rect 5520 11885 5525 11915
rect 5555 11885 5685 11915
rect 5715 11885 5845 11915
rect 5875 11885 6005 11915
rect 6035 11885 6165 11915
rect 6195 11885 6325 11915
rect 6355 11885 6485 11915
rect 6515 11885 6645 11915
rect 6675 11885 6805 11915
rect 6835 11885 6965 11915
rect 6995 11885 7125 11915
rect 7155 11885 7285 11915
rect 7315 11885 7320 11915
rect 5520 11880 7320 11885
rect 7360 11915 7720 11920
rect 7360 11885 7365 11915
rect 7395 11885 7525 11915
rect 7555 11885 7685 11915
rect 7715 11885 7720 11915
rect 7360 11880 7720 11885
rect 5520 11835 7320 11840
rect 5520 11805 5525 11835
rect 5555 11805 5685 11835
rect 5715 11805 5845 11835
rect 5875 11805 6005 11835
rect 6035 11805 6165 11835
rect 6195 11805 6325 11835
rect 6355 11805 6485 11835
rect 6515 11805 6645 11835
rect 6675 11805 6805 11835
rect 6835 11805 6965 11835
rect 6995 11805 7125 11835
rect 7155 11805 7285 11835
rect 7315 11805 7320 11835
rect 5520 11800 7320 11805
rect 7360 11835 7720 11840
rect 7360 11805 7365 11835
rect 7395 11805 7525 11835
rect 7555 11805 7685 11835
rect 7715 11805 7720 11835
rect 7360 11800 7720 11805
rect 5520 11755 7320 11760
rect 5520 11725 5525 11755
rect 5555 11725 5685 11755
rect 5715 11725 5845 11755
rect 5875 11725 6005 11755
rect 6035 11725 6165 11755
rect 6195 11725 6325 11755
rect 6355 11725 6485 11755
rect 6515 11725 6645 11755
rect 6675 11725 6805 11755
rect 6835 11725 6965 11755
rect 6995 11725 7125 11755
rect 7155 11725 7285 11755
rect 7315 11725 7320 11755
rect 5520 11720 7320 11725
rect 7360 11755 7720 11760
rect 7360 11725 7365 11755
rect 7395 11725 7525 11755
rect 7555 11725 7685 11755
rect 7715 11725 7720 11755
rect 7360 11720 7720 11725
rect 5520 11675 7320 11680
rect 5520 11645 5525 11675
rect 5555 11645 5685 11675
rect 5715 11645 5845 11675
rect 5875 11645 6005 11675
rect 6035 11645 6165 11675
rect 6195 11645 6325 11675
rect 6355 11645 6485 11675
rect 6515 11645 6645 11675
rect 6675 11645 6805 11675
rect 6835 11645 6965 11675
rect 6995 11645 7125 11675
rect 7155 11645 7285 11675
rect 7315 11645 7320 11675
rect 5520 11640 7320 11645
rect 7360 11675 7720 11680
rect 7360 11645 7365 11675
rect 7395 11645 7525 11675
rect 7555 11645 7685 11675
rect 7715 11645 7720 11675
rect 7360 11640 7720 11645
rect 5520 11595 7320 11600
rect 5520 11565 5525 11595
rect 5555 11565 5685 11595
rect 5715 11565 5845 11595
rect 5875 11565 6005 11595
rect 6035 11565 6165 11595
rect 6195 11565 6325 11595
rect 6355 11565 6485 11595
rect 6515 11565 6645 11595
rect 6675 11565 6805 11595
rect 6835 11565 6965 11595
rect 6995 11565 7125 11595
rect 7155 11565 7285 11595
rect 7315 11565 7320 11595
rect 5520 11560 7320 11565
rect 7360 11595 7720 11600
rect 7360 11565 7365 11595
rect 7395 11565 7525 11595
rect 7555 11565 7685 11595
rect 7715 11565 7720 11595
rect 7360 11560 7720 11565
rect 5520 11515 7320 11520
rect 5520 11485 5525 11515
rect 5555 11485 5685 11515
rect 5715 11485 5845 11515
rect 5875 11485 6005 11515
rect 6035 11485 6165 11515
rect 6195 11485 6325 11515
rect 6355 11485 6485 11515
rect 6515 11485 6645 11515
rect 6675 11485 6805 11515
rect 6835 11485 6965 11515
rect 6995 11485 7125 11515
rect 7155 11485 7285 11515
rect 7315 11485 7320 11515
rect 5520 11480 7320 11485
rect 7360 11515 7720 11520
rect 7360 11485 7365 11515
rect 7395 11485 7525 11515
rect 7555 11485 7685 11515
rect 7715 11485 7720 11515
rect 7360 11480 7720 11485
rect 5520 11435 7320 11440
rect 5520 11405 5525 11435
rect 5555 11405 5685 11435
rect 5715 11405 5845 11435
rect 5875 11405 6005 11435
rect 6035 11405 6165 11435
rect 6195 11405 6325 11435
rect 6355 11405 6485 11435
rect 6515 11405 6645 11435
rect 6675 11405 6805 11435
rect 6835 11405 6965 11435
rect 6995 11405 7125 11435
rect 7155 11405 7285 11435
rect 7315 11405 7320 11435
rect 5520 11400 7320 11405
rect 7360 11435 7720 11440
rect 7360 11405 7365 11435
rect 7395 11405 7525 11435
rect 7555 11405 7685 11435
rect 7715 11405 7720 11435
rect 7360 11400 7720 11405
rect 5520 11355 7320 11360
rect 5520 11325 5525 11355
rect 5555 11325 5685 11355
rect 5715 11325 5845 11355
rect 5875 11325 6005 11355
rect 6035 11325 6165 11355
rect 6195 11325 6325 11355
rect 6355 11325 6485 11355
rect 6515 11325 6645 11355
rect 6675 11325 6805 11355
rect 6835 11325 6965 11355
rect 6995 11325 7125 11355
rect 7155 11325 7285 11355
rect 7315 11325 7320 11355
rect 5520 11320 7320 11325
rect 7360 11355 7720 11360
rect 7360 11325 7365 11355
rect 7395 11325 7525 11355
rect 7555 11325 7685 11355
rect 7715 11325 7720 11355
rect 7360 11320 7720 11325
rect 5480 11275 7240 11280
rect 5480 11245 7205 11275
rect 7235 11245 7240 11275
rect 5480 11240 7240 11245
rect 7360 11275 7720 11280
rect 7360 11245 7365 11275
rect 7395 11245 7525 11275
rect 7555 11245 7685 11275
rect 7715 11245 7720 11275
rect 7360 11240 7720 11245
rect 5520 11195 7320 11200
rect 5520 11165 5525 11195
rect 5555 11165 5685 11195
rect 5715 11165 5845 11195
rect 5875 11165 6005 11195
rect 6035 11165 6165 11195
rect 6195 11165 6325 11195
rect 6355 11165 6485 11195
rect 6515 11165 6645 11195
rect 6675 11165 6805 11195
rect 6835 11165 6965 11195
rect 6995 11165 7125 11195
rect 7155 11165 7285 11195
rect 7315 11165 7320 11195
rect 5520 11160 7320 11165
rect 7360 11195 7720 11200
rect 7360 11165 7365 11195
rect 7395 11165 7525 11195
rect 7555 11165 7685 11195
rect 7715 11165 7720 11195
rect 7360 11160 7720 11165
rect 5520 11115 7320 11120
rect 5520 11085 5525 11115
rect 5555 11085 5685 11115
rect 5715 11085 5845 11115
rect 5875 11085 6005 11115
rect 6035 11085 6165 11115
rect 6195 11085 6325 11115
rect 6355 11085 6485 11115
rect 6515 11085 6645 11115
rect 6675 11085 6805 11115
rect 6835 11085 6965 11115
rect 6995 11085 7125 11115
rect 7155 11085 7285 11115
rect 7315 11085 7320 11115
rect 5520 11080 7320 11085
rect 7360 11115 7720 11120
rect 7360 11085 7365 11115
rect 7395 11085 7525 11115
rect 7555 11085 7685 11115
rect 7715 11085 7720 11115
rect 7360 11080 7720 11085
rect 5520 11035 7320 11040
rect 5520 11005 5525 11035
rect 5555 11005 5685 11035
rect 5715 11005 5845 11035
rect 5875 11005 6005 11035
rect 6035 11005 6165 11035
rect 6195 11005 6325 11035
rect 6355 11005 6485 11035
rect 6515 11005 6645 11035
rect 6675 11005 6805 11035
rect 6835 11005 6965 11035
rect 6995 11005 7125 11035
rect 7155 11005 7285 11035
rect 7315 11005 7320 11035
rect 5520 11000 7320 11005
rect 7360 11035 7720 11040
rect 7360 11005 7365 11035
rect 7395 11005 7525 11035
rect 7555 11005 7685 11035
rect 7715 11005 7720 11035
rect 7360 11000 7720 11005
rect 5480 10955 7240 10960
rect 5480 10925 7205 10955
rect 7235 10925 7240 10955
rect 5480 10920 7240 10925
rect 7360 10955 7720 10960
rect 7360 10925 7365 10955
rect 7395 10925 7525 10955
rect 7555 10925 7685 10955
rect 7715 10925 7720 10955
rect 7360 10920 7720 10925
rect 5480 10875 7320 10880
rect 5480 10845 5525 10875
rect 5555 10845 5685 10875
rect 5715 10845 5845 10875
rect 5875 10845 6005 10875
rect 6035 10845 6165 10875
rect 6195 10845 6325 10875
rect 6355 10845 6485 10875
rect 6515 10845 6645 10875
rect 6675 10845 6805 10875
rect 6835 10845 6965 10875
rect 6995 10845 7125 10875
rect 7155 10845 7285 10875
rect 7315 10845 7320 10875
rect 5480 10840 7320 10845
rect 7360 10875 7720 10880
rect 7360 10845 7365 10875
rect 7395 10845 7525 10875
rect 7555 10845 7685 10875
rect 7715 10845 7720 10875
rect 7360 10840 7720 10845
rect 5480 10795 7080 10800
rect 5480 10765 7045 10795
rect 7075 10765 7080 10795
rect 5480 10760 7080 10765
rect 7120 10795 7320 10800
rect 7120 10765 7125 10795
rect 7155 10765 7285 10795
rect 7315 10765 7320 10795
rect 7120 10760 7320 10765
rect 7360 10795 7720 10800
rect 7360 10765 7365 10795
rect 7395 10765 7525 10795
rect 7555 10765 7685 10795
rect 7715 10765 7720 10795
rect 7360 10760 7720 10765
rect 5520 10715 7320 10720
rect 5520 10685 5525 10715
rect 5555 10685 5685 10715
rect 5715 10685 5845 10715
rect 5875 10685 6005 10715
rect 6035 10685 6165 10715
rect 6195 10685 6325 10715
rect 6355 10685 6485 10715
rect 6515 10685 6645 10715
rect 6675 10685 6805 10715
rect 6835 10685 6965 10715
rect 6995 10685 7125 10715
rect 7155 10685 7285 10715
rect 7315 10685 7320 10715
rect 5520 10680 7320 10685
rect 7360 10715 7720 10720
rect 7360 10685 7365 10715
rect 7395 10685 7525 10715
rect 7555 10685 7685 10715
rect 7715 10685 7720 10715
rect 7360 10680 7720 10685
rect 5520 10635 7320 10640
rect 5520 10605 5525 10635
rect 5555 10605 5685 10635
rect 5715 10605 5845 10635
rect 5875 10605 6005 10635
rect 6035 10605 6165 10635
rect 6195 10605 6325 10635
rect 6355 10605 6485 10635
rect 6515 10605 6645 10635
rect 6675 10605 6805 10635
rect 6835 10605 6965 10635
rect 6995 10605 7125 10635
rect 7155 10605 7285 10635
rect 7315 10605 7320 10635
rect 5520 10600 7320 10605
rect 7360 10635 7720 10640
rect 7360 10605 7365 10635
rect 7395 10605 7525 10635
rect 7555 10605 7685 10635
rect 7715 10605 7720 10635
rect 7360 10600 7720 10605
rect 5480 10555 7080 10560
rect 5480 10525 7045 10555
rect 7075 10525 7080 10555
rect 5480 10520 7080 10525
rect 7120 10555 7320 10560
rect 7120 10525 7125 10555
rect 7155 10525 7285 10555
rect 7315 10525 7320 10555
rect 7120 10520 7320 10525
rect 7360 10555 7720 10560
rect 7360 10525 7365 10555
rect 7395 10525 7525 10555
rect 7555 10525 7685 10555
rect 7715 10525 7720 10555
rect 7360 10520 7720 10525
rect 5520 10475 7320 10480
rect 5520 10445 5525 10475
rect 5555 10445 5685 10475
rect 5715 10445 5845 10475
rect 5875 10445 6005 10475
rect 6035 10445 6165 10475
rect 6195 10445 6325 10475
rect 6355 10445 6485 10475
rect 6515 10445 6645 10475
rect 6675 10445 6805 10475
rect 6835 10445 6965 10475
rect 6995 10445 7125 10475
rect 7155 10445 7285 10475
rect 7315 10445 7320 10475
rect 5520 10440 7320 10445
rect 7360 10475 7720 10480
rect 7360 10445 7365 10475
rect 7395 10445 7525 10475
rect 7555 10445 7685 10475
rect 7715 10445 7720 10475
rect 7360 10440 7720 10445
rect 5480 10395 6920 10400
rect 5480 10365 6885 10395
rect 6915 10365 6920 10395
rect 5480 10360 6920 10365
rect 6960 10395 7320 10400
rect 6960 10365 6965 10395
rect 6995 10365 7125 10395
rect 7155 10365 7285 10395
rect 7315 10365 7320 10395
rect 6960 10360 7320 10365
rect 7360 10395 7720 10400
rect 7360 10365 7365 10395
rect 7395 10365 7525 10395
rect 7555 10365 7685 10395
rect 7715 10365 7720 10395
rect 7360 10360 7720 10365
rect 5520 10315 7320 10320
rect 5520 10285 5525 10315
rect 5555 10285 5685 10315
rect 5715 10285 5845 10315
rect 5875 10285 6005 10315
rect 6035 10285 6165 10315
rect 6195 10285 6325 10315
rect 6355 10285 6485 10315
rect 6515 10285 6645 10315
rect 6675 10285 6805 10315
rect 6835 10285 6965 10315
rect 6995 10285 7125 10315
rect 7155 10285 7285 10315
rect 7315 10285 7320 10315
rect 5520 10280 7320 10285
rect 7360 10315 7720 10320
rect 7360 10285 7365 10315
rect 7395 10285 7525 10315
rect 7555 10285 7685 10315
rect 7715 10285 7720 10315
rect 7360 10280 7720 10285
rect 5520 10235 7320 10240
rect 5520 10205 5525 10235
rect 5555 10205 5685 10235
rect 5715 10205 5845 10235
rect 5875 10205 6005 10235
rect 6035 10205 6165 10235
rect 6195 10205 6325 10235
rect 6355 10205 6485 10235
rect 6515 10205 6645 10235
rect 6675 10205 6805 10235
rect 6835 10205 6965 10235
rect 6995 10205 7125 10235
rect 7155 10205 7285 10235
rect 7315 10205 7320 10235
rect 5520 10200 7320 10205
rect 7360 10235 7720 10240
rect 7360 10205 7365 10235
rect 7395 10205 7525 10235
rect 7555 10205 7685 10235
rect 7715 10205 7720 10235
rect 7360 10200 7720 10205
rect 5520 10155 7320 10160
rect 5520 10125 5525 10155
rect 5555 10125 5685 10155
rect 5715 10125 5845 10155
rect 5875 10125 6005 10155
rect 6035 10125 6165 10155
rect 6195 10125 6325 10155
rect 6355 10125 6485 10155
rect 6515 10125 6645 10155
rect 6675 10125 6805 10155
rect 6835 10125 6965 10155
rect 6995 10125 7125 10155
rect 7155 10125 7285 10155
rect 7315 10125 7320 10155
rect 5520 10120 7320 10125
rect 7360 10155 7720 10160
rect 7360 10125 7365 10155
rect 7395 10125 7525 10155
rect 7555 10125 7685 10155
rect 7715 10125 7720 10155
rect 7360 10120 7720 10125
rect 5520 10075 7320 10080
rect 5520 10045 5525 10075
rect 5555 10045 5685 10075
rect 5715 10045 5845 10075
rect 5875 10045 6005 10075
rect 6035 10045 6165 10075
rect 6195 10045 6325 10075
rect 6355 10045 6485 10075
rect 6515 10045 6645 10075
rect 6675 10045 6805 10075
rect 6835 10045 6965 10075
rect 6995 10045 7125 10075
rect 7155 10045 7285 10075
rect 7315 10045 7320 10075
rect 5520 10040 7320 10045
rect 7360 10075 7720 10080
rect 7360 10045 7365 10075
rect 7395 10045 7525 10075
rect 7555 10045 7685 10075
rect 7715 10045 7720 10075
rect 7360 10040 7720 10045
rect 5520 9995 7320 10000
rect 5520 9965 5525 9995
rect 5555 9965 5685 9995
rect 5715 9965 5845 9995
rect 5875 9965 6005 9995
rect 6035 9965 6165 9995
rect 6195 9965 6325 9995
rect 6355 9965 6485 9995
rect 6515 9965 6645 9995
rect 6675 9965 6805 9995
rect 6835 9965 6965 9995
rect 6995 9965 7125 9995
rect 7155 9965 7285 9995
rect 7315 9965 7320 9995
rect 5520 9960 7320 9965
rect 7360 9995 7720 10000
rect 7360 9965 7365 9995
rect 7395 9965 7525 9995
rect 7555 9965 7685 9995
rect 7715 9965 7720 9995
rect 7360 9960 7720 9965
rect 5520 9915 7320 9920
rect 5520 9885 5525 9915
rect 5555 9885 5685 9915
rect 5715 9885 5845 9915
rect 5875 9885 6005 9915
rect 6035 9885 6165 9915
rect 6195 9885 6325 9915
rect 6355 9885 6485 9915
rect 6515 9885 6645 9915
rect 6675 9885 6805 9915
rect 6835 9885 6965 9915
rect 6995 9885 7125 9915
rect 7155 9885 7285 9915
rect 7315 9885 7320 9915
rect 5520 9880 7320 9885
rect 7360 9915 7720 9920
rect 7360 9885 7365 9915
rect 7395 9885 7525 9915
rect 7555 9885 7685 9915
rect 7715 9885 7720 9915
rect 7360 9880 7720 9885
rect 5520 9835 7320 9840
rect 5520 9805 5525 9835
rect 5555 9805 5685 9835
rect 5715 9805 5845 9835
rect 5875 9805 6005 9835
rect 6035 9805 6165 9835
rect 6195 9805 6325 9835
rect 6355 9805 6485 9835
rect 6515 9805 6645 9835
rect 6675 9805 6805 9835
rect 6835 9805 6965 9835
rect 6995 9805 7125 9835
rect 7155 9805 7285 9835
rect 7315 9805 7320 9835
rect 5520 9800 7320 9805
rect 7360 9835 7720 9840
rect 7360 9805 7365 9835
rect 7395 9805 7525 9835
rect 7555 9805 7685 9835
rect 7715 9805 7720 9835
rect 7360 9800 7720 9805
rect 5520 9755 7320 9760
rect 5520 9725 5525 9755
rect 5555 9725 5685 9755
rect 5715 9725 5845 9755
rect 5875 9725 6005 9755
rect 6035 9725 6165 9755
rect 6195 9725 6325 9755
rect 6355 9725 6485 9755
rect 6515 9725 6645 9755
rect 6675 9725 6805 9755
rect 6835 9725 6965 9755
rect 6995 9725 7125 9755
rect 7155 9725 7285 9755
rect 7315 9725 7320 9755
rect 5520 9720 7320 9725
rect 7360 9755 7720 9760
rect 7360 9725 7365 9755
rect 7395 9725 7525 9755
rect 7555 9725 7685 9755
rect 7715 9725 7720 9755
rect 7360 9720 7720 9725
rect 5520 9675 7320 9680
rect 5520 9645 5525 9675
rect 5555 9645 5685 9675
rect 5715 9645 5845 9675
rect 5875 9645 6005 9675
rect 6035 9645 6165 9675
rect 6195 9645 6325 9675
rect 6355 9645 6485 9675
rect 6515 9645 6645 9675
rect 6675 9645 6805 9675
rect 6835 9645 6965 9675
rect 6995 9645 7125 9675
rect 7155 9645 7285 9675
rect 7315 9645 7320 9675
rect 5520 9640 7320 9645
rect 7360 9675 7720 9680
rect 7360 9645 7365 9675
rect 7395 9645 7525 9675
rect 7555 9645 7685 9675
rect 7715 9645 7720 9675
rect 7360 9640 7720 9645
rect 5520 9595 7320 9600
rect 5520 9565 5525 9595
rect 5555 9565 5685 9595
rect 5715 9565 5845 9595
rect 5875 9565 6005 9595
rect 6035 9565 6165 9595
rect 6195 9565 6325 9595
rect 6355 9565 6485 9595
rect 6515 9565 6645 9595
rect 6675 9565 6805 9595
rect 6835 9565 6965 9595
rect 6995 9565 7125 9595
rect 7155 9565 7285 9595
rect 7315 9565 7320 9595
rect 5520 9560 7320 9565
rect 7360 9595 7720 9600
rect 7360 9565 7365 9595
rect 7395 9565 7525 9595
rect 7555 9565 7685 9595
rect 7715 9565 7720 9595
rect 7360 9560 7720 9565
rect 5520 9515 7320 9520
rect 5520 9485 5525 9515
rect 5555 9485 5685 9515
rect 5715 9485 5845 9515
rect 5875 9485 6005 9515
rect 6035 9485 6165 9515
rect 6195 9485 6325 9515
rect 6355 9485 6485 9515
rect 6515 9485 6645 9515
rect 6675 9485 6805 9515
rect 6835 9485 6965 9515
rect 6995 9485 7125 9515
rect 7155 9485 7285 9515
rect 7315 9485 7320 9515
rect 5520 9480 7320 9485
rect 7360 9515 7720 9520
rect 7360 9485 7365 9515
rect 7395 9485 7525 9515
rect 7555 9485 7685 9515
rect 7715 9485 7720 9515
rect 7360 9480 7720 9485
rect 5520 9435 7320 9440
rect 5520 9405 5525 9435
rect 5555 9405 5685 9435
rect 5715 9405 5845 9435
rect 5875 9405 6005 9435
rect 6035 9405 6165 9435
rect 6195 9405 6325 9435
rect 6355 9405 6485 9435
rect 6515 9405 6645 9435
rect 6675 9405 6805 9435
rect 6835 9405 6965 9435
rect 6995 9405 7125 9435
rect 7155 9405 7285 9435
rect 7315 9405 7320 9435
rect 5520 9400 7320 9405
rect 7360 9435 7720 9440
rect 7360 9405 7365 9435
rect 7395 9405 7525 9435
rect 7555 9405 7685 9435
rect 7715 9405 7720 9435
rect 7360 9400 7720 9405
rect 5520 9355 7320 9360
rect 5520 9325 5525 9355
rect 5555 9325 5685 9355
rect 5715 9325 5845 9355
rect 5875 9325 6005 9355
rect 6035 9325 6165 9355
rect 6195 9325 6325 9355
rect 6355 9325 6485 9355
rect 6515 9325 6645 9355
rect 6675 9325 6805 9355
rect 6835 9325 6965 9355
rect 6995 9325 7125 9355
rect 7155 9325 7285 9355
rect 7315 9325 7320 9355
rect 5520 9320 7320 9325
rect 7360 9355 7720 9360
rect 7360 9325 7365 9355
rect 7395 9325 7525 9355
rect 7555 9325 7685 9355
rect 7715 9325 7720 9355
rect 7360 9320 7720 9325
rect 5520 9275 7320 9280
rect 5520 9245 5525 9275
rect 5555 9245 5685 9275
rect 5715 9245 5845 9275
rect 5875 9245 6005 9275
rect 6035 9245 6165 9275
rect 6195 9245 6325 9275
rect 6355 9245 6485 9275
rect 6515 9245 6645 9275
rect 6675 9245 6805 9275
rect 6835 9245 6965 9275
rect 6995 9245 7125 9275
rect 7155 9245 7285 9275
rect 7315 9245 7320 9275
rect 5520 9240 7320 9245
rect 7360 9275 7720 9280
rect 7360 9245 7365 9275
rect 7395 9245 7525 9275
rect 7555 9245 7685 9275
rect 7715 9245 7720 9275
rect 7360 9240 7720 9245
rect 5480 9195 7240 9200
rect 5480 9165 7205 9195
rect 7235 9165 7240 9195
rect 5480 9160 7240 9165
rect 7360 9195 7720 9200
rect 7360 9165 7365 9195
rect 7395 9165 7525 9195
rect 7555 9165 7685 9195
rect 7715 9165 7720 9195
rect 7360 9160 7720 9165
rect 5520 9115 7320 9120
rect 5520 9085 5525 9115
rect 5555 9085 5685 9115
rect 5715 9085 5845 9115
rect 5875 9085 6005 9115
rect 6035 9085 6165 9115
rect 6195 9085 6325 9115
rect 6355 9085 6485 9115
rect 6515 9085 6645 9115
rect 6675 9085 6805 9115
rect 6835 9085 6965 9115
rect 6995 9085 7125 9115
rect 7155 9085 7285 9115
rect 7315 9085 7320 9115
rect 5520 9080 7320 9085
rect 7360 9115 7720 9120
rect 7360 9085 7365 9115
rect 7395 9085 7525 9115
rect 7555 9085 7685 9115
rect 7715 9085 7720 9115
rect 7360 9080 7720 9085
rect 5520 9035 7320 9040
rect 5520 9005 5525 9035
rect 5555 9005 5685 9035
rect 5715 9005 5845 9035
rect 5875 9005 6005 9035
rect 6035 9005 6165 9035
rect 6195 9005 6325 9035
rect 6355 9005 6485 9035
rect 6515 9005 6645 9035
rect 6675 9005 6805 9035
rect 6835 9005 6965 9035
rect 6995 9005 7125 9035
rect 7155 9005 7285 9035
rect 7315 9005 7320 9035
rect 5520 9000 7320 9005
rect 7360 9035 7720 9040
rect 7360 9005 7365 9035
rect 7395 9005 7525 9035
rect 7555 9005 7685 9035
rect 7715 9005 7720 9035
rect 7360 9000 7720 9005
rect 5520 8955 7320 8960
rect 5520 8925 5525 8955
rect 5555 8925 5685 8955
rect 5715 8925 5845 8955
rect 5875 8925 6005 8955
rect 6035 8925 6165 8955
rect 6195 8925 6325 8955
rect 6355 8925 6485 8955
rect 6515 8925 6645 8955
rect 6675 8925 6805 8955
rect 6835 8925 6965 8955
rect 6995 8925 7125 8955
rect 7155 8925 7285 8955
rect 7315 8925 7320 8955
rect 5520 8920 7320 8925
rect 7360 8955 7720 8960
rect 7360 8925 7365 8955
rect 7395 8925 7525 8955
rect 7555 8925 7685 8955
rect 7715 8925 7720 8955
rect 7360 8920 7720 8925
rect 5480 8875 7640 8880
rect 5480 8845 7605 8875
rect 7635 8845 7640 8875
rect 5480 8840 7640 8845
rect 5480 8795 7720 8800
rect 5480 8765 7365 8795
rect 7395 8765 7525 8795
rect 7555 8765 7685 8795
rect 7715 8765 7720 8795
rect 5480 8760 7720 8765
rect 5480 8715 7480 8720
rect 5480 8685 7445 8715
rect 7475 8685 7480 8715
rect 5480 8680 7480 8685
rect 5520 8635 7320 8640
rect 5520 8605 5525 8635
rect 5555 8605 5685 8635
rect 5715 8605 5845 8635
rect 5875 8605 6005 8635
rect 6035 8605 6165 8635
rect 6195 8605 6325 8635
rect 6355 8605 6485 8635
rect 6515 8605 6645 8635
rect 6675 8605 6805 8635
rect 6835 8605 6965 8635
rect 6995 8605 7125 8635
rect 7155 8605 7285 8635
rect 7315 8605 7320 8635
rect 5520 8600 7320 8605
rect 7360 8635 7720 8640
rect 7360 8605 7365 8635
rect 7395 8605 7525 8635
rect 7555 8605 7685 8635
rect 7715 8605 7720 8635
rect 7360 8600 7720 8605
rect 5520 8555 7320 8560
rect 5520 8525 5525 8555
rect 5555 8525 5685 8555
rect 5715 8525 5845 8555
rect 5875 8525 6005 8555
rect 6035 8525 6165 8555
rect 6195 8525 6325 8555
rect 6355 8525 6485 8555
rect 6515 8525 6645 8555
rect 6675 8525 6805 8555
rect 6835 8525 6965 8555
rect 6995 8525 7125 8555
rect 7155 8525 7285 8555
rect 7315 8525 7320 8555
rect 5520 8520 7320 8525
rect 7360 8555 7720 8560
rect 7360 8525 7365 8555
rect 7395 8525 7525 8555
rect 7555 8525 7685 8555
rect 7715 8525 7720 8555
rect 7360 8520 7720 8525
rect 5480 8475 7080 8480
rect 5480 8445 7045 8475
rect 7075 8445 7080 8475
rect 5480 8440 7080 8445
rect 7120 8475 7320 8480
rect 7120 8445 7125 8475
rect 7155 8445 7285 8475
rect 7315 8445 7320 8475
rect 7120 8440 7320 8445
rect 7360 8475 7720 8480
rect 7360 8445 7365 8475
rect 7395 8445 7525 8475
rect 7555 8445 7685 8475
rect 7715 8445 7720 8475
rect 7360 8440 7720 8445
rect 5520 8395 7320 8400
rect 5520 8365 5525 8395
rect 5555 8365 5685 8395
rect 5715 8365 5845 8395
rect 5875 8365 6005 8395
rect 6035 8365 6165 8395
rect 6195 8365 6325 8395
rect 6355 8365 6485 8395
rect 6515 8365 6645 8395
rect 6675 8365 6805 8395
rect 6835 8365 6965 8395
rect 6995 8365 7125 8395
rect 7155 8365 7285 8395
rect 7315 8365 7320 8395
rect 5520 8360 7320 8365
rect 7360 8395 7720 8400
rect 7360 8365 7365 8395
rect 7395 8365 7525 8395
rect 7555 8365 7685 8395
rect 7715 8365 7720 8395
rect 7360 8360 7720 8365
rect 5480 8315 6760 8320
rect 5480 8285 6725 8315
rect 6755 8285 6760 8315
rect 5480 8280 6760 8285
rect 6800 8315 7320 8320
rect 6800 8285 6805 8315
rect 6835 8285 6965 8315
rect 6995 8285 7125 8315
rect 7155 8285 7285 8315
rect 7315 8285 7320 8315
rect 6800 8280 7320 8285
rect 7360 8315 7720 8320
rect 7360 8285 7365 8315
rect 7395 8285 7525 8315
rect 7555 8285 7685 8315
rect 7715 8285 7720 8315
rect 7360 8280 7720 8285
rect 5520 8235 7320 8240
rect 5520 8205 5525 8235
rect 5555 8205 5685 8235
rect 5715 8205 5845 8235
rect 5875 8205 6005 8235
rect 6035 8205 6165 8235
rect 6195 8205 6325 8235
rect 6355 8205 6485 8235
rect 6515 8205 6645 8235
rect 6675 8205 6805 8235
rect 6835 8205 6965 8235
rect 6995 8205 7125 8235
rect 7155 8205 7285 8235
rect 7315 8205 7320 8235
rect 5520 8200 7320 8205
rect 7360 8235 7720 8240
rect 7360 8205 7365 8235
rect 7395 8205 7525 8235
rect 7555 8205 7685 8235
rect 7715 8205 7720 8235
rect 7360 8200 7720 8205
rect 5520 8155 7320 8160
rect 5520 8125 5525 8155
rect 5555 8125 5685 8155
rect 5715 8125 5845 8155
rect 5875 8125 6005 8155
rect 6035 8125 6165 8155
rect 6195 8125 6325 8155
rect 6355 8125 6485 8155
rect 6515 8125 6645 8155
rect 6675 8125 6805 8155
rect 6835 8125 6965 8155
rect 6995 8125 7125 8155
rect 7155 8125 7285 8155
rect 7315 8125 7320 8155
rect 5520 8120 7320 8125
rect 7360 8155 7720 8160
rect 7360 8125 7365 8155
rect 7395 8125 7525 8155
rect 7555 8125 7685 8155
rect 7715 8125 7720 8155
rect 7360 8120 7720 8125
rect 5520 8075 7320 8080
rect 5520 8045 5525 8075
rect 5555 8045 5685 8075
rect 5715 8045 5845 8075
rect 5875 8045 6005 8075
rect 6035 8045 6165 8075
rect 6195 8045 6325 8075
rect 6355 8045 6485 8075
rect 6515 8045 6645 8075
rect 6675 8045 6805 8075
rect 6835 8045 6965 8075
rect 6995 8045 7125 8075
rect 7155 8045 7285 8075
rect 7315 8045 7320 8075
rect 5520 8040 7320 8045
rect 7360 8075 7720 8080
rect 7360 8045 7365 8075
rect 7395 8045 7525 8075
rect 7555 8045 7685 8075
rect 7715 8045 7720 8075
rect 7360 8040 7720 8045
rect 5520 7995 7320 8000
rect 5520 7965 5525 7995
rect 5555 7965 5685 7995
rect 5715 7965 5845 7995
rect 5875 7965 6005 7995
rect 6035 7965 6165 7995
rect 6195 7965 6325 7995
rect 6355 7965 6485 7995
rect 6515 7965 6645 7995
rect 6675 7965 6805 7995
rect 6835 7965 6965 7995
rect 6995 7965 7125 7995
rect 7155 7965 7285 7995
rect 7315 7965 7320 7995
rect 5520 7960 7320 7965
rect 7360 7995 7720 8000
rect 7360 7965 7365 7995
rect 7395 7965 7525 7995
rect 7555 7965 7685 7995
rect 7715 7965 7720 7995
rect 7360 7960 7720 7965
rect 5520 7915 7320 7920
rect 5520 7885 5525 7915
rect 5555 7885 5685 7915
rect 5715 7885 5845 7915
rect 5875 7885 6005 7915
rect 6035 7885 6165 7915
rect 6195 7885 6325 7915
rect 6355 7885 6485 7915
rect 6515 7885 6645 7915
rect 6675 7885 6805 7915
rect 6835 7885 6965 7915
rect 6995 7885 7125 7915
rect 7155 7885 7285 7915
rect 7315 7885 7320 7915
rect 5520 7880 7320 7885
rect 7360 7915 7720 7920
rect 7360 7885 7365 7915
rect 7395 7885 7525 7915
rect 7555 7885 7685 7915
rect 7715 7885 7720 7915
rect 7360 7880 7720 7885
rect 5520 7835 7320 7840
rect 5520 7805 5525 7835
rect 5555 7805 5685 7835
rect 5715 7805 5845 7835
rect 5875 7805 6005 7835
rect 6035 7805 6165 7835
rect 6195 7805 6325 7835
rect 6355 7805 6485 7835
rect 6515 7805 6645 7835
rect 6675 7805 6805 7835
rect 6835 7805 6965 7835
rect 6995 7805 7125 7835
rect 7155 7805 7285 7835
rect 7315 7805 7320 7835
rect 5520 7800 7320 7805
rect 7360 7835 7720 7840
rect 7360 7805 7365 7835
rect 7395 7805 7525 7835
rect 7555 7805 7685 7835
rect 7715 7805 7720 7835
rect 7360 7800 7720 7805
rect 5520 7755 7320 7760
rect 5520 7725 5525 7755
rect 5555 7725 5685 7755
rect 5715 7725 5845 7755
rect 5875 7725 6005 7755
rect 6035 7725 6165 7755
rect 6195 7725 6325 7755
rect 6355 7725 6485 7755
rect 6515 7725 6645 7755
rect 6675 7725 6805 7755
rect 6835 7725 6965 7755
rect 6995 7725 7125 7755
rect 7155 7725 7285 7755
rect 7315 7725 7320 7755
rect 5520 7720 7320 7725
rect 7360 7755 7720 7760
rect 7360 7725 7365 7755
rect 7395 7725 7525 7755
rect 7555 7725 7685 7755
rect 7715 7725 7720 7755
rect 7360 7720 7720 7725
rect 5520 7675 7320 7680
rect 5520 7645 5525 7675
rect 5555 7645 5685 7675
rect 5715 7645 5845 7675
rect 5875 7645 6005 7675
rect 6035 7645 6165 7675
rect 6195 7645 6325 7675
rect 6355 7645 6485 7675
rect 6515 7645 6645 7675
rect 6675 7645 6805 7675
rect 6835 7645 6965 7675
rect 6995 7645 7125 7675
rect 7155 7645 7285 7675
rect 7315 7645 7320 7675
rect 5520 7640 7320 7645
rect 7360 7675 7720 7680
rect 7360 7645 7365 7675
rect 7395 7645 7525 7675
rect 7555 7645 7685 7675
rect 7715 7645 7720 7675
rect 7360 7640 7720 7645
rect 5520 7595 7320 7600
rect 5520 7565 5525 7595
rect 5555 7565 5685 7595
rect 5715 7565 5845 7595
rect 5875 7565 6005 7595
rect 6035 7565 6165 7595
rect 6195 7565 6325 7595
rect 6355 7565 6485 7595
rect 6515 7565 6645 7595
rect 6675 7565 6805 7595
rect 6835 7565 6965 7595
rect 6995 7565 7125 7595
rect 7155 7565 7285 7595
rect 7315 7565 7320 7595
rect 5520 7560 7320 7565
rect 7360 7595 7720 7600
rect 7360 7565 7365 7595
rect 7395 7565 7525 7595
rect 7555 7565 7685 7595
rect 7715 7565 7720 7595
rect 7360 7560 7720 7565
rect 5520 7515 7320 7520
rect 5520 7485 5525 7515
rect 5555 7485 5685 7515
rect 5715 7485 5845 7515
rect 5875 7485 6005 7515
rect 6035 7485 6165 7515
rect 6195 7485 6325 7515
rect 6355 7485 6485 7515
rect 6515 7485 6645 7515
rect 6675 7485 6805 7515
rect 6835 7485 6965 7515
rect 6995 7485 7125 7515
rect 7155 7485 7285 7515
rect 7315 7485 7320 7515
rect 5520 7480 7320 7485
rect 7360 7515 7720 7520
rect 7360 7485 7365 7515
rect 7395 7485 7525 7515
rect 7555 7485 7685 7515
rect 7715 7485 7720 7515
rect 7360 7480 7720 7485
rect 5520 7435 7320 7440
rect 5520 7405 5525 7435
rect 5555 7405 5685 7435
rect 5715 7405 5845 7435
rect 5875 7405 6005 7435
rect 6035 7405 6165 7435
rect 6195 7405 6325 7435
rect 6355 7405 6485 7435
rect 6515 7405 6645 7435
rect 6675 7405 6805 7435
rect 6835 7405 6965 7435
rect 6995 7405 7125 7435
rect 7155 7405 7285 7435
rect 7315 7405 7320 7435
rect 5520 7400 7320 7405
rect 7360 7435 7720 7440
rect 7360 7405 7365 7435
rect 7395 7405 7525 7435
rect 7555 7405 7685 7435
rect 7715 7405 7720 7435
rect 7360 7400 7720 7405
rect 5520 7355 7320 7360
rect 5520 7325 5525 7355
rect 5555 7325 5685 7355
rect 5715 7325 5845 7355
rect 5875 7325 6005 7355
rect 6035 7325 6165 7355
rect 6195 7325 6325 7355
rect 6355 7325 6485 7355
rect 6515 7325 6645 7355
rect 6675 7325 6805 7355
rect 6835 7325 6965 7355
rect 6995 7325 7125 7355
rect 7155 7325 7285 7355
rect 7315 7325 7320 7355
rect 5520 7320 7320 7325
rect 7360 7355 7720 7360
rect 7360 7325 7365 7355
rect 7395 7325 7525 7355
rect 7555 7325 7685 7355
rect 7715 7325 7720 7355
rect 7360 7320 7720 7325
rect 5520 7275 7320 7280
rect 5520 7245 5525 7275
rect 5555 7245 5685 7275
rect 5715 7245 5845 7275
rect 5875 7245 6005 7275
rect 6035 7245 6165 7275
rect 6195 7245 6325 7275
rect 6355 7245 6485 7275
rect 6515 7245 6645 7275
rect 6675 7245 6805 7275
rect 6835 7245 6965 7275
rect 6995 7245 7125 7275
rect 7155 7245 7285 7275
rect 7315 7245 7320 7275
rect 5520 7240 7320 7245
rect 7360 7275 7720 7280
rect 7360 7245 7365 7275
rect 7395 7245 7525 7275
rect 7555 7245 7685 7275
rect 7715 7245 7720 7275
rect 7360 7240 7720 7245
rect 5520 7195 7320 7200
rect 5520 7165 5525 7195
rect 5555 7165 5685 7195
rect 5715 7165 5845 7195
rect 5875 7165 6005 7195
rect 6035 7165 6165 7195
rect 6195 7165 6325 7195
rect 6355 7165 6485 7195
rect 6515 7165 6645 7195
rect 6675 7165 6805 7195
rect 6835 7165 6965 7195
rect 6995 7165 7125 7195
rect 7155 7165 7285 7195
rect 7315 7165 7320 7195
rect 5520 7160 7320 7165
rect 7360 7195 7720 7200
rect 7360 7165 7365 7195
rect 7395 7165 7525 7195
rect 7555 7165 7685 7195
rect 7715 7165 7720 7195
rect 7360 7160 7720 7165
rect 5480 7115 6120 7120
rect 5480 7085 6085 7115
rect 6115 7085 6120 7115
rect 5480 7080 6120 7085
rect 6160 7115 7320 7120
rect 6160 7085 6165 7115
rect 6195 7085 6325 7115
rect 6355 7085 6485 7115
rect 6515 7085 6645 7115
rect 6675 7085 6805 7115
rect 6835 7085 6965 7115
rect 6995 7085 7125 7115
rect 7155 7085 7285 7115
rect 7315 7085 7320 7115
rect 6160 7080 7320 7085
rect 7360 7115 7720 7120
rect 7360 7085 7365 7115
rect 7395 7085 7525 7115
rect 7555 7085 7685 7115
rect 7715 7085 7720 7115
rect 7360 7080 7720 7085
rect 5520 7035 7320 7040
rect 5520 7005 5525 7035
rect 5555 7005 5685 7035
rect 5715 7005 5845 7035
rect 5875 7005 6005 7035
rect 6035 7005 6165 7035
rect 6195 7005 6325 7035
rect 6355 7005 6485 7035
rect 6515 7005 6645 7035
rect 6675 7005 6805 7035
rect 6835 7005 6965 7035
rect 6995 7005 7125 7035
rect 7155 7005 7285 7035
rect 7315 7005 7320 7035
rect 5520 7000 7320 7005
rect 7360 7035 7720 7040
rect 7360 7005 7365 7035
rect 7395 7005 7525 7035
rect 7555 7005 7685 7035
rect 7715 7005 7720 7035
rect 7360 7000 7720 7005
rect 5520 6955 7320 6960
rect 5520 6925 5525 6955
rect 5555 6925 5685 6955
rect 5715 6925 5845 6955
rect 5875 6925 6005 6955
rect 6035 6925 6165 6955
rect 6195 6925 6325 6955
rect 6355 6925 6485 6955
rect 6515 6925 6645 6955
rect 6675 6925 6805 6955
rect 6835 6925 6965 6955
rect 6995 6925 7125 6955
rect 7155 6925 7285 6955
rect 7315 6925 7320 6955
rect 5520 6920 7320 6925
rect 7360 6955 7720 6960
rect 7360 6925 7365 6955
rect 7395 6925 7525 6955
rect 7555 6925 7685 6955
rect 7715 6925 7720 6955
rect 7360 6920 7720 6925
rect 5480 6875 6280 6880
rect 5480 6845 6245 6875
rect 6275 6845 6280 6875
rect 5480 6840 6280 6845
rect 6320 6875 7320 6880
rect 6320 6845 6325 6875
rect 6355 6845 6485 6875
rect 6515 6845 6645 6875
rect 6675 6845 6805 6875
rect 6835 6845 6965 6875
rect 6995 6845 7125 6875
rect 7155 6845 7285 6875
rect 7315 6845 7320 6875
rect 6320 6840 7320 6845
rect 7360 6875 7720 6880
rect 7360 6845 7365 6875
rect 7395 6845 7525 6875
rect 7555 6845 7685 6875
rect 7715 6845 7720 6875
rect 7360 6840 7720 6845
rect 5520 6795 7320 6800
rect 5520 6765 5525 6795
rect 5555 6765 5685 6795
rect 5715 6765 5845 6795
rect 5875 6765 6005 6795
rect 6035 6765 6165 6795
rect 6195 6765 6325 6795
rect 6355 6765 6485 6795
rect 6515 6765 6645 6795
rect 6675 6765 6805 6795
rect 6835 6765 6965 6795
rect 6995 6765 7125 6795
rect 7155 6765 7285 6795
rect 7315 6765 7320 6795
rect 5520 6760 7320 6765
rect 7360 6795 7720 6800
rect 7360 6765 7365 6795
rect 7395 6765 7525 6795
rect 7555 6765 7685 6795
rect 7715 6765 7720 6795
rect 7360 6760 7720 6765
rect 5520 6715 7320 6720
rect 5520 6685 5525 6715
rect 5555 6685 5685 6715
rect 5715 6685 5845 6715
rect 5875 6685 6005 6715
rect 6035 6685 6165 6715
rect 6195 6685 6325 6715
rect 6355 6685 6485 6715
rect 6515 6685 6645 6715
rect 6675 6685 6805 6715
rect 6835 6685 6965 6715
rect 6995 6685 7125 6715
rect 7155 6685 7285 6715
rect 7315 6685 7320 6715
rect 5520 6680 7320 6685
rect 7360 6715 7720 6720
rect 7360 6685 7365 6715
rect 7395 6685 7525 6715
rect 7555 6685 7685 6715
rect 7715 6685 7720 6715
rect 7360 6680 7720 6685
rect 5520 6635 7320 6640
rect 5520 6605 5525 6635
rect 5555 6605 5685 6635
rect 5715 6605 5845 6635
rect 5875 6605 6005 6635
rect 6035 6605 6165 6635
rect 6195 6605 6325 6635
rect 6355 6605 6485 6635
rect 6515 6605 6645 6635
rect 6675 6605 6805 6635
rect 6835 6605 6965 6635
rect 6995 6605 7125 6635
rect 7155 6605 7285 6635
rect 7315 6605 7320 6635
rect 5520 6600 7320 6605
rect 7360 6635 7720 6640
rect 7360 6605 7365 6635
rect 7395 6605 7525 6635
rect 7555 6605 7685 6635
rect 7715 6605 7720 6635
rect 7360 6600 7720 6605
rect 5520 6555 7320 6560
rect 5520 6525 5525 6555
rect 5555 6525 5685 6555
rect 5715 6525 5845 6555
rect 5875 6525 6005 6555
rect 6035 6525 6165 6555
rect 6195 6525 6325 6555
rect 6355 6525 6485 6555
rect 6515 6525 6645 6555
rect 6675 6525 6805 6555
rect 6835 6525 6965 6555
rect 6995 6525 7125 6555
rect 7155 6525 7285 6555
rect 7315 6525 7320 6555
rect 5520 6520 7320 6525
rect 7360 6555 7720 6560
rect 7360 6525 7365 6555
rect 7395 6525 7525 6555
rect 7555 6525 7685 6555
rect 7715 6525 7720 6555
rect 7360 6520 7720 6525
rect 5520 6475 7320 6480
rect 5520 6445 5525 6475
rect 5555 6445 5685 6475
rect 5715 6445 5845 6475
rect 5875 6445 6005 6475
rect 6035 6445 6165 6475
rect 6195 6445 6325 6475
rect 6355 6445 6485 6475
rect 6515 6445 6645 6475
rect 6675 6445 6805 6475
rect 6835 6445 6965 6475
rect 6995 6445 7125 6475
rect 7155 6445 7285 6475
rect 7315 6445 7320 6475
rect 5520 6440 7320 6445
rect 7360 6475 7720 6480
rect 7360 6445 7365 6475
rect 7395 6445 7525 6475
rect 7555 6445 7685 6475
rect 7715 6445 7720 6475
rect 7360 6440 7720 6445
rect 5480 6395 6600 6400
rect 5480 6365 6565 6395
rect 6595 6365 6600 6395
rect 5480 6360 6600 6365
rect 6640 6395 7320 6400
rect 6640 6365 6645 6395
rect 6675 6365 6805 6395
rect 6835 6365 6965 6395
rect 6995 6365 7125 6395
rect 7155 6365 7285 6395
rect 7315 6365 7320 6395
rect 6640 6360 7320 6365
rect 7360 6395 7720 6400
rect 7360 6365 7365 6395
rect 7395 6365 7525 6395
rect 7555 6365 7685 6395
rect 7715 6365 7720 6395
rect 7360 6360 7720 6365
rect 5520 6315 7320 6320
rect 5520 6285 5525 6315
rect 5555 6285 5685 6315
rect 5715 6285 5845 6315
rect 5875 6285 6005 6315
rect 6035 6285 6165 6315
rect 6195 6285 6325 6315
rect 6355 6285 6485 6315
rect 6515 6285 6645 6315
rect 6675 6285 6805 6315
rect 6835 6285 6965 6315
rect 6995 6285 7125 6315
rect 7155 6285 7285 6315
rect 7315 6285 7320 6315
rect 5520 6280 7320 6285
rect 7360 6315 7720 6320
rect 7360 6285 7365 6315
rect 7395 6285 7525 6315
rect 7555 6285 7685 6315
rect 7715 6285 7720 6315
rect 7360 6280 7720 6285
rect 5520 6235 7320 6240
rect 5520 6205 5525 6235
rect 5555 6205 5685 6235
rect 5715 6205 5845 6235
rect 5875 6205 6005 6235
rect 6035 6205 6165 6235
rect 6195 6205 6325 6235
rect 6355 6205 6485 6235
rect 6515 6205 6645 6235
rect 6675 6205 6805 6235
rect 6835 6205 6965 6235
rect 6995 6205 7125 6235
rect 7155 6205 7285 6235
rect 7315 6205 7320 6235
rect 5520 6200 7320 6205
rect 7360 6235 7720 6240
rect 7360 6205 7365 6235
rect 7395 6205 7525 6235
rect 7555 6205 7685 6235
rect 7715 6205 7720 6235
rect 7360 6200 7720 6205
rect 5520 6155 7320 6160
rect 5520 6125 5525 6155
rect 5555 6125 5685 6155
rect 5715 6125 5845 6155
rect 5875 6125 6005 6155
rect 6035 6125 6165 6155
rect 6195 6125 6325 6155
rect 6355 6125 6485 6155
rect 6515 6125 6645 6155
rect 6675 6125 6805 6155
rect 6835 6125 6965 6155
rect 6995 6125 7125 6155
rect 7155 6125 7285 6155
rect 7315 6125 7320 6155
rect 5520 6120 7320 6125
rect 7360 6155 7720 6160
rect 7360 6125 7365 6155
rect 7395 6125 7525 6155
rect 7555 6125 7685 6155
rect 7715 6125 7720 6155
rect 7360 6120 7720 6125
rect 5480 6075 7080 6080
rect 5480 6045 7045 6075
rect 7075 6045 7080 6075
rect 5480 6040 7080 6045
rect 7120 6075 7320 6080
rect 7120 6045 7125 6075
rect 7155 6045 7285 6075
rect 7315 6045 7320 6075
rect 7120 6040 7320 6045
rect 7360 6075 7720 6080
rect 7360 6045 7365 6075
rect 7395 6045 7525 6075
rect 7555 6045 7685 6075
rect 7715 6045 7720 6075
rect 7360 6040 7720 6045
rect 5520 5995 7320 6000
rect 5520 5965 5525 5995
rect 5555 5965 5685 5995
rect 5715 5965 5845 5995
rect 5875 5965 6005 5995
rect 6035 5965 6165 5995
rect 6195 5965 6325 5995
rect 6355 5965 6485 5995
rect 6515 5965 6645 5995
rect 6675 5965 6805 5995
rect 6835 5965 6965 5995
rect 6995 5965 7125 5995
rect 7155 5965 7285 5995
rect 7315 5965 7320 5995
rect 5520 5960 7320 5965
rect 7360 5995 7720 6000
rect 7360 5965 7365 5995
rect 7395 5965 7525 5995
rect 7555 5965 7685 5995
rect 7715 5965 7720 5995
rect 7360 5960 7720 5965
rect 5480 5915 6920 5920
rect 5480 5885 6885 5915
rect 6915 5885 6920 5915
rect 5480 5880 6920 5885
rect 6960 5915 7320 5920
rect 6960 5885 6965 5915
rect 6995 5885 7125 5915
rect 7155 5885 7285 5915
rect 7315 5885 7320 5915
rect 6960 5880 7320 5885
rect 7360 5915 7720 5920
rect 7360 5885 7365 5915
rect 7395 5885 7525 5915
rect 7555 5885 7685 5915
rect 7715 5885 7720 5915
rect 7360 5880 7720 5885
rect 5520 5835 7320 5840
rect 5520 5805 5525 5835
rect 5555 5805 5685 5835
rect 5715 5805 5845 5835
rect 5875 5805 6005 5835
rect 6035 5805 6165 5835
rect 6195 5805 6325 5835
rect 6355 5805 6485 5835
rect 6515 5805 6645 5835
rect 6675 5805 6805 5835
rect 6835 5805 6965 5835
rect 6995 5805 7125 5835
rect 7155 5805 7285 5835
rect 7315 5805 7320 5835
rect 5520 5800 7320 5805
rect 7360 5835 7720 5840
rect 7360 5805 7365 5835
rect 7395 5805 7525 5835
rect 7555 5805 7685 5835
rect 7715 5805 7720 5835
rect 7360 5800 7720 5805
rect 5520 5755 7320 5760
rect 5520 5725 5525 5755
rect 5555 5725 5685 5755
rect 5715 5725 5845 5755
rect 5875 5725 6005 5755
rect 6035 5725 6165 5755
rect 6195 5725 6325 5755
rect 6355 5725 6485 5755
rect 6515 5725 6645 5755
rect 6675 5725 6805 5755
rect 6835 5725 6965 5755
rect 6995 5725 7125 5755
rect 7155 5725 7285 5755
rect 7315 5725 7320 5755
rect 5520 5720 7320 5725
rect 7360 5755 7720 5760
rect 7360 5725 7365 5755
rect 7395 5725 7525 5755
rect 7555 5725 7685 5755
rect 7715 5725 7720 5755
rect 7360 5720 7720 5725
rect 5520 5675 7320 5680
rect 5520 5645 5525 5675
rect 5555 5645 5685 5675
rect 5715 5645 5845 5675
rect 5875 5645 6005 5675
rect 6035 5645 6165 5675
rect 6195 5645 6325 5675
rect 6355 5645 6485 5675
rect 6515 5645 6645 5675
rect 6675 5645 6805 5675
rect 6835 5645 6965 5675
rect 6995 5645 7125 5675
rect 7155 5645 7285 5675
rect 7315 5645 7320 5675
rect 5520 5640 7320 5645
rect 7360 5675 7720 5680
rect 7360 5645 7365 5675
rect 7395 5645 7525 5675
rect 7555 5645 7685 5675
rect 7715 5645 7720 5675
rect 7360 5640 7720 5645
rect 5520 5595 7320 5600
rect 5520 5565 5525 5595
rect 5555 5565 5685 5595
rect 5715 5565 5845 5595
rect 5875 5565 6005 5595
rect 6035 5565 6165 5595
rect 6195 5565 6325 5595
rect 6355 5565 6485 5595
rect 6515 5565 6645 5595
rect 6675 5565 6805 5595
rect 6835 5565 6965 5595
rect 6995 5565 7125 5595
rect 7155 5565 7285 5595
rect 7315 5565 7320 5595
rect 5520 5560 7320 5565
rect 7360 5595 7720 5600
rect 7360 5565 7365 5595
rect 7395 5565 7525 5595
rect 7555 5565 7685 5595
rect 7715 5565 7720 5595
rect 7360 5560 7720 5565
rect 5520 5515 7320 5520
rect 5520 5485 5525 5515
rect 5555 5485 5685 5515
rect 5715 5485 5845 5515
rect 5875 5485 6005 5515
rect 6035 5485 6165 5515
rect 6195 5485 6325 5515
rect 6355 5485 6485 5515
rect 6515 5485 6645 5515
rect 6675 5485 6805 5515
rect 6835 5485 6965 5515
rect 6995 5485 7125 5515
rect 7155 5485 7285 5515
rect 7315 5485 7320 5515
rect 5520 5480 7320 5485
rect 7360 5515 7720 5520
rect 7360 5485 7365 5515
rect 7395 5485 7525 5515
rect 7555 5485 7685 5515
rect 7715 5485 7720 5515
rect 7360 5480 7720 5485
rect 5520 5435 7320 5440
rect 5520 5405 5525 5435
rect 5555 5405 5685 5435
rect 5715 5405 5845 5435
rect 5875 5405 6005 5435
rect 6035 5405 6165 5435
rect 6195 5405 6325 5435
rect 6355 5405 6485 5435
rect 6515 5405 6645 5435
rect 6675 5405 6805 5435
rect 6835 5405 6965 5435
rect 6995 5405 7125 5435
rect 7155 5405 7285 5435
rect 7315 5405 7320 5435
rect 5520 5400 7320 5405
rect 7360 5435 7720 5440
rect 7360 5405 7365 5435
rect 7395 5405 7525 5435
rect 7555 5405 7685 5435
rect 7715 5405 7720 5435
rect 7360 5400 7720 5405
rect 5520 5355 7320 5360
rect 5520 5325 5525 5355
rect 5555 5325 5685 5355
rect 5715 5325 5845 5355
rect 5875 5325 6005 5355
rect 6035 5325 6165 5355
rect 6195 5325 6325 5355
rect 6355 5325 6485 5355
rect 6515 5325 6645 5355
rect 6675 5325 6805 5355
rect 6835 5325 6965 5355
rect 6995 5325 7125 5355
rect 7155 5325 7285 5355
rect 7315 5325 7320 5355
rect 5520 5320 7320 5325
rect 7360 5355 7720 5360
rect 7360 5325 7365 5355
rect 7395 5325 7525 5355
rect 7555 5325 7685 5355
rect 7715 5325 7720 5355
rect 7360 5320 7720 5325
rect 5520 5275 7320 5280
rect 5520 5245 5525 5275
rect 5555 5245 5685 5275
rect 5715 5245 5845 5275
rect 5875 5245 6005 5275
rect 6035 5245 6165 5275
rect 6195 5245 6325 5275
rect 6355 5245 6485 5275
rect 6515 5245 6645 5275
rect 6675 5245 6805 5275
rect 6835 5245 6965 5275
rect 6995 5245 7125 5275
rect 7155 5245 7285 5275
rect 7315 5245 7320 5275
rect 5520 5240 7320 5245
rect 7360 5275 7720 5280
rect 7360 5245 7365 5275
rect 7395 5245 7525 5275
rect 7555 5245 7685 5275
rect 7715 5245 7720 5275
rect 7360 5240 7720 5245
rect 5520 5195 7320 5200
rect 5520 5165 5525 5195
rect 5555 5165 5685 5195
rect 5715 5165 5845 5195
rect 5875 5165 6005 5195
rect 6035 5165 6165 5195
rect 6195 5165 6325 5195
rect 6355 5165 6485 5195
rect 6515 5165 6645 5195
rect 6675 5165 6805 5195
rect 6835 5165 6965 5195
rect 6995 5165 7125 5195
rect 7155 5165 7285 5195
rect 7315 5165 7320 5195
rect 5520 5160 7320 5165
rect 7360 5195 7720 5200
rect 7360 5165 7365 5195
rect 7395 5165 7525 5195
rect 7555 5165 7685 5195
rect 7715 5165 7720 5195
rect 7360 5160 7720 5165
rect 5520 5115 7320 5120
rect 5520 5085 5525 5115
rect 5555 5085 5685 5115
rect 5715 5085 5845 5115
rect 5875 5085 6005 5115
rect 6035 5085 6165 5115
rect 6195 5085 6325 5115
rect 6355 5085 6485 5115
rect 6515 5085 6645 5115
rect 6675 5085 6805 5115
rect 6835 5085 6965 5115
rect 6995 5085 7125 5115
rect 7155 5085 7285 5115
rect 7315 5085 7320 5115
rect 5520 5080 7320 5085
rect 7360 5115 7720 5120
rect 7360 5085 7365 5115
rect 7395 5085 7525 5115
rect 7555 5085 7685 5115
rect 7715 5085 7720 5115
rect 7360 5080 7720 5085
rect 5520 5035 7320 5040
rect 5520 5005 5525 5035
rect 5555 5005 5685 5035
rect 5715 5005 5845 5035
rect 5875 5005 6005 5035
rect 6035 5005 6165 5035
rect 6195 5005 6325 5035
rect 6355 5005 6485 5035
rect 6515 5005 6645 5035
rect 6675 5005 6805 5035
rect 6835 5005 6965 5035
rect 6995 5005 7125 5035
rect 7155 5005 7285 5035
rect 7315 5005 7320 5035
rect 5520 5000 7320 5005
rect 7360 5035 7720 5040
rect 7360 5005 7365 5035
rect 7395 5005 7525 5035
rect 7555 5005 7685 5035
rect 7715 5005 7720 5035
rect 7360 5000 7720 5005
rect 5520 4955 7320 4960
rect 5520 4925 5525 4955
rect 5555 4925 5685 4955
rect 5715 4925 5845 4955
rect 5875 4925 6005 4955
rect 6035 4925 6165 4955
rect 6195 4925 6325 4955
rect 6355 4925 6485 4955
rect 6515 4925 6645 4955
rect 6675 4925 6805 4955
rect 6835 4925 6965 4955
rect 6995 4925 7125 4955
rect 7155 4925 7285 4955
rect 7315 4925 7320 4955
rect 5520 4920 7320 4925
rect 7360 4955 7720 4960
rect 7360 4925 7365 4955
rect 7395 4925 7525 4955
rect 7555 4925 7685 4955
rect 7715 4925 7720 4955
rect 7360 4920 7720 4925
rect 5520 4875 7320 4880
rect 5520 4845 5525 4875
rect 5555 4845 5685 4875
rect 5715 4845 5845 4875
rect 5875 4845 6005 4875
rect 6035 4845 6165 4875
rect 6195 4845 6325 4875
rect 6355 4845 6485 4875
rect 6515 4845 6645 4875
rect 6675 4845 6805 4875
rect 6835 4845 6965 4875
rect 6995 4845 7125 4875
rect 7155 4845 7285 4875
rect 7315 4845 7320 4875
rect 5520 4840 7320 4845
rect 7360 4875 7720 4880
rect 7360 4845 7365 4875
rect 7395 4845 7525 4875
rect 7555 4845 7685 4875
rect 7715 4845 7720 4875
rect 7360 4840 7720 4845
rect 5520 4795 7320 4800
rect 5520 4765 5525 4795
rect 5555 4765 5685 4795
rect 5715 4765 5845 4795
rect 5875 4765 6005 4795
rect 6035 4765 6165 4795
rect 6195 4765 6325 4795
rect 6355 4765 6485 4795
rect 6515 4765 6645 4795
rect 6675 4765 6805 4795
rect 6835 4765 6965 4795
rect 6995 4765 7125 4795
rect 7155 4765 7285 4795
rect 7315 4765 7320 4795
rect 5520 4760 7320 4765
rect 7360 4795 7720 4800
rect 7360 4765 7365 4795
rect 7395 4765 7525 4795
rect 7555 4765 7685 4795
rect 7715 4765 7720 4795
rect 7360 4760 7720 4765
rect 5480 4715 6120 4720
rect 5480 4685 6085 4715
rect 6115 4685 6120 4715
rect 5480 4680 6120 4685
rect 6160 4715 7320 4720
rect 6160 4685 6165 4715
rect 6195 4685 6325 4715
rect 6355 4685 6485 4715
rect 6515 4685 6645 4715
rect 6675 4685 6805 4715
rect 6835 4685 6965 4715
rect 6995 4685 7125 4715
rect 7155 4685 7285 4715
rect 7315 4685 7320 4715
rect 6160 4680 7320 4685
rect 7360 4715 7720 4720
rect 7360 4685 7365 4715
rect 7395 4685 7525 4715
rect 7555 4685 7685 4715
rect 7715 4685 7720 4715
rect 7360 4680 7720 4685
rect 5520 4635 7320 4640
rect 5520 4605 5525 4635
rect 5555 4605 5685 4635
rect 5715 4605 5845 4635
rect 5875 4605 6005 4635
rect 6035 4605 6165 4635
rect 6195 4605 6325 4635
rect 6355 4605 6485 4635
rect 6515 4605 6645 4635
rect 6675 4605 6805 4635
rect 6835 4605 6965 4635
rect 6995 4605 7125 4635
rect 7155 4605 7285 4635
rect 7315 4605 7320 4635
rect 5520 4600 7320 4605
rect 7360 4635 7720 4640
rect 7360 4605 7365 4635
rect 7395 4605 7525 4635
rect 7555 4605 7685 4635
rect 7715 4605 7720 4635
rect 7360 4600 7720 4605
rect 5520 4555 7320 4560
rect 5520 4525 5525 4555
rect 5555 4525 5685 4555
rect 5715 4525 5845 4555
rect 5875 4525 6005 4555
rect 6035 4525 6165 4555
rect 6195 4525 6325 4555
rect 6355 4525 6485 4555
rect 6515 4525 6645 4555
rect 6675 4525 6805 4555
rect 6835 4525 6965 4555
rect 6995 4525 7125 4555
rect 7155 4525 7285 4555
rect 7315 4525 7320 4555
rect 5520 4520 7320 4525
rect 7360 4555 7720 4560
rect 7360 4525 7365 4555
rect 7395 4525 7525 4555
rect 7555 4525 7685 4555
rect 7715 4525 7720 4555
rect 7360 4520 7720 4525
rect 5480 4475 6280 4480
rect 5480 4445 6245 4475
rect 6275 4445 6280 4475
rect 5480 4440 6280 4445
rect 6320 4475 7320 4480
rect 6320 4445 6325 4475
rect 6355 4445 6485 4475
rect 6515 4445 6645 4475
rect 6675 4445 6805 4475
rect 6835 4445 6965 4475
rect 6995 4445 7125 4475
rect 7155 4445 7285 4475
rect 7315 4445 7320 4475
rect 6320 4440 7320 4445
rect 7360 4475 7720 4480
rect 7360 4445 7365 4475
rect 7395 4445 7525 4475
rect 7555 4445 7685 4475
rect 7715 4445 7720 4475
rect 7360 4440 7720 4445
rect 5520 4395 7320 4400
rect 5520 4365 5525 4395
rect 5555 4365 5685 4395
rect 5715 4365 5845 4395
rect 5875 4365 6005 4395
rect 6035 4365 6165 4395
rect 6195 4365 6325 4395
rect 6355 4365 6485 4395
rect 6515 4365 6645 4395
rect 6675 4365 6805 4395
rect 6835 4365 6965 4395
rect 6995 4365 7125 4395
rect 7155 4365 7285 4395
rect 7315 4365 7320 4395
rect 5520 4360 7320 4365
rect 7360 4395 7720 4400
rect 7360 4365 7365 4395
rect 7395 4365 7525 4395
rect 7555 4365 7685 4395
rect 7715 4365 7720 4395
rect 7360 4360 7720 4365
rect 5520 4315 7320 4320
rect 5520 4285 5525 4315
rect 5555 4285 5685 4315
rect 5715 4285 5845 4315
rect 5875 4285 6005 4315
rect 6035 4285 6165 4315
rect 6195 4285 6325 4315
rect 6355 4285 6485 4315
rect 6515 4285 6645 4315
rect 6675 4285 6805 4315
rect 6835 4285 6965 4315
rect 6995 4285 7125 4315
rect 7155 4285 7285 4315
rect 7315 4285 7320 4315
rect 5520 4280 7320 4285
rect 7360 4315 7720 4320
rect 7360 4285 7365 4315
rect 7395 4285 7525 4315
rect 7555 4285 7685 4315
rect 7715 4285 7720 4315
rect 7360 4280 7720 4285
rect 5520 4235 7320 4240
rect 5520 4205 5525 4235
rect 5555 4205 5685 4235
rect 5715 4205 5845 4235
rect 5875 4205 6005 4235
rect 6035 4205 6165 4235
rect 6195 4205 6325 4235
rect 6355 4205 6485 4235
rect 6515 4205 6645 4235
rect 6675 4205 6805 4235
rect 6835 4205 6965 4235
rect 6995 4205 7125 4235
rect 7155 4205 7285 4235
rect 7315 4205 7320 4235
rect 5520 4200 7320 4205
rect 7360 4235 7720 4240
rect 7360 4205 7365 4235
rect 7395 4205 7525 4235
rect 7555 4205 7685 4235
rect 7715 4205 7720 4235
rect 7360 4200 7720 4205
rect 5520 4155 7320 4160
rect 5520 4125 5525 4155
rect 5555 4125 5685 4155
rect 5715 4125 5845 4155
rect 5875 4125 6005 4155
rect 6035 4125 6165 4155
rect 6195 4125 6325 4155
rect 6355 4125 6485 4155
rect 6515 4125 6645 4155
rect 6675 4125 6805 4155
rect 6835 4125 6965 4155
rect 6995 4125 7125 4155
rect 7155 4125 7285 4155
rect 7315 4125 7320 4155
rect 5520 4120 7320 4125
rect 7360 4155 7720 4160
rect 7360 4125 7365 4155
rect 7395 4125 7525 4155
rect 7555 4125 7685 4155
rect 7715 4125 7720 4155
rect 7360 4120 7720 4125
rect 5520 4075 7320 4080
rect 5520 4045 5525 4075
rect 5555 4045 5685 4075
rect 5715 4045 5845 4075
rect 5875 4045 6005 4075
rect 6035 4045 6165 4075
rect 6195 4045 6325 4075
rect 6355 4045 6485 4075
rect 6515 4045 6645 4075
rect 6675 4045 6805 4075
rect 6835 4045 6965 4075
rect 6995 4045 7125 4075
rect 7155 4045 7285 4075
rect 7315 4045 7320 4075
rect 5520 4040 7320 4045
rect 7360 4075 7720 4080
rect 7360 4045 7365 4075
rect 7395 4045 7525 4075
rect 7555 4045 7685 4075
rect 7715 4045 7720 4075
rect 7360 4040 7720 4045
rect 5480 3995 6440 4000
rect 5480 3965 6405 3995
rect 6435 3965 6440 3995
rect 5480 3960 6440 3965
rect 6480 3995 7320 4000
rect 6480 3965 6485 3995
rect 6515 3965 6645 3995
rect 6675 3965 6805 3995
rect 6835 3965 6965 3995
rect 6995 3965 7125 3995
rect 7155 3965 7285 3995
rect 7315 3965 7320 3995
rect 6480 3960 7320 3965
rect 7360 3995 7720 4000
rect 7360 3965 7365 3995
rect 7395 3965 7525 3995
rect 7555 3965 7685 3995
rect 7715 3965 7720 3995
rect 7360 3960 7720 3965
rect 5520 3915 7320 3920
rect 5520 3885 5525 3915
rect 5555 3885 5685 3915
rect 5715 3885 5845 3915
rect 5875 3885 6005 3915
rect 6035 3885 6165 3915
rect 6195 3885 6325 3915
rect 6355 3885 6485 3915
rect 6515 3885 6645 3915
rect 6675 3885 6805 3915
rect 6835 3885 6965 3915
rect 6995 3885 7125 3915
rect 7155 3885 7285 3915
rect 7315 3885 7320 3915
rect 5520 3880 7320 3885
rect 7360 3915 7720 3920
rect 7360 3885 7365 3915
rect 7395 3885 7525 3915
rect 7555 3885 7685 3915
rect 7715 3885 7720 3915
rect 7360 3880 7720 3885
rect 5520 3835 7320 3840
rect 5520 3805 5525 3835
rect 5555 3805 5685 3835
rect 5715 3805 5845 3835
rect 5875 3805 6005 3835
rect 6035 3805 6165 3835
rect 6195 3805 6325 3835
rect 6355 3805 6485 3835
rect 6515 3805 6645 3835
rect 6675 3805 6805 3835
rect 6835 3805 6965 3835
rect 6995 3805 7125 3835
rect 7155 3805 7285 3835
rect 7315 3805 7320 3835
rect 5520 3800 7320 3805
rect 7360 3835 7720 3840
rect 7360 3805 7365 3835
rect 7395 3805 7525 3835
rect 7555 3805 7685 3835
rect 7715 3805 7720 3835
rect 7360 3800 7720 3805
rect 5520 3755 7320 3760
rect 5520 3725 5525 3755
rect 5555 3725 5685 3755
rect 5715 3725 5845 3755
rect 5875 3725 6005 3755
rect 6035 3725 6165 3755
rect 6195 3725 6325 3755
rect 6355 3725 6485 3755
rect 6515 3725 6645 3755
rect 6675 3725 6805 3755
rect 6835 3725 6965 3755
rect 6995 3725 7125 3755
rect 7155 3725 7285 3755
rect 7315 3725 7320 3755
rect 5520 3720 7320 3725
rect 7360 3755 7720 3760
rect 7360 3725 7365 3755
rect 7395 3725 7525 3755
rect 7555 3725 7685 3755
rect 7715 3725 7720 3755
rect 7360 3720 7720 3725
rect 5480 3675 7080 3680
rect 5480 3645 7045 3675
rect 7075 3645 7080 3675
rect 5480 3640 7080 3645
rect 7120 3675 7320 3680
rect 7120 3645 7125 3675
rect 7155 3645 7285 3675
rect 7315 3645 7320 3675
rect 7120 3640 7320 3645
rect 7360 3675 7720 3680
rect 7360 3645 7365 3675
rect 7395 3645 7525 3675
rect 7555 3645 7685 3675
rect 7715 3645 7720 3675
rect 7360 3640 7720 3645
rect 5520 3595 7320 3600
rect 5520 3565 5525 3595
rect 5555 3565 5685 3595
rect 5715 3565 5845 3595
rect 5875 3565 6005 3595
rect 6035 3565 6165 3595
rect 6195 3565 6325 3595
rect 6355 3565 6485 3595
rect 6515 3565 6645 3595
rect 6675 3565 6805 3595
rect 6835 3565 6965 3595
rect 6995 3565 7125 3595
rect 7155 3565 7285 3595
rect 7315 3565 7320 3595
rect 5520 3560 7320 3565
rect 7360 3595 7720 3600
rect 7360 3565 7365 3595
rect 7395 3565 7525 3595
rect 7555 3565 7685 3595
rect 7715 3565 7720 3595
rect 7360 3560 7720 3565
rect 5480 3515 6760 3520
rect 5480 3485 6725 3515
rect 6755 3485 6760 3515
rect 5480 3480 6760 3485
rect 6800 3515 7320 3520
rect 6800 3485 6805 3515
rect 6835 3485 6965 3515
rect 6995 3485 7125 3515
rect 7155 3485 7285 3515
rect 7315 3485 7320 3515
rect 6800 3480 7320 3485
rect 7360 3515 7720 3520
rect 7360 3485 7365 3515
rect 7395 3485 7525 3515
rect 7555 3485 7685 3515
rect 7715 3485 7720 3515
rect 7360 3480 7720 3485
rect 5520 3435 7320 3440
rect 5520 3405 5525 3435
rect 5555 3405 5685 3435
rect 5715 3405 5845 3435
rect 5875 3405 6005 3435
rect 6035 3405 6165 3435
rect 6195 3405 6325 3435
rect 6355 3405 6485 3435
rect 6515 3405 6645 3435
rect 6675 3405 6805 3435
rect 6835 3405 6965 3435
rect 6995 3405 7125 3435
rect 7155 3405 7285 3435
rect 7315 3405 7320 3435
rect 5520 3400 7320 3405
rect 7360 3435 7720 3440
rect 7360 3405 7365 3435
rect 7395 3405 7525 3435
rect 7555 3405 7685 3435
rect 7715 3405 7720 3435
rect 7360 3400 7720 3405
rect 5520 3355 7320 3360
rect 5520 3325 5525 3355
rect 5555 3325 5685 3355
rect 5715 3325 5845 3355
rect 5875 3325 6005 3355
rect 6035 3325 6165 3355
rect 6195 3325 6325 3355
rect 6355 3325 6485 3355
rect 6515 3325 6645 3355
rect 6675 3325 6805 3355
rect 6835 3325 6965 3355
rect 6995 3325 7125 3355
rect 7155 3325 7285 3355
rect 7315 3325 7320 3355
rect 5520 3320 7320 3325
rect 7360 3355 7720 3360
rect 7360 3325 7365 3355
rect 7395 3325 7525 3355
rect 7555 3325 7685 3355
rect 7715 3325 7720 3355
rect 7360 3320 7720 3325
rect 5520 3275 7320 3280
rect 5520 3245 5525 3275
rect 5555 3245 5685 3275
rect 5715 3245 5845 3275
rect 5875 3245 6005 3275
rect 6035 3245 6165 3275
rect 6195 3245 6325 3275
rect 6355 3245 6485 3275
rect 6515 3245 6645 3275
rect 6675 3245 6805 3275
rect 6835 3245 6965 3275
rect 6995 3245 7125 3275
rect 7155 3245 7285 3275
rect 7315 3245 7320 3275
rect 5520 3240 7320 3245
rect 7360 3275 7720 3280
rect 7360 3245 7365 3275
rect 7395 3245 7525 3275
rect 7555 3245 7685 3275
rect 7715 3245 7720 3275
rect 7360 3240 7720 3245
rect 5520 3195 7320 3200
rect 5520 3165 5525 3195
rect 5555 3165 5685 3195
rect 5715 3165 5845 3195
rect 5875 3165 6005 3195
rect 6035 3165 6165 3195
rect 6195 3165 6325 3195
rect 6355 3165 6485 3195
rect 6515 3165 6645 3195
rect 6675 3165 6805 3195
rect 6835 3165 6965 3195
rect 6995 3165 7125 3195
rect 7155 3165 7285 3195
rect 7315 3165 7320 3195
rect 5520 3160 7320 3165
rect 7360 3195 7720 3200
rect 7360 3165 7365 3195
rect 7395 3165 7525 3195
rect 7555 3165 7685 3195
rect 7715 3165 7720 3195
rect 7360 3160 7720 3165
rect 5520 3115 7320 3120
rect 5520 3085 5525 3115
rect 5555 3085 5685 3115
rect 5715 3085 5845 3115
rect 5875 3085 6005 3115
rect 6035 3085 6165 3115
rect 6195 3085 6325 3115
rect 6355 3085 6485 3115
rect 6515 3085 6645 3115
rect 6675 3085 6805 3115
rect 6835 3085 6965 3115
rect 6995 3085 7125 3115
rect 7155 3085 7285 3115
rect 7315 3085 7320 3115
rect 5520 3080 7320 3085
rect 7360 3115 7720 3120
rect 7360 3085 7365 3115
rect 7395 3085 7525 3115
rect 7555 3085 7685 3115
rect 7715 3085 7720 3115
rect 7360 3080 7720 3085
rect 5520 3035 7320 3040
rect 5520 3005 5525 3035
rect 5555 3005 5685 3035
rect 5715 3005 5845 3035
rect 5875 3005 6005 3035
rect 6035 3005 6165 3035
rect 6195 3005 6325 3035
rect 6355 3005 6485 3035
rect 6515 3005 6645 3035
rect 6675 3005 6805 3035
rect 6835 3005 6965 3035
rect 6995 3005 7125 3035
rect 7155 3005 7285 3035
rect 7315 3005 7320 3035
rect 5520 3000 7320 3005
rect 7360 3035 7720 3040
rect 7360 3005 7365 3035
rect 7395 3005 7525 3035
rect 7555 3005 7685 3035
rect 7715 3005 7720 3035
rect 7360 3000 7720 3005
rect 5520 2955 7320 2960
rect 5520 2925 5525 2955
rect 5555 2925 5685 2955
rect 5715 2925 5845 2955
rect 5875 2925 6005 2955
rect 6035 2925 6165 2955
rect 6195 2925 6325 2955
rect 6355 2925 6485 2955
rect 6515 2925 6645 2955
rect 6675 2925 6805 2955
rect 6835 2925 6965 2955
rect 6995 2925 7125 2955
rect 7155 2925 7285 2955
rect 7315 2925 7320 2955
rect 5520 2920 7320 2925
rect 7360 2955 7720 2960
rect 7360 2925 7365 2955
rect 7395 2925 7525 2955
rect 7555 2925 7685 2955
rect 7715 2925 7720 2955
rect 7360 2920 7720 2925
rect 5520 2875 7320 2880
rect 5520 2845 5525 2875
rect 5555 2845 5685 2875
rect 5715 2845 5845 2875
rect 5875 2845 6005 2875
rect 6035 2845 6165 2875
rect 6195 2845 6325 2875
rect 6355 2845 6485 2875
rect 6515 2845 6645 2875
rect 6675 2845 6805 2875
rect 6835 2845 6965 2875
rect 6995 2845 7125 2875
rect 7155 2845 7285 2875
rect 7315 2845 7320 2875
rect 5520 2840 7320 2845
rect 7360 2875 7720 2880
rect 7360 2845 7365 2875
rect 7395 2845 7525 2875
rect 7555 2845 7685 2875
rect 7715 2845 7720 2875
rect 7360 2840 7720 2845
rect 5520 2795 7320 2800
rect 5520 2765 5525 2795
rect 5555 2765 5685 2795
rect 5715 2765 5845 2795
rect 5875 2765 6005 2795
rect 6035 2765 6165 2795
rect 6195 2765 6325 2795
rect 6355 2765 6485 2795
rect 6515 2765 6645 2795
rect 6675 2765 6805 2795
rect 6835 2765 6965 2795
rect 6995 2765 7125 2795
rect 7155 2765 7285 2795
rect 7315 2765 7320 2795
rect 5520 2760 7320 2765
rect 7360 2795 7720 2800
rect 7360 2765 7365 2795
rect 7395 2765 7525 2795
rect 7555 2765 7685 2795
rect 7715 2765 7720 2795
rect 7360 2760 7720 2765
rect 5520 2715 7320 2720
rect 5520 2685 5525 2715
rect 5555 2685 5685 2715
rect 5715 2685 5845 2715
rect 5875 2685 6005 2715
rect 6035 2685 6165 2715
rect 6195 2685 6325 2715
rect 6355 2685 6485 2715
rect 6515 2685 6645 2715
rect 6675 2685 6805 2715
rect 6835 2685 6965 2715
rect 6995 2685 7125 2715
rect 7155 2685 7285 2715
rect 7315 2685 7320 2715
rect 5520 2680 7320 2685
rect 7360 2715 7720 2720
rect 7360 2685 7365 2715
rect 7395 2685 7525 2715
rect 7555 2685 7685 2715
rect 7715 2685 7720 2715
rect 7360 2680 7720 2685
rect 5520 2635 7320 2640
rect 5520 2605 5525 2635
rect 5555 2605 5685 2635
rect 5715 2605 5845 2635
rect 5875 2605 6005 2635
rect 6035 2605 6165 2635
rect 6195 2605 6325 2635
rect 6355 2605 6485 2635
rect 6515 2605 6645 2635
rect 6675 2605 6805 2635
rect 6835 2605 6965 2635
rect 6995 2605 7125 2635
rect 7155 2605 7285 2635
rect 7315 2605 7320 2635
rect 5520 2600 7320 2605
rect 7360 2635 7720 2640
rect 7360 2605 7365 2635
rect 7395 2605 7525 2635
rect 7555 2605 7685 2635
rect 7715 2605 7720 2635
rect 7360 2600 7720 2605
rect 5520 2555 7320 2560
rect 5520 2525 5525 2555
rect 5555 2525 5685 2555
rect 5715 2525 5845 2555
rect 5875 2525 6005 2555
rect 6035 2525 6165 2555
rect 6195 2525 6325 2555
rect 6355 2525 6485 2555
rect 6515 2525 6645 2555
rect 6675 2525 6805 2555
rect 6835 2525 6965 2555
rect 6995 2525 7125 2555
rect 7155 2525 7285 2555
rect 7315 2525 7320 2555
rect 5520 2520 7320 2525
rect 7360 2555 7720 2560
rect 7360 2525 7365 2555
rect 7395 2525 7525 2555
rect 7555 2525 7685 2555
rect 7715 2525 7720 2555
rect 7360 2520 7720 2525
rect 5520 2475 7320 2480
rect 5520 2445 5525 2475
rect 5555 2445 5685 2475
rect 5715 2445 5845 2475
rect 5875 2445 6005 2475
rect 6035 2445 6165 2475
rect 6195 2445 6325 2475
rect 6355 2445 6485 2475
rect 6515 2445 6645 2475
rect 6675 2445 6805 2475
rect 6835 2445 6965 2475
rect 6995 2445 7125 2475
rect 7155 2445 7285 2475
rect 7315 2445 7320 2475
rect 5520 2440 7320 2445
rect 7360 2475 7720 2480
rect 7360 2445 7365 2475
rect 7395 2445 7525 2475
rect 7555 2445 7685 2475
rect 7715 2445 7720 2475
rect 7360 2440 7720 2445
rect 5520 2395 7320 2400
rect 5520 2365 5525 2395
rect 5555 2365 5685 2395
rect 5715 2365 5845 2395
rect 5875 2365 6005 2395
rect 6035 2365 6165 2395
rect 6195 2365 6325 2395
rect 6355 2365 6485 2395
rect 6515 2365 6645 2395
rect 6675 2365 6805 2395
rect 6835 2365 6965 2395
rect 6995 2365 7125 2395
rect 7155 2365 7285 2395
rect 7315 2365 7320 2395
rect 5520 2360 7320 2365
rect 7360 2395 7720 2400
rect 7360 2365 7365 2395
rect 7395 2365 7525 2395
rect 7555 2365 7685 2395
rect 7715 2365 7720 2395
rect 7360 2360 7720 2365
rect 5480 2315 6120 2320
rect 5480 2285 6085 2315
rect 6115 2285 6120 2315
rect 5480 2280 6120 2285
rect 6160 2315 7320 2320
rect 6160 2285 6165 2315
rect 6195 2285 6325 2315
rect 6355 2285 6485 2315
rect 6515 2285 6645 2315
rect 6675 2285 6805 2315
rect 6835 2285 6965 2315
rect 6995 2285 7125 2315
rect 7155 2285 7285 2315
rect 7315 2285 7320 2315
rect 6160 2280 7320 2285
rect 7360 2315 7720 2320
rect 7360 2285 7365 2315
rect 7395 2285 7525 2315
rect 7555 2285 7685 2315
rect 7715 2285 7720 2315
rect 7360 2280 7720 2285
rect 5520 2235 7320 2240
rect 5520 2205 5525 2235
rect 5555 2205 5685 2235
rect 5715 2205 5845 2235
rect 5875 2205 6005 2235
rect 6035 2205 6165 2235
rect 6195 2205 6325 2235
rect 6355 2205 6485 2235
rect 6515 2205 6645 2235
rect 6675 2205 6805 2235
rect 6835 2205 6965 2235
rect 6995 2205 7125 2235
rect 7155 2205 7285 2235
rect 7315 2205 7320 2235
rect 5520 2200 7320 2205
rect 7360 2235 7720 2240
rect 7360 2205 7365 2235
rect 7395 2205 7525 2235
rect 7555 2205 7685 2235
rect 7715 2205 7720 2235
rect 7360 2200 7720 2205
rect 5520 2155 7320 2160
rect 5520 2125 5525 2155
rect 5555 2125 5685 2155
rect 5715 2125 5845 2155
rect 5875 2125 6005 2155
rect 6035 2125 6165 2155
rect 6195 2125 6325 2155
rect 6355 2125 6485 2155
rect 6515 2125 6645 2155
rect 6675 2125 6805 2155
rect 6835 2125 6965 2155
rect 6995 2125 7125 2155
rect 7155 2125 7285 2155
rect 7315 2125 7320 2155
rect 5520 2120 7320 2125
rect 7360 2155 7720 2160
rect 7360 2125 7365 2155
rect 7395 2125 7525 2155
rect 7555 2125 7685 2155
rect 7715 2125 7720 2155
rect 7360 2120 7720 2125
rect 5520 2075 7320 2080
rect 5520 2045 5525 2075
rect 5555 2045 5685 2075
rect 5715 2045 5845 2075
rect 5875 2045 6005 2075
rect 6035 2045 6165 2075
rect 6195 2045 6325 2075
rect 6355 2045 6485 2075
rect 6515 2045 6645 2075
rect 6675 2045 6805 2075
rect 6835 2045 6965 2075
rect 6995 2045 7125 2075
rect 7155 2045 7285 2075
rect 7315 2045 7320 2075
rect 5520 2040 7320 2045
rect 7360 2075 7720 2080
rect 7360 2045 7365 2075
rect 7395 2045 7525 2075
rect 7555 2045 7685 2075
rect 7715 2045 7720 2075
rect 7360 2040 7720 2045
rect 5520 1995 7320 2000
rect 5520 1965 5525 1995
rect 5555 1965 5685 1995
rect 5715 1965 5845 1995
rect 5875 1965 6005 1995
rect 6035 1965 6165 1995
rect 6195 1965 6325 1995
rect 6355 1965 6485 1995
rect 6515 1965 6645 1995
rect 6675 1965 6805 1995
rect 6835 1965 6965 1995
rect 6995 1965 7125 1995
rect 7155 1965 7285 1995
rect 7315 1965 7320 1995
rect 5520 1960 7320 1965
rect 7360 1995 7720 2000
rect 7360 1965 7365 1995
rect 7395 1965 7525 1995
rect 7555 1965 7685 1995
rect 7715 1965 7720 1995
rect 7360 1960 7720 1965
rect 5520 1915 7320 1920
rect 5520 1885 5525 1915
rect 5555 1885 5685 1915
rect 5715 1885 5845 1915
rect 5875 1885 6005 1915
rect 6035 1885 6165 1915
rect 6195 1885 6325 1915
rect 6355 1885 6485 1915
rect 6515 1885 6645 1915
rect 6675 1885 6805 1915
rect 6835 1885 6965 1915
rect 6995 1885 7125 1915
rect 7155 1885 7285 1915
rect 7315 1885 7320 1915
rect 5520 1880 7320 1885
rect 7360 1915 7720 1920
rect 7360 1885 7365 1915
rect 7395 1885 7525 1915
rect 7555 1885 7685 1915
rect 7715 1885 7720 1915
rect 7360 1880 7720 1885
rect 5520 1835 7320 1840
rect 5520 1805 5525 1835
rect 5555 1805 5685 1835
rect 5715 1805 5845 1835
rect 5875 1805 6005 1835
rect 6035 1805 6165 1835
rect 6195 1805 6325 1835
rect 6355 1805 6485 1835
rect 6515 1805 6645 1835
rect 6675 1805 6805 1835
rect 6835 1805 6965 1835
rect 6995 1805 7125 1835
rect 7155 1805 7285 1835
rect 7315 1805 7320 1835
rect 5520 1800 7320 1805
rect 7360 1835 7720 1840
rect 7360 1805 7365 1835
rect 7395 1805 7525 1835
rect 7555 1805 7685 1835
rect 7715 1805 7720 1835
rect 7360 1800 7720 1805
rect 5520 1755 7320 1760
rect 5520 1725 5525 1755
rect 5555 1725 5685 1755
rect 5715 1725 5845 1755
rect 5875 1725 6005 1755
rect 6035 1725 6165 1755
rect 6195 1725 6325 1755
rect 6355 1725 6485 1755
rect 6515 1725 6645 1755
rect 6675 1725 6805 1755
rect 6835 1725 6965 1755
rect 6995 1725 7125 1755
rect 7155 1725 7285 1755
rect 7315 1725 7320 1755
rect 5520 1720 7320 1725
rect 7360 1755 7720 1760
rect 7360 1725 7365 1755
rect 7395 1725 7525 1755
rect 7555 1725 7685 1755
rect 7715 1725 7720 1755
rect 7360 1720 7720 1725
rect 5520 1675 7320 1680
rect 5520 1645 5525 1675
rect 5555 1645 5685 1675
rect 5715 1645 5845 1675
rect 5875 1645 6005 1675
rect 6035 1645 6165 1675
rect 6195 1645 6325 1675
rect 6355 1645 6485 1675
rect 6515 1645 6645 1675
rect 6675 1645 6805 1675
rect 6835 1645 6965 1675
rect 6995 1645 7125 1675
rect 7155 1645 7285 1675
rect 7315 1645 7320 1675
rect 5520 1640 7320 1645
rect 7360 1675 7720 1680
rect 7360 1645 7365 1675
rect 7395 1645 7525 1675
rect 7555 1645 7685 1675
rect 7715 1645 7720 1675
rect 7360 1640 7720 1645
rect 5480 1595 5960 1600
rect 5480 1565 5925 1595
rect 5955 1565 5960 1595
rect 5480 1560 5960 1565
rect 6000 1595 7320 1600
rect 6000 1565 6005 1595
rect 6035 1565 6165 1595
rect 6195 1565 6325 1595
rect 6355 1565 6485 1595
rect 6515 1565 6645 1595
rect 6675 1565 6805 1595
rect 6835 1565 6965 1595
rect 6995 1565 7125 1595
rect 7155 1565 7285 1595
rect 7315 1565 7320 1595
rect 6000 1560 7320 1565
rect 7360 1595 7720 1600
rect 7360 1565 7365 1595
rect 7395 1565 7525 1595
rect 7555 1565 7685 1595
rect 7715 1565 7720 1595
rect 7360 1560 7720 1565
rect 5520 1515 7320 1520
rect 5520 1485 5525 1515
rect 5555 1485 5685 1515
rect 5715 1485 5845 1515
rect 5875 1485 6005 1515
rect 6035 1485 6165 1515
rect 6195 1485 6325 1515
rect 6355 1485 6485 1515
rect 6515 1485 6645 1515
rect 6675 1485 6805 1515
rect 6835 1485 6965 1515
rect 6995 1485 7125 1515
rect 7155 1485 7285 1515
rect 7315 1485 7320 1515
rect 5520 1480 7320 1485
rect 7360 1515 7720 1520
rect 7360 1485 7365 1515
rect 7395 1485 7525 1515
rect 7555 1485 7685 1515
rect 7715 1485 7720 1515
rect 7360 1480 7720 1485
rect 5520 1435 7320 1440
rect 5520 1405 5525 1435
rect 5555 1405 5685 1435
rect 5715 1405 5845 1435
rect 5875 1405 6005 1435
rect 6035 1405 6165 1435
rect 6195 1405 6325 1435
rect 6355 1405 6485 1435
rect 6515 1405 6645 1435
rect 6675 1405 6805 1435
rect 6835 1405 6965 1435
rect 6995 1405 7125 1435
rect 7155 1405 7285 1435
rect 7315 1405 7320 1435
rect 5520 1400 7320 1405
rect 7360 1435 7720 1440
rect 7360 1405 7365 1435
rect 7395 1405 7525 1435
rect 7555 1405 7685 1435
rect 7715 1405 7720 1435
rect 7360 1400 7720 1405
rect 5520 1355 7320 1360
rect 5520 1325 5525 1355
rect 5555 1325 5685 1355
rect 5715 1325 5845 1355
rect 5875 1325 6005 1355
rect 6035 1325 6165 1355
rect 6195 1325 6325 1355
rect 6355 1325 6485 1355
rect 6515 1325 6645 1355
rect 6675 1325 6805 1355
rect 6835 1325 6965 1355
rect 6995 1325 7125 1355
rect 7155 1325 7285 1355
rect 7315 1325 7320 1355
rect 5520 1320 7320 1325
rect 7360 1355 7720 1360
rect 7360 1325 7365 1355
rect 7395 1325 7525 1355
rect 7555 1325 7685 1355
rect 7715 1325 7720 1355
rect 7360 1320 7720 1325
rect 5480 1275 5640 1280
rect 5480 1245 5605 1275
rect 5635 1245 5640 1275
rect 5480 1240 5640 1245
rect 5680 1275 7320 1280
rect 5680 1245 5685 1275
rect 5715 1245 5845 1275
rect 5875 1245 6005 1275
rect 6035 1245 6165 1275
rect 6195 1245 6325 1275
rect 6355 1245 6485 1275
rect 6515 1245 6645 1275
rect 6675 1245 6805 1275
rect 6835 1245 6965 1275
rect 6995 1245 7125 1275
rect 7155 1245 7285 1275
rect 7315 1245 7320 1275
rect 5680 1240 7320 1245
rect 7360 1275 7720 1280
rect 7360 1245 7365 1275
rect 7395 1245 7525 1275
rect 7555 1245 7685 1275
rect 7715 1245 7720 1275
rect 7360 1240 7720 1245
rect 5520 1195 7320 1200
rect 5520 1165 5525 1195
rect 5555 1165 5685 1195
rect 5715 1165 5845 1195
rect 5875 1165 6005 1195
rect 6035 1165 6165 1195
rect 6195 1165 6325 1195
rect 6355 1165 6485 1195
rect 6515 1165 6645 1195
rect 6675 1165 6805 1195
rect 6835 1165 6965 1195
rect 6995 1165 7125 1195
rect 7155 1165 7285 1195
rect 7315 1165 7320 1195
rect 5520 1160 7320 1165
rect 7360 1195 7720 1200
rect 7360 1165 7365 1195
rect 7395 1165 7525 1195
rect 7555 1165 7685 1195
rect 7715 1165 7720 1195
rect 7360 1160 7720 1165
rect 5520 1115 7320 1120
rect 5520 1085 5525 1115
rect 5555 1085 5685 1115
rect 5715 1085 5845 1115
rect 5875 1085 6005 1115
rect 6035 1085 6165 1115
rect 6195 1085 6325 1115
rect 6355 1085 6485 1115
rect 6515 1085 6645 1115
rect 6675 1085 6805 1115
rect 6835 1085 6965 1115
rect 6995 1085 7125 1115
rect 7155 1085 7285 1115
rect 7315 1085 7320 1115
rect 5520 1080 7320 1085
rect 7360 1115 7720 1120
rect 7360 1085 7365 1115
rect 7395 1085 7525 1115
rect 7555 1085 7685 1115
rect 7715 1085 7720 1115
rect 7360 1080 7720 1085
rect 5520 1035 7320 1040
rect 5520 1005 5525 1035
rect 5555 1005 5685 1035
rect 5715 1005 5845 1035
rect 5875 1005 6005 1035
rect 6035 1005 6165 1035
rect 6195 1005 6325 1035
rect 6355 1005 6485 1035
rect 6515 1005 6645 1035
rect 6675 1005 6805 1035
rect 6835 1005 6965 1035
rect 6995 1005 7125 1035
rect 7155 1005 7285 1035
rect 7315 1005 7320 1035
rect 5520 1000 7320 1005
rect 7360 1035 7720 1040
rect 7360 1005 7365 1035
rect 7395 1005 7525 1035
rect 7555 1005 7685 1035
rect 7715 1005 7720 1035
rect 7360 1000 7720 1005
rect 5520 955 7320 960
rect 5520 925 5525 955
rect 5555 925 5685 955
rect 5715 925 5845 955
rect 5875 925 6005 955
rect 6035 925 6165 955
rect 6195 925 6325 955
rect 6355 925 6485 955
rect 6515 925 6645 955
rect 6675 925 6805 955
rect 6835 925 6965 955
rect 6995 925 7125 955
rect 7155 925 7285 955
rect 7315 925 7320 955
rect 5520 920 7320 925
rect 7360 955 7720 960
rect 7360 925 7365 955
rect 7395 925 7525 955
rect 7555 925 7685 955
rect 7715 925 7720 955
rect 7360 920 7720 925
rect 5520 875 7320 880
rect 5520 845 5525 875
rect 5555 845 5685 875
rect 5715 845 5845 875
rect 5875 845 6005 875
rect 6035 845 6165 875
rect 6195 845 6325 875
rect 6355 845 6485 875
rect 6515 845 6645 875
rect 6675 845 6805 875
rect 6835 845 6965 875
rect 6995 845 7125 875
rect 7155 845 7285 875
rect 7315 845 7320 875
rect 5520 840 7320 845
rect 7360 875 7720 880
rect 7360 845 7365 875
rect 7395 845 7525 875
rect 7555 845 7685 875
rect 7715 845 7720 875
rect 7360 840 7720 845
rect 5520 795 7320 800
rect 5520 765 5525 795
rect 5555 765 5685 795
rect 5715 765 5845 795
rect 5875 765 6005 795
rect 6035 765 6165 795
rect 6195 765 6325 795
rect 6355 765 6485 795
rect 6515 765 6645 795
rect 6675 765 6805 795
rect 6835 765 6965 795
rect 6995 765 7125 795
rect 7155 765 7285 795
rect 7315 765 7320 795
rect 5520 760 7320 765
rect 7360 795 7720 800
rect 7360 765 7365 795
rect 7395 765 7525 795
rect 7555 765 7685 795
rect 7715 765 7720 795
rect 7360 760 7720 765
rect 5480 715 5800 720
rect 5480 685 5765 715
rect 5795 685 5800 715
rect 5480 680 5800 685
rect 5840 715 7320 720
rect 5840 685 5845 715
rect 5875 685 6005 715
rect 6035 685 6165 715
rect 6195 685 6325 715
rect 6355 685 6485 715
rect 6515 685 6645 715
rect 6675 685 6805 715
rect 6835 685 6965 715
rect 6995 685 7125 715
rect 7155 685 7285 715
rect 7315 685 7320 715
rect 5840 680 7320 685
rect 7360 715 7720 720
rect 7360 685 7365 715
rect 7395 685 7525 715
rect 7555 685 7685 715
rect 7715 685 7720 715
rect 7360 680 7720 685
rect 5520 595 7320 600
rect 5520 565 5525 595
rect 5555 565 5685 595
rect 5715 565 5845 595
rect 5875 565 6005 595
rect 6035 565 6165 595
rect 6195 565 6325 595
rect 6355 565 6485 595
rect 6515 565 6645 595
rect 6675 565 6805 595
rect 6835 565 6965 595
rect 6995 565 7125 595
rect 7155 565 7285 595
rect 7315 565 7320 595
rect 5520 560 7320 565
rect 7360 595 7720 600
rect 7360 565 7365 595
rect 7395 565 7525 595
rect 7555 565 7685 595
rect 7715 565 7720 595
rect 7360 560 7720 565
rect 5520 515 7320 520
rect 5520 485 5525 515
rect 5555 485 5685 515
rect 5715 485 5845 515
rect 5875 485 6005 515
rect 6035 485 6165 515
rect 6195 485 6325 515
rect 6355 485 6485 515
rect 6515 485 6645 515
rect 6675 485 6805 515
rect 6835 485 6965 515
rect 6995 485 7125 515
rect 7155 485 7285 515
rect 7315 485 7320 515
rect 5520 480 7320 485
rect 7360 515 7720 520
rect 7360 485 7365 515
rect 7395 485 7525 515
rect 7555 485 7685 515
rect 7715 485 7720 515
rect 7360 480 7720 485
rect 5480 435 5640 440
rect 5480 405 5605 435
rect 5635 405 5640 435
rect 5480 400 5640 405
rect 5680 435 7320 440
rect 5680 405 5685 435
rect 5715 405 5845 435
rect 5875 405 6005 435
rect 6035 405 6165 435
rect 6195 405 6325 435
rect 6355 405 6485 435
rect 6515 405 6645 435
rect 6675 405 6805 435
rect 6835 405 6965 435
rect 6995 405 7125 435
rect 7155 405 7285 435
rect 7315 405 7320 435
rect 5680 400 7320 405
rect 7360 435 7720 440
rect 7360 405 7365 435
rect 7395 405 7525 435
rect 7555 405 7685 435
rect 7715 405 7720 435
rect 7360 400 7720 405
rect 5520 355 7320 360
rect 5520 325 5525 355
rect 5555 325 5685 355
rect 5715 325 5845 355
rect 5875 325 6005 355
rect 6035 325 6165 355
rect 6195 325 6325 355
rect 6355 325 6485 355
rect 6515 325 6645 355
rect 6675 325 6805 355
rect 6835 325 6965 355
rect 6995 325 7125 355
rect 7155 325 7285 355
rect 7315 325 7320 355
rect 5520 320 7320 325
rect 7360 355 7720 360
rect 7360 325 7365 355
rect 7395 325 7525 355
rect 7555 325 7685 355
rect 7715 325 7720 355
rect 7360 320 7720 325
rect 5520 275 7320 280
rect 5520 245 5525 275
rect 5555 245 5685 275
rect 5715 245 5845 275
rect 5875 245 6005 275
rect 6035 245 6165 275
rect 6195 245 6325 275
rect 6355 245 6485 275
rect 6515 245 6645 275
rect 6675 245 6805 275
rect 6835 245 6965 275
rect 6995 245 7125 275
rect 7155 245 7285 275
rect 7315 245 7320 275
rect 5520 240 7320 245
rect 7360 275 7720 280
rect 7360 245 7365 275
rect 7395 245 7525 275
rect 7555 245 7685 275
rect 7715 245 7720 275
rect 7360 240 7720 245
rect 5520 195 7320 200
rect 5520 165 5525 195
rect 5555 165 5685 195
rect 5715 165 5845 195
rect 5875 165 6005 195
rect 6035 165 6165 195
rect 6195 165 6325 195
rect 6355 165 6485 195
rect 6515 165 6645 195
rect 6675 165 6805 195
rect 6835 165 6965 195
rect 6995 165 7125 195
rect 7155 165 7285 195
rect 7315 165 7320 195
rect 5520 160 7320 165
rect 7360 195 7720 200
rect 7360 165 7365 195
rect 7395 165 7525 195
rect 7555 165 7685 195
rect 7715 165 7720 195
rect 7360 160 7720 165
rect 5520 115 7320 120
rect 5520 85 5525 115
rect 5555 85 5685 115
rect 5715 85 5845 115
rect 5875 85 6005 115
rect 6035 85 6165 115
rect 6195 85 6325 115
rect 6355 85 6485 115
rect 6515 85 6645 115
rect 6675 85 6805 115
rect 6835 85 6965 115
rect 6995 85 7125 115
rect 7155 85 7285 115
rect 7315 85 7320 115
rect 5520 80 7320 85
rect 7360 115 7720 120
rect 7360 85 7365 115
rect 7395 85 7525 115
rect 7555 85 7685 115
rect 7715 85 7720 115
rect 7360 80 7720 85
rect 5520 35 7320 40
rect 5520 5 5525 35
rect 5555 5 5685 35
rect 5715 5 5845 35
rect 5875 5 6005 35
rect 6035 5 6165 35
rect 6195 5 6325 35
rect 6355 5 6485 35
rect 6515 5 6645 35
rect 6675 5 6805 35
rect 6835 5 6965 35
rect 6995 5 7125 35
rect 7155 5 7285 35
rect 7315 5 7320 35
rect 5520 0 7320 5
rect 7360 35 7720 40
rect 7360 5 7365 35
rect 7395 5 7525 35
rect 7555 5 7685 35
rect 7715 5 7720 35
rect 7360 0 7720 5
<< via2 >>
rect 5525 16565 5555 16595
rect 5685 16565 5715 16595
rect 5845 16565 5875 16595
rect 6005 16565 6035 16595
rect 6165 16565 6195 16595
rect 6325 16565 6355 16595
rect 6485 16565 6515 16595
rect 6645 16565 6675 16595
rect 6805 16565 6835 16595
rect 6965 16565 6995 16595
rect 7125 16565 7155 16595
rect 7285 16565 7315 16595
rect 7365 16565 7395 16595
rect 7525 16565 7555 16595
rect 7685 16565 7715 16595
rect 5525 16485 5555 16515
rect 5685 16485 5715 16515
rect 5845 16485 5875 16515
rect 6005 16485 6035 16515
rect 6165 16485 6195 16515
rect 6325 16485 6355 16515
rect 6485 16485 6515 16515
rect 6645 16485 6675 16515
rect 6805 16485 6835 16515
rect 6965 16485 6995 16515
rect 7125 16485 7155 16515
rect 7285 16485 7315 16515
rect 7365 16485 7395 16515
rect 7525 16485 7555 16515
rect 7685 16485 7715 16515
rect 5525 16405 5555 16435
rect 5685 16405 5715 16435
rect 5845 16405 5875 16435
rect 6005 16405 6035 16435
rect 6165 16405 6195 16435
rect 6325 16405 6355 16435
rect 6485 16405 6515 16435
rect 6645 16405 6675 16435
rect 6805 16405 6835 16435
rect 6965 16405 6995 16435
rect 7125 16405 7155 16435
rect 7285 16405 7315 16435
rect 7365 16405 7395 16435
rect 7525 16405 7555 16435
rect 7685 16405 7715 16435
rect 5525 16325 5555 16355
rect 5685 16325 5715 16355
rect 5845 16325 5875 16355
rect 6005 16325 6035 16355
rect 6165 16325 6195 16355
rect 6325 16325 6355 16355
rect 6485 16325 6515 16355
rect 6645 16325 6675 16355
rect 6805 16325 6835 16355
rect 6965 16325 6995 16355
rect 7125 16325 7155 16355
rect 7285 16325 7315 16355
rect 7365 16325 7395 16355
rect 7525 16325 7555 16355
rect 7685 16325 7715 16355
rect 5525 16245 5555 16275
rect 5685 16245 5715 16275
rect 5845 16245 5875 16275
rect 6005 16245 6035 16275
rect 6165 16245 6195 16275
rect 6325 16245 6355 16275
rect 6485 16245 6515 16275
rect 6645 16245 6675 16275
rect 6805 16245 6835 16275
rect 6965 16245 6995 16275
rect 7125 16245 7155 16275
rect 7285 16245 7315 16275
rect 7365 16245 7395 16275
rect 7525 16245 7555 16275
rect 7685 16245 7715 16275
rect 5525 16165 5555 16195
rect 5685 16165 5715 16195
rect 5845 16165 5875 16195
rect 6005 16165 6035 16195
rect 6165 16165 6195 16195
rect 6325 16165 6355 16195
rect 6485 16165 6515 16195
rect 6645 16165 6675 16195
rect 6805 16165 6835 16195
rect 6965 16165 6995 16195
rect 7125 16165 7155 16195
rect 7285 16165 7315 16195
rect 7365 16165 7395 16195
rect 7525 16165 7555 16195
rect 7685 16165 7715 16195
rect 5525 16085 5555 16115
rect 5685 16085 5715 16115
rect 5845 16085 5875 16115
rect 6005 16085 6035 16115
rect 6165 16085 6195 16115
rect 6325 16085 6355 16115
rect 6485 16085 6515 16115
rect 6645 16085 6675 16115
rect 6805 16085 6835 16115
rect 6965 16085 6995 16115
rect 7125 16085 7155 16115
rect 7285 16085 7315 16115
rect 7365 16085 7395 16115
rect 7525 16085 7555 16115
rect 7685 16085 7715 16115
rect 5525 16005 5555 16035
rect 5685 16005 5715 16035
rect 5845 16005 5875 16035
rect 6005 16005 6035 16035
rect 6165 16005 6195 16035
rect 6325 16005 6355 16035
rect 6485 16005 6515 16035
rect 6645 16005 6675 16035
rect 6805 16005 6835 16035
rect 6965 16005 6995 16035
rect 7125 16005 7155 16035
rect 7285 16005 7315 16035
rect 7365 16005 7395 16035
rect 7525 16005 7555 16035
rect 7685 16005 7715 16035
rect 5525 15925 5555 15955
rect 5685 15925 5715 15955
rect 5845 15925 5875 15955
rect 6005 15925 6035 15955
rect 6165 15925 6195 15955
rect 6325 15925 6355 15955
rect 6485 15925 6515 15955
rect 6645 15925 6675 15955
rect 6805 15925 6835 15955
rect 6965 15925 6995 15955
rect 7125 15925 7155 15955
rect 7285 15925 7315 15955
rect 7365 15925 7395 15955
rect 7525 15925 7555 15955
rect 7685 15925 7715 15955
rect 7365 15845 7395 15875
rect 7525 15845 7555 15875
rect 7685 15845 7715 15875
rect 7605 15765 7635 15795
rect 7365 15685 7395 15715
rect 7525 15685 7555 15715
rect 7685 15685 7715 15715
rect 7445 15605 7475 15635
rect 7365 15525 7395 15555
rect 7525 15525 7555 15555
rect 7685 15525 7715 15555
rect 5525 15405 5555 15435
rect 5685 15405 5715 15435
rect 5845 15405 5875 15435
rect 6005 15405 6035 15435
rect 6165 15405 6195 15435
rect 6325 15405 6355 15435
rect 6485 15405 6515 15435
rect 6645 15405 6675 15435
rect 6805 15405 6835 15435
rect 6965 15405 6995 15435
rect 7125 15405 7155 15435
rect 7285 15405 7315 15435
rect 7365 15405 7395 15435
rect 7525 15405 7555 15435
rect 7685 15405 7715 15435
rect 5525 15325 5555 15355
rect 5685 15325 5715 15355
rect 5845 15325 5875 15355
rect 6005 15325 6035 15355
rect 6165 15325 6195 15355
rect 6325 15325 6355 15355
rect 6485 15325 6515 15355
rect 6645 15325 6675 15355
rect 6805 15325 6835 15355
rect 6965 15325 6995 15355
rect 7125 15325 7155 15355
rect 7285 15325 7315 15355
rect 7365 15325 7395 15355
rect 7525 15325 7555 15355
rect 7685 15325 7715 15355
rect 5525 15245 5555 15275
rect 5685 15245 5715 15275
rect 5845 15245 5875 15275
rect 6005 15245 6035 15275
rect 6165 15245 6195 15275
rect 6325 15245 6355 15275
rect 6485 15245 6515 15275
rect 6645 15245 6675 15275
rect 6805 15245 6835 15275
rect 6965 15245 6995 15275
rect 7125 15245 7155 15275
rect 7285 15245 7315 15275
rect 7365 15245 7395 15275
rect 7525 15245 7555 15275
rect 7685 15245 7715 15275
rect 5525 15165 5555 15195
rect 5685 15165 5715 15195
rect 5845 15165 5875 15195
rect 6005 15165 6035 15195
rect 6165 15165 6195 15195
rect 6325 15165 6355 15195
rect 6485 15165 6515 15195
rect 6645 15165 6675 15195
rect 6805 15165 6835 15195
rect 6965 15165 6995 15195
rect 7125 15165 7155 15195
rect 7285 15165 7315 15195
rect 7365 15165 7395 15195
rect 7525 15165 7555 15195
rect 7685 15165 7715 15195
rect 5525 15085 5555 15115
rect 5685 15085 5715 15115
rect 5845 15085 5875 15115
rect 6005 15085 6035 15115
rect 6165 15085 6195 15115
rect 6325 15085 6355 15115
rect 6485 15085 6515 15115
rect 6645 15085 6675 15115
rect 6805 15085 6835 15115
rect 6965 15085 6995 15115
rect 7125 15085 7155 15115
rect 7285 15085 7315 15115
rect 7365 15085 7395 15115
rect 7525 15085 7555 15115
rect 7685 15085 7715 15115
rect 6085 15005 6115 15035
rect 6165 15005 6195 15035
rect 6325 15005 6355 15035
rect 6485 15005 6515 15035
rect 6645 15005 6675 15035
rect 6805 15005 6835 15035
rect 6965 15005 6995 15035
rect 7125 15005 7155 15035
rect 7285 15005 7315 15035
rect 7365 15005 7395 15035
rect 7525 15005 7555 15035
rect 7685 15005 7715 15035
rect 5525 14925 5555 14955
rect 5685 14925 5715 14955
rect 5845 14925 5875 14955
rect 6005 14925 6035 14955
rect 6165 14925 6195 14955
rect 6325 14925 6355 14955
rect 6485 14925 6515 14955
rect 6645 14925 6675 14955
rect 6805 14925 6835 14955
rect 6965 14925 6995 14955
rect 7125 14925 7155 14955
rect 7285 14925 7315 14955
rect 7365 14925 7395 14955
rect 7525 14925 7555 14955
rect 7685 14925 7715 14955
rect 5525 14845 5555 14875
rect 5685 14845 5715 14875
rect 5845 14845 5875 14875
rect 6005 14845 6035 14875
rect 6165 14845 6195 14875
rect 6325 14845 6355 14875
rect 6485 14845 6515 14875
rect 6645 14845 6675 14875
rect 6805 14845 6835 14875
rect 6965 14845 6995 14875
rect 7125 14845 7155 14875
rect 7285 14845 7315 14875
rect 7365 14845 7395 14875
rect 7525 14845 7555 14875
rect 7685 14845 7715 14875
rect 5525 14765 5555 14795
rect 5685 14765 5715 14795
rect 5845 14765 5875 14795
rect 6005 14765 6035 14795
rect 6165 14765 6195 14795
rect 6325 14765 6355 14795
rect 6485 14765 6515 14795
rect 6645 14765 6675 14795
rect 6805 14765 6835 14795
rect 6965 14765 6995 14795
rect 7125 14765 7155 14795
rect 7285 14765 7315 14795
rect 7365 14765 7395 14795
rect 7525 14765 7555 14795
rect 7685 14765 7715 14795
rect 5525 14685 5555 14715
rect 5685 14685 5715 14715
rect 5845 14685 5875 14715
rect 6005 14685 6035 14715
rect 6165 14685 6195 14715
rect 6325 14685 6355 14715
rect 6485 14685 6515 14715
rect 6645 14685 6675 14715
rect 6805 14685 6835 14715
rect 6965 14685 6995 14715
rect 7125 14685 7155 14715
rect 7285 14685 7315 14715
rect 7365 14685 7395 14715
rect 7525 14685 7555 14715
rect 7685 14685 7715 14715
rect 5925 14605 5955 14635
rect 6005 14605 6035 14635
rect 6165 14605 6195 14635
rect 6325 14605 6355 14635
rect 6485 14605 6515 14635
rect 6645 14605 6675 14635
rect 6805 14605 6835 14635
rect 6965 14605 6995 14635
rect 7125 14605 7155 14635
rect 7285 14605 7315 14635
rect 7365 14605 7395 14635
rect 7525 14605 7555 14635
rect 7685 14605 7715 14635
rect 5525 14525 5555 14555
rect 5685 14525 5715 14555
rect 5845 14525 5875 14555
rect 6005 14525 6035 14555
rect 6165 14525 6195 14555
rect 6325 14525 6355 14555
rect 6485 14525 6515 14555
rect 6645 14525 6675 14555
rect 6805 14525 6835 14555
rect 6965 14525 6995 14555
rect 7125 14525 7155 14555
rect 7285 14525 7315 14555
rect 7365 14525 7395 14555
rect 7525 14525 7555 14555
rect 7685 14525 7715 14555
rect 5525 14445 5555 14475
rect 5685 14445 5715 14475
rect 5845 14445 5875 14475
rect 6005 14445 6035 14475
rect 6165 14445 6195 14475
rect 6325 14445 6355 14475
rect 6485 14445 6515 14475
rect 6645 14445 6675 14475
rect 6805 14445 6835 14475
rect 6965 14445 6995 14475
rect 7125 14445 7155 14475
rect 7285 14445 7315 14475
rect 7365 14445 7395 14475
rect 7525 14445 7555 14475
rect 7685 14445 7715 14475
rect 6965 14365 6995 14395
rect 7125 14365 7155 14395
rect 7285 14365 7315 14395
rect 7365 14365 7395 14395
rect 7525 14365 7555 14395
rect 7685 14365 7715 14395
rect 7205 14285 7235 14315
rect 7365 14285 7395 14315
rect 7525 14285 7555 14315
rect 7685 14285 7715 14315
rect 6965 14205 6995 14235
rect 7125 14205 7155 14235
rect 7285 14205 7315 14235
rect 7365 14205 7395 14235
rect 7525 14205 7555 14235
rect 7685 14205 7715 14235
rect 7045 14125 7075 14155
rect 7365 14125 7395 14155
rect 7525 14125 7555 14155
rect 7685 14125 7715 14155
rect 6965 14045 6995 14075
rect 7125 14045 7155 14075
rect 7285 14045 7315 14075
rect 7365 14045 7395 14075
rect 7525 14045 7555 14075
rect 7685 14045 7715 14075
rect 5525 13965 5555 13995
rect 5685 13965 5715 13995
rect 5845 13965 5875 13995
rect 6005 13965 6035 13995
rect 6165 13965 6195 13995
rect 6325 13965 6355 13995
rect 6485 13965 6515 13995
rect 6645 13965 6675 13995
rect 6805 13965 6835 13995
rect 6965 13965 6995 13995
rect 7125 13965 7155 13995
rect 7285 13965 7315 13995
rect 7365 13965 7395 13995
rect 7525 13965 7555 13995
rect 7685 13965 7715 13995
rect 5765 13885 5795 13915
rect 5845 13845 5875 13875
rect 6005 13845 6035 13875
rect 6165 13845 6195 13875
rect 6325 13845 6355 13875
rect 6485 13845 6515 13875
rect 6645 13845 6675 13875
rect 6805 13845 6835 13875
rect 6965 13845 6995 13875
rect 7125 13845 7155 13875
rect 7285 13845 7315 13875
rect 7365 13845 7395 13875
rect 7525 13845 7555 13875
rect 7685 13845 7715 13875
rect 5525 13765 5555 13795
rect 5685 13765 5715 13795
rect 5845 13765 5875 13795
rect 6005 13765 6035 13795
rect 6165 13765 6195 13795
rect 6325 13765 6355 13795
rect 6485 13765 6515 13795
rect 6645 13765 6675 13795
rect 6805 13765 6835 13795
rect 6965 13765 6995 13795
rect 7125 13765 7155 13795
rect 7285 13765 7315 13795
rect 7365 13765 7395 13795
rect 7525 13765 7555 13795
rect 7685 13765 7715 13795
rect 5525 13685 5555 13715
rect 5685 13685 5715 13715
rect 5845 13685 5875 13715
rect 6005 13685 6035 13715
rect 6165 13685 6195 13715
rect 6325 13685 6355 13715
rect 6485 13685 6515 13715
rect 6645 13685 6675 13715
rect 6805 13685 6835 13715
rect 6965 13685 6995 13715
rect 7125 13685 7155 13715
rect 7285 13685 7315 13715
rect 7365 13685 7395 13715
rect 7525 13685 7555 13715
rect 7685 13685 7715 13715
rect 5525 13605 5555 13635
rect 5685 13605 5715 13635
rect 5845 13605 5875 13635
rect 6005 13605 6035 13635
rect 6165 13605 6195 13635
rect 6325 13605 6355 13635
rect 6485 13605 6515 13635
rect 6645 13605 6675 13635
rect 6805 13605 6835 13635
rect 6965 13605 6995 13635
rect 7125 13605 7155 13635
rect 7285 13605 7315 13635
rect 7365 13605 7395 13635
rect 7525 13605 7555 13635
rect 7685 13605 7715 13635
rect 6085 13525 6115 13555
rect 6165 13525 6195 13555
rect 6325 13525 6355 13555
rect 6485 13525 6515 13555
rect 6645 13525 6675 13555
rect 6805 13525 6835 13555
rect 6965 13525 6995 13555
rect 7125 13525 7155 13555
rect 7285 13525 7315 13555
rect 7365 13525 7395 13555
rect 7525 13525 7555 13555
rect 7685 13525 7715 13555
rect 5525 13445 5555 13475
rect 5685 13445 5715 13475
rect 5845 13445 5875 13475
rect 6005 13445 6035 13475
rect 6165 13445 6195 13475
rect 6325 13445 6355 13475
rect 6485 13445 6515 13475
rect 6645 13445 6675 13475
rect 6805 13445 6835 13475
rect 6965 13445 6995 13475
rect 7125 13445 7155 13475
rect 7285 13445 7315 13475
rect 7365 13445 7395 13475
rect 7525 13445 7555 13475
rect 7685 13445 7715 13475
rect 5525 13365 5555 13395
rect 5685 13365 5715 13395
rect 5845 13365 5875 13395
rect 6005 13365 6035 13395
rect 6165 13365 6195 13395
rect 6325 13365 6355 13395
rect 6485 13365 6515 13395
rect 6645 13365 6675 13395
rect 6805 13365 6835 13395
rect 6965 13365 6995 13395
rect 7125 13365 7155 13395
rect 7285 13365 7315 13395
rect 7365 13365 7395 13395
rect 7525 13365 7555 13395
rect 7685 13365 7715 13395
rect 5525 13285 5555 13315
rect 5685 13285 5715 13315
rect 5845 13285 5875 13315
rect 6005 13285 6035 13315
rect 6165 13285 6195 13315
rect 6325 13285 6355 13315
rect 6485 13285 6515 13315
rect 6645 13285 6675 13315
rect 6805 13285 6835 13315
rect 6965 13285 6995 13315
rect 7125 13285 7155 13315
rect 7285 13285 7315 13315
rect 7365 13285 7395 13315
rect 7525 13285 7555 13315
rect 7685 13285 7715 13315
rect 5525 13205 5555 13235
rect 5685 13205 5715 13235
rect 5845 13205 5875 13235
rect 6005 13205 6035 13235
rect 6165 13205 6195 13235
rect 6325 13205 6355 13235
rect 6485 13205 6515 13235
rect 6645 13205 6675 13235
rect 6805 13205 6835 13235
rect 6965 13205 6995 13235
rect 7125 13205 7155 13235
rect 7285 13205 7315 13235
rect 7365 13205 7395 13235
rect 7525 13205 7555 13235
rect 7685 13205 7715 13235
rect 5925 13125 5955 13155
rect 6005 13125 6035 13155
rect 6165 13125 6195 13155
rect 6325 13125 6355 13155
rect 6485 13125 6515 13155
rect 6645 13125 6675 13155
rect 6805 13125 6835 13155
rect 6965 13125 6995 13155
rect 7125 13125 7155 13155
rect 7285 13125 7315 13155
rect 7365 13125 7395 13155
rect 7525 13125 7555 13155
rect 7685 13125 7715 13155
rect 5525 13045 5555 13075
rect 5685 13045 5715 13075
rect 5845 13045 5875 13075
rect 6005 13045 6035 13075
rect 6165 13045 6195 13075
rect 6325 13045 6355 13075
rect 6485 13045 6515 13075
rect 6645 13045 6675 13075
rect 6805 13045 6835 13075
rect 6965 13045 6995 13075
rect 7125 13045 7155 13075
rect 7285 13045 7315 13075
rect 7365 13045 7395 13075
rect 7525 13045 7555 13075
rect 7685 13045 7715 13075
rect 5525 12965 5555 12995
rect 5685 12965 5715 12995
rect 5845 12965 5875 12995
rect 6005 12965 6035 12995
rect 6165 12965 6195 12995
rect 6325 12965 6355 12995
rect 6485 12965 6515 12995
rect 6645 12965 6675 12995
rect 6805 12965 6835 12995
rect 6965 12965 6995 12995
rect 7125 12965 7155 12995
rect 7285 12965 7315 12995
rect 7365 12965 7395 12995
rect 7525 12965 7555 12995
rect 7685 12965 7715 12995
rect 7365 12885 7395 12915
rect 7525 12885 7555 12915
rect 7685 12885 7715 12915
rect 7605 12805 7635 12835
rect 7365 12725 7395 12755
rect 7525 12725 7555 12755
rect 7685 12725 7715 12755
rect 7445 12645 7475 12675
rect 7365 12565 7395 12595
rect 7525 12565 7555 12595
rect 7685 12565 7715 12595
rect 5525 12485 5555 12515
rect 5685 12485 5715 12515
rect 5845 12485 5875 12515
rect 6005 12485 6035 12515
rect 6165 12485 6195 12515
rect 6325 12485 6355 12515
rect 6485 12485 6515 12515
rect 6645 12485 6675 12515
rect 6805 12485 6835 12515
rect 6965 12485 6995 12515
rect 7125 12485 7155 12515
rect 7285 12485 7315 12515
rect 7365 12445 7395 12475
rect 7525 12445 7555 12475
rect 7685 12445 7715 12475
rect 5765 12405 5795 12435
rect 5845 12405 5875 12435
rect 6005 12405 6035 12435
rect 6165 12405 6195 12435
rect 6325 12405 6355 12435
rect 6485 12405 6515 12435
rect 6645 12405 6675 12435
rect 6805 12405 6835 12435
rect 6965 12405 6995 12435
rect 7125 12405 7155 12435
rect 7285 12405 7315 12435
rect 7365 12365 7395 12395
rect 7525 12365 7555 12395
rect 7685 12365 7715 12395
rect 5525 12285 5555 12315
rect 5685 12285 5715 12315
rect 5845 12285 5875 12315
rect 6005 12285 6035 12315
rect 6165 12285 6195 12315
rect 6325 12285 6355 12315
rect 6485 12285 6515 12315
rect 6645 12285 6675 12315
rect 6805 12285 6835 12315
rect 6965 12285 6995 12315
rect 7125 12285 7155 12315
rect 7285 12285 7315 12315
rect 7365 12285 7395 12315
rect 7525 12285 7555 12315
rect 7685 12285 7715 12315
rect 5525 12205 5555 12235
rect 5685 12205 5715 12235
rect 5845 12205 5875 12235
rect 6005 12205 6035 12235
rect 6165 12205 6195 12235
rect 6325 12205 6355 12235
rect 6485 12205 6515 12235
rect 6645 12205 6675 12235
rect 6805 12205 6835 12235
rect 6965 12205 6995 12235
rect 7125 12205 7155 12235
rect 7285 12205 7315 12235
rect 7365 12205 7395 12235
rect 7525 12205 7555 12235
rect 7685 12205 7715 12235
rect 5525 12125 5555 12155
rect 5685 12125 5715 12155
rect 5845 12125 5875 12155
rect 6005 12125 6035 12155
rect 6165 12125 6195 12155
rect 6325 12125 6355 12155
rect 6485 12125 6515 12155
rect 6645 12125 6675 12155
rect 6805 12125 6835 12155
rect 6965 12125 6995 12155
rect 7125 12125 7155 12155
rect 7285 12125 7315 12155
rect 7365 12125 7395 12155
rect 7525 12125 7555 12155
rect 7685 12125 7715 12155
rect 5525 12045 5555 12075
rect 5685 12045 5715 12075
rect 5845 12045 5875 12075
rect 6005 12045 6035 12075
rect 6165 12045 6195 12075
rect 6325 12045 6355 12075
rect 6485 12045 6515 12075
rect 6645 12045 6675 12075
rect 6805 12045 6835 12075
rect 6965 12045 6995 12075
rect 7125 12045 7155 12075
rect 7285 12045 7315 12075
rect 7365 12045 7395 12075
rect 7525 12045 7555 12075
rect 7685 12045 7715 12075
rect 5525 11965 5555 11995
rect 5685 11965 5715 11995
rect 5845 11965 5875 11995
rect 6005 11965 6035 11995
rect 6165 11965 6195 11995
rect 6325 11965 6355 11995
rect 6485 11965 6515 11995
rect 6645 11965 6675 11995
rect 6805 11965 6835 11995
rect 6965 11965 6995 11995
rect 7125 11965 7155 11995
rect 7285 11965 7315 11995
rect 7365 11965 7395 11995
rect 7525 11965 7555 11995
rect 7685 11965 7715 11995
rect 5525 11885 5555 11915
rect 5685 11885 5715 11915
rect 5845 11885 5875 11915
rect 6005 11885 6035 11915
rect 6165 11885 6195 11915
rect 6325 11885 6355 11915
rect 6485 11885 6515 11915
rect 6645 11885 6675 11915
rect 6805 11885 6835 11915
rect 6965 11885 6995 11915
rect 7125 11885 7155 11915
rect 7285 11885 7315 11915
rect 7365 11885 7395 11915
rect 7525 11885 7555 11915
rect 7685 11885 7715 11915
rect 5525 11805 5555 11835
rect 5685 11805 5715 11835
rect 5845 11805 5875 11835
rect 6005 11805 6035 11835
rect 6165 11805 6195 11835
rect 6325 11805 6355 11835
rect 6485 11805 6515 11835
rect 6645 11805 6675 11835
rect 6805 11805 6835 11835
rect 6965 11805 6995 11835
rect 7125 11805 7155 11835
rect 7285 11805 7315 11835
rect 7365 11805 7395 11835
rect 7525 11805 7555 11835
rect 7685 11805 7715 11835
rect 5525 11725 5555 11755
rect 5685 11725 5715 11755
rect 5845 11725 5875 11755
rect 6005 11725 6035 11755
rect 6165 11725 6195 11755
rect 6325 11725 6355 11755
rect 6485 11725 6515 11755
rect 6645 11725 6675 11755
rect 6805 11725 6835 11755
rect 6965 11725 6995 11755
rect 7125 11725 7155 11755
rect 7285 11725 7315 11755
rect 7365 11725 7395 11755
rect 7525 11725 7555 11755
rect 7685 11725 7715 11755
rect 5525 11645 5555 11675
rect 5685 11645 5715 11675
rect 5845 11645 5875 11675
rect 6005 11645 6035 11675
rect 6165 11645 6195 11675
rect 6325 11645 6355 11675
rect 6485 11645 6515 11675
rect 6645 11645 6675 11675
rect 6805 11645 6835 11675
rect 6965 11645 6995 11675
rect 7125 11645 7155 11675
rect 7285 11645 7315 11675
rect 7365 11645 7395 11675
rect 7525 11645 7555 11675
rect 7685 11645 7715 11675
rect 5525 11565 5555 11595
rect 5685 11565 5715 11595
rect 5845 11565 5875 11595
rect 6005 11565 6035 11595
rect 6165 11565 6195 11595
rect 6325 11565 6355 11595
rect 6485 11565 6515 11595
rect 6645 11565 6675 11595
rect 6805 11565 6835 11595
rect 6965 11565 6995 11595
rect 7125 11565 7155 11595
rect 7285 11565 7315 11595
rect 7365 11565 7395 11595
rect 7525 11565 7555 11595
rect 7685 11565 7715 11595
rect 5525 11485 5555 11515
rect 5685 11485 5715 11515
rect 5845 11485 5875 11515
rect 6005 11485 6035 11515
rect 6165 11485 6195 11515
rect 6325 11485 6355 11515
rect 6485 11485 6515 11515
rect 6645 11485 6675 11515
rect 6805 11485 6835 11515
rect 6965 11485 6995 11515
rect 7125 11485 7155 11515
rect 7285 11485 7315 11515
rect 7365 11485 7395 11515
rect 7525 11485 7555 11515
rect 7685 11485 7715 11515
rect 5525 11405 5555 11435
rect 5685 11405 5715 11435
rect 5845 11405 5875 11435
rect 6005 11405 6035 11435
rect 6165 11405 6195 11435
rect 6325 11405 6355 11435
rect 6485 11405 6515 11435
rect 6645 11405 6675 11435
rect 6805 11405 6835 11435
rect 6965 11405 6995 11435
rect 7125 11405 7155 11435
rect 7285 11405 7315 11435
rect 7365 11405 7395 11435
rect 7525 11405 7555 11435
rect 7685 11405 7715 11435
rect 5525 11325 5555 11355
rect 5685 11325 5715 11355
rect 5845 11325 5875 11355
rect 6005 11325 6035 11355
rect 6165 11325 6195 11355
rect 6325 11325 6355 11355
rect 6485 11325 6515 11355
rect 6645 11325 6675 11355
rect 6805 11325 6835 11355
rect 6965 11325 6995 11355
rect 7125 11325 7155 11355
rect 7285 11325 7315 11355
rect 7365 11325 7395 11355
rect 7525 11325 7555 11355
rect 7685 11325 7715 11355
rect 7205 11245 7235 11275
rect 7365 11245 7395 11275
rect 7525 11245 7555 11275
rect 7685 11245 7715 11275
rect 5525 11165 5555 11195
rect 5685 11165 5715 11195
rect 5845 11165 5875 11195
rect 6005 11165 6035 11195
rect 6165 11165 6195 11195
rect 6325 11165 6355 11195
rect 6485 11165 6515 11195
rect 6645 11165 6675 11195
rect 6805 11165 6835 11195
rect 6965 11165 6995 11195
rect 7125 11165 7155 11195
rect 7285 11165 7315 11195
rect 7365 11165 7395 11195
rect 7525 11165 7555 11195
rect 7685 11165 7715 11195
rect 5525 11085 5555 11115
rect 5685 11085 5715 11115
rect 5845 11085 5875 11115
rect 6005 11085 6035 11115
rect 6165 11085 6195 11115
rect 6325 11085 6355 11115
rect 6485 11085 6515 11115
rect 6645 11085 6675 11115
rect 6805 11085 6835 11115
rect 6965 11085 6995 11115
rect 7125 11085 7155 11115
rect 7285 11085 7315 11115
rect 7365 11085 7395 11115
rect 7525 11085 7555 11115
rect 7685 11085 7715 11115
rect 5525 11005 5555 11035
rect 5685 11005 5715 11035
rect 5845 11005 5875 11035
rect 6005 11005 6035 11035
rect 6165 11005 6195 11035
rect 6325 11005 6355 11035
rect 6485 11005 6515 11035
rect 6645 11005 6675 11035
rect 6805 11005 6835 11035
rect 6965 11005 6995 11035
rect 7125 11005 7155 11035
rect 7285 11005 7315 11035
rect 7365 11005 7395 11035
rect 7525 11005 7555 11035
rect 7685 11005 7715 11035
rect 7205 10925 7235 10955
rect 7365 10925 7395 10955
rect 7525 10925 7555 10955
rect 7685 10925 7715 10955
rect 5525 10845 5555 10875
rect 5685 10845 5715 10875
rect 5845 10845 5875 10875
rect 6005 10845 6035 10875
rect 6165 10845 6195 10875
rect 6325 10845 6355 10875
rect 6485 10845 6515 10875
rect 6645 10845 6675 10875
rect 6805 10845 6835 10875
rect 6965 10845 6995 10875
rect 7125 10845 7155 10875
rect 7285 10845 7315 10875
rect 7365 10845 7395 10875
rect 7525 10845 7555 10875
rect 7685 10845 7715 10875
rect 7045 10765 7075 10795
rect 7125 10765 7155 10795
rect 7285 10765 7315 10795
rect 7365 10765 7395 10795
rect 7525 10765 7555 10795
rect 7685 10765 7715 10795
rect 5525 10685 5555 10715
rect 5685 10685 5715 10715
rect 5845 10685 5875 10715
rect 6005 10685 6035 10715
rect 6165 10685 6195 10715
rect 6325 10685 6355 10715
rect 6485 10685 6515 10715
rect 6645 10685 6675 10715
rect 6805 10685 6835 10715
rect 6965 10685 6995 10715
rect 7125 10685 7155 10715
rect 7285 10685 7315 10715
rect 7365 10685 7395 10715
rect 7525 10685 7555 10715
rect 7685 10685 7715 10715
rect 5525 10605 5555 10635
rect 5685 10605 5715 10635
rect 5845 10605 5875 10635
rect 6005 10605 6035 10635
rect 6165 10605 6195 10635
rect 6325 10605 6355 10635
rect 6485 10605 6515 10635
rect 6645 10605 6675 10635
rect 6805 10605 6835 10635
rect 6965 10605 6995 10635
rect 7125 10605 7155 10635
rect 7285 10605 7315 10635
rect 7365 10605 7395 10635
rect 7525 10605 7555 10635
rect 7685 10605 7715 10635
rect 7045 10525 7075 10555
rect 7125 10525 7155 10555
rect 7285 10525 7315 10555
rect 7365 10525 7395 10555
rect 7525 10525 7555 10555
rect 7685 10525 7715 10555
rect 5525 10445 5555 10475
rect 5685 10445 5715 10475
rect 5845 10445 5875 10475
rect 6005 10445 6035 10475
rect 6165 10445 6195 10475
rect 6325 10445 6355 10475
rect 6485 10445 6515 10475
rect 6645 10445 6675 10475
rect 6805 10445 6835 10475
rect 6965 10445 6995 10475
rect 7125 10445 7155 10475
rect 7285 10445 7315 10475
rect 7365 10445 7395 10475
rect 7525 10445 7555 10475
rect 7685 10445 7715 10475
rect 6885 10365 6915 10395
rect 6965 10365 6995 10395
rect 7125 10365 7155 10395
rect 7285 10365 7315 10395
rect 7365 10365 7395 10395
rect 7525 10365 7555 10395
rect 7685 10365 7715 10395
rect 5525 10285 5555 10315
rect 5685 10285 5715 10315
rect 5845 10285 5875 10315
rect 6005 10285 6035 10315
rect 6165 10285 6195 10315
rect 6325 10285 6355 10315
rect 6485 10285 6515 10315
rect 6645 10285 6675 10315
rect 6805 10285 6835 10315
rect 6965 10285 6995 10315
rect 7125 10285 7155 10315
rect 7285 10285 7315 10315
rect 7365 10285 7395 10315
rect 7525 10285 7555 10315
rect 7685 10285 7715 10315
rect 5525 10205 5555 10235
rect 5685 10205 5715 10235
rect 5845 10205 5875 10235
rect 6005 10205 6035 10235
rect 6165 10205 6195 10235
rect 6325 10205 6355 10235
rect 6485 10205 6515 10235
rect 6645 10205 6675 10235
rect 6805 10205 6835 10235
rect 6965 10205 6995 10235
rect 7125 10205 7155 10235
rect 7285 10205 7315 10235
rect 7365 10205 7395 10235
rect 7525 10205 7555 10235
rect 7685 10205 7715 10235
rect 5525 10125 5555 10155
rect 5685 10125 5715 10155
rect 5845 10125 5875 10155
rect 6005 10125 6035 10155
rect 6165 10125 6195 10155
rect 6325 10125 6355 10155
rect 6485 10125 6515 10155
rect 6645 10125 6675 10155
rect 6805 10125 6835 10155
rect 6965 10125 6995 10155
rect 7125 10125 7155 10155
rect 7285 10125 7315 10155
rect 7365 10125 7395 10155
rect 7525 10125 7555 10155
rect 7685 10125 7715 10155
rect 5525 10045 5555 10075
rect 5685 10045 5715 10075
rect 5845 10045 5875 10075
rect 6005 10045 6035 10075
rect 6165 10045 6195 10075
rect 6325 10045 6355 10075
rect 6485 10045 6515 10075
rect 6645 10045 6675 10075
rect 6805 10045 6835 10075
rect 6965 10045 6995 10075
rect 7125 10045 7155 10075
rect 7285 10045 7315 10075
rect 7365 10045 7395 10075
rect 7525 10045 7555 10075
rect 7685 10045 7715 10075
rect 5525 9965 5555 9995
rect 5685 9965 5715 9995
rect 5845 9965 5875 9995
rect 6005 9965 6035 9995
rect 6165 9965 6195 9995
rect 6325 9965 6355 9995
rect 6485 9965 6515 9995
rect 6645 9965 6675 9995
rect 6805 9965 6835 9995
rect 6965 9965 6995 9995
rect 7125 9965 7155 9995
rect 7285 9965 7315 9995
rect 7365 9965 7395 9995
rect 7525 9965 7555 9995
rect 7685 9965 7715 9995
rect 5525 9885 5555 9915
rect 5685 9885 5715 9915
rect 5845 9885 5875 9915
rect 6005 9885 6035 9915
rect 6165 9885 6195 9915
rect 6325 9885 6355 9915
rect 6485 9885 6515 9915
rect 6645 9885 6675 9915
rect 6805 9885 6835 9915
rect 6965 9885 6995 9915
rect 7125 9885 7155 9915
rect 7285 9885 7315 9915
rect 7365 9885 7395 9915
rect 7525 9885 7555 9915
rect 7685 9885 7715 9915
rect 5525 9805 5555 9835
rect 5685 9805 5715 9835
rect 5845 9805 5875 9835
rect 6005 9805 6035 9835
rect 6165 9805 6195 9835
rect 6325 9805 6355 9835
rect 6485 9805 6515 9835
rect 6645 9805 6675 9835
rect 6805 9805 6835 9835
rect 6965 9805 6995 9835
rect 7125 9805 7155 9835
rect 7285 9805 7315 9835
rect 7365 9805 7395 9835
rect 7525 9805 7555 9835
rect 7685 9805 7715 9835
rect 5525 9725 5555 9755
rect 5685 9725 5715 9755
rect 5845 9725 5875 9755
rect 6005 9725 6035 9755
rect 6165 9725 6195 9755
rect 6325 9725 6355 9755
rect 6485 9725 6515 9755
rect 6645 9725 6675 9755
rect 6805 9725 6835 9755
rect 6965 9725 6995 9755
rect 7125 9725 7155 9755
rect 7285 9725 7315 9755
rect 7365 9725 7395 9755
rect 7525 9725 7555 9755
rect 7685 9725 7715 9755
rect 5525 9645 5555 9675
rect 5685 9645 5715 9675
rect 5845 9645 5875 9675
rect 6005 9645 6035 9675
rect 6165 9645 6195 9675
rect 6325 9645 6355 9675
rect 6485 9645 6515 9675
rect 6645 9645 6675 9675
rect 6805 9645 6835 9675
rect 6965 9645 6995 9675
rect 7125 9645 7155 9675
rect 7285 9645 7315 9675
rect 7365 9645 7395 9675
rect 7525 9645 7555 9675
rect 7685 9645 7715 9675
rect 5525 9565 5555 9595
rect 5685 9565 5715 9595
rect 5845 9565 5875 9595
rect 6005 9565 6035 9595
rect 6165 9565 6195 9595
rect 6325 9565 6355 9595
rect 6485 9565 6515 9595
rect 6645 9565 6675 9595
rect 6805 9565 6835 9595
rect 6965 9565 6995 9595
rect 7125 9565 7155 9595
rect 7285 9565 7315 9595
rect 7365 9565 7395 9595
rect 7525 9565 7555 9595
rect 7685 9565 7715 9595
rect 5525 9485 5555 9515
rect 5685 9485 5715 9515
rect 5845 9485 5875 9515
rect 6005 9485 6035 9515
rect 6165 9485 6195 9515
rect 6325 9485 6355 9515
rect 6485 9485 6515 9515
rect 6645 9485 6675 9515
rect 6805 9485 6835 9515
rect 6965 9485 6995 9515
rect 7125 9485 7155 9515
rect 7285 9485 7315 9515
rect 7365 9485 7395 9515
rect 7525 9485 7555 9515
rect 7685 9485 7715 9515
rect 5525 9405 5555 9435
rect 5685 9405 5715 9435
rect 5845 9405 5875 9435
rect 6005 9405 6035 9435
rect 6165 9405 6195 9435
rect 6325 9405 6355 9435
rect 6485 9405 6515 9435
rect 6645 9405 6675 9435
rect 6805 9405 6835 9435
rect 6965 9405 6995 9435
rect 7125 9405 7155 9435
rect 7285 9405 7315 9435
rect 7365 9405 7395 9435
rect 7525 9405 7555 9435
rect 7685 9405 7715 9435
rect 5525 9325 5555 9355
rect 5685 9325 5715 9355
rect 5845 9325 5875 9355
rect 6005 9325 6035 9355
rect 6165 9325 6195 9355
rect 6325 9325 6355 9355
rect 6485 9325 6515 9355
rect 6645 9325 6675 9355
rect 6805 9325 6835 9355
rect 6965 9325 6995 9355
rect 7125 9325 7155 9355
rect 7285 9325 7315 9355
rect 7365 9325 7395 9355
rect 7525 9325 7555 9355
rect 7685 9325 7715 9355
rect 5525 9245 5555 9275
rect 5685 9245 5715 9275
rect 5845 9245 5875 9275
rect 6005 9245 6035 9275
rect 6165 9245 6195 9275
rect 6325 9245 6355 9275
rect 6485 9245 6515 9275
rect 6645 9245 6675 9275
rect 6805 9245 6835 9275
rect 6965 9245 6995 9275
rect 7125 9245 7155 9275
rect 7285 9245 7315 9275
rect 7365 9245 7395 9275
rect 7525 9245 7555 9275
rect 7685 9245 7715 9275
rect 7205 9165 7235 9195
rect 7365 9165 7395 9195
rect 7525 9165 7555 9195
rect 7685 9165 7715 9195
rect 5525 9085 5555 9115
rect 5685 9085 5715 9115
rect 5845 9085 5875 9115
rect 6005 9085 6035 9115
rect 6165 9085 6195 9115
rect 6325 9085 6355 9115
rect 6485 9085 6515 9115
rect 6645 9085 6675 9115
rect 6805 9085 6835 9115
rect 6965 9085 6995 9115
rect 7125 9085 7155 9115
rect 7285 9085 7315 9115
rect 7365 9085 7395 9115
rect 7525 9085 7555 9115
rect 7685 9085 7715 9115
rect 5525 9005 5555 9035
rect 5685 9005 5715 9035
rect 5845 9005 5875 9035
rect 6005 9005 6035 9035
rect 6165 9005 6195 9035
rect 6325 9005 6355 9035
rect 6485 9005 6515 9035
rect 6645 9005 6675 9035
rect 6805 9005 6835 9035
rect 6965 9005 6995 9035
rect 7125 9005 7155 9035
rect 7285 9005 7315 9035
rect 7365 9005 7395 9035
rect 7525 9005 7555 9035
rect 7685 9005 7715 9035
rect 5525 8925 5555 8955
rect 5685 8925 5715 8955
rect 5845 8925 5875 8955
rect 6005 8925 6035 8955
rect 6165 8925 6195 8955
rect 6325 8925 6355 8955
rect 6485 8925 6515 8955
rect 6645 8925 6675 8955
rect 6805 8925 6835 8955
rect 6965 8925 6995 8955
rect 7125 8925 7155 8955
rect 7285 8925 7315 8955
rect 7365 8925 7395 8955
rect 7525 8925 7555 8955
rect 7685 8925 7715 8955
rect 7605 8845 7635 8875
rect 7365 8765 7395 8795
rect 7525 8765 7555 8795
rect 7685 8765 7715 8795
rect 7445 8685 7475 8715
rect 5525 8605 5555 8635
rect 5685 8605 5715 8635
rect 5845 8605 5875 8635
rect 6005 8605 6035 8635
rect 6165 8605 6195 8635
rect 6325 8605 6355 8635
rect 6485 8605 6515 8635
rect 6645 8605 6675 8635
rect 6805 8605 6835 8635
rect 6965 8605 6995 8635
rect 7125 8605 7155 8635
rect 7285 8605 7315 8635
rect 7365 8605 7395 8635
rect 7525 8605 7555 8635
rect 7685 8605 7715 8635
rect 5525 8525 5555 8555
rect 5685 8525 5715 8555
rect 5845 8525 5875 8555
rect 6005 8525 6035 8555
rect 6165 8525 6195 8555
rect 6325 8525 6355 8555
rect 6485 8525 6515 8555
rect 6645 8525 6675 8555
rect 6805 8525 6835 8555
rect 6965 8525 6995 8555
rect 7125 8525 7155 8555
rect 7285 8525 7315 8555
rect 7365 8525 7395 8555
rect 7525 8525 7555 8555
rect 7685 8525 7715 8555
rect 7045 8445 7075 8475
rect 7125 8445 7155 8475
rect 7285 8445 7315 8475
rect 7365 8445 7395 8475
rect 7525 8445 7555 8475
rect 7685 8445 7715 8475
rect 5525 8365 5555 8395
rect 5685 8365 5715 8395
rect 5845 8365 5875 8395
rect 6005 8365 6035 8395
rect 6165 8365 6195 8395
rect 6325 8365 6355 8395
rect 6485 8365 6515 8395
rect 6645 8365 6675 8395
rect 6805 8365 6835 8395
rect 6965 8365 6995 8395
rect 7125 8365 7155 8395
rect 7285 8365 7315 8395
rect 7365 8365 7395 8395
rect 7525 8365 7555 8395
rect 7685 8365 7715 8395
rect 6725 8285 6755 8315
rect 6805 8285 6835 8315
rect 6965 8285 6995 8315
rect 7125 8285 7155 8315
rect 7285 8285 7315 8315
rect 7365 8285 7395 8315
rect 7525 8285 7555 8315
rect 7685 8285 7715 8315
rect 5525 8205 5555 8235
rect 5685 8205 5715 8235
rect 5845 8205 5875 8235
rect 6005 8205 6035 8235
rect 6165 8205 6195 8235
rect 6325 8205 6355 8235
rect 6485 8205 6515 8235
rect 6645 8205 6675 8235
rect 6805 8205 6835 8235
rect 6965 8205 6995 8235
rect 7125 8205 7155 8235
rect 7285 8205 7315 8235
rect 7365 8205 7395 8235
rect 7525 8205 7555 8235
rect 7685 8205 7715 8235
rect 5525 8125 5555 8155
rect 5685 8125 5715 8155
rect 5845 8125 5875 8155
rect 6005 8125 6035 8155
rect 6165 8125 6195 8155
rect 6325 8125 6355 8155
rect 6485 8125 6515 8155
rect 6645 8125 6675 8155
rect 6805 8125 6835 8155
rect 6965 8125 6995 8155
rect 7125 8125 7155 8155
rect 7285 8125 7315 8155
rect 7365 8125 7395 8155
rect 7525 8125 7555 8155
rect 7685 8125 7715 8155
rect 5525 8045 5555 8075
rect 5685 8045 5715 8075
rect 5845 8045 5875 8075
rect 6005 8045 6035 8075
rect 6165 8045 6195 8075
rect 6325 8045 6355 8075
rect 6485 8045 6515 8075
rect 6645 8045 6675 8075
rect 6805 8045 6835 8075
rect 6965 8045 6995 8075
rect 7125 8045 7155 8075
rect 7285 8045 7315 8075
rect 7365 8045 7395 8075
rect 7525 8045 7555 8075
rect 7685 8045 7715 8075
rect 5525 7965 5555 7995
rect 5685 7965 5715 7995
rect 5845 7965 5875 7995
rect 6005 7965 6035 7995
rect 6165 7965 6195 7995
rect 6325 7965 6355 7995
rect 6485 7965 6515 7995
rect 6645 7965 6675 7995
rect 6805 7965 6835 7995
rect 6965 7965 6995 7995
rect 7125 7965 7155 7995
rect 7285 7965 7315 7995
rect 7365 7965 7395 7995
rect 7525 7965 7555 7995
rect 7685 7965 7715 7995
rect 5525 7885 5555 7915
rect 5685 7885 5715 7915
rect 5845 7885 5875 7915
rect 6005 7885 6035 7915
rect 6165 7885 6195 7915
rect 6325 7885 6355 7915
rect 6485 7885 6515 7915
rect 6645 7885 6675 7915
rect 6805 7885 6835 7915
rect 6965 7885 6995 7915
rect 7125 7885 7155 7915
rect 7285 7885 7315 7915
rect 7365 7885 7395 7915
rect 7525 7885 7555 7915
rect 7685 7885 7715 7915
rect 5525 7805 5555 7835
rect 5685 7805 5715 7835
rect 5845 7805 5875 7835
rect 6005 7805 6035 7835
rect 6165 7805 6195 7835
rect 6325 7805 6355 7835
rect 6485 7805 6515 7835
rect 6645 7805 6675 7835
rect 6805 7805 6835 7835
rect 6965 7805 6995 7835
rect 7125 7805 7155 7835
rect 7285 7805 7315 7835
rect 7365 7805 7395 7835
rect 7525 7805 7555 7835
rect 7685 7805 7715 7835
rect 5525 7725 5555 7755
rect 5685 7725 5715 7755
rect 5845 7725 5875 7755
rect 6005 7725 6035 7755
rect 6165 7725 6195 7755
rect 6325 7725 6355 7755
rect 6485 7725 6515 7755
rect 6645 7725 6675 7755
rect 6805 7725 6835 7755
rect 6965 7725 6995 7755
rect 7125 7725 7155 7755
rect 7285 7725 7315 7755
rect 7365 7725 7395 7755
rect 7525 7725 7555 7755
rect 7685 7725 7715 7755
rect 5525 7645 5555 7675
rect 5685 7645 5715 7675
rect 5845 7645 5875 7675
rect 6005 7645 6035 7675
rect 6165 7645 6195 7675
rect 6325 7645 6355 7675
rect 6485 7645 6515 7675
rect 6645 7645 6675 7675
rect 6805 7645 6835 7675
rect 6965 7645 6995 7675
rect 7125 7645 7155 7675
rect 7285 7645 7315 7675
rect 7365 7645 7395 7675
rect 7525 7645 7555 7675
rect 7685 7645 7715 7675
rect 5525 7565 5555 7595
rect 5685 7565 5715 7595
rect 5845 7565 5875 7595
rect 6005 7565 6035 7595
rect 6165 7565 6195 7595
rect 6325 7565 6355 7595
rect 6485 7565 6515 7595
rect 6645 7565 6675 7595
rect 6805 7565 6835 7595
rect 6965 7565 6995 7595
rect 7125 7565 7155 7595
rect 7285 7565 7315 7595
rect 7365 7565 7395 7595
rect 7525 7565 7555 7595
rect 7685 7565 7715 7595
rect 5525 7485 5555 7515
rect 5685 7485 5715 7515
rect 5845 7485 5875 7515
rect 6005 7485 6035 7515
rect 6165 7485 6195 7515
rect 6325 7485 6355 7515
rect 6485 7485 6515 7515
rect 6645 7485 6675 7515
rect 6805 7485 6835 7515
rect 6965 7485 6995 7515
rect 7125 7485 7155 7515
rect 7285 7485 7315 7515
rect 7365 7485 7395 7515
rect 7525 7485 7555 7515
rect 7685 7485 7715 7515
rect 5525 7405 5555 7435
rect 5685 7405 5715 7435
rect 5845 7405 5875 7435
rect 6005 7405 6035 7435
rect 6165 7405 6195 7435
rect 6325 7405 6355 7435
rect 6485 7405 6515 7435
rect 6645 7405 6675 7435
rect 6805 7405 6835 7435
rect 6965 7405 6995 7435
rect 7125 7405 7155 7435
rect 7285 7405 7315 7435
rect 7365 7405 7395 7435
rect 7525 7405 7555 7435
rect 7685 7405 7715 7435
rect 5525 7325 5555 7355
rect 5685 7325 5715 7355
rect 5845 7325 5875 7355
rect 6005 7325 6035 7355
rect 6165 7325 6195 7355
rect 6325 7325 6355 7355
rect 6485 7325 6515 7355
rect 6645 7325 6675 7355
rect 6805 7325 6835 7355
rect 6965 7325 6995 7355
rect 7125 7325 7155 7355
rect 7285 7325 7315 7355
rect 7365 7325 7395 7355
rect 7525 7325 7555 7355
rect 7685 7325 7715 7355
rect 5525 7245 5555 7275
rect 5685 7245 5715 7275
rect 5845 7245 5875 7275
rect 6005 7245 6035 7275
rect 6165 7245 6195 7275
rect 6325 7245 6355 7275
rect 6485 7245 6515 7275
rect 6645 7245 6675 7275
rect 6805 7245 6835 7275
rect 6965 7245 6995 7275
rect 7125 7245 7155 7275
rect 7285 7245 7315 7275
rect 7365 7245 7395 7275
rect 7525 7245 7555 7275
rect 7685 7245 7715 7275
rect 5525 7165 5555 7195
rect 5685 7165 5715 7195
rect 5845 7165 5875 7195
rect 6005 7165 6035 7195
rect 6165 7165 6195 7195
rect 6325 7165 6355 7195
rect 6485 7165 6515 7195
rect 6645 7165 6675 7195
rect 6805 7165 6835 7195
rect 6965 7165 6995 7195
rect 7125 7165 7155 7195
rect 7285 7165 7315 7195
rect 7365 7165 7395 7195
rect 7525 7165 7555 7195
rect 7685 7165 7715 7195
rect 6085 7085 6115 7115
rect 6165 7085 6195 7115
rect 6325 7085 6355 7115
rect 6485 7085 6515 7115
rect 6645 7085 6675 7115
rect 6805 7085 6835 7115
rect 6965 7085 6995 7115
rect 7125 7085 7155 7115
rect 7285 7085 7315 7115
rect 7365 7085 7395 7115
rect 7525 7085 7555 7115
rect 7685 7085 7715 7115
rect 5525 7005 5555 7035
rect 5685 7005 5715 7035
rect 5845 7005 5875 7035
rect 6005 7005 6035 7035
rect 6165 7005 6195 7035
rect 6325 7005 6355 7035
rect 6485 7005 6515 7035
rect 6645 7005 6675 7035
rect 6805 7005 6835 7035
rect 6965 7005 6995 7035
rect 7125 7005 7155 7035
rect 7285 7005 7315 7035
rect 7365 7005 7395 7035
rect 7525 7005 7555 7035
rect 7685 7005 7715 7035
rect 5525 6925 5555 6955
rect 5685 6925 5715 6955
rect 5845 6925 5875 6955
rect 6005 6925 6035 6955
rect 6165 6925 6195 6955
rect 6325 6925 6355 6955
rect 6485 6925 6515 6955
rect 6645 6925 6675 6955
rect 6805 6925 6835 6955
rect 6965 6925 6995 6955
rect 7125 6925 7155 6955
rect 7285 6925 7315 6955
rect 7365 6925 7395 6955
rect 7525 6925 7555 6955
rect 7685 6925 7715 6955
rect 6245 6845 6275 6875
rect 6325 6845 6355 6875
rect 6485 6845 6515 6875
rect 6645 6845 6675 6875
rect 6805 6845 6835 6875
rect 6965 6845 6995 6875
rect 7125 6845 7155 6875
rect 7285 6845 7315 6875
rect 7365 6845 7395 6875
rect 7525 6845 7555 6875
rect 7685 6845 7715 6875
rect 5525 6765 5555 6795
rect 5685 6765 5715 6795
rect 5845 6765 5875 6795
rect 6005 6765 6035 6795
rect 6165 6765 6195 6795
rect 6325 6765 6355 6795
rect 6485 6765 6515 6795
rect 6645 6765 6675 6795
rect 6805 6765 6835 6795
rect 6965 6765 6995 6795
rect 7125 6765 7155 6795
rect 7285 6765 7315 6795
rect 7365 6765 7395 6795
rect 7525 6765 7555 6795
rect 7685 6765 7715 6795
rect 5525 6685 5555 6715
rect 5685 6685 5715 6715
rect 5845 6685 5875 6715
rect 6005 6685 6035 6715
rect 6165 6685 6195 6715
rect 6325 6685 6355 6715
rect 6485 6685 6515 6715
rect 6645 6685 6675 6715
rect 6805 6685 6835 6715
rect 6965 6685 6995 6715
rect 7125 6685 7155 6715
rect 7285 6685 7315 6715
rect 7365 6685 7395 6715
rect 7525 6685 7555 6715
rect 7685 6685 7715 6715
rect 5525 6605 5555 6635
rect 5685 6605 5715 6635
rect 5845 6605 5875 6635
rect 6005 6605 6035 6635
rect 6165 6605 6195 6635
rect 6325 6605 6355 6635
rect 6485 6605 6515 6635
rect 6645 6605 6675 6635
rect 6805 6605 6835 6635
rect 6965 6605 6995 6635
rect 7125 6605 7155 6635
rect 7285 6605 7315 6635
rect 7365 6605 7395 6635
rect 7525 6605 7555 6635
rect 7685 6605 7715 6635
rect 5525 6525 5555 6555
rect 5685 6525 5715 6555
rect 5845 6525 5875 6555
rect 6005 6525 6035 6555
rect 6165 6525 6195 6555
rect 6325 6525 6355 6555
rect 6485 6525 6515 6555
rect 6645 6525 6675 6555
rect 6805 6525 6835 6555
rect 6965 6525 6995 6555
rect 7125 6525 7155 6555
rect 7285 6525 7315 6555
rect 7365 6525 7395 6555
rect 7525 6525 7555 6555
rect 7685 6525 7715 6555
rect 5525 6445 5555 6475
rect 5685 6445 5715 6475
rect 5845 6445 5875 6475
rect 6005 6445 6035 6475
rect 6165 6445 6195 6475
rect 6325 6445 6355 6475
rect 6485 6445 6515 6475
rect 6645 6445 6675 6475
rect 6805 6445 6835 6475
rect 6965 6445 6995 6475
rect 7125 6445 7155 6475
rect 7285 6445 7315 6475
rect 7365 6445 7395 6475
rect 7525 6445 7555 6475
rect 7685 6445 7715 6475
rect 6565 6365 6595 6395
rect 6645 6365 6675 6395
rect 6805 6365 6835 6395
rect 6965 6365 6995 6395
rect 7125 6365 7155 6395
rect 7285 6365 7315 6395
rect 7365 6365 7395 6395
rect 7525 6365 7555 6395
rect 7685 6365 7715 6395
rect 5525 6285 5555 6315
rect 5685 6285 5715 6315
rect 5845 6285 5875 6315
rect 6005 6285 6035 6315
rect 6165 6285 6195 6315
rect 6325 6285 6355 6315
rect 6485 6285 6515 6315
rect 6645 6285 6675 6315
rect 6805 6285 6835 6315
rect 6965 6285 6995 6315
rect 7125 6285 7155 6315
rect 7285 6285 7315 6315
rect 7365 6285 7395 6315
rect 7525 6285 7555 6315
rect 7685 6285 7715 6315
rect 5525 6205 5555 6235
rect 5685 6205 5715 6235
rect 5845 6205 5875 6235
rect 6005 6205 6035 6235
rect 6165 6205 6195 6235
rect 6325 6205 6355 6235
rect 6485 6205 6515 6235
rect 6645 6205 6675 6235
rect 6805 6205 6835 6235
rect 6965 6205 6995 6235
rect 7125 6205 7155 6235
rect 7285 6205 7315 6235
rect 7365 6205 7395 6235
rect 7525 6205 7555 6235
rect 7685 6205 7715 6235
rect 5525 6125 5555 6155
rect 5685 6125 5715 6155
rect 5845 6125 5875 6155
rect 6005 6125 6035 6155
rect 6165 6125 6195 6155
rect 6325 6125 6355 6155
rect 6485 6125 6515 6155
rect 6645 6125 6675 6155
rect 6805 6125 6835 6155
rect 6965 6125 6995 6155
rect 7125 6125 7155 6155
rect 7285 6125 7315 6155
rect 7365 6125 7395 6155
rect 7525 6125 7555 6155
rect 7685 6125 7715 6155
rect 7045 6045 7075 6075
rect 7125 6045 7155 6075
rect 7285 6045 7315 6075
rect 7365 6045 7395 6075
rect 7525 6045 7555 6075
rect 7685 6045 7715 6075
rect 5525 5965 5555 5995
rect 5685 5965 5715 5995
rect 5845 5965 5875 5995
rect 6005 5965 6035 5995
rect 6165 5965 6195 5995
rect 6325 5965 6355 5995
rect 6485 5965 6515 5995
rect 6645 5965 6675 5995
rect 6805 5965 6835 5995
rect 6965 5965 6995 5995
rect 7125 5965 7155 5995
rect 7285 5965 7315 5995
rect 7365 5965 7395 5995
rect 7525 5965 7555 5995
rect 7685 5965 7715 5995
rect 6885 5885 6915 5915
rect 6965 5885 6995 5915
rect 7125 5885 7155 5915
rect 7285 5885 7315 5915
rect 7365 5885 7395 5915
rect 7525 5885 7555 5915
rect 7685 5885 7715 5915
rect 5525 5805 5555 5835
rect 5685 5805 5715 5835
rect 5845 5805 5875 5835
rect 6005 5805 6035 5835
rect 6165 5805 6195 5835
rect 6325 5805 6355 5835
rect 6485 5805 6515 5835
rect 6645 5805 6675 5835
rect 6805 5805 6835 5835
rect 6965 5805 6995 5835
rect 7125 5805 7155 5835
rect 7285 5805 7315 5835
rect 7365 5805 7395 5835
rect 7525 5805 7555 5835
rect 7685 5805 7715 5835
rect 5525 5725 5555 5755
rect 5685 5725 5715 5755
rect 5845 5725 5875 5755
rect 6005 5725 6035 5755
rect 6165 5725 6195 5755
rect 6325 5725 6355 5755
rect 6485 5725 6515 5755
rect 6645 5725 6675 5755
rect 6805 5725 6835 5755
rect 6965 5725 6995 5755
rect 7125 5725 7155 5755
rect 7285 5725 7315 5755
rect 7365 5725 7395 5755
rect 7525 5725 7555 5755
rect 7685 5725 7715 5755
rect 5525 5645 5555 5675
rect 5685 5645 5715 5675
rect 5845 5645 5875 5675
rect 6005 5645 6035 5675
rect 6165 5645 6195 5675
rect 6325 5645 6355 5675
rect 6485 5645 6515 5675
rect 6645 5645 6675 5675
rect 6805 5645 6835 5675
rect 6965 5645 6995 5675
rect 7125 5645 7155 5675
rect 7285 5645 7315 5675
rect 7365 5645 7395 5675
rect 7525 5645 7555 5675
rect 7685 5645 7715 5675
rect 5525 5565 5555 5595
rect 5685 5565 5715 5595
rect 5845 5565 5875 5595
rect 6005 5565 6035 5595
rect 6165 5565 6195 5595
rect 6325 5565 6355 5595
rect 6485 5565 6515 5595
rect 6645 5565 6675 5595
rect 6805 5565 6835 5595
rect 6965 5565 6995 5595
rect 7125 5565 7155 5595
rect 7285 5565 7315 5595
rect 7365 5565 7395 5595
rect 7525 5565 7555 5595
rect 7685 5565 7715 5595
rect 5525 5485 5555 5515
rect 5685 5485 5715 5515
rect 5845 5485 5875 5515
rect 6005 5485 6035 5515
rect 6165 5485 6195 5515
rect 6325 5485 6355 5515
rect 6485 5485 6515 5515
rect 6645 5485 6675 5515
rect 6805 5485 6835 5515
rect 6965 5485 6995 5515
rect 7125 5485 7155 5515
rect 7285 5485 7315 5515
rect 7365 5485 7395 5515
rect 7525 5485 7555 5515
rect 7685 5485 7715 5515
rect 5525 5405 5555 5435
rect 5685 5405 5715 5435
rect 5845 5405 5875 5435
rect 6005 5405 6035 5435
rect 6165 5405 6195 5435
rect 6325 5405 6355 5435
rect 6485 5405 6515 5435
rect 6645 5405 6675 5435
rect 6805 5405 6835 5435
rect 6965 5405 6995 5435
rect 7125 5405 7155 5435
rect 7285 5405 7315 5435
rect 7365 5405 7395 5435
rect 7525 5405 7555 5435
rect 7685 5405 7715 5435
rect 5525 5325 5555 5355
rect 5685 5325 5715 5355
rect 5845 5325 5875 5355
rect 6005 5325 6035 5355
rect 6165 5325 6195 5355
rect 6325 5325 6355 5355
rect 6485 5325 6515 5355
rect 6645 5325 6675 5355
rect 6805 5325 6835 5355
rect 6965 5325 6995 5355
rect 7125 5325 7155 5355
rect 7285 5325 7315 5355
rect 7365 5325 7395 5355
rect 7525 5325 7555 5355
rect 7685 5325 7715 5355
rect 5525 5245 5555 5275
rect 5685 5245 5715 5275
rect 5845 5245 5875 5275
rect 6005 5245 6035 5275
rect 6165 5245 6195 5275
rect 6325 5245 6355 5275
rect 6485 5245 6515 5275
rect 6645 5245 6675 5275
rect 6805 5245 6835 5275
rect 6965 5245 6995 5275
rect 7125 5245 7155 5275
rect 7285 5245 7315 5275
rect 7365 5245 7395 5275
rect 7525 5245 7555 5275
rect 7685 5245 7715 5275
rect 5525 5165 5555 5195
rect 5685 5165 5715 5195
rect 5845 5165 5875 5195
rect 6005 5165 6035 5195
rect 6165 5165 6195 5195
rect 6325 5165 6355 5195
rect 6485 5165 6515 5195
rect 6645 5165 6675 5195
rect 6805 5165 6835 5195
rect 6965 5165 6995 5195
rect 7125 5165 7155 5195
rect 7285 5165 7315 5195
rect 7365 5165 7395 5195
rect 7525 5165 7555 5195
rect 7685 5165 7715 5195
rect 5525 5085 5555 5115
rect 5685 5085 5715 5115
rect 5845 5085 5875 5115
rect 6005 5085 6035 5115
rect 6165 5085 6195 5115
rect 6325 5085 6355 5115
rect 6485 5085 6515 5115
rect 6645 5085 6675 5115
rect 6805 5085 6835 5115
rect 6965 5085 6995 5115
rect 7125 5085 7155 5115
rect 7285 5085 7315 5115
rect 7365 5085 7395 5115
rect 7525 5085 7555 5115
rect 7685 5085 7715 5115
rect 5525 5005 5555 5035
rect 5685 5005 5715 5035
rect 5845 5005 5875 5035
rect 6005 5005 6035 5035
rect 6165 5005 6195 5035
rect 6325 5005 6355 5035
rect 6485 5005 6515 5035
rect 6645 5005 6675 5035
rect 6805 5005 6835 5035
rect 6965 5005 6995 5035
rect 7125 5005 7155 5035
rect 7285 5005 7315 5035
rect 7365 5005 7395 5035
rect 7525 5005 7555 5035
rect 7685 5005 7715 5035
rect 5525 4925 5555 4955
rect 5685 4925 5715 4955
rect 5845 4925 5875 4955
rect 6005 4925 6035 4955
rect 6165 4925 6195 4955
rect 6325 4925 6355 4955
rect 6485 4925 6515 4955
rect 6645 4925 6675 4955
rect 6805 4925 6835 4955
rect 6965 4925 6995 4955
rect 7125 4925 7155 4955
rect 7285 4925 7315 4955
rect 7365 4925 7395 4955
rect 7525 4925 7555 4955
rect 7685 4925 7715 4955
rect 5525 4845 5555 4875
rect 5685 4845 5715 4875
rect 5845 4845 5875 4875
rect 6005 4845 6035 4875
rect 6165 4845 6195 4875
rect 6325 4845 6355 4875
rect 6485 4845 6515 4875
rect 6645 4845 6675 4875
rect 6805 4845 6835 4875
rect 6965 4845 6995 4875
rect 7125 4845 7155 4875
rect 7285 4845 7315 4875
rect 7365 4845 7395 4875
rect 7525 4845 7555 4875
rect 7685 4845 7715 4875
rect 5525 4765 5555 4795
rect 5685 4765 5715 4795
rect 5845 4765 5875 4795
rect 6005 4765 6035 4795
rect 6165 4765 6195 4795
rect 6325 4765 6355 4795
rect 6485 4765 6515 4795
rect 6645 4765 6675 4795
rect 6805 4765 6835 4795
rect 6965 4765 6995 4795
rect 7125 4765 7155 4795
rect 7285 4765 7315 4795
rect 7365 4765 7395 4795
rect 7525 4765 7555 4795
rect 7685 4765 7715 4795
rect 6085 4685 6115 4715
rect 6165 4685 6195 4715
rect 6325 4685 6355 4715
rect 6485 4685 6515 4715
rect 6645 4685 6675 4715
rect 6805 4685 6835 4715
rect 6965 4685 6995 4715
rect 7125 4685 7155 4715
rect 7285 4685 7315 4715
rect 7365 4685 7395 4715
rect 7525 4685 7555 4715
rect 7685 4685 7715 4715
rect 5525 4605 5555 4635
rect 5685 4605 5715 4635
rect 5845 4605 5875 4635
rect 6005 4605 6035 4635
rect 6165 4605 6195 4635
rect 6325 4605 6355 4635
rect 6485 4605 6515 4635
rect 6645 4605 6675 4635
rect 6805 4605 6835 4635
rect 6965 4605 6995 4635
rect 7125 4605 7155 4635
rect 7285 4605 7315 4635
rect 7365 4605 7395 4635
rect 7525 4605 7555 4635
rect 7685 4605 7715 4635
rect 5525 4525 5555 4555
rect 5685 4525 5715 4555
rect 5845 4525 5875 4555
rect 6005 4525 6035 4555
rect 6165 4525 6195 4555
rect 6325 4525 6355 4555
rect 6485 4525 6515 4555
rect 6645 4525 6675 4555
rect 6805 4525 6835 4555
rect 6965 4525 6995 4555
rect 7125 4525 7155 4555
rect 7285 4525 7315 4555
rect 7365 4525 7395 4555
rect 7525 4525 7555 4555
rect 7685 4525 7715 4555
rect 6245 4445 6275 4475
rect 6325 4445 6355 4475
rect 6485 4445 6515 4475
rect 6645 4445 6675 4475
rect 6805 4445 6835 4475
rect 6965 4445 6995 4475
rect 7125 4445 7155 4475
rect 7285 4445 7315 4475
rect 7365 4445 7395 4475
rect 7525 4445 7555 4475
rect 7685 4445 7715 4475
rect 5525 4365 5555 4395
rect 5685 4365 5715 4395
rect 5845 4365 5875 4395
rect 6005 4365 6035 4395
rect 6165 4365 6195 4395
rect 6325 4365 6355 4395
rect 6485 4365 6515 4395
rect 6645 4365 6675 4395
rect 6805 4365 6835 4395
rect 6965 4365 6995 4395
rect 7125 4365 7155 4395
rect 7285 4365 7315 4395
rect 7365 4365 7395 4395
rect 7525 4365 7555 4395
rect 7685 4365 7715 4395
rect 5525 4285 5555 4315
rect 5685 4285 5715 4315
rect 5845 4285 5875 4315
rect 6005 4285 6035 4315
rect 6165 4285 6195 4315
rect 6325 4285 6355 4315
rect 6485 4285 6515 4315
rect 6645 4285 6675 4315
rect 6805 4285 6835 4315
rect 6965 4285 6995 4315
rect 7125 4285 7155 4315
rect 7285 4285 7315 4315
rect 7365 4285 7395 4315
rect 7525 4285 7555 4315
rect 7685 4285 7715 4315
rect 5525 4205 5555 4235
rect 5685 4205 5715 4235
rect 5845 4205 5875 4235
rect 6005 4205 6035 4235
rect 6165 4205 6195 4235
rect 6325 4205 6355 4235
rect 6485 4205 6515 4235
rect 6645 4205 6675 4235
rect 6805 4205 6835 4235
rect 6965 4205 6995 4235
rect 7125 4205 7155 4235
rect 7285 4205 7315 4235
rect 7365 4205 7395 4235
rect 7525 4205 7555 4235
rect 7685 4205 7715 4235
rect 5525 4125 5555 4155
rect 5685 4125 5715 4155
rect 5845 4125 5875 4155
rect 6005 4125 6035 4155
rect 6165 4125 6195 4155
rect 6325 4125 6355 4155
rect 6485 4125 6515 4155
rect 6645 4125 6675 4155
rect 6805 4125 6835 4155
rect 6965 4125 6995 4155
rect 7125 4125 7155 4155
rect 7285 4125 7315 4155
rect 7365 4125 7395 4155
rect 7525 4125 7555 4155
rect 7685 4125 7715 4155
rect 5525 4045 5555 4075
rect 5685 4045 5715 4075
rect 5845 4045 5875 4075
rect 6005 4045 6035 4075
rect 6165 4045 6195 4075
rect 6325 4045 6355 4075
rect 6485 4045 6515 4075
rect 6645 4045 6675 4075
rect 6805 4045 6835 4075
rect 6965 4045 6995 4075
rect 7125 4045 7155 4075
rect 7285 4045 7315 4075
rect 7365 4045 7395 4075
rect 7525 4045 7555 4075
rect 7685 4045 7715 4075
rect 6405 3965 6435 3995
rect 6485 3965 6515 3995
rect 6645 3965 6675 3995
rect 6805 3965 6835 3995
rect 6965 3965 6995 3995
rect 7125 3965 7155 3995
rect 7285 3965 7315 3995
rect 7365 3965 7395 3995
rect 7525 3965 7555 3995
rect 7685 3965 7715 3995
rect 5525 3885 5555 3915
rect 5685 3885 5715 3915
rect 5845 3885 5875 3915
rect 6005 3885 6035 3915
rect 6165 3885 6195 3915
rect 6325 3885 6355 3915
rect 6485 3885 6515 3915
rect 6645 3885 6675 3915
rect 6805 3885 6835 3915
rect 6965 3885 6995 3915
rect 7125 3885 7155 3915
rect 7285 3885 7315 3915
rect 7365 3885 7395 3915
rect 7525 3885 7555 3915
rect 7685 3885 7715 3915
rect 5525 3805 5555 3835
rect 5685 3805 5715 3835
rect 5845 3805 5875 3835
rect 6005 3805 6035 3835
rect 6165 3805 6195 3835
rect 6325 3805 6355 3835
rect 6485 3805 6515 3835
rect 6645 3805 6675 3835
rect 6805 3805 6835 3835
rect 6965 3805 6995 3835
rect 7125 3805 7155 3835
rect 7285 3805 7315 3835
rect 7365 3805 7395 3835
rect 7525 3805 7555 3835
rect 7685 3805 7715 3835
rect 5525 3725 5555 3755
rect 5685 3725 5715 3755
rect 5845 3725 5875 3755
rect 6005 3725 6035 3755
rect 6165 3725 6195 3755
rect 6325 3725 6355 3755
rect 6485 3725 6515 3755
rect 6645 3725 6675 3755
rect 6805 3725 6835 3755
rect 6965 3725 6995 3755
rect 7125 3725 7155 3755
rect 7285 3725 7315 3755
rect 7365 3725 7395 3755
rect 7525 3725 7555 3755
rect 7685 3725 7715 3755
rect 7045 3645 7075 3675
rect 7125 3645 7155 3675
rect 7285 3645 7315 3675
rect 7365 3645 7395 3675
rect 7525 3645 7555 3675
rect 7685 3645 7715 3675
rect 5525 3565 5555 3595
rect 5685 3565 5715 3595
rect 5845 3565 5875 3595
rect 6005 3565 6035 3595
rect 6165 3565 6195 3595
rect 6325 3565 6355 3595
rect 6485 3565 6515 3595
rect 6645 3565 6675 3595
rect 6805 3565 6835 3595
rect 6965 3565 6995 3595
rect 7125 3565 7155 3595
rect 7285 3565 7315 3595
rect 7365 3565 7395 3595
rect 7525 3565 7555 3595
rect 7685 3565 7715 3595
rect 6725 3485 6755 3515
rect 6805 3485 6835 3515
rect 6965 3485 6995 3515
rect 7125 3485 7155 3515
rect 7285 3485 7315 3515
rect 7365 3485 7395 3515
rect 7525 3485 7555 3515
rect 7685 3485 7715 3515
rect 5525 3405 5555 3435
rect 5685 3405 5715 3435
rect 5845 3405 5875 3435
rect 6005 3405 6035 3435
rect 6165 3405 6195 3435
rect 6325 3405 6355 3435
rect 6485 3405 6515 3435
rect 6645 3405 6675 3435
rect 6805 3405 6835 3435
rect 6965 3405 6995 3435
rect 7125 3405 7155 3435
rect 7285 3405 7315 3435
rect 7365 3405 7395 3435
rect 7525 3405 7555 3435
rect 7685 3405 7715 3435
rect 5525 3325 5555 3355
rect 5685 3325 5715 3355
rect 5845 3325 5875 3355
rect 6005 3325 6035 3355
rect 6165 3325 6195 3355
rect 6325 3325 6355 3355
rect 6485 3325 6515 3355
rect 6645 3325 6675 3355
rect 6805 3325 6835 3355
rect 6965 3325 6995 3355
rect 7125 3325 7155 3355
rect 7285 3325 7315 3355
rect 7365 3325 7395 3355
rect 7525 3325 7555 3355
rect 7685 3325 7715 3355
rect 5525 3245 5555 3275
rect 5685 3245 5715 3275
rect 5845 3245 5875 3275
rect 6005 3245 6035 3275
rect 6165 3245 6195 3275
rect 6325 3245 6355 3275
rect 6485 3245 6515 3275
rect 6645 3245 6675 3275
rect 6805 3245 6835 3275
rect 6965 3245 6995 3275
rect 7125 3245 7155 3275
rect 7285 3245 7315 3275
rect 7365 3245 7395 3275
rect 7525 3245 7555 3275
rect 7685 3245 7715 3275
rect 5525 3165 5555 3195
rect 5685 3165 5715 3195
rect 5845 3165 5875 3195
rect 6005 3165 6035 3195
rect 6165 3165 6195 3195
rect 6325 3165 6355 3195
rect 6485 3165 6515 3195
rect 6645 3165 6675 3195
rect 6805 3165 6835 3195
rect 6965 3165 6995 3195
rect 7125 3165 7155 3195
rect 7285 3165 7315 3195
rect 7365 3165 7395 3195
rect 7525 3165 7555 3195
rect 7685 3165 7715 3195
rect 5525 3085 5555 3115
rect 5685 3085 5715 3115
rect 5845 3085 5875 3115
rect 6005 3085 6035 3115
rect 6165 3085 6195 3115
rect 6325 3085 6355 3115
rect 6485 3085 6515 3115
rect 6645 3085 6675 3115
rect 6805 3085 6835 3115
rect 6965 3085 6995 3115
rect 7125 3085 7155 3115
rect 7285 3085 7315 3115
rect 7365 3085 7395 3115
rect 7525 3085 7555 3115
rect 7685 3085 7715 3115
rect 5525 3005 5555 3035
rect 5685 3005 5715 3035
rect 5845 3005 5875 3035
rect 6005 3005 6035 3035
rect 6165 3005 6195 3035
rect 6325 3005 6355 3035
rect 6485 3005 6515 3035
rect 6645 3005 6675 3035
rect 6805 3005 6835 3035
rect 6965 3005 6995 3035
rect 7125 3005 7155 3035
rect 7285 3005 7315 3035
rect 7365 3005 7395 3035
rect 7525 3005 7555 3035
rect 7685 3005 7715 3035
rect 5525 2925 5555 2955
rect 5685 2925 5715 2955
rect 5845 2925 5875 2955
rect 6005 2925 6035 2955
rect 6165 2925 6195 2955
rect 6325 2925 6355 2955
rect 6485 2925 6515 2955
rect 6645 2925 6675 2955
rect 6805 2925 6835 2955
rect 6965 2925 6995 2955
rect 7125 2925 7155 2955
rect 7285 2925 7315 2955
rect 7365 2925 7395 2955
rect 7525 2925 7555 2955
rect 7685 2925 7715 2955
rect 5525 2845 5555 2875
rect 5685 2845 5715 2875
rect 5845 2845 5875 2875
rect 6005 2845 6035 2875
rect 6165 2845 6195 2875
rect 6325 2845 6355 2875
rect 6485 2845 6515 2875
rect 6645 2845 6675 2875
rect 6805 2845 6835 2875
rect 6965 2845 6995 2875
rect 7125 2845 7155 2875
rect 7285 2845 7315 2875
rect 7365 2845 7395 2875
rect 7525 2845 7555 2875
rect 7685 2845 7715 2875
rect 5525 2765 5555 2795
rect 5685 2765 5715 2795
rect 5845 2765 5875 2795
rect 6005 2765 6035 2795
rect 6165 2765 6195 2795
rect 6325 2765 6355 2795
rect 6485 2765 6515 2795
rect 6645 2765 6675 2795
rect 6805 2765 6835 2795
rect 6965 2765 6995 2795
rect 7125 2765 7155 2795
rect 7285 2765 7315 2795
rect 7365 2765 7395 2795
rect 7525 2765 7555 2795
rect 7685 2765 7715 2795
rect 5525 2685 5555 2715
rect 5685 2685 5715 2715
rect 5845 2685 5875 2715
rect 6005 2685 6035 2715
rect 6165 2685 6195 2715
rect 6325 2685 6355 2715
rect 6485 2685 6515 2715
rect 6645 2685 6675 2715
rect 6805 2685 6835 2715
rect 6965 2685 6995 2715
rect 7125 2685 7155 2715
rect 7285 2685 7315 2715
rect 7365 2685 7395 2715
rect 7525 2685 7555 2715
rect 7685 2685 7715 2715
rect 5525 2605 5555 2635
rect 5685 2605 5715 2635
rect 5845 2605 5875 2635
rect 6005 2605 6035 2635
rect 6165 2605 6195 2635
rect 6325 2605 6355 2635
rect 6485 2605 6515 2635
rect 6645 2605 6675 2635
rect 6805 2605 6835 2635
rect 6965 2605 6995 2635
rect 7125 2605 7155 2635
rect 7285 2605 7315 2635
rect 7365 2605 7395 2635
rect 7525 2605 7555 2635
rect 7685 2605 7715 2635
rect 5525 2525 5555 2555
rect 5685 2525 5715 2555
rect 5845 2525 5875 2555
rect 6005 2525 6035 2555
rect 6165 2525 6195 2555
rect 6325 2525 6355 2555
rect 6485 2525 6515 2555
rect 6645 2525 6675 2555
rect 6805 2525 6835 2555
rect 6965 2525 6995 2555
rect 7125 2525 7155 2555
rect 7285 2525 7315 2555
rect 7365 2525 7395 2555
rect 7525 2525 7555 2555
rect 7685 2525 7715 2555
rect 5525 2445 5555 2475
rect 5685 2445 5715 2475
rect 5845 2445 5875 2475
rect 6005 2445 6035 2475
rect 6165 2445 6195 2475
rect 6325 2445 6355 2475
rect 6485 2445 6515 2475
rect 6645 2445 6675 2475
rect 6805 2445 6835 2475
rect 6965 2445 6995 2475
rect 7125 2445 7155 2475
rect 7285 2445 7315 2475
rect 7365 2445 7395 2475
rect 7525 2445 7555 2475
rect 7685 2445 7715 2475
rect 5525 2365 5555 2395
rect 5685 2365 5715 2395
rect 5845 2365 5875 2395
rect 6005 2365 6035 2395
rect 6165 2365 6195 2395
rect 6325 2365 6355 2395
rect 6485 2365 6515 2395
rect 6645 2365 6675 2395
rect 6805 2365 6835 2395
rect 6965 2365 6995 2395
rect 7125 2365 7155 2395
rect 7285 2365 7315 2395
rect 7365 2365 7395 2395
rect 7525 2365 7555 2395
rect 7685 2365 7715 2395
rect 6085 2285 6115 2315
rect 6165 2285 6195 2315
rect 6325 2285 6355 2315
rect 6485 2285 6515 2315
rect 6645 2285 6675 2315
rect 6805 2285 6835 2315
rect 6965 2285 6995 2315
rect 7125 2285 7155 2315
rect 7285 2285 7315 2315
rect 7365 2285 7395 2315
rect 7525 2285 7555 2315
rect 7685 2285 7715 2315
rect 5525 2205 5555 2235
rect 5685 2205 5715 2235
rect 5845 2205 5875 2235
rect 6005 2205 6035 2235
rect 6165 2205 6195 2235
rect 6325 2205 6355 2235
rect 6485 2205 6515 2235
rect 6645 2205 6675 2235
rect 6805 2205 6835 2235
rect 6965 2205 6995 2235
rect 7125 2205 7155 2235
rect 7285 2205 7315 2235
rect 7365 2205 7395 2235
rect 7525 2205 7555 2235
rect 7685 2205 7715 2235
rect 5525 2125 5555 2155
rect 5685 2125 5715 2155
rect 5845 2125 5875 2155
rect 6005 2125 6035 2155
rect 6165 2125 6195 2155
rect 6325 2125 6355 2155
rect 6485 2125 6515 2155
rect 6645 2125 6675 2155
rect 6805 2125 6835 2155
rect 6965 2125 6995 2155
rect 7125 2125 7155 2155
rect 7285 2125 7315 2155
rect 7365 2125 7395 2155
rect 7525 2125 7555 2155
rect 7685 2125 7715 2155
rect 5525 2045 5555 2075
rect 5685 2045 5715 2075
rect 5845 2045 5875 2075
rect 6005 2045 6035 2075
rect 6165 2045 6195 2075
rect 6325 2045 6355 2075
rect 6485 2045 6515 2075
rect 6645 2045 6675 2075
rect 6805 2045 6835 2075
rect 6965 2045 6995 2075
rect 7125 2045 7155 2075
rect 7285 2045 7315 2075
rect 7365 2045 7395 2075
rect 7525 2045 7555 2075
rect 7685 2045 7715 2075
rect 5525 1965 5555 1995
rect 5685 1965 5715 1995
rect 5845 1965 5875 1995
rect 6005 1965 6035 1995
rect 6165 1965 6195 1995
rect 6325 1965 6355 1995
rect 6485 1965 6515 1995
rect 6645 1965 6675 1995
rect 6805 1965 6835 1995
rect 6965 1965 6995 1995
rect 7125 1965 7155 1995
rect 7285 1965 7315 1995
rect 7365 1965 7395 1995
rect 7525 1965 7555 1995
rect 7685 1965 7715 1995
rect 5525 1885 5555 1915
rect 5685 1885 5715 1915
rect 5845 1885 5875 1915
rect 6005 1885 6035 1915
rect 6165 1885 6195 1915
rect 6325 1885 6355 1915
rect 6485 1885 6515 1915
rect 6645 1885 6675 1915
rect 6805 1885 6835 1915
rect 6965 1885 6995 1915
rect 7125 1885 7155 1915
rect 7285 1885 7315 1915
rect 7365 1885 7395 1915
rect 7525 1885 7555 1915
rect 7685 1885 7715 1915
rect 5525 1805 5555 1835
rect 5685 1805 5715 1835
rect 5845 1805 5875 1835
rect 6005 1805 6035 1835
rect 6165 1805 6195 1835
rect 6325 1805 6355 1835
rect 6485 1805 6515 1835
rect 6645 1805 6675 1835
rect 6805 1805 6835 1835
rect 6965 1805 6995 1835
rect 7125 1805 7155 1835
rect 7285 1805 7315 1835
rect 7365 1805 7395 1835
rect 7525 1805 7555 1835
rect 7685 1805 7715 1835
rect 5525 1725 5555 1755
rect 5685 1725 5715 1755
rect 5845 1725 5875 1755
rect 6005 1725 6035 1755
rect 6165 1725 6195 1755
rect 6325 1725 6355 1755
rect 6485 1725 6515 1755
rect 6645 1725 6675 1755
rect 6805 1725 6835 1755
rect 6965 1725 6995 1755
rect 7125 1725 7155 1755
rect 7285 1725 7315 1755
rect 7365 1725 7395 1755
rect 7525 1725 7555 1755
rect 7685 1725 7715 1755
rect 5525 1645 5555 1675
rect 5685 1645 5715 1675
rect 5845 1645 5875 1675
rect 6005 1645 6035 1675
rect 6165 1645 6195 1675
rect 6325 1645 6355 1675
rect 6485 1645 6515 1675
rect 6645 1645 6675 1675
rect 6805 1645 6835 1675
rect 6965 1645 6995 1675
rect 7125 1645 7155 1675
rect 7285 1645 7315 1675
rect 7365 1645 7395 1675
rect 7525 1645 7555 1675
rect 7685 1645 7715 1675
rect 5925 1565 5955 1595
rect 6005 1565 6035 1595
rect 6165 1565 6195 1595
rect 6325 1565 6355 1595
rect 6485 1565 6515 1595
rect 6645 1565 6675 1595
rect 6805 1565 6835 1595
rect 6965 1565 6995 1595
rect 7125 1565 7155 1595
rect 7285 1565 7315 1595
rect 7365 1565 7395 1595
rect 7525 1565 7555 1595
rect 7685 1565 7715 1595
rect 5525 1485 5555 1515
rect 5685 1485 5715 1515
rect 5845 1485 5875 1515
rect 6005 1485 6035 1515
rect 6165 1485 6195 1515
rect 6325 1485 6355 1515
rect 6485 1485 6515 1515
rect 6645 1485 6675 1515
rect 6805 1485 6835 1515
rect 6965 1485 6995 1515
rect 7125 1485 7155 1515
rect 7285 1485 7315 1515
rect 7365 1485 7395 1515
rect 7525 1485 7555 1515
rect 7685 1485 7715 1515
rect 5525 1405 5555 1435
rect 5685 1405 5715 1435
rect 5845 1405 5875 1435
rect 6005 1405 6035 1435
rect 6165 1405 6195 1435
rect 6325 1405 6355 1435
rect 6485 1405 6515 1435
rect 6645 1405 6675 1435
rect 6805 1405 6835 1435
rect 6965 1405 6995 1435
rect 7125 1405 7155 1435
rect 7285 1405 7315 1435
rect 7365 1405 7395 1435
rect 7525 1405 7555 1435
rect 7685 1405 7715 1435
rect 5525 1325 5555 1355
rect 5685 1325 5715 1355
rect 5845 1325 5875 1355
rect 6005 1325 6035 1355
rect 6165 1325 6195 1355
rect 6325 1325 6355 1355
rect 6485 1325 6515 1355
rect 6645 1325 6675 1355
rect 6805 1325 6835 1355
rect 6965 1325 6995 1355
rect 7125 1325 7155 1355
rect 7285 1325 7315 1355
rect 7365 1325 7395 1355
rect 7525 1325 7555 1355
rect 7685 1325 7715 1355
rect 5605 1245 5635 1275
rect 5685 1245 5715 1275
rect 5845 1245 5875 1275
rect 6005 1245 6035 1275
rect 6165 1245 6195 1275
rect 6325 1245 6355 1275
rect 6485 1245 6515 1275
rect 6645 1245 6675 1275
rect 6805 1245 6835 1275
rect 6965 1245 6995 1275
rect 7125 1245 7155 1275
rect 7285 1245 7315 1275
rect 7365 1245 7395 1275
rect 7525 1245 7555 1275
rect 7685 1245 7715 1275
rect 5525 1165 5555 1195
rect 5685 1165 5715 1195
rect 5845 1165 5875 1195
rect 6005 1165 6035 1195
rect 6165 1165 6195 1195
rect 6325 1165 6355 1195
rect 6485 1165 6515 1195
rect 6645 1165 6675 1195
rect 6805 1165 6835 1195
rect 6965 1165 6995 1195
rect 7125 1165 7155 1195
rect 7285 1165 7315 1195
rect 7365 1165 7395 1195
rect 7525 1165 7555 1195
rect 7685 1165 7715 1195
rect 5525 1085 5555 1115
rect 5685 1085 5715 1115
rect 5845 1085 5875 1115
rect 6005 1085 6035 1115
rect 6165 1085 6195 1115
rect 6325 1085 6355 1115
rect 6485 1085 6515 1115
rect 6645 1085 6675 1115
rect 6805 1085 6835 1115
rect 6965 1085 6995 1115
rect 7125 1085 7155 1115
rect 7285 1085 7315 1115
rect 7365 1085 7395 1115
rect 7525 1085 7555 1115
rect 7685 1085 7715 1115
rect 5525 1005 5555 1035
rect 5685 1005 5715 1035
rect 5845 1005 5875 1035
rect 6005 1005 6035 1035
rect 6165 1005 6195 1035
rect 6325 1005 6355 1035
rect 6485 1005 6515 1035
rect 6645 1005 6675 1035
rect 6805 1005 6835 1035
rect 6965 1005 6995 1035
rect 7125 1005 7155 1035
rect 7285 1005 7315 1035
rect 7365 1005 7395 1035
rect 7525 1005 7555 1035
rect 7685 1005 7715 1035
rect 5525 925 5555 955
rect 5685 925 5715 955
rect 5845 925 5875 955
rect 6005 925 6035 955
rect 6165 925 6195 955
rect 6325 925 6355 955
rect 6485 925 6515 955
rect 6645 925 6675 955
rect 6805 925 6835 955
rect 6965 925 6995 955
rect 7125 925 7155 955
rect 7285 925 7315 955
rect 7365 925 7395 955
rect 7525 925 7555 955
rect 7685 925 7715 955
rect 5525 845 5555 875
rect 5685 845 5715 875
rect 5845 845 5875 875
rect 6005 845 6035 875
rect 6165 845 6195 875
rect 6325 845 6355 875
rect 6485 845 6515 875
rect 6645 845 6675 875
rect 6805 845 6835 875
rect 6965 845 6995 875
rect 7125 845 7155 875
rect 7285 845 7315 875
rect 7365 845 7395 875
rect 7525 845 7555 875
rect 7685 845 7715 875
rect 5525 765 5555 795
rect 5685 765 5715 795
rect 5845 765 5875 795
rect 6005 765 6035 795
rect 6165 765 6195 795
rect 6325 765 6355 795
rect 6485 765 6515 795
rect 6645 765 6675 795
rect 6805 765 6835 795
rect 6965 765 6995 795
rect 7125 765 7155 795
rect 7285 765 7315 795
rect 7365 765 7395 795
rect 7525 765 7555 795
rect 7685 765 7715 795
rect 5765 685 5795 715
rect 5845 685 5875 715
rect 6005 685 6035 715
rect 6165 685 6195 715
rect 6325 685 6355 715
rect 6485 685 6515 715
rect 6645 685 6675 715
rect 6805 685 6835 715
rect 6965 685 6995 715
rect 7125 685 7155 715
rect 7285 685 7315 715
rect 7365 685 7395 715
rect 7525 685 7555 715
rect 7685 685 7715 715
rect 5525 565 5555 595
rect 5685 565 5715 595
rect 5845 565 5875 595
rect 6005 565 6035 595
rect 6165 565 6195 595
rect 6325 565 6355 595
rect 6485 565 6515 595
rect 6645 565 6675 595
rect 6805 565 6835 595
rect 6965 565 6995 595
rect 7125 565 7155 595
rect 7285 565 7315 595
rect 7365 565 7395 595
rect 7525 565 7555 595
rect 7685 565 7715 595
rect 5525 485 5555 515
rect 5685 485 5715 515
rect 5845 485 5875 515
rect 6005 485 6035 515
rect 6165 485 6195 515
rect 6325 485 6355 515
rect 6485 485 6515 515
rect 6645 485 6675 515
rect 6805 485 6835 515
rect 6965 485 6995 515
rect 7125 485 7155 515
rect 7285 485 7315 515
rect 7365 485 7395 515
rect 7525 485 7555 515
rect 7685 485 7715 515
rect 5605 405 5635 435
rect 5685 405 5715 435
rect 5845 405 5875 435
rect 6005 405 6035 435
rect 6165 405 6195 435
rect 6325 405 6355 435
rect 6485 405 6515 435
rect 6645 405 6675 435
rect 6805 405 6835 435
rect 6965 405 6995 435
rect 7125 405 7155 435
rect 7285 405 7315 435
rect 7365 405 7395 435
rect 7525 405 7555 435
rect 7685 405 7715 435
rect 5525 325 5555 355
rect 5685 325 5715 355
rect 5845 325 5875 355
rect 6005 325 6035 355
rect 6165 325 6195 355
rect 6325 325 6355 355
rect 6485 325 6515 355
rect 6645 325 6675 355
rect 6805 325 6835 355
rect 6965 325 6995 355
rect 7125 325 7155 355
rect 7285 325 7315 355
rect 7365 325 7395 355
rect 7525 325 7555 355
rect 7685 325 7715 355
rect 5525 245 5555 275
rect 5685 245 5715 275
rect 5845 245 5875 275
rect 6005 245 6035 275
rect 6165 245 6195 275
rect 6325 245 6355 275
rect 6485 245 6515 275
rect 6645 245 6675 275
rect 6805 245 6835 275
rect 6965 245 6995 275
rect 7125 245 7155 275
rect 7285 245 7315 275
rect 7365 245 7395 275
rect 7525 245 7555 275
rect 7685 245 7715 275
rect 5525 165 5555 195
rect 5685 165 5715 195
rect 5845 165 5875 195
rect 6005 165 6035 195
rect 6165 165 6195 195
rect 6325 165 6355 195
rect 6485 165 6515 195
rect 6645 165 6675 195
rect 6805 165 6835 195
rect 6965 165 6995 195
rect 7125 165 7155 195
rect 7285 165 7315 195
rect 7365 165 7395 195
rect 7525 165 7555 195
rect 7685 165 7715 195
rect 5525 85 5555 115
rect 5685 85 5715 115
rect 5845 85 5875 115
rect 6005 85 6035 115
rect 6165 85 6195 115
rect 6325 85 6355 115
rect 6485 85 6515 115
rect 6645 85 6675 115
rect 6805 85 6835 115
rect 6965 85 6995 115
rect 7125 85 7155 115
rect 7285 85 7315 115
rect 7365 85 7395 115
rect 7525 85 7555 115
rect 7685 85 7715 115
rect 5525 5 5555 35
rect 5685 5 5715 35
rect 5845 5 5875 35
rect 6005 5 6035 35
rect 6165 5 6195 35
rect 6325 5 6355 35
rect 6485 5 6515 35
rect 6645 5 6675 35
rect 6805 5 6835 35
rect 6965 5 6995 35
rect 7125 5 7155 35
rect 7285 5 7315 35
rect 7365 5 7395 35
rect 7525 5 7555 35
rect 7685 5 7715 35
<< metal3 >>
rect 7360 19716 7400 19720
rect 7360 19684 7364 19716
rect 7396 19684 7400 19716
rect 560 19636 1640 19640
rect 560 19604 564 19636
rect 1636 19604 1640 19636
rect 560 18520 1640 19604
rect 1680 19636 2760 19640
rect 1680 19604 1684 19636
rect 2756 19604 2760 19636
rect 1680 18520 2760 19604
rect 2800 19636 3880 19640
rect 2800 19604 2804 19636
rect 3876 19604 3880 19636
rect 2800 18520 3880 19604
rect 3920 19636 5000 19640
rect 3920 19604 3924 19636
rect 4996 19604 5000 19636
rect 3920 18520 5000 19604
rect 5040 19636 6120 19640
rect 5040 19604 5044 19636
rect 6116 19604 6120 19636
rect 5040 18520 6120 19604
rect 6160 19636 7240 19640
rect 6160 19604 6164 19636
rect 7236 19604 7240 19636
rect 6160 18520 7240 19604
rect 560 18480 7240 18520
rect 560 18400 7240 18440
rect 560 17316 1640 18400
rect 560 17284 564 17316
rect 1636 17284 1640 17316
rect 560 17280 1640 17284
rect 1680 17316 2760 18400
rect 1680 17284 1684 17316
rect 2756 17284 2760 17316
rect 1680 17280 2760 17284
rect 2800 17316 3880 18400
rect 2800 17284 2804 17316
rect 3876 17284 3880 17316
rect 2800 17280 3880 17284
rect 3920 17316 5000 18400
rect 3920 17284 3924 17316
rect 4996 17284 5000 17316
rect 3920 17280 5000 17284
rect 5040 17316 6120 18400
rect 5040 17284 5044 17316
rect 6116 17284 6120 17316
rect 5040 17280 6120 17284
rect 6160 17316 7240 18400
rect 6160 17284 6164 17316
rect 7236 17284 7240 17316
rect 6160 17280 7240 17284
rect 7280 17156 7320 19680
rect 7280 17124 7284 17156
rect 7316 17124 7320 17156
rect 5520 16836 5560 16840
rect 5520 16644 5524 16836
rect 5556 16644 5560 16836
rect 5520 16596 5560 16644
rect 5680 16836 5720 16840
rect 5680 16644 5684 16836
rect 5716 16644 5720 16836
rect 5520 16564 5524 16596
rect 5556 16564 5560 16596
rect 5520 16516 5560 16564
rect 5520 16484 5524 16516
rect 5556 16484 5560 16516
rect 5520 16436 5560 16484
rect 5520 16404 5524 16436
rect 5556 16404 5560 16436
rect 5520 16356 5560 16404
rect 5520 16324 5524 16356
rect 5556 16324 5560 16356
rect 5520 16276 5560 16324
rect 5520 16244 5524 16276
rect 5556 16244 5560 16276
rect 5520 16196 5560 16244
rect 5520 16164 5524 16196
rect 5556 16164 5560 16196
rect 5520 16116 5560 16164
rect 5520 16084 5524 16116
rect 5556 16084 5560 16116
rect 5520 16036 5560 16084
rect 5520 16004 5524 16036
rect 5556 16004 5560 16036
rect 5520 15956 5560 16004
rect 5520 15924 5524 15956
rect 5556 15924 5560 15956
rect 5520 15436 5560 15924
rect 5520 15404 5524 15436
rect 5556 15404 5560 15436
rect 5520 15356 5560 15404
rect 5520 15324 5524 15356
rect 5556 15324 5560 15356
rect 5520 15276 5560 15324
rect 5520 15244 5524 15276
rect 5556 15244 5560 15276
rect 5520 15196 5560 15244
rect 5520 15164 5524 15196
rect 5556 15164 5560 15196
rect 5520 15116 5560 15164
rect 5520 15084 5524 15116
rect 5556 15084 5560 15116
rect 5520 14956 5560 15084
rect 5520 14924 5524 14956
rect 5556 14924 5560 14956
rect 5520 14876 5560 14924
rect 5520 14844 5524 14876
rect 5556 14844 5560 14876
rect 5520 14796 5560 14844
rect 5520 14764 5524 14796
rect 5556 14764 5560 14796
rect 5520 14716 5560 14764
rect 5520 14684 5524 14716
rect 5556 14684 5560 14716
rect 5520 14556 5560 14684
rect 5520 14524 5524 14556
rect 5556 14524 5560 14556
rect 5520 14476 5560 14524
rect 5520 14444 5524 14476
rect 5556 14444 5560 14476
rect 5520 13996 5560 14444
rect 5520 13964 5524 13996
rect 5556 13964 5560 13996
rect 5520 13796 5560 13964
rect 5520 13764 5524 13796
rect 5556 13764 5560 13796
rect 5520 13716 5560 13764
rect 5520 13684 5524 13716
rect 5556 13684 5560 13716
rect 5520 13636 5560 13684
rect 5520 13604 5524 13636
rect 5556 13604 5560 13636
rect 5520 13476 5560 13604
rect 5520 13444 5524 13476
rect 5556 13444 5560 13476
rect 5520 13396 5560 13444
rect 5520 13364 5524 13396
rect 5556 13364 5560 13396
rect 5520 13316 5560 13364
rect 5520 13284 5524 13316
rect 5556 13284 5560 13316
rect 5520 13236 5560 13284
rect 5520 13204 5524 13236
rect 5556 13204 5560 13236
rect 5520 13076 5560 13204
rect 5520 13044 5524 13076
rect 5556 13044 5560 13076
rect 5520 12996 5560 13044
rect 5520 12964 5524 12996
rect 5556 12964 5560 12996
rect 5520 12516 5560 12964
rect 5520 12484 5524 12516
rect 5556 12484 5560 12516
rect 5520 12316 5560 12484
rect 5520 12284 5524 12316
rect 5556 12284 5560 12316
rect 5520 12236 5560 12284
rect 5520 12204 5524 12236
rect 5556 12204 5560 12236
rect 5520 12156 5560 12204
rect 5520 12124 5524 12156
rect 5556 12124 5560 12156
rect 5520 12076 5560 12124
rect 5520 12044 5524 12076
rect 5556 12044 5560 12076
rect 5520 11996 5560 12044
rect 5520 11964 5524 11996
rect 5556 11964 5560 11996
rect 5520 11916 5560 11964
rect 5520 11884 5524 11916
rect 5556 11884 5560 11916
rect 5520 11836 5560 11884
rect 5520 11804 5524 11836
rect 5556 11804 5560 11836
rect 5520 11756 5560 11804
rect 5520 11724 5524 11756
rect 5556 11724 5560 11756
rect 5520 11676 5560 11724
rect 5520 11644 5524 11676
rect 5556 11644 5560 11676
rect 5520 11596 5560 11644
rect 5520 11564 5524 11596
rect 5556 11564 5560 11596
rect 5520 11516 5560 11564
rect 5520 11484 5524 11516
rect 5556 11484 5560 11516
rect 5520 11436 5560 11484
rect 5520 11404 5524 11436
rect 5556 11404 5560 11436
rect 5520 11356 5560 11404
rect 5520 11324 5524 11356
rect 5556 11324 5560 11356
rect 5520 11196 5560 11324
rect 5520 11164 5524 11196
rect 5556 11164 5560 11196
rect 5520 11116 5560 11164
rect 5520 11084 5524 11116
rect 5556 11084 5560 11116
rect 5520 11036 5560 11084
rect 5520 11004 5524 11036
rect 5556 11004 5560 11036
rect 5520 10876 5560 11004
rect 5520 10844 5524 10876
rect 5556 10844 5560 10876
rect 5520 10716 5560 10844
rect 5520 10684 5524 10716
rect 5556 10684 5560 10716
rect 5520 10636 5560 10684
rect 5520 10604 5524 10636
rect 5556 10604 5560 10636
rect 5520 10476 5560 10604
rect 5520 10444 5524 10476
rect 5556 10444 5560 10476
rect 5520 10316 5560 10444
rect 5520 10284 5524 10316
rect 5556 10284 5560 10316
rect 5520 10236 5560 10284
rect 5520 10204 5524 10236
rect 5556 10204 5560 10236
rect 5520 10156 5560 10204
rect 5520 10124 5524 10156
rect 5556 10124 5560 10156
rect 5520 10076 5560 10124
rect 5520 10044 5524 10076
rect 5556 10044 5560 10076
rect 5520 9996 5560 10044
rect 5520 9964 5524 9996
rect 5556 9964 5560 9996
rect 5520 9916 5560 9964
rect 5520 9884 5524 9916
rect 5556 9884 5560 9916
rect 5520 9836 5560 9884
rect 5520 9804 5524 9836
rect 5556 9804 5560 9836
rect 5520 9756 5560 9804
rect 5520 9724 5524 9756
rect 5556 9724 5560 9756
rect 5520 9676 5560 9724
rect 5520 9644 5524 9676
rect 5556 9644 5560 9676
rect 5520 9596 5560 9644
rect 5520 9564 5524 9596
rect 5556 9564 5560 9596
rect 5520 9516 5560 9564
rect 5520 9484 5524 9516
rect 5556 9484 5560 9516
rect 5520 9436 5560 9484
rect 5520 9404 5524 9436
rect 5556 9404 5560 9436
rect 5520 9356 5560 9404
rect 5520 9324 5524 9356
rect 5556 9324 5560 9356
rect 5520 9276 5560 9324
rect 5520 9244 5524 9276
rect 5556 9244 5560 9276
rect 5520 9116 5560 9244
rect 5520 9084 5524 9116
rect 5556 9084 5560 9116
rect 5520 9036 5560 9084
rect 5520 9004 5524 9036
rect 5556 9004 5560 9036
rect 5520 8956 5560 9004
rect 5520 8924 5524 8956
rect 5556 8924 5560 8956
rect 5520 8636 5560 8924
rect 5520 8604 5524 8636
rect 5556 8604 5560 8636
rect 5520 8556 5560 8604
rect 5520 8524 5524 8556
rect 5556 8524 5560 8556
rect 5520 8396 5560 8524
rect 5520 8364 5524 8396
rect 5556 8364 5560 8396
rect 5520 8236 5560 8364
rect 5520 8204 5524 8236
rect 5556 8204 5560 8236
rect 5520 8156 5560 8204
rect 5520 8124 5524 8156
rect 5556 8124 5560 8156
rect 5520 8076 5560 8124
rect 5520 8044 5524 8076
rect 5556 8044 5560 8076
rect 5520 7996 5560 8044
rect 5520 7964 5524 7996
rect 5556 7964 5560 7996
rect 5520 7916 5560 7964
rect 5520 7884 5524 7916
rect 5556 7884 5560 7916
rect 5520 7836 5560 7884
rect 5520 7804 5524 7836
rect 5556 7804 5560 7836
rect 5520 7756 5560 7804
rect 5520 7724 5524 7756
rect 5556 7724 5560 7756
rect 5520 7676 5560 7724
rect 5520 7644 5524 7676
rect 5556 7644 5560 7676
rect 5520 7596 5560 7644
rect 5520 7564 5524 7596
rect 5556 7564 5560 7596
rect 5520 7516 5560 7564
rect 5520 7484 5524 7516
rect 5556 7484 5560 7516
rect 5520 7436 5560 7484
rect 5520 7404 5524 7436
rect 5556 7404 5560 7436
rect 5520 7356 5560 7404
rect 5520 7324 5524 7356
rect 5556 7324 5560 7356
rect 5520 7276 5560 7324
rect 5520 7244 5524 7276
rect 5556 7244 5560 7276
rect 5520 7196 5560 7244
rect 5520 7164 5524 7196
rect 5556 7164 5560 7196
rect 5520 7036 5560 7164
rect 5520 7004 5524 7036
rect 5556 7004 5560 7036
rect 5520 6956 5560 7004
rect 5520 6924 5524 6956
rect 5556 6924 5560 6956
rect 5520 6796 5560 6924
rect 5520 6764 5524 6796
rect 5556 6764 5560 6796
rect 5520 6716 5560 6764
rect 5520 6684 5524 6716
rect 5556 6684 5560 6716
rect 5520 6636 5560 6684
rect 5520 6604 5524 6636
rect 5556 6604 5560 6636
rect 5520 6556 5560 6604
rect 5520 6524 5524 6556
rect 5556 6524 5560 6556
rect 5520 6476 5560 6524
rect 5520 6444 5524 6476
rect 5556 6444 5560 6476
rect 5520 6316 5560 6444
rect 5520 6284 5524 6316
rect 5556 6284 5560 6316
rect 5520 6236 5560 6284
rect 5520 6204 5524 6236
rect 5556 6204 5560 6236
rect 5520 6156 5560 6204
rect 5520 6124 5524 6156
rect 5556 6124 5560 6156
rect 5520 5996 5560 6124
rect 5520 5964 5524 5996
rect 5556 5964 5560 5996
rect 5520 5836 5560 5964
rect 5520 5804 5524 5836
rect 5556 5804 5560 5836
rect 5520 5756 5560 5804
rect 5520 5724 5524 5756
rect 5556 5724 5560 5756
rect 5520 5676 5560 5724
rect 5520 5644 5524 5676
rect 5556 5644 5560 5676
rect 5520 5596 5560 5644
rect 5520 5564 5524 5596
rect 5556 5564 5560 5596
rect 5520 5516 5560 5564
rect 5520 5484 5524 5516
rect 5556 5484 5560 5516
rect 5520 5436 5560 5484
rect 5520 5404 5524 5436
rect 5556 5404 5560 5436
rect 5520 5356 5560 5404
rect 5520 5324 5524 5356
rect 5556 5324 5560 5356
rect 5520 5276 5560 5324
rect 5520 5244 5524 5276
rect 5556 5244 5560 5276
rect 5520 5196 5560 5244
rect 5520 5164 5524 5196
rect 5556 5164 5560 5196
rect 5520 5116 5560 5164
rect 5520 5084 5524 5116
rect 5556 5084 5560 5116
rect 5520 5036 5560 5084
rect 5520 5004 5524 5036
rect 5556 5004 5560 5036
rect 5520 4956 5560 5004
rect 5520 4924 5524 4956
rect 5556 4924 5560 4956
rect 5520 4876 5560 4924
rect 5520 4844 5524 4876
rect 5556 4844 5560 4876
rect 5520 4796 5560 4844
rect 5520 4764 5524 4796
rect 5556 4764 5560 4796
rect 5520 4636 5560 4764
rect 5520 4604 5524 4636
rect 5556 4604 5560 4636
rect 5520 4556 5560 4604
rect 5520 4524 5524 4556
rect 5556 4524 5560 4556
rect 5520 4396 5560 4524
rect 5520 4364 5524 4396
rect 5556 4364 5560 4396
rect 5520 4316 5560 4364
rect 5520 4284 5524 4316
rect 5556 4284 5560 4316
rect 5520 4236 5560 4284
rect 5520 4204 5524 4236
rect 5556 4204 5560 4236
rect 5520 4156 5560 4204
rect 5520 4124 5524 4156
rect 5556 4124 5560 4156
rect 5520 4076 5560 4124
rect 5520 4044 5524 4076
rect 5556 4044 5560 4076
rect 5520 3916 5560 4044
rect 5520 3884 5524 3916
rect 5556 3884 5560 3916
rect 5520 3836 5560 3884
rect 5520 3804 5524 3836
rect 5556 3804 5560 3836
rect 5520 3756 5560 3804
rect 5520 3724 5524 3756
rect 5556 3724 5560 3756
rect 5520 3596 5560 3724
rect 5520 3564 5524 3596
rect 5556 3564 5560 3596
rect 5520 3436 5560 3564
rect 5520 3404 5524 3436
rect 5556 3404 5560 3436
rect 5520 3356 5560 3404
rect 5520 3324 5524 3356
rect 5556 3324 5560 3356
rect 5520 3276 5560 3324
rect 5520 3244 5524 3276
rect 5556 3244 5560 3276
rect 5520 3196 5560 3244
rect 5520 3164 5524 3196
rect 5556 3164 5560 3196
rect 5520 3116 5560 3164
rect 5520 3084 5524 3116
rect 5556 3084 5560 3116
rect 5520 3036 5560 3084
rect 5520 3004 5524 3036
rect 5556 3004 5560 3036
rect 5520 2956 5560 3004
rect 5520 2924 5524 2956
rect 5556 2924 5560 2956
rect 5520 2876 5560 2924
rect 5520 2844 5524 2876
rect 5556 2844 5560 2876
rect 5520 2796 5560 2844
rect 5520 2764 5524 2796
rect 5556 2764 5560 2796
rect 5520 2716 5560 2764
rect 5520 2684 5524 2716
rect 5556 2684 5560 2716
rect 5520 2636 5560 2684
rect 5520 2604 5524 2636
rect 5556 2604 5560 2636
rect 5520 2556 5560 2604
rect 5520 2524 5524 2556
rect 5556 2524 5560 2556
rect 5520 2476 5560 2524
rect 5520 2444 5524 2476
rect 5556 2444 5560 2476
rect 5520 2396 5560 2444
rect 5520 2364 5524 2396
rect 5556 2364 5560 2396
rect 5520 2236 5560 2364
rect 5520 2204 5524 2236
rect 5556 2204 5560 2236
rect 5520 2156 5560 2204
rect 5520 2124 5524 2156
rect 5556 2124 5560 2156
rect 5520 2076 5560 2124
rect 5520 2044 5524 2076
rect 5556 2044 5560 2076
rect 5520 1996 5560 2044
rect 5520 1964 5524 1996
rect 5556 1964 5560 1996
rect 5520 1916 5560 1964
rect 5520 1884 5524 1916
rect 5556 1884 5560 1916
rect 5520 1836 5560 1884
rect 5520 1804 5524 1836
rect 5556 1804 5560 1836
rect 5520 1756 5560 1804
rect 5520 1724 5524 1756
rect 5556 1724 5560 1756
rect 5520 1676 5560 1724
rect 5520 1644 5524 1676
rect 5556 1644 5560 1676
rect 5520 1516 5560 1644
rect 5520 1484 5524 1516
rect 5556 1484 5560 1516
rect 5520 1436 5560 1484
rect 5520 1404 5524 1436
rect 5556 1404 5560 1436
rect 5520 1356 5560 1404
rect 5520 1324 5524 1356
rect 5556 1324 5560 1356
rect 5520 1196 5560 1324
rect 5520 1164 5524 1196
rect 5556 1164 5560 1196
rect 5520 1116 5560 1164
rect 5520 1084 5524 1116
rect 5556 1084 5560 1116
rect 5520 1036 5560 1084
rect 5520 1004 5524 1036
rect 5556 1004 5560 1036
rect 5520 956 5560 1004
rect 5520 924 5524 956
rect 5556 924 5560 956
rect 5520 876 5560 924
rect 5520 844 5524 876
rect 5556 844 5560 876
rect 5520 796 5560 844
rect 5520 764 5524 796
rect 5556 764 5560 796
rect 5520 596 5560 764
rect 5520 564 5524 596
rect 5556 564 5560 596
rect 5520 516 5560 564
rect 5520 484 5524 516
rect 5556 484 5560 516
rect 5520 356 5560 484
rect 5520 324 5524 356
rect 5556 324 5560 356
rect 5520 276 5560 324
rect 5520 244 5524 276
rect 5556 244 5560 276
rect 5520 196 5560 244
rect 5520 164 5524 196
rect 5556 164 5560 196
rect 5520 116 5560 164
rect 5520 84 5524 116
rect 5556 84 5560 116
rect 5520 36 5560 84
rect 5520 4 5524 36
rect 5556 4 5560 36
rect 5520 -40 5560 4
rect 5600 1275 5640 16640
rect 5600 1245 5605 1275
rect 5635 1245 5640 1275
rect 5600 435 5640 1245
rect 5600 405 5605 435
rect 5635 405 5640 435
rect 5600 -40 5640 405
rect 5680 16596 5720 16644
rect 5840 16836 5880 16840
rect 5840 16644 5844 16836
rect 5876 16644 5880 16836
rect 5680 16564 5684 16596
rect 5716 16564 5720 16596
rect 5680 16516 5720 16564
rect 5680 16484 5684 16516
rect 5716 16484 5720 16516
rect 5680 16436 5720 16484
rect 5680 16404 5684 16436
rect 5716 16404 5720 16436
rect 5680 16356 5720 16404
rect 5680 16324 5684 16356
rect 5716 16324 5720 16356
rect 5680 16276 5720 16324
rect 5680 16244 5684 16276
rect 5716 16244 5720 16276
rect 5680 16196 5720 16244
rect 5680 16164 5684 16196
rect 5716 16164 5720 16196
rect 5680 16116 5720 16164
rect 5680 16084 5684 16116
rect 5716 16084 5720 16116
rect 5680 16036 5720 16084
rect 5680 16004 5684 16036
rect 5716 16004 5720 16036
rect 5680 15956 5720 16004
rect 5680 15924 5684 15956
rect 5716 15924 5720 15956
rect 5680 15436 5720 15924
rect 5680 15404 5684 15436
rect 5716 15404 5720 15436
rect 5680 15356 5720 15404
rect 5680 15324 5684 15356
rect 5716 15324 5720 15356
rect 5680 15276 5720 15324
rect 5680 15244 5684 15276
rect 5716 15244 5720 15276
rect 5680 15196 5720 15244
rect 5680 15164 5684 15196
rect 5716 15164 5720 15196
rect 5680 15116 5720 15164
rect 5680 15084 5684 15116
rect 5716 15084 5720 15116
rect 5680 14956 5720 15084
rect 5680 14924 5684 14956
rect 5716 14924 5720 14956
rect 5680 14876 5720 14924
rect 5680 14844 5684 14876
rect 5716 14844 5720 14876
rect 5680 14796 5720 14844
rect 5680 14764 5684 14796
rect 5716 14764 5720 14796
rect 5680 14716 5720 14764
rect 5680 14684 5684 14716
rect 5716 14684 5720 14716
rect 5680 14556 5720 14684
rect 5680 14524 5684 14556
rect 5716 14524 5720 14556
rect 5680 14476 5720 14524
rect 5680 14444 5684 14476
rect 5716 14444 5720 14476
rect 5680 13996 5720 14444
rect 5680 13964 5684 13996
rect 5716 13964 5720 13996
rect 5680 13796 5720 13964
rect 5680 13764 5684 13796
rect 5716 13764 5720 13796
rect 5680 13716 5720 13764
rect 5680 13684 5684 13716
rect 5716 13684 5720 13716
rect 5680 13636 5720 13684
rect 5680 13604 5684 13636
rect 5716 13604 5720 13636
rect 5680 13476 5720 13604
rect 5680 13444 5684 13476
rect 5716 13444 5720 13476
rect 5680 13396 5720 13444
rect 5680 13364 5684 13396
rect 5716 13364 5720 13396
rect 5680 13316 5720 13364
rect 5680 13284 5684 13316
rect 5716 13284 5720 13316
rect 5680 13236 5720 13284
rect 5680 13204 5684 13236
rect 5716 13204 5720 13236
rect 5680 13076 5720 13204
rect 5680 13044 5684 13076
rect 5716 13044 5720 13076
rect 5680 12996 5720 13044
rect 5680 12964 5684 12996
rect 5716 12964 5720 12996
rect 5680 12516 5720 12964
rect 5680 12484 5684 12516
rect 5716 12484 5720 12516
rect 5680 12316 5720 12484
rect 5680 12284 5684 12316
rect 5716 12284 5720 12316
rect 5680 12236 5720 12284
rect 5680 12204 5684 12236
rect 5716 12204 5720 12236
rect 5680 12156 5720 12204
rect 5680 12124 5684 12156
rect 5716 12124 5720 12156
rect 5680 12076 5720 12124
rect 5680 12044 5684 12076
rect 5716 12044 5720 12076
rect 5680 11996 5720 12044
rect 5680 11964 5684 11996
rect 5716 11964 5720 11996
rect 5680 11916 5720 11964
rect 5680 11884 5684 11916
rect 5716 11884 5720 11916
rect 5680 11836 5720 11884
rect 5680 11804 5684 11836
rect 5716 11804 5720 11836
rect 5680 11756 5720 11804
rect 5680 11724 5684 11756
rect 5716 11724 5720 11756
rect 5680 11676 5720 11724
rect 5680 11644 5684 11676
rect 5716 11644 5720 11676
rect 5680 11596 5720 11644
rect 5680 11564 5684 11596
rect 5716 11564 5720 11596
rect 5680 11516 5720 11564
rect 5680 11484 5684 11516
rect 5716 11484 5720 11516
rect 5680 11436 5720 11484
rect 5680 11404 5684 11436
rect 5716 11404 5720 11436
rect 5680 11356 5720 11404
rect 5680 11324 5684 11356
rect 5716 11324 5720 11356
rect 5680 11196 5720 11324
rect 5680 11164 5684 11196
rect 5716 11164 5720 11196
rect 5680 11116 5720 11164
rect 5680 11084 5684 11116
rect 5716 11084 5720 11116
rect 5680 11036 5720 11084
rect 5680 11004 5684 11036
rect 5716 11004 5720 11036
rect 5680 10876 5720 11004
rect 5680 10844 5684 10876
rect 5716 10844 5720 10876
rect 5680 10716 5720 10844
rect 5680 10684 5684 10716
rect 5716 10684 5720 10716
rect 5680 10636 5720 10684
rect 5680 10604 5684 10636
rect 5716 10604 5720 10636
rect 5680 10476 5720 10604
rect 5680 10444 5684 10476
rect 5716 10444 5720 10476
rect 5680 10316 5720 10444
rect 5680 10284 5684 10316
rect 5716 10284 5720 10316
rect 5680 10236 5720 10284
rect 5680 10204 5684 10236
rect 5716 10204 5720 10236
rect 5680 10156 5720 10204
rect 5680 10124 5684 10156
rect 5716 10124 5720 10156
rect 5680 10076 5720 10124
rect 5680 10044 5684 10076
rect 5716 10044 5720 10076
rect 5680 9996 5720 10044
rect 5680 9964 5684 9996
rect 5716 9964 5720 9996
rect 5680 9916 5720 9964
rect 5680 9884 5684 9916
rect 5716 9884 5720 9916
rect 5680 9836 5720 9884
rect 5680 9804 5684 9836
rect 5716 9804 5720 9836
rect 5680 9756 5720 9804
rect 5680 9724 5684 9756
rect 5716 9724 5720 9756
rect 5680 9676 5720 9724
rect 5680 9644 5684 9676
rect 5716 9644 5720 9676
rect 5680 9596 5720 9644
rect 5680 9564 5684 9596
rect 5716 9564 5720 9596
rect 5680 9516 5720 9564
rect 5680 9484 5684 9516
rect 5716 9484 5720 9516
rect 5680 9436 5720 9484
rect 5680 9404 5684 9436
rect 5716 9404 5720 9436
rect 5680 9356 5720 9404
rect 5680 9324 5684 9356
rect 5716 9324 5720 9356
rect 5680 9276 5720 9324
rect 5680 9244 5684 9276
rect 5716 9244 5720 9276
rect 5680 9116 5720 9244
rect 5680 9084 5684 9116
rect 5716 9084 5720 9116
rect 5680 9036 5720 9084
rect 5680 9004 5684 9036
rect 5716 9004 5720 9036
rect 5680 8956 5720 9004
rect 5680 8924 5684 8956
rect 5716 8924 5720 8956
rect 5680 8636 5720 8924
rect 5680 8604 5684 8636
rect 5716 8604 5720 8636
rect 5680 8556 5720 8604
rect 5680 8524 5684 8556
rect 5716 8524 5720 8556
rect 5680 8396 5720 8524
rect 5680 8364 5684 8396
rect 5716 8364 5720 8396
rect 5680 8236 5720 8364
rect 5680 8204 5684 8236
rect 5716 8204 5720 8236
rect 5680 8156 5720 8204
rect 5680 8124 5684 8156
rect 5716 8124 5720 8156
rect 5680 8076 5720 8124
rect 5680 8044 5684 8076
rect 5716 8044 5720 8076
rect 5680 7996 5720 8044
rect 5680 7964 5684 7996
rect 5716 7964 5720 7996
rect 5680 7916 5720 7964
rect 5680 7884 5684 7916
rect 5716 7884 5720 7916
rect 5680 7836 5720 7884
rect 5680 7804 5684 7836
rect 5716 7804 5720 7836
rect 5680 7756 5720 7804
rect 5680 7724 5684 7756
rect 5716 7724 5720 7756
rect 5680 7676 5720 7724
rect 5680 7644 5684 7676
rect 5716 7644 5720 7676
rect 5680 7596 5720 7644
rect 5680 7564 5684 7596
rect 5716 7564 5720 7596
rect 5680 7516 5720 7564
rect 5680 7484 5684 7516
rect 5716 7484 5720 7516
rect 5680 7436 5720 7484
rect 5680 7404 5684 7436
rect 5716 7404 5720 7436
rect 5680 7356 5720 7404
rect 5680 7324 5684 7356
rect 5716 7324 5720 7356
rect 5680 7276 5720 7324
rect 5680 7244 5684 7276
rect 5716 7244 5720 7276
rect 5680 7196 5720 7244
rect 5680 7164 5684 7196
rect 5716 7164 5720 7196
rect 5680 7036 5720 7164
rect 5680 7004 5684 7036
rect 5716 7004 5720 7036
rect 5680 6956 5720 7004
rect 5680 6924 5684 6956
rect 5716 6924 5720 6956
rect 5680 6796 5720 6924
rect 5680 6764 5684 6796
rect 5716 6764 5720 6796
rect 5680 6716 5720 6764
rect 5680 6684 5684 6716
rect 5716 6684 5720 6716
rect 5680 6636 5720 6684
rect 5680 6604 5684 6636
rect 5716 6604 5720 6636
rect 5680 6556 5720 6604
rect 5680 6524 5684 6556
rect 5716 6524 5720 6556
rect 5680 6476 5720 6524
rect 5680 6444 5684 6476
rect 5716 6444 5720 6476
rect 5680 6316 5720 6444
rect 5680 6284 5684 6316
rect 5716 6284 5720 6316
rect 5680 6236 5720 6284
rect 5680 6204 5684 6236
rect 5716 6204 5720 6236
rect 5680 6156 5720 6204
rect 5680 6124 5684 6156
rect 5716 6124 5720 6156
rect 5680 5996 5720 6124
rect 5680 5964 5684 5996
rect 5716 5964 5720 5996
rect 5680 5836 5720 5964
rect 5680 5804 5684 5836
rect 5716 5804 5720 5836
rect 5680 5756 5720 5804
rect 5680 5724 5684 5756
rect 5716 5724 5720 5756
rect 5680 5676 5720 5724
rect 5680 5644 5684 5676
rect 5716 5644 5720 5676
rect 5680 5596 5720 5644
rect 5680 5564 5684 5596
rect 5716 5564 5720 5596
rect 5680 5516 5720 5564
rect 5680 5484 5684 5516
rect 5716 5484 5720 5516
rect 5680 5436 5720 5484
rect 5680 5404 5684 5436
rect 5716 5404 5720 5436
rect 5680 5356 5720 5404
rect 5680 5324 5684 5356
rect 5716 5324 5720 5356
rect 5680 5276 5720 5324
rect 5680 5244 5684 5276
rect 5716 5244 5720 5276
rect 5680 5196 5720 5244
rect 5680 5164 5684 5196
rect 5716 5164 5720 5196
rect 5680 5116 5720 5164
rect 5680 5084 5684 5116
rect 5716 5084 5720 5116
rect 5680 5036 5720 5084
rect 5680 5004 5684 5036
rect 5716 5004 5720 5036
rect 5680 4956 5720 5004
rect 5680 4924 5684 4956
rect 5716 4924 5720 4956
rect 5680 4876 5720 4924
rect 5680 4844 5684 4876
rect 5716 4844 5720 4876
rect 5680 4796 5720 4844
rect 5680 4764 5684 4796
rect 5716 4764 5720 4796
rect 5680 4636 5720 4764
rect 5680 4604 5684 4636
rect 5716 4604 5720 4636
rect 5680 4556 5720 4604
rect 5680 4524 5684 4556
rect 5716 4524 5720 4556
rect 5680 4396 5720 4524
rect 5680 4364 5684 4396
rect 5716 4364 5720 4396
rect 5680 4316 5720 4364
rect 5680 4284 5684 4316
rect 5716 4284 5720 4316
rect 5680 4236 5720 4284
rect 5680 4204 5684 4236
rect 5716 4204 5720 4236
rect 5680 4156 5720 4204
rect 5680 4124 5684 4156
rect 5716 4124 5720 4156
rect 5680 4076 5720 4124
rect 5680 4044 5684 4076
rect 5716 4044 5720 4076
rect 5680 3916 5720 4044
rect 5680 3884 5684 3916
rect 5716 3884 5720 3916
rect 5680 3836 5720 3884
rect 5680 3804 5684 3836
rect 5716 3804 5720 3836
rect 5680 3756 5720 3804
rect 5680 3724 5684 3756
rect 5716 3724 5720 3756
rect 5680 3596 5720 3724
rect 5680 3564 5684 3596
rect 5716 3564 5720 3596
rect 5680 3436 5720 3564
rect 5680 3404 5684 3436
rect 5716 3404 5720 3436
rect 5680 3356 5720 3404
rect 5680 3324 5684 3356
rect 5716 3324 5720 3356
rect 5680 3276 5720 3324
rect 5680 3244 5684 3276
rect 5716 3244 5720 3276
rect 5680 3196 5720 3244
rect 5680 3164 5684 3196
rect 5716 3164 5720 3196
rect 5680 3116 5720 3164
rect 5680 3084 5684 3116
rect 5716 3084 5720 3116
rect 5680 3036 5720 3084
rect 5680 3004 5684 3036
rect 5716 3004 5720 3036
rect 5680 2956 5720 3004
rect 5680 2924 5684 2956
rect 5716 2924 5720 2956
rect 5680 2876 5720 2924
rect 5680 2844 5684 2876
rect 5716 2844 5720 2876
rect 5680 2796 5720 2844
rect 5680 2764 5684 2796
rect 5716 2764 5720 2796
rect 5680 2716 5720 2764
rect 5680 2684 5684 2716
rect 5716 2684 5720 2716
rect 5680 2636 5720 2684
rect 5680 2604 5684 2636
rect 5716 2604 5720 2636
rect 5680 2556 5720 2604
rect 5680 2524 5684 2556
rect 5716 2524 5720 2556
rect 5680 2476 5720 2524
rect 5680 2444 5684 2476
rect 5716 2444 5720 2476
rect 5680 2396 5720 2444
rect 5680 2364 5684 2396
rect 5716 2364 5720 2396
rect 5680 2236 5720 2364
rect 5680 2204 5684 2236
rect 5716 2204 5720 2236
rect 5680 2156 5720 2204
rect 5680 2124 5684 2156
rect 5716 2124 5720 2156
rect 5680 2076 5720 2124
rect 5680 2044 5684 2076
rect 5716 2044 5720 2076
rect 5680 1996 5720 2044
rect 5680 1964 5684 1996
rect 5716 1964 5720 1996
rect 5680 1916 5720 1964
rect 5680 1884 5684 1916
rect 5716 1884 5720 1916
rect 5680 1836 5720 1884
rect 5680 1804 5684 1836
rect 5716 1804 5720 1836
rect 5680 1756 5720 1804
rect 5680 1724 5684 1756
rect 5716 1724 5720 1756
rect 5680 1676 5720 1724
rect 5680 1644 5684 1676
rect 5716 1644 5720 1676
rect 5680 1516 5720 1644
rect 5680 1484 5684 1516
rect 5716 1484 5720 1516
rect 5680 1436 5720 1484
rect 5680 1404 5684 1436
rect 5716 1404 5720 1436
rect 5680 1356 5720 1404
rect 5680 1324 5684 1356
rect 5716 1324 5720 1356
rect 5680 1276 5720 1324
rect 5680 1244 5684 1276
rect 5716 1244 5720 1276
rect 5680 1196 5720 1244
rect 5680 1164 5684 1196
rect 5716 1164 5720 1196
rect 5680 1116 5720 1164
rect 5680 1084 5684 1116
rect 5716 1084 5720 1116
rect 5680 1036 5720 1084
rect 5680 1004 5684 1036
rect 5716 1004 5720 1036
rect 5680 956 5720 1004
rect 5680 924 5684 956
rect 5716 924 5720 956
rect 5680 876 5720 924
rect 5680 844 5684 876
rect 5716 844 5720 876
rect 5680 796 5720 844
rect 5680 764 5684 796
rect 5716 764 5720 796
rect 5680 596 5720 764
rect 5680 564 5684 596
rect 5716 564 5720 596
rect 5680 516 5720 564
rect 5680 484 5684 516
rect 5716 484 5720 516
rect 5680 436 5720 484
rect 5680 404 5684 436
rect 5716 404 5720 436
rect 5680 356 5720 404
rect 5680 324 5684 356
rect 5716 324 5720 356
rect 5680 276 5720 324
rect 5680 244 5684 276
rect 5716 244 5720 276
rect 5680 196 5720 244
rect 5680 164 5684 196
rect 5716 164 5720 196
rect 5680 116 5720 164
rect 5680 84 5684 116
rect 5716 84 5720 116
rect 5680 36 5720 84
rect 5680 4 5684 36
rect 5716 4 5720 36
rect 5680 -40 5720 4
rect 5760 13915 5800 16640
rect 5760 13885 5765 13915
rect 5795 13885 5800 13915
rect 5760 12435 5800 13885
rect 5760 12405 5765 12435
rect 5795 12405 5800 12435
rect 5760 715 5800 12405
rect 5760 685 5765 715
rect 5795 685 5800 715
rect 5760 -40 5800 685
rect 5840 16596 5880 16644
rect 6000 16836 6040 16840
rect 6000 16644 6004 16836
rect 6036 16644 6040 16836
rect 5840 16564 5844 16596
rect 5876 16564 5880 16596
rect 5840 16516 5880 16564
rect 5840 16484 5844 16516
rect 5876 16484 5880 16516
rect 5840 16436 5880 16484
rect 5840 16404 5844 16436
rect 5876 16404 5880 16436
rect 5840 16356 5880 16404
rect 5840 16324 5844 16356
rect 5876 16324 5880 16356
rect 5840 16276 5880 16324
rect 5840 16244 5844 16276
rect 5876 16244 5880 16276
rect 5840 16196 5880 16244
rect 5840 16164 5844 16196
rect 5876 16164 5880 16196
rect 5840 16116 5880 16164
rect 5840 16084 5844 16116
rect 5876 16084 5880 16116
rect 5840 16036 5880 16084
rect 5840 16004 5844 16036
rect 5876 16004 5880 16036
rect 5840 15956 5880 16004
rect 5840 15924 5844 15956
rect 5876 15924 5880 15956
rect 5840 15436 5880 15924
rect 5840 15404 5844 15436
rect 5876 15404 5880 15436
rect 5840 15356 5880 15404
rect 5840 15324 5844 15356
rect 5876 15324 5880 15356
rect 5840 15276 5880 15324
rect 5840 15244 5844 15276
rect 5876 15244 5880 15276
rect 5840 15196 5880 15244
rect 5840 15164 5844 15196
rect 5876 15164 5880 15196
rect 5840 15116 5880 15164
rect 5840 15084 5844 15116
rect 5876 15084 5880 15116
rect 5840 14956 5880 15084
rect 5840 14924 5844 14956
rect 5876 14924 5880 14956
rect 5840 14876 5880 14924
rect 5840 14844 5844 14876
rect 5876 14844 5880 14876
rect 5840 14796 5880 14844
rect 5840 14764 5844 14796
rect 5876 14764 5880 14796
rect 5840 14716 5880 14764
rect 5840 14684 5844 14716
rect 5876 14684 5880 14716
rect 5840 14556 5880 14684
rect 5840 14524 5844 14556
rect 5876 14524 5880 14556
rect 5840 14476 5880 14524
rect 5840 14444 5844 14476
rect 5876 14444 5880 14476
rect 5840 13996 5880 14444
rect 5840 13964 5844 13996
rect 5876 13964 5880 13996
rect 5840 13876 5880 13964
rect 5840 13844 5844 13876
rect 5876 13844 5880 13876
rect 5840 13796 5880 13844
rect 5840 13764 5844 13796
rect 5876 13764 5880 13796
rect 5840 13716 5880 13764
rect 5840 13684 5844 13716
rect 5876 13684 5880 13716
rect 5840 13636 5880 13684
rect 5840 13604 5844 13636
rect 5876 13604 5880 13636
rect 5840 13476 5880 13604
rect 5840 13444 5844 13476
rect 5876 13444 5880 13476
rect 5840 13396 5880 13444
rect 5840 13364 5844 13396
rect 5876 13364 5880 13396
rect 5840 13316 5880 13364
rect 5840 13284 5844 13316
rect 5876 13284 5880 13316
rect 5840 13236 5880 13284
rect 5840 13204 5844 13236
rect 5876 13204 5880 13236
rect 5840 13076 5880 13204
rect 5840 13044 5844 13076
rect 5876 13044 5880 13076
rect 5840 12996 5880 13044
rect 5840 12964 5844 12996
rect 5876 12964 5880 12996
rect 5840 12516 5880 12964
rect 5840 12484 5844 12516
rect 5876 12484 5880 12516
rect 5840 12436 5880 12484
rect 5840 12404 5844 12436
rect 5876 12404 5880 12436
rect 5840 12316 5880 12404
rect 5840 12284 5844 12316
rect 5876 12284 5880 12316
rect 5840 12236 5880 12284
rect 5840 12204 5844 12236
rect 5876 12204 5880 12236
rect 5840 12156 5880 12204
rect 5840 12124 5844 12156
rect 5876 12124 5880 12156
rect 5840 12076 5880 12124
rect 5840 12044 5844 12076
rect 5876 12044 5880 12076
rect 5840 11996 5880 12044
rect 5840 11964 5844 11996
rect 5876 11964 5880 11996
rect 5840 11916 5880 11964
rect 5840 11884 5844 11916
rect 5876 11884 5880 11916
rect 5840 11836 5880 11884
rect 5840 11804 5844 11836
rect 5876 11804 5880 11836
rect 5840 11756 5880 11804
rect 5840 11724 5844 11756
rect 5876 11724 5880 11756
rect 5840 11676 5880 11724
rect 5840 11644 5844 11676
rect 5876 11644 5880 11676
rect 5840 11596 5880 11644
rect 5840 11564 5844 11596
rect 5876 11564 5880 11596
rect 5840 11516 5880 11564
rect 5840 11484 5844 11516
rect 5876 11484 5880 11516
rect 5840 11436 5880 11484
rect 5840 11404 5844 11436
rect 5876 11404 5880 11436
rect 5840 11356 5880 11404
rect 5840 11324 5844 11356
rect 5876 11324 5880 11356
rect 5840 11196 5880 11324
rect 5840 11164 5844 11196
rect 5876 11164 5880 11196
rect 5840 11116 5880 11164
rect 5840 11084 5844 11116
rect 5876 11084 5880 11116
rect 5840 11036 5880 11084
rect 5840 11004 5844 11036
rect 5876 11004 5880 11036
rect 5840 10876 5880 11004
rect 5840 10844 5844 10876
rect 5876 10844 5880 10876
rect 5840 10716 5880 10844
rect 5840 10684 5844 10716
rect 5876 10684 5880 10716
rect 5840 10636 5880 10684
rect 5840 10604 5844 10636
rect 5876 10604 5880 10636
rect 5840 10476 5880 10604
rect 5840 10444 5844 10476
rect 5876 10444 5880 10476
rect 5840 10316 5880 10444
rect 5840 10284 5844 10316
rect 5876 10284 5880 10316
rect 5840 10236 5880 10284
rect 5840 10204 5844 10236
rect 5876 10204 5880 10236
rect 5840 10156 5880 10204
rect 5840 10124 5844 10156
rect 5876 10124 5880 10156
rect 5840 10076 5880 10124
rect 5840 10044 5844 10076
rect 5876 10044 5880 10076
rect 5840 9996 5880 10044
rect 5840 9964 5844 9996
rect 5876 9964 5880 9996
rect 5840 9916 5880 9964
rect 5840 9884 5844 9916
rect 5876 9884 5880 9916
rect 5840 9836 5880 9884
rect 5840 9804 5844 9836
rect 5876 9804 5880 9836
rect 5840 9756 5880 9804
rect 5840 9724 5844 9756
rect 5876 9724 5880 9756
rect 5840 9676 5880 9724
rect 5840 9644 5844 9676
rect 5876 9644 5880 9676
rect 5840 9596 5880 9644
rect 5840 9564 5844 9596
rect 5876 9564 5880 9596
rect 5840 9516 5880 9564
rect 5840 9484 5844 9516
rect 5876 9484 5880 9516
rect 5840 9436 5880 9484
rect 5840 9404 5844 9436
rect 5876 9404 5880 9436
rect 5840 9356 5880 9404
rect 5840 9324 5844 9356
rect 5876 9324 5880 9356
rect 5840 9276 5880 9324
rect 5840 9244 5844 9276
rect 5876 9244 5880 9276
rect 5840 9116 5880 9244
rect 5840 9084 5844 9116
rect 5876 9084 5880 9116
rect 5840 9036 5880 9084
rect 5840 9004 5844 9036
rect 5876 9004 5880 9036
rect 5840 8956 5880 9004
rect 5840 8924 5844 8956
rect 5876 8924 5880 8956
rect 5840 8636 5880 8924
rect 5840 8604 5844 8636
rect 5876 8604 5880 8636
rect 5840 8556 5880 8604
rect 5840 8524 5844 8556
rect 5876 8524 5880 8556
rect 5840 8396 5880 8524
rect 5840 8364 5844 8396
rect 5876 8364 5880 8396
rect 5840 8236 5880 8364
rect 5840 8204 5844 8236
rect 5876 8204 5880 8236
rect 5840 8156 5880 8204
rect 5840 8124 5844 8156
rect 5876 8124 5880 8156
rect 5840 8076 5880 8124
rect 5840 8044 5844 8076
rect 5876 8044 5880 8076
rect 5840 7996 5880 8044
rect 5840 7964 5844 7996
rect 5876 7964 5880 7996
rect 5840 7916 5880 7964
rect 5840 7884 5844 7916
rect 5876 7884 5880 7916
rect 5840 7836 5880 7884
rect 5840 7804 5844 7836
rect 5876 7804 5880 7836
rect 5840 7756 5880 7804
rect 5840 7724 5844 7756
rect 5876 7724 5880 7756
rect 5840 7676 5880 7724
rect 5840 7644 5844 7676
rect 5876 7644 5880 7676
rect 5840 7596 5880 7644
rect 5840 7564 5844 7596
rect 5876 7564 5880 7596
rect 5840 7516 5880 7564
rect 5840 7484 5844 7516
rect 5876 7484 5880 7516
rect 5840 7436 5880 7484
rect 5840 7404 5844 7436
rect 5876 7404 5880 7436
rect 5840 7356 5880 7404
rect 5840 7324 5844 7356
rect 5876 7324 5880 7356
rect 5840 7276 5880 7324
rect 5840 7244 5844 7276
rect 5876 7244 5880 7276
rect 5840 7196 5880 7244
rect 5840 7164 5844 7196
rect 5876 7164 5880 7196
rect 5840 7036 5880 7164
rect 5840 7004 5844 7036
rect 5876 7004 5880 7036
rect 5840 6956 5880 7004
rect 5840 6924 5844 6956
rect 5876 6924 5880 6956
rect 5840 6796 5880 6924
rect 5840 6764 5844 6796
rect 5876 6764 5880 6796
rect 5840 6716 5880 6764
rect 5840 6684 5844 6716
rect 5876 6684 5880 6716
rect 5840 6636 5880 6684
rect 5840 6604 5844 6636
rect 5876 6604 5880 6636
rect 5840 6556 5880 6604
rect 5840 6524 5844 6556
rect 5876 6524 5880 6556
rect 5840 6476 5880 6524
rect 5840 6444 5844 6476
rect 5876 6444 5880 6476
rect 5840 6316 5880 6444
rect 5840 6284 5844 6316
rect 5876 6284 5880 6316
rect 5840 6236 5880 6284
rect 5840 6204 5844 6236
rect 5876 6204 5880 6236
rect 5840 6156 5880 6204
rect 5840 6124 5844 6156
rect 5876 6124 5880 6156
rect 5840 5996 5880 6124
rect 5840 5964 5844 5996
rect 5876 5964 5880 5996
rect 5840 5836 5880 5964
rect 5840 5804 5844 5836
rect 5876 5804 5880 5836
rect 5840 5756 5880 5804
rect 5840 5724 5844 5756
rect 5876 5724 5880 5756
rect 5840 5676 5880 5724
rect 5840 5644 5844 5676
rect 5876 5644 5880 5676
rect 5840 5596 5880 5644
rect 5840 5564 5844 5596
rect 5876 5564 5880 5596
rect 5840 5516 5880 5564
rect 5840 5484 5844 5516
rect 5876 5484 5880 5516
rect 5840 5436 5880 5484
rect 5840 5404 5844 5436
rect 5876 5404 5880 5436
rect 5840 5356 5880 5404
rect 5840 5324 5844 5356
rect 5876 5324 5880 5356
rect 5840 5276 5880 5324
rect 5840 5244 5844 5276
rect 5876 5244 5880 5276
rect 5840 5196 5880 5244
rect 5840 5164 5844 5196
rect 5876 5164 5880 5196
rect 5840 5116 5880 5164
rect 5840 5084 5844 5116
rect 5876 5084 5880 5116
rect 5840 5036 5880 5084
rect 5840 5004 5844 5036
rect 5876 5004 5880 5036
rect 5840 4956 5880 5004
rect 5840 4924 5844 4956
rect 5876 4924 5880 4956
rect 5840 4876 5880 4924
rect 5840 4844 5844 4876
rect 5876 4844 5880 4876
rect 5840 4796 5880 4844
rect 5840 4764 5844 4796
rect 5876 4764 5880 4796
rect 5840 4636 5880 4764
rect 5840 4604 5844 4636
rect 5876 4604 5880 4636
rect 5840 4556 5880 4604
rect 5840 4524 5844 4556
rect 5876 4524 5880 4556
rect 5840 4396 5880 4524
rect 5840 4364 5844 4396
rect 5876 4364 5880 4396
rect 5840 4316 5880 4364
rect 5840 4284 5844 4316
rect 5876 4284 5880 4316
rect 5840 4236 5880 4284
rect 5840 4204 5844 4236
rect 5876 4204 5880 4236
rect 5840 4156 5880 4204
rect 5840 4124 5844 4156
rect 5876 4124 5880 4156
rect 5840 4076 5880 4124
rect 5840 4044 5844 4076
rect 5876 4044 5880 4076
rect 5840 3916 5880 4044
rect 5840 3884 5844 3916
rect 5876 3884 5880 3916
rect 5840 3836 5880 3884
rect 5840 3804 5844 3836
rect 5876 3804 5880 3836
rect 5840 3756 5880 3804
rect 5840 3724 5844 3756
rect 5876 3724 5880 3756
rect 5840 3596 5880 3724
rect 5840 3564 5844 3596
rect 5876 3564 5880 3596
rect 5840 3436 5880 3564
rect 5840 3404 5844 3436
rect 5876 3404 5880 3436
rect 5840 3356 5880 3404
rect 5840 3324 5844 3356
rect 5876 3324 5880 3356
rect 5840 3276 5880 3324
rect 5840 3244 5844 3276
rect 5876 3244 5880 3276
rect 5840 3196 5880 3244
rect 5840 3164 5844 3196
rect 5876 3164 5880 3196
rect 5840 3116 5880 3164
rect 5840 3084 5844 3116
rect 5876 3084 5880 3116
rect 5840 3036 5880 3084
rect 5840 3004 5844 3036
rect 5876 3004 5880 3036
rect 5840 2956 5880 3004
rect 5840 2924 5844 2956
rect 5876 2924 5880 2956
rect 5840 2876 5880 2924
rect 5840 2844 5844 2876
rect 5876 2844 5880 2876
rect 5840 2796 5880 2844
rect 5840 2764 5844 2796
rect 5876 2764 5880 2796
rect 5840 2716 5880 2764
rect 5840 2684 5844 2716
rect 5876 2684 5880 2716
rect 5840 2636 5880 2684
rect 5840 2604 5844 2636
rect 5876 2604 5880 2636
rect 5840 2556 5880 2604
rect 5840 2524 5844 2556
rect 5876 2524 5880 2556
rect 5840 2476 5880 2524
rect 5840 2444 5844 2476
rect 5876 2444 5880 2476
rect 5840 2396 5880 2444
rect 5840 2364 5844 2396
rect 5876 2364 5880 2396
rect 5840 2236 5880 2364
rect 5840 2204 5844 2236
rect 5876 2204 5880 2236
rect 5840 2156 5880 2204
rect 5840 2124 5844 2156
rect 5876 2124 5880 2156
rect 5840 2076 5880 2124
rect 5840 2044 5844 2076
rect 5876 2044 5880 2076
rect 5840 1996 5880 2044
rect 5840 1964 5844 1996
rect 5876 1964 5880 1996
rect 5840 1916 5880 1964
rect 5840 1884 5844 1916
rect 5876 1884 5880 1916
rect 5840 1836 5880 1884
rect 5840 1804 5844 1836
rect 5876 1804 5880 1836
rect 5840 1756 5880 1804
rect 5840 1724 5844 1756
rect 5876 1724 5880 1756
rect 5840 1676 5880 1724
rect 5840 1644 5844 1676
rect 5876 1644 5880 1676
rect 5840 1516 5880 1644
rect 5840 1484 5844 1516
rect 5876 1484 5880 1516
rect 5840 1436 5880 1484
rect 5840 1404 5844 1436
rect 5876 1404 5880 1436
rect 5840 1356 5880 1404
rect 5840 1324 5844 1356
rect 5876 1324 5880 1356
rect 5840 1276 5880 1324
rect 5840 1244 5844 1276
rect 5876 1244 5880 1276
rect 5840 1196 5880 1244
rect 5840 1164 5844 1196
rect 5876 1164 5880 1196
rect 5840 1116 5880 1164
rect 5840 1084 5844 1116
rect 5876 1084 5880 1116
rect 5840 1036 5880 1084
rect 5840 1004 5844 1036
rect 5876 1004 5880 1036
rect 5840 956 5880 1004
rect 5840 924 5844 956
rect 5876 924 5880 956
rect 5840 876 5880 924
rect 5840 844 5844 876
rect 5876 844 5880 876
rect 5840 796 5880 844
rect 5840 764 5844 796
rect 5876 764 5880 796
rect 5840 716 5880 764
rect 5840 684 5844 716
rect 5876 684 5880 716
rect 5840 596 5880 684
rect 5840 564 5844 596
rect 5876 564 5880 596
rect 5840 516 5880 564
rect 5840 484 5844 516
rect 5876 484 5880 516
rect 5840 436 5880 484
rect 5840 404 5844 436
rect 5876 404 5880 436
rect 5840 356 5880 404
rect 5840 324 5844 356
rect 5876 324 5880 356
rect 5840 276 5880 324
rect 5840 244 5844 276
rect 5876 244 5880 276
rect 5840 196 5880 244
rect 5840 164 5844 196
rect 5876 164 5880 196
rect 5840 116 5880 164
rect 5840 84 5844 116
rect 5876 84 5880 116
rect 5840 36 5880 84
rect 5840 4 5844 36
rect 5876 4 5880 36
rect 5840 -40 5880 4
rect 5920 14635 5960 16640
rect 5920 14605 5925 14635
rect 5955 14605 5960 14635
rect 5920 13155 5960 14605
rect 5920 13125 5925 13155
rect 5955 13125 5960 13155
rect 5920 1595 5960 13125
rect 5920 1565 5925 1595
rect 5955 1565 5960 1595
rect 5920 -40 5960 1565
rect 6000 16596 6040 16644
rect 6160 16836 6200 16840
rect 6160 16644 6164 16836
rect 6196 16644 6200 16836
rect 6000 16564 6004 16596
rect 6036 16564 6040 16596
rect 6000 16516 6040 16564
rect 6000 16484 6004 16516
rect 6036 16484 6040 16516
rect 6000 16436 6040 16484
rect 6000 16404 6004 16436
rect 6036 16404 6040 16436
rect 6000 16356 6040 16404
rect 6000 16324 6004 16356
rect 6036 16324 6040 16356
rect 6000 16276 6040 16324
rect 6000 16244 6004 16276
rect 6036 16244 6040 16276
rect 6000 16196 6040 16244
rect 6000 16164 6004 16196
rect 6036 16164 6040 16196
rect 6000 16116 6040 16164
rect 6000 16084 6004 16116
rect 6036 16084 6040 16116
rect 6000 16036 6040 16084
rect 6000 16004 6004 16036
rect 6036 16004 6040 16036
rect 6000 15956 6040 16004
rect 6000 15924 6004 15956
rect 6036 15924 6040 15956
rect 6000 15436 6040 15924
rect 6000 15404 6004 15436
rect 6036 15404 6040 15436
rect 6000 15356 6040 15404
rect 6000 15324 6004 15356
rect 6036 15324 6040 15356
rect 6000 15276 6040 15324
rect 6000 15244 6004 15276
rect 6036 15244 6040 15276
rect 6000 15196 6040 15244
rect 6000 15164 6004 15196
rect 6036 15164 6040 15196
rect 6000 15116 6040 15164
rect 6000 15084 6004 15116
rect 6036 15084 6040 15116
rect 6000 14956 6040 15084
rect 6000 14924 6004 14956
rect 6036 14924 6040 14956
rect 6000 14876 6040 14924
rect 6000 14844 6004 14876
rect 6036 14844 6040 14876
rect 6000 14796 6040 14844
rect 6000 14764 6004 14796
rect 6036 14764 6040 14796
rect 6000 14716 6040 14764
rect 6000 14684 6004 14716
rect 6036 14684 6040 14716
rect 6000 14636 6040 14684
rect 6000 14604 6004 14636
rect 6036 14604 6040 14636
rect 6000 14556 6040 14604
rect 6000 14524 6004 14556
rect 6036 14524 6040 14556
rect 6000 14476 6040 14524
rect 6000 14444 6004 14476
rect 6036 14444 6040 14476
rect 6000 13996 6040 14444
rect 6000 13964 6004 13996
rect 6036 13964 6040 13996
rect 6000 13876 6040 13964
rect 6000 13844 6004 13876
rect 6036 13844 6040 13876
rect 6000 13796 6040 13844
rect 6000 13764 6004 13796
rect 6036 13764 6040 13796
rect 6000 13716 6040 13764
rect 6000 13684 6004 13716
rect 6036 13684 6040 13716
rect 6000 13636 6040 13684
rect 6000 13604 6004 13636
rect 6036 13604 6040 13636
rect 6000 13476 6040 13604
rect 6000 13444 6004 13476
rect 6036 13444 6040 13476
rect 6000 13396 6040 13444
rect 6000 13364 6004 13396
rect 6036 13364 6040 13396
rect 6000 13316 6040 13364
rect 6000 13284 6004 13316
rect 6036 13284 6040 13316
rect 6000 13236 6040 13284
rect 6000 13204 6004 13236
rect 6036 13204 6040 13236
rect 6000 13156 6040 13204
rect 6000 13124 6004 13156
rect 6036 13124 6040 13156
rect 6000 13076 6040 13124
rect 6000 13044 6004 13076
rect 6036 13044 6040 13076
rect 6000 12996 6040 13044
rect 6000 12964 6004 12996
rect 6036 12964 6040 12996
rect 6000 12516 6040 12964
rect 6000 12484 6004 12516
rect 6036 12484 6040 12516
rect 6000 12436 6040 12484
rect 6000 12404 6004 12436
rect 6036 12404 6040 12436
rect 6000 12316 6040 12404
rect 6000 12284 6004 12316
rect 6036 12284 6040 12316
rect 6000 12236 6040 12284
rect 6000 12204 6004 12236
rect 6036 12204 6040 12236
rect 6000 12156 6040 12204
rect 6000 12124 6004 12156
rect 6036 12124 6040 12156
rect 6000 12076 6040 12124
rect 6000 12044 6004 12076
rect 6036 12044 6040 12076
rect 6000 11996 6040 12044
rect 6000 11964 6004 11996
rect 6036 11964 6040 11996
rect 6000 11916 6040 11964
rect 6000 11884 6004 11916
rect 6036 11884 6040 11916
rect 6000 11836 6040 11884
rect 6000 11804 6004 11836
rect 6036 11804 6040 11836
rect 6000 11756 6040 11804
rect 6000 11724 6004 11756
rect 6036 11724 6040 11756
rect 6000 11676 6040 11724
rect 6000 11644 6004 11676
rect 6036 11644 6040 11676
rect 6000 11596 6040 11644
rect 6000 11564 6004 11596
rect 6036 11564 6040 11596
rect 6000 11516 6040 11564
rect 6000 11484 6004 11516
rect 6036 11484 6040 11516
rect 6000 11436 6040 11484
rect 6000 11404 6004 11436
rect 6036 11404 6040 11436
rect 6000 11356 6040 11404
rect 6000 11324 6004 11356
rect 6036 11324 6040 11356
rect 6000 11196 6040 11324
rect 6000 11164 6004 11196
rect 6036 11164 6040 11196
rect 6000 11116 6040 11164
rect 6000 11084 6004 11116
rect 6036 11084 6040 11116
rect 6000 11036 6040 11084
rect 6000 11004 6004 11036
rect 6036 11004 6040 11036
rect 6000 10876 6040 11004
rect 6000 10844 6004 10876
rect 6036 10844 6040 10876
rect 6000 10716 6040 10844
rect 6000 10684 6004 10716
rect 6036 10684 6040 10716
rect 6000 10636 6040 10684
rect 6000 10604 6004 10636
rect 6036 10604 6040 10636
rect 6000 10476 6040 10604
rect 6000 10444 6004 10476
rect 6036 10444 6040 10476
rect 6000 10316 6040 10444
rect 6000 10284 6004 10316
rect 6036 10284 6040 10316
rect 6000 10236 6040 10284
rect 6000 10204 6004 10236
rect 6036 10204 6040 10236
rect 6000 10156 6040 10204
rect 6000 10124 6004 10156
rect 6036 10124 6040 10156
rect 6000 10076 6040 10124
rect 6000 10044 6004 10076
rect 6036 10044 6040 10076
rect 6000 9996 6040 10044
rect 6000 9964 6004 9996
rect 6036 9964 6040 9996
rect 6000 9916 6040 9964
rect 6000 9884 6004 9916
rect 6036 9884 6040 9916
rect 6000 9836 6040 9884
rect 6000 9804 6004 9836
rect 6036 9804 6040 9836
rect 6000 9756 6040 9804
rect 6000 9724 6004 9756
rect 6036 9724 6040 9756
rect 6000 9676 6040 9724
rect 6000 9644 6004 9676
rect 6036 9644 6040 9676
rect 6000 9596 6040 9644
rect 6000 9564 6004 9596
rect 6036 9564 6040 9596
rect 6000 9516 6040 9564
rect 6000 9484 6004 9516
rect 6036 9484 6040 9516
rect 6000 9436 6040 9484
rect 6000 9404 6004 9436
rect 6036 9404 6040 9436
rect 6000 9356 6040 9404
rect 6000 9324 6004 9356
rect 6036 9324 6040 9356
rect 6000 9276 6040 9324
rect 6000 9244 6004 9276
rect 6036 9244 6040 9276
rect 6000 9116 6040 9244
rect 6000 9084 6004 9116
rect 6036 9084 6040 9116
rect 6000 9036 6040 9084
rect 6000 9004 6004 9036
rect 6036 9004 6040 9036
rect 6000 8956 6040 9004
rect 6000 8924 6004 8956
rect 6036 8924 6040 8956
rect 6000 8636 6040 8924
rect 6000 8604 6004 8636
rect 6036 8604 6040 8636
rect 6000 8556 6040 8604
rect 6000 8524 6004 8556
rect 6036 8524 6040 8556
rect 6000 8396 6040 8524
rect 6000 8364 6004 8396
rect 6036 8364 6040 8396
rect 6000 8236 6040 8364
rect 6000 8204 6004 8236
rect 6036 8204 6040 8236
rect 6000 8156 6040 8204
rect 6000 8124 6004 8156
rect 6036 8124 6040 8156
rect 6000 8076 6040 8124
rect 6000 8044 6004 8076
rect 6036 8044 6040 8076
rect 6000 7996 6040 8044
rect 6000 7964 6004 7996
rect 6036 7964 6040 7996
rect 6000 7916 6040 7964
rect 6000 7884 6004 7916
rect 6036 7884 6040 7916
rect 6000 7836 6040 7884
rect 6000 7804 6004 7836
rect 6036 7804 6040 7836
rect 6000 7756 6040 7804
rect 6000 7724 6004 7756
rect 6036 7724 6040 7756
rect 6000 7676 6040 7724
rect 6000 7644 6004 7676
rect 6036 7644 6040 7676
rect 6000 7596 6040 7644
rect 6000 7564 6004 7596
rect 6036 7564 6040 7596
rect 6000 7516 6040 7564
rect 6000 7484 6004 7516
rect 6036 7484 6040 7516
rect 6000 7436 6040 7484
rect 6000 7404 6004 7436
rect 6036 7404 6040 7436
rect 6000 7356 6040 7404
rect 6000 7324 6004 7356
rect 6036 7324 6040 7356
rect 6000 7276 6040 7324
rect 6000 7244 6004 7276
rect 6036 7244 6040 7276
rect 6000 7196 6040 7244
rect 6000 7164 6004 7196
rect 6036 7164 6040 7196
rect 6000 7036 6040 7164
rect 6000 7004 6004 7036
rect 6036 7004 6040 7036
rect 6000 6956 6040 7004
rect 6000 6924 6004 6956
rect 6036 6924 6040 6956
rect 6000 6796 6040 6924
rect 6000 6764 6004 6796
rect 6036 6764 6040 6796
rect 6000 6716 6040 6764
rect 6000 6684 6004 6716
rect 6036 6684 6040 6716
rect 6000 6636 6040 6684
rect 6000 6604 6004 6636
rect 6036 6604 6040 6636
rect 6000 6556 6040 6604
rect 6000 6524 6004 6556
rect 6036 6524 6040 6556
rect 6000 6476 6040 6524
rect 6000 6444 6004 6476
rect 6036 6444 6040 6476
rect 6000 6316 6040 6444
rect 6000 6284 6004 6316
rect 6036 6284 6040 6316
rect 6000 6236 6040 6284
rect 6000 6204 6004 6236
rect 6036 6204 6040 6236
rect 6000 6156 6040 6204
rect 6000 6124 6004 6156
rect 6036 6124 6040 6156
rect 6000 5996 6040 6124
rect 6000 5964 6004 5996
rect 6036 5964 6040 5996
rect 6000 5836 6040 5964
rect 6000 5804 6004 5836
rect 6036 5804 6040 5836
rect 6000 5756 6040 5804
rect 6000 5724 6004 5756
rect 6036 5724 6040 5756
rect 6000 5676 6040 5724
rect 6000 5644 6004 5676
rect 6036 5644 6040 5676
rect 6000 5596 6040 5644
rect 6000 5564 6004 5596
rect 6036 5564 6040 5596
rect 6000 5516 6040 5564
rect 6000 5484 6004 5516
rect 6036 5484 6040 5516
rect 6000 5436 6040 5484
rect 6000 5404 6004 5436
rect 6036 5404 6040 5436
rect 6000 5356 6040 5404
rect 6000 5324 6004 5356
rect 6036 5324 6040 5356
rect 6000 5276 6040 5324
rect 6000 5244 6004 5276
rect 6036 5244 6040 5276
rect 6000 5196 6040 5244
rect 6000 5164 6004 5196
rect 6036 5164 6040 5196
rect 6000 5116 6040 5164
rect 6000 5084 6004 5116
rect 6036 5084 6040 5116
rect 6000 5036 6040 5084
rect 6000 5004 6004 5036
rect 6036 5004 6040 5036
rect 6000 4956 6040 5004
rect 6000 4924 6004 4956
rect 6036 4924 6040 4956
rect 6000 4876 6040 4924
rect 6000 4844 6004 4876
rect 6036 4844 6040 4876
rect 6000 4796 6040 4844
rect 6000 4764 6004 4796
rect 6036 4764 6040 4796
rect 6000 4636 6040 4764
rect 6000 4604 6004 4636
rect 6036 4604 6040 4636
rect 6000 4556 6040 4604
rect 6000 4524 6004 4556
rect 6036 4524 6040 4556
rect 6000 4396 6040 4524
rect 6000 4364 6004 4396
rect 6036 4364 6040 4396
rect 6000 4316 6040 4364
rect 6000 4284 6004 4316
rect 6036 4284 6040 4316
rect 6000 4236 6040 4284
rect 6000 4204 6004 4236
rect 6036 4204 6040 4236
rect 6000 4156 6040 4204
rect 6000 4124 6004 4156
rect 6036 4124 6040 4156
rect 6000 4076 6040 4124
rect 6000 4044 6004 4076
rect 6036 4044 6040 4076
rect 6000 3916 6040 4044
rect 6000 3884 6004 3916
rect 6036 3884 6040 3916
rect 6000 3836 6040 3884
rect 6000 3804 6004 3836
rect 6036 3804 6040 3836
rect 6000 3756 6040 3804
rect 6000 3724 6004 3756
rect 6036 3724 6040 3756
rect 6000 3596 6040 3724
rect 6000 3564 6004 3596
rect 6036 3564 6040 3596
rect 6000 3436 6040 3564
rect 6000 3404 6004 3436
rect 6036 3404 6040 3436
rect 6000 3356 6040 3404
rect 6000 3324 6004 3356
rect 6036 3324 6040 3356
rect 6000 3276 6040 3324
rect 6000 3244 6004 3276
rect 6036 3244 6040 3276
rect 6000 3196 6040 3244
rect 6000 3164 6004 3196
rect 6036 3164 6040 3196
rect 6000 3116 6040 3164
rect 6000 3084 6004 3116
rect 6036 3084 6040 3116
rect 6000 3036 6040 3084
rect 6000 3004 6004 3036
rect 6036 3004 6040 3036
rect 6000 2956 6040 3004
rect 6000 2924 6004 2956
rect 6036 2924 6040 2956
rect 6000 2876 6040 2924
rect 6000 2844 6004 2876
rect 6036 2844 6040 2876
rect 6000 2796 6040 2844
rect 6000 2764 6004 2796
rect 6036 2764 6040 2796
rect 6000 2716 6040 2764
rect 6000 2684 6004 2716
rect 6036 2684 6040 2716
rect 6000 2636 6040 2684
rect 6000 2604 6004 2636
rect 6036 2604 6040 2636
rect 6000 2556 6040 2604
rect 6000 2524 6004 2556
rect 6036 2524 6040 2556
rect 6000 2476 6040 2524
rect 6000 2444 6004 2476
rect 6036 2444 6040 2476
rect 6000 2396 6040 2444
rect 6000 2364 6004 2396
rect 6036 2364 6040 2396
rect 6000 2236 6040 2364
rect 6000 2204 6004 2236
rect 6036 2204 6040 2236
rect 6000 2156 6040 2204
rect 6000 2124 6004 2156
rect 6036 2124 6040 2156
rect 6000 2076 6040 2124
rect 6000 2044 6004 2076
rect 6036 2044 6040 2076
rect 6000 1996 6040 2044
rect 6000 1964 6004 1996
rect 6036 1964 6040 1996
rect 6000 1916 6040 1964
rect 6000 1884 6004 1916
rect 6036 1884 6040 1916
rect 6000 1836 6040 1884
rect 6000 1804 6004 1836
rect 6036 1804 6040 1836
rect 6000 1756 6040 1804
rect 6000 1724 6004 1756
rect 6036 1724 6040 1756
rect 6000 1676 6040 1724
rect 6000 1644 6004 1676
rect 6036 1644 6040 1676
rect 6000 1596 6040 1644
rect 6000 1564 6004 1596
rect 6036 1564 6040 1596
rect 6000 1516 6040 1564
rect 6000 1484 6004 1516
rect 6036 1484 6040 1516
rect 6000 1436 6040 1484
rect 6000 1404 6004 1436
rect 6036 1404 6040 1436
rect 6000 1356 6040 1404
rect 6000 1324 6004 1356
rect 6036 1324 6040 1356
rect 6000 1276 6040 1324
rect 6000 1244 6004 1276
rect 6036 1244 6040 1276
rect 6000 1196 6040 1244
rect 6000 1164 6004 1196
rect 6036 1164 6040 1196
rect 6000 1116 6040 1164
rect 6000 1084 6004 1116
rect 6036 1084 6040 1116
rect 6000 1036 6040 1084
rect 6000 1004 6004 1036
rect 6036 1004 6040 1036
rect 6000 956 6040 1004
rect 6000 924 6004 956
rect 6036 924 6040 956
rect 6000 876 6040 924
rect 6000 844 6004 876
rect 6036 844 6040 876
rect 6000 796 6040 844
rect 6000 764 6004 796
rect 6036 764 6040 796
rect 6000 716 6040 764
rect 6000 684 6004 716
rect 6036 684 6040 716
rect 6000 596 6040 684
rect 6000 564 6004 596
rect 6036 564 6040 596
rect 6000 516 6040 564
rect 6000 484 6004 516
rect 6036 484 6040 516
rect 6000 436 6040 484
rect 6000 404 6004 436
rect 6036 404 6040 436
rect 6000 356 6040 404
rect 6000 324 6004 356
rect 6036 324 6040 356
rect 6000 276 6040 324
rect 6000 244 6004 276
rect 6036 244 6040 276
rect 6000 196 6040 244
rect 6000 164 6004 196
rect 6036 164 6040 196
rect 6000 116 6040 164
rect 6000 84 6004 116
rect 6036 84 6040 116
rect 6000 36 6040 84
rect 6000 4 6004 36
rect 6036 4 6040 36
rect 6000 -40 6040 4
rect 6080 15035 6120 16640
rect 6080 15005 6085 15035
rect 6115 15005 6120 15035
rect 6080 13555 6120 15005
rect 6080 13525 6085 13555
rect 6115 13525 6120 13555
rect 6080 7115 6120 13525
rect 6080 7085 6085 7115
rect 6115 7085 6120 7115
rect 6080 4715 6120 7085
rect 6080 4685 6085 4715
rect 6115 4685 6120 4715
rect 6080 2315 6120 4685
rect 6080 2285 6085 2315
rect 6115 2285 6120 2315
rect 6080 -40 6120 2285
rect 6160 16596 6200 16644
rect 6320 16836 6360 16840
rect 6320 16644 6324 16836
rect 6356 16644 6360 16836
rect 6160 16564 6164 16596
rect 6196 16564 6200 16596
rect 6160 16516 6200 16564
rect 6160 16484 6164 16516
rect 6196 16484 6200 16516
rect 6160 16436 6200 16484
rect 6160 16404 6164 16436
rect 6196 16404 6200 16436
rect 6160 16356 6200 16404
rect 6160 16324 6164 16356
rect 6196 16324 6200 16356
rect 6160 16276 6200 16324
rect 6160 16244 6164 16276
rect 6196 16244 6200 16276
rect 6160 16196 6200 16244
rect 6160 16164 6164 16196
rect 6196 16164 6200 16196
rect 6160 16116 6200 16164
rect 6160 16084 6164 16116
rect 6196 16084 6200 16116
rect 6160 16036 6200 16084
rect 6160 16004 6164 16036
rect 6196 16004 6200 16036
rect 6160 15956 6200 16004
rect 6160 15924 6164 15956
rect 6196 15924 6200 15956
rect 6160 15436 6200 15924
rect 6160 15404 6164 15436
rect 6196 15404 6200 15436
rect 6160 15356 6200 15404
rect 6160 15324 6164 15356
rect 6196 15324 6200 15356
rect 6160 15276 6200 15324
rect 6160 15244 6164 15276
rect 6196 15244 6200 15276
rect 6160 15196 6200 15244
rect 6160 15164 6164 15196
rect 6196 15164 6200 15196
rect 6160 15116 6200 15164
rect 6160 15084 6164 15116
rect 6196 15084 6200 15116
rect 6160 15036 6200 15084
rect 6160 15004 6164 15036
rect 6196 15004 6200 15036
rect 6160 14956 6200 15004
rect 6160 14924 6164 14956
rect 6196 14924 6200 14956
rect 6160 14876 6200 14924
rect 6160 14844 6164 14876
rect 6196 14844 6200 14876
rect 6160 14796 6200 14844
rect 6160 14764 6164 14796
rect 6196 14764 6200 14796
rect 6160 14716 6200 14764
rect 6160 14684 6164 14716
rect 6196 14684 6200 14716
rect 6160 14636 6200 14684
rect 6160 14604 6164 14636
rect 6196 14604 6200 14636
rect 6160 14556 6200 14604
rect 6160 14524 6164 14556
rect 6196 14524 6200 14556
rect 6160 14476 6200 14524
rect 6160 14444 6164 14476
rect 6196 14444 6200 14476
rect 6160 13996 6200 14444
rect 6160 13964 6164 13996
rect 6196 13964 6200 13996
rect 6160 13876 6200 13964
rect 6160 13844 6164 13876
rect 6196 13844 6200 13876
rect 6160 13796 6200 13844
rect 6160 13764 6164 13796
rect 6196 13764 6200 13796
rect 6160 13716 6200 13764
rect 6160 13684 6164 13716
rect 6196 13684 6200 13716
rect 6160 13636 6200 13684
rect 6160 13604 6164 13636
rect 6196 13604 6200 13636
rect 6160 13556 6200 13604
rect 6160 13524 6164 13556
rect 6196 13524 6200 13556
rect 6160 13476 6200 13524
rect 6160 13444 6164 13476
rect 6196 13444 6200 13476
rect 6160 13396 6200 13444
rect 6160 13364 6164 13396
rect 6196 13364 6200 13396
rect 6160 13316 6200 13364
rect 6160 13284 6164 13316
rect 6196 13284 6200 13316
rect 6160 13236 6200 13284
rect 6160 13204 6164 13236
rect 6196 13204 6200 13236
rect 6160 13156 6200 13204
rect 6160 13124 6164 13156
rect 6196 13124 6200 13156
rect 6160 13076 6200 13124
rect 6160 13044 6164 13076
rect 6196 13044 6200 13076
rect 6160 12996 6200 13044
rect 6160 12964 6164 12996
rect 6196 12964 6200 12996
rect 6160 12516 6200 12964
rect 6160 12484 6164 12516
rect 6196 12484 6200 12516
rect 6160 12436 6200 12484
rect 6160 12404 6164 12436
rect 6196 12404 6200 12436
rect 6160 12316 6200 12404
rect 6160 12284 6164 12316
rect 6196 12284 6200 12316
rect 6160 12236 6200 12284
rect 6160 12204 6164 12236
rect 6196 12204 6200 12236
rect 6160 12156 6200 12204
rect 6160 12124 6164 12156
rect 6196 12124 6200 12156
rect 6160 12076 6200 12124
rect 6160 12044 6164 12076
rect 6196 12044 6200 12076
rect 6160 11996 6200 12044
rect 6160 11964 6164 11996
rect 6196 11964 6200 11996
rect 6160 11916 6200 11964
rect 6160 11884 6164 11916
rect 6196 11884 6200 11916
rect 6160 11836 6200 11884
rect 6160 11804 6164 11836
rect 6196 11804 6200 11836
rect 6160 11756 6200 11804
rect 6160 11724 6164 11756
rect 6196 11724 6200 11756
rect 6160 11676 6200 11724
rect 6160 11644 6164 11676
rect 6196 11644 6200 11676
rect 6160 11596 6200 11644
rect 6160 11564 6164 11596
rect 6196 11564 6200 11596
rect 6160 11516 6200 11564
rect 6160 11484 6164 11516
rect 6196 11484 6200 11516
rect 6160 11436 6200 11484
rect 6160 11404 6164 11436
rect 6196 11404 6200 11436
rect 6160 11356 6200 11404
rect 6160 11324 6164 11356
rect 6196 11324 6200 11356
rect 6160 11196 6200 11324
rect 6160 11164 6164 11196
rect 6196 11164 6200 11196
rect 6160 11116 6200 11164
rect 6160 11084 6164 11116
rect 6196 11084 6200 11116
rect 6160 11036 6200 11084
rect 6160 11004 6164 11036
rect 6196 11004 6200 11036
rect 6160 10876 6200 11004
rect 6160 10844 6164 10876
rect 6196 10844 6200 10876
rect 6160 10716 6200 10844
rect 6160 10684 6164 10716
rect 6196 10684 6200 10716
rect 6160 10636 6200 10684
rect 6160 10604 6164 10636
rect 6196 10604 6200 10636
rect 6160 10476 6200 10604
rect 6160 10444 6164 10476
rect 6196 10444 6200 10476
rect 6160 10316 6200 10444
rect 6160 10284 6164 10316
rect 6196 10284 6200 10316
rect 6160 10236 6200 10284
rect 6160 10204 6164 10236
rect 6196 10204 6200 10236
rect 6160 10156 6200 10204
rect 6160 10124 6164 10156
rect 6196 10124 6200 10156
rect 6160 10076 6200 10124
rect 6160 10044 6164 10076
rect 6196 10044 6200 10076
rect 6160 9996 6200 10044
rect 6160 9964 6164 9996
rect 6196 9964 6200 9996
rect 6160 9916 6200 9964
rect 6160 9884 6164 9916
rect 6196 9884 6200 9916
rect 6160 9836 6200 9884
rect 6160 9804 6164 9836
rect 6196 9804 6200 9836
rect 6160 9756 6200 9804
rect 6160 9724 6164 9756
rect 6196 9724 6200 9756
rect 6160 9676 6200 9724
rect 6160 9644 6164 9676
rect 6196 9644 6200 9676
rect 6160 9596 6200 9644
rect 6160 9564 6164 9596
rect 6196 9564 6200 9596
rect 6160 9516 6200 9564
rect 6160 9484 6164 9516
rect 6196 9484 6200 9516
rect 6160 9436 6200 9484
rect 6160 9404 6164 9436
rect 6196 9404 6200 9436
rect 6160 9356 6200 9404
rect 6160 9324 6164 9356
rect 6196 9324 6200 9356
rect 6160 9276 6200 9324
rect 6160 9244 6164 9276
rect 6196 9244 6200 9276
rect 6160 9116 6200 9244
rect 6160 9084 6164 9116
rect 6196 9084 6200 9116
rect 6160 9036 6200 9084
rect 6160 9004 6164 9036
rect 6196 9004 6200 9036
rect 6160 8956 6200 9004
rect 6160 8924 6164 8956
rect 6196 8924 6200 8956
rect 6160 8636 6200 8924
rect 6160 8604 6164 8636
rect 6196 8604 6200 8636
rect 6160 8556 6200 8604
rect 6160 8524 6164 8556
rect 6196 8524 6200 8556
rect 6160 8396 6200 8524
rect 6160 8364 6164 8396
rect 6196 8364 6200 8396
rect 6160 8236 6200 8364
rect 6160 8204 6164 8236
rect 6196 8204 6200 8236
rect 6160 8156 6200 8204
rect 6160 8124 6164 8156
rect 6196 8124 6200 8156
rect 6160 8076 6200 8124
rect 6160 8044 6164 8076
rect 6196 8044 6200 8076
rect 6160 7996 6200 8044
rect 6160 7964 6164 7996
rect 6196 7964 6200 7996
rect 6160 7916 6200 7964
rect 6160 7884 6164 7916
rect 6196 7884 6200 7916
rect 6160 7836 6200 7884
rect 6160 7804 6164 7836
rect 6196 7804 6200 7836
rect 6160 7756 6200 7804
rect 6160 7724 6164 7756
rect 6196 7724 6200 7756
rect 6160 7676 6200 7724
rect 6160 7644 6164 7676
rect 6196 7644 6200 7676
rect 6160 7596 6200 7644
rect 6160 7564 6164 7596
rect 6196 7564 6200 7596
rect 6160 7516 6200 7564
rect 6160 7484 6164 7516
rect 6196 7484 6200 7516
rect 6160 7436 6200 7484
rect 6160 7404 6164 7436
rect 6196 7404 6200 7436
rect 6160 7356 6200 7404
rect 6160 7324 6164 7356
rect 6196 7324 6200 7356
rect 6160 7276 6200 7324
rect 6160 7244 6164 7276
rect 6196 7244 6200 7276
rect 6160 7196 6200 7244
rect 6160 7164 6164 7196
rect 6196 7164 6200 7196
rect 6160 7116 6200 7164
rect 6160 7084 6164 7116
rect 6196 7084 6200 7116
rect 6160 7036 6200 7084
rect 6160 7004 6164 7036
rect 6196 7004 6200 7036
rect 6160 6956 6200 7004
rect 6160 6924 6164 6956
rect 6196 6924 6200 6956
rect 6160 6796 6200 6924
rect 6160 6764 6164 6796
rect 6196 6764 6200 6796
rect 6160 6716 6200 6764
rect 6160 6684 6164 6716
rect 6196 6684 6200 6716
rect 6160 6636 6200 6684
rect 6160 6604 6164 6636
rect 6196 6604 6200 6636
rect 6160 6556 6200 6604
rect 6160 6524 6164 6556
rect 6196 6524 6200 6556
rect 6160 6476 6200 6524
rect 6160 6444 6164 6476
rect 6196 6444 6200 6476
rect 6160 6316 6200 6444
rect 6160 6284 6164 6316
rect 6196 6284 6200 6316
rect 6160 6236 6200 6284
rect 6160 6204 6164 6236
rect 6196 6204 6200 6236
rect 6160 6156 6200 6204
rect 6160 6124 6164 6156
rect 6196 6124 6200 6156
rect 6160 5996 6200 6124
rect 6160 5964 6164 5996
rect 6196 5964 6200 5996
rect 6160 5836 6200 5964
rect 6160 5804 6164 5836
rect 6196 5804 6200 5836
rect 6160 5756 6200 5804
rect 6160 5724 6164 5756
rect 6196 5724 6200 5756
rect 6160 5676 6200 5724
rect 6160 5644 6164 5676
rect 6196 5644 6200 5676
rect 6160 5596 6200 5644
rect 6160 5564 6164 5596
rect 6196 5564 6200 5596
rect 6160 5516 6200 5564
rect 6160 5484 6164 5516
rect 6196 5484 6200 5516
rect 6160 5436 6200 5484
rect 6160 5404 6164 5436
rect 6196 5404 6200 5436
rect 6160 5356 6200 5404
rect 6160 5324 6164 5356
rect 6196 5324 6200 5356
rect 6160 5276 6200 5324
rect 6160 5244 6164 5276
rect 6196 5244 6200 5276
rect 6160 5196 6200 5244
rect 6160 5164 6164 5196
rect 6196 5164 6200 5196
rect 6160 5116 6200 5164
rect 6160 5084 6164 5116
rect 6196 5084 6200 5116
rect 6160 5036 6200 5084
rect 6160 5004 6164 5036
rect 6196 5004 6200 5036
rect 6160 4956 6200 5004
rect 6160 4924 6164 4956
rect 6196 4924 6200 4956
rect 6160 4876 6200 4924
rect 6160 4844 6164 4876
rect 6196 4844 6200 4876
rect 6160 4796 6200 4844
rect 6160 4764 6164 4796
rect 6196 4764 6200 4796
rect 6160 4716 6200 4764
rect 6160 4684 6164 4716
rect 6196 4684 6200 4716
rect 6160 4636 6200 4684
rect 6160 4604 6164 4636
rect 6196 4604 6200 4636
rect 6160 4556 6200 4604
rect 6160 4524 6164 4556
rect 6196 4524 6200 4556
rect 6160 4396 6200 4524
rect 6160 4364 6164 4396
rect 6196 4364 6200 4396
rect 6160 4316 6200 4364
rect 6160 4284 6164 4316
rect 6196 4284 6200 4316
rect 6160 4236 6200 4284
rect 6160 4204 6164 4236
rect 6196 4204 6200 4236
rect 6160 4156 6200 4204
rect 6160 4124 6164 4156
rect 6196 4124 6200 4156
rect 6160 4076 6200 4124
rect 6160 4044 6164 4076
rect 6196 4044 6200 4076
rect 6160 3916 6200 4044
rect 6160 3884 6164 3916
rect 6196 3884 6200 3916
rect 6160 3836 6200 3884
rect 6160 3804 6164 3836
rect 6196 3804 6200 3836
rect 6160 3756 6200 3804
rect 6160 3724 6164 3756
rect 6196 3724 6200 3756
rect 6160 3596 6200 3724
rect 6160 3564 6164 3596
rect 6196 3564 6200 3596
rect 6160 3436 6200 3564
rect 6160 3404 6164 3436
rect 6196 3404 6200 3436
rect 6160 3356 6200 3404
rect 6160 3324 6164 3356
rect 6196 3324 6200 3356
rect 6160 3276 6200 3324
rect 6160 3244 6164 3276
rect 6196 3244 6200 3276
rect 6160 3196 6200 3244
rect 6160 3164 6164 3196
rect 6196 3164 6200 3196
rect 6160 3116 6200 3164
rect 6160 3084 6164 3116
rect 6196 3084 6200 3116
rect 6160 3036 6200 3084
rect 6160 3004 6164 3036
rect 6196 3004 6200 3036
rect 6160 2956 6200 3004
rect 6160 2924 6164 2956
rect 6196 2924 6200 2956
rect 6160 2876 6200 2924
rect 6160 2844 6164 2876
rect 6196 2844 6200 2876
rect 6160 2796 6200 2844
rect 6160 2764 6164 2796
rect 6196 2764 6200 2796
rect 6160 2716 6200 2764
rect 6160 2684 6164 2716
rect 6196 2684 6200 2716
rect 6160 2636 6200 2684
rect 6160 2604 6164 2636
rect 6196 2604 6200 2636
rect 6160 2556 6200 2604
rect 6160 2524 6164 2556
rect 6196 2524 6200 2556
rect 6160 2476 6200 2524
rect 6160 2444 6164 2476
rect 6196 2444 6200 2476
rect 6160 2396 6200 2444
rect 6160 2364 6164 2396
rect 6196 2364 6200 2396
rect 6160 2316 6200 2364
rect 6160 2284 6164 2316
rect 6196 2284 6200 2316
rect 6160 2236 6200 2284
rect 6160 2204 6164 2236
rect 6196 2204 6200 2236
rect 6160 2156 6200 2204
rect 6160 2124 6164 2156
rect 6196 2124 6200 2156
rect 6160 2076 6200 2124
rect 6160 2044 6164 2076
rect 6196 2044 6200 2076
rect 6160 1996 6200 2044
rect 6160 1964 6164 1996
rect 6196 1964 6200 1996
rect 6160 1916 6200 1964
rect 6160 1884 6164 1916
rect 6196 1884 6200 1916
rect 6160 1836 6200 1884
rect 6160 1804 6164 1836
rect 6196 1804 6200 1836
rect 6160 1756 6200 1804
rect 6160 1724 6164 1756
rect 6196 1724 6200 1756
rect 6160 1676 6200 1724
rect 6160 1644 6164 1676
rect 6196 1644 6200 1676
rect 6160 1596 6200 1644
rect 6160 1564 6164 1596
rect 6196 1564 6200 1596
rect 6160 1516 6200 1564
rect 6160 1484 6164 1516
rect 6196 1484 6200 1516
rect 6160 1436 6200 1484
rect 6160 1404 6164 1436
rect 6196 1404 6200 1436
rect 6160 1356 6200 1404
rect 6160 1324 6164 1356
rect 6196 1324 6200 1356
rect 6160 1276 6200 1324
rect 6160 1244 6164 1276
rect 6196 1244 6200 1276
rect 6160 1196 6200 1244
rect 6160 1164 6164 1196
rect 6196 1164 6200 1196
rect 6160 1116 6200 1164
rect 6160 1084 6164 1116
rect 6196 1084 6200 1116
rect 6160 1036 6200 1084
rect 6160 1004 6164 1036
rect 6196 1004 6200 1036
rect 6160 956 6200 1004
rect 6160 924 6164 956
rect 6196 924 6200 956
rect 6160 876 6200 924
rect 6160 844 6164 876
rect 6196 844 6200 876
rect 6160 796 6200 844
rect 6160 764 6164 796
rect 6196 764 6200 796
rect 6160 716 6200 764
rect 6160 684 6164 716
rect 6196 684 6200 716
rect 6160 596 6200 684
rect 6160 564 6164 596
rect 6196 564 6200 596
rect 6160 516 6200 564
rect 6160 484 6164 516
rect 6196 484 6200 516
rect 6160 436 6200 484
rect 6160 404 6164 436
rect 6196 404 6200 436
rect 6160 356 6200 404
rect 6160 324 6164 356
rect 6196 324 6200 356
rect 6160 276 6200 324
rect 6160 244 6164 276
rect 6196 244 6200 276
rect 6160 196 6200 244
rect 6160 164 6164 196
rect 6196 164 6200 196
rect 6160 116 6200 164
rect 6160 84 6164 116
rect 6196 84 6200 116
rect 6160 36 6200 84
rect 6160 4 6164 36
rect 6196 4 6200 36
rect 6160 -40 6200 4
rect 6240 6875 6280 16640
rect 6240 6845 6245 6875
rect 6275 6845 6280 6875
rect 6240 4475 6280 6845
rect 6240 4445 6245 4475
rect 6275 4445 6280 4475
rect 6240 -40 6280 4445
rect 6320 16596 6360 16644
rect 6480 16836 6520 16840
rect 6480 16644 6484 16836
rect 6516 16644 6520 16836
rect 6320 16564 6324 16596
rect 6356 16564 6360 16596
rect 6320 16516 6360 16564
rect 6320 16484 6324 16516
rect 6356 16484 6360 16516
rect 6320 16436 6360 16484
rect 6320 16404 6324 16436
rect 6356 16404 6360 16436
rect 6320 16356 6360 16404
rect 6320 16324 6324 16356
rect 6356 16324 6360 16356
rect 6320 16276 6360 16324
rect 6320 16244 6324 16276
rect 6356 16244 6360 16276
rect 6320 16196 6360 16244
rect 6320 16164 6324 16196
rect 6356 16164 6360 16196
rect 6320 16116 6360 16164
rect 6320 16084 6324 16116
rect 6356 16084 6360 16116
rect 6320 16036 6360 16084
rect 6320 16004 6324 16036
rect 6356 16004 6360 16036
rect 6320 15956 6360 16004
rect 6320 15924 6324 15956
rect 6356 15924 6360 15956
rect 6320 15436 6360 15924
rect 6320 15404 6324 15436
rect 6356 15404 6360 15436
rect 6320 15356 6360 15404
rect 6320 15324 6324 15356
rect 6356 15324 6360 15356
rect 6320 15276 6360 15324
rect 6320 15244 6324 15276
rect 6356 15244 6360 15276
rect 6320 15196 6360 15244
rect 6320 15164 6324 15196
rect 6356 15164 6360 15196
rect 6320 15116 6360 15164
rect 6320 15084 6324 15116
rect 6356 15084 6360 15116
rect 6320 15036 6360 15084
rect 6320 15004 6324 15036
rect 6356 15004 6360 15036
rect 6320 14956 6360 15004
rect 6320 14924 6324 14956
rect 6356 14924 6360 14956
rect 6320 14876 6360 14924
rect 6320 14844 6324 14876
rect 6356 14844 6360 14876
rect 6320 14796 6360 14844
rect 6320 14764 6324 14796
rect 6356 14764 6360 14796
rect 6320 14716 6360 14764
rect 6320 14684 6324 14716
rect 6356 14684 6360 14716
rect 6320 14636 6360 14684
rect 6320 14604 6324 14636
rect 6356 14604 6360 14636
rect 6320 14556 6360 14604
rect 6320 14524 6324 14556
rect 6356 14524 6360 14556
rect 6320 14476 6360 14524
rect 6320 14444 6324 14476
rect 6356 14444 6360 14476
rect 6320 13996 6360 14444
rect 6320 13964 6324 13996
rect 6356 13964 6360 13996
rect 6320 13876 6360 13964
rect 6320 13844 6324 13876
rect 6356 13844 6360 13876
rect 6320 13796 6360 13844
rect 6320 13764 6324 13796
rect 6356 13764 6360 13796
rect 6320 13716 6360 13764
rect 6320 13684 6324 13716
rect 6356 13684 6360 13716
rect 6320 13636 6360 13684
rect 6320 13604 6324 13636
rect 6356 13604 6360 13636
rect 6320 13556 6360 13604
rect 6320 13524 6324 13556
rect 6356 13524 6360 13556
rect 6320 13476 6360 13524
rect 6320 13444 6324 13476
rect 6356 13444 6360 13476
rect 6320 13396 6360 13444
rect 6320 13364 6324 13396
rect 6356 13364 6360 13396
rect 6320 13316 6360 13364
rect 6320 13284 6324 13316
rect 6356 13284 6360 13316
rect 6320 13236 6360 13284
rect 6320 13204 6324 13236
rect 6356 13204 6360 13236
rect 6320 13156 6360 13204
rect 6320 13124 6324 13156
rect 6356 13124 6360 13156
rect 6320 13076 6360 13124
rect 6320 13044 6324 13076
rect 6356 13044 6360 13076
rect 6320 12996 6360 13044
rect 6320 12964 6324 12996
rect 6356 12964 6360 12996
rect 6320 12516 6360 12964
rect 6320 12484 6324 12516
rect 6356 12484 6360 12516
rect 6320 12436 6360 12484
rect 6320 12404 6324 12436
rect 6356 12404 6360 12436
rect 6320 12316 6360 12404
rect 6320 12284 6324 12316
rect 6356 12284 6360 12316
rect 6320 12236 6360 12284
rect 6320 12204 6324 12236
rect 6356 12204 6360 12236
rect 6320 12156 6360 12204
rect 6320 12124 6324 12156
rect 6356 12124 6360 12156
rect 6320 12076 6360 12124
rect 6320 12044 6324 12076
rect 6356 12044 6360 12076
rect 6320 11996 6360 12044
rect 6320 11964 6324 11996
rect 6356 11964 6360 11996
rect 6320 11916 6360 11964
rect 6320 11884 6324 11916
rect 6356 11884 6360 11916
rect 6320 11836 6360 11884
rect 6320 11804 6324 11836
rect 6356 11804 6360 11836
rect 6320 11756 6360 11804
rect 6320 11724 6324 11756
rect 6356 11724 6360 11756
rect 6320 11676 6360 11724
rect 6320 11644 6324 11676
rect 6356 11644 6360 11676
rect 6320 11596 6360 11644
rect 6320 11564 6324 11596
rect 6356 11564 6360 11596
rect 6320 11516 6360 11564
rect 6320 11484 6324 11516
rect 6356 11484 6360 11516
rect 6320 11436 6360 11484
rect 6320 11404 6324 11436
rect 6356 11404 6360 11436
rect 6320 11356 6360 11404
rect 6320 11324 6324 11356
rect 6356 11324 6360 11356
rect 6320 11196 6360 11324
rect 6320 11164 6324 11196
rect 6356 11164 6360 11196
rect 6320 11116 6360 11164
rect 6320 11084 6324 11116
rect 6356 11084 6360 11116
rect 6320 11036 6360 11084
rect 6320 11004 6324 11036
rect 6356 11004 6360 11036
rect 6320 10876 6360 11004
rect 6320 10844 6324 10876
rect 6356 10844 6360 10876
rect 6320 10716 6360 10844
rect 6320 10684 6324 10716
rect 6356 10684 6360 10716
rect 6320 10636 6360 10684
rect 6320 10604 6324 10636
rect 6356 10604 6360 10636
rect 6320 10476 6360 10604
rect 6320 10444 6324 10476
rect 6356 10444 6360 10476
rect 6320 10316 6360 10444
rect 6320 10284 6324 10316
rect 6356 10284 6360 10316
rect 6320 10236 6360 10284
rect 6320 10204 6324 10236
rect 6356 10204 6360 10236
rect 6320 10156 6360 10204
rect 6320 10124 6324 10156
rect 6356 10124 6360 10156
rect 6320 10076 6360 10124
rect 6320 10044 6324 10076
rect 6356 10044 6360 10076
rect 6320 9996 6360 10044
rect 6320 9964 6324 9996
rect 6356 9964 6360 9996
rect 6320 9916 6360 9964
rect 6320 9884 6324 9916
rect 6356 9884 6360 9916
rect 6320 9836 6360 9884
rect 6320 9804 6324 9836
rect 6356 9804 6360 9836
rect 6320 9756 6360 9804
rect 6320 9724 6324 9756
rect 6356 9724 6360 9756
rect 6320 9676 6360 9724
rect 6320 9644 6324 9676
rect 6356 9644 6360 9676
rect 6320 9596 6360 9644
rect 6320 9564 6324 9596
rect 6356 9564 6360 9596
rect 6320 9516 6360 9564
rect 6320 9484 6324 9516
rect 6356 9484 6360 9516
rect 6320 9436 6360 9484
rect 6320 9404 6324 9436
rect 6356 9404 6360 9436
rect 6320 9356 6360 9404
rect 6320 9324 6324 9356
rect 6356 9324 6360 9356
rect 6320 9276 6360 9324
rect 6320 9244 6324 9276
rect 6356 9244 6360 9276
rect 6320 9116 6360 9244
rect 6320 9084 6324 9116
rect 6356 9084 6360 9116
rect 6320 9036 6360 9084
rect 6320 9004 6324 9036
rect 6356 9004 6360 9036
rect 6320 8956 6360 9004
rect 6320 8924 6324 8956
rect 6356 8924 6360 8956
rect 6320 8636 6360 8924
rect 6320 8604 6324 8636
rect 6356 8604 6360 8636
rect 6320 8556 6360 8604
rect 6320 8524 6324 8556
rect 6356 8524 6360 8556
rect 6320 8396 6360 8524
rect 6320 8364 6324 8396
rect 6356 8364 6360 8396
rect 6320 8236 6360 8364
rect 6320 8204 6324 8236
rect 6356 8204 6360 8236
rect 6320 8156 6360 8204
rect 6320 8124 6324 8156
rect 6356 8124 6360 8156
rect 6320 8076 6360 8124
rect 6320 8044 6324 8076
rect 6356 8044 6360 8076
rect 6320 7996 6360 8044
rect 6320 7964 6324 7996
rect 6356 7964 6360 7996
rect 6320 7916 6360 7964
rect 6320 7884 6324 7916
rect 6356 7884 6360 7916
rect 6320 7836 6360 7884
rect 6320 7804 6324 7836
rect 6356 7804 6360 7836
rect 6320 7756 6360 7804
rect 6320 7724 6324 7756
rect 6356 7724 6360 7756
rect 6320 7676 6360 7724
rect 6320 7644 6324 7676
rect 6356 7644 6360 7676
rect 6320 7596 6360 7644
rect 6320 7564 6324 7596
rect 6356 7564 6360 7596
rect 6320 7516 6360 7564
rect 6320 7484 6324 7516
rect 6356 7484 6360 7516
rect 6320 7436 6360 7484
rect 6320 7404 6324 7436
rect 6356 7404 6360 7436
rect 6320 7356 6360 7404
rect 6320 7324 6324 7356
rect 6356 7324 6360 7356
rect 6320 7276 6360 7324
rect 6320 7244 6324 7276
rect 6356 7244 6360 7276
rect 6320 7196 6360 7244
rect 6320 7164 6324 7196
rect 6356 7164 6360 7196
rect 6320 7116 6360 7164
rect 6320 7084 6324 7116
rect 6356 7084 6360 7116
rect 6320 7036 6360 7084
rect 6320 7004 6324 7036
rect 6356 7004 6360 7036
rect 6320 6956 6360 7004
rect 6320 6924 6324 6956
rect 6356 6924 6360 6956
rect 6320 6876 6360 6924
rect 6320 6844 6324 6876
rect 6356 6844 6360 6876
rect 6320 6796 6360 6844
rect 6320 6764 6324 6796
rect 6356 6764 6360 6796
rect 6320 6716 6360 6764
rect 6320 6684 6324 6716
rect 6356 6684 6360 6716
rect 6320 6636 6360 6684
rect 6320 6604 6324 6636
rect 6356 6604 6360 6636
rect 6320 6556 6360 6604
rect 6320 6524 6324 6556
rect 6356 6524 6360 6556
rect 6320 6476 6360 6524
rect 6320 6444 6324 6476
rect 6356 6444 6360 6476
rect 6320 6316 6360 6444
rect 6320 6284 6324 6316
rect 6356 6284 6360 6316
rect 6320 6236 6360 6284
rect 6320 6204 6324 6236
rect 6356 6204 6360 6236
rect 6320 6156 6360 6204
rect 6320 6124 6324 6156
rect 6356 6124 6360 6156
rect 6320 5996 6360 6124
rect 6320 5964 6324 5996
rect 6356 5964 6360 5996
rect 6320 5836 6360 5964
rect 6320 5804 6324 5836
rect 6356 5804 6360 5836
rect 6320 5756 6360 5804
rect 6320 5724 6324 5756
rect 6356 5724 6360 5756
rect 6320 5676 6360 5724
rect 6320 5644 6324 5676
rect 6356 5644 6360 5676
rect 6320 5596 6360 5644
rect 6320 5564 6324 5596
rect 6356 5564 6360 5596
rect 6320 5516 6360 5564
rect 6320 5484 6324 5516
rect 6356 5484 6360 5516
rect 6320 5436 6360 5484
rect 6320 5404 6324 5436
rect 6356 5404 6360 5436
rect 6320 5356 6360 5404
rect 6320 5324 6324 5356
rect 6356 5324 6360 5356
rect 6320 5276 6360 5324
rect 6320 5244 6324 5276
rect 6356 5244 6360 5276
rect 6320 5196 6360 5244
rect 6320 5164 6324 5196
rect 6356 5164 6360 5196
rect 6320 5116 6360 5164
rect 6320 5084 6324 5116
rect 6356 5084 6360 5116
rect 6320 5036 6360 5084
rect 6320 5004 6324 5036
rect 6356 5004 6360 5036
rect 6320 4956 6360 5004
rect 6320 4924 6324 4956
rect 6356 4924 6360 4956
rect 6320 4876 6360 4924
rect 6320 4844 6324 4876
rect 6356 4844 6360 4876
rect 6320 4796 6360 4844
rect 6320 4764 6324 4796
rect 6356 4764 6360 4796
rect 6320 4716 6360 4764
rect 6320 4684 6324 4716
rect 6356 4684 6360 4716
rect 6320 4636 6360 4684
rect 6320 4604 6324 4636
rect 6356 4604 6360 4636
rect 6320 4556 6360 4604
rect 6320 4524 6324 4556
rect 6356 4524 6360 4556
rect 6320 4476 6360 4524
rect 6320 4444 6324 4476
rect 6356 4444 6360 4476
rect 6320 4396 6360 4444
rect 6320 4364 6324 4396
rect 6356 4364 6360 4396
rect 6320 4316 6360 4364
rect 6320 4284 6324 4316
rect 6356 4284 6360 4316
rect 6320 4236 6360 4284
rect 6320 4204 6324 4236
rect 6356 4204 6360 4236
rect 6320 4156 6360 4204
rect 6320 4124 6324 4156
rect 6356 4124 6360 4156
rect 6320 4076 6360 4124
rect 6320 4044 6324 4076
rect 6356 4044 6360 4076
rect 6320 3916 6360 4044
rect 6320 3884 6324 3916
rect 6356 3884 6360 3916
rect 6320 3836 6360 3884
rect 6320 3804 6324 3836
rect 6356 3804 6360 3836
rect 6320 3756 6360 3804
rect 6320 3724 6324 3756
rect 6356 3724 6360 3756
rect 6320 3596 6360 3724
rect 6320 3564 6324 3596
rect 6356 3564 6360 3596
rect 6320 3436 6360 3564
rect 6320 3404 6324 3436
rect 6356 3404 6360 3436
rect 6320 3356 6360 3404
rect 6320 3324 6324 3356
rect 6356 3324 6360 3356
rect 6320 3276 6360 3324
rect 6320 3244 6324 3276
rect 6356 3244 6360 3276
rect 6320 3196 6360 3244
rect 6320 3164 6324 3196
rect 6356 3164 6360 3196
rect 6320 3116 6360 3164
rect 6320 3084 6324 3116
rect 6356 3084 6360 3116
rect 6320 3036 6360 3084
rect 6320 3004 6324 3036
rect 6356 3004 6360 3036
rect 6320 2956 6360 3004
rect 6320 2924 6324 2956
rect 6356 2924 6360 2956
rect 6320 2876 6360 2924
rect 6320 2844 6324 2876
rect 6356 2844 6360 2876
rect 6320 2796 6360 2844
rect 6320 2764 6324 2796
rect 6356 2764 6360 2796
rect 6320 2716 6360 2764
rect 6320 2684 6324 2716
rect 6356 2684 6360 2716
rect 6320 2636 6360 2684
rect 6320 2604 6324 2636
rect 6356 2604 6360 2636
rect 6320 2556 6360 2604
rect 6320 2524 6324 2556
rect 6356 2524 6360 2556
rect 6320 2476 6360 2524
rect 6320 2444 6324 2476
rect 6356 2444 6360 2476
rect 6320 2396 6360 2444
rect 6320 2364 6324 2396
rect 6356 2364 6360 2396
rect 6320 2316 6360 2364
rect 6320 2284 6324 2316
rect 6356 2284 6360 2316
rect 6320 2236 6360 2284
rect 6320 2204 6324 2236
rect 6356 2204 6360 2236
rect 6320 2156 6360 2204
rect 6320 2124 6324 2156
rect 6356 2124 6360 2156
rect 6320 2076 6360 2124
rect 6320 2044 6324 2076
rect 6356 2044 6360 2076
rect 6320 1996 6360 2044
rect 6320 1964 6324 1996
rect 6356 1964 6360 1996
rect 6320 1916 6360 1964
rect 6320 1884 6324 1916
rect 6356 1884 6360 1916
rect 6320 1836 6360 1884
rect 6320 1804 6324 1836
rect 6356 1804 6360 1836
rect 6320 1756 6360 1804
rect 6320 1724 6324 1756
rect 6356 1724 6360 1756
rect 6320 1676 6360 1724
rect 6320 1644 6324 1676
rect 6356 1644 6360 1676
rect 6320 1596 6360 1644
rect 6320 1564 6324 1596
rect 6356 1564 6360 1596
rect 6320 1516 6360 1564
rect 6320 1484 6324 1516
rect 6356 1484 6360 1516
rect 6320 1436 6360 1484
rect 6320 1404 6324 1436
rect 6356 1404 6360 1436
rect 6320 1356 6360 1404
rect 6320 1324 6324 1356
rect 6356 1324 6360 1356
rect 6320 1276 6360 1324
rect 6320 1244 6324 1276
rect 6356 1244 6360 1276
rect 6320 1196 6360 1244
rect 6320 1164 6324 1196
rect 6356 1164 6360 1196
rect 6320 1116 6360 1164
rect 6320 1084 6324 1116
rect 6356 1084 6360 1116
rect 6320 1036 6360 1084
rect 6320 1004 6324 1036
rect 6356 1004 6360 1036
rect 6320 956 6360 1004
rect 6320 924 6324 956
rect 6356 924 6360 956
rect 6320 876 6360 924
rect 6320 844 6324 876
rect 6356 844 6360 876
rect 6320 796 6360 844
rect 6320 764 6324 796
rect 6356 764 6360 796
rect 6320 716 6360 764
rect 6320 684 6324 716
rect 6356 684 6360 716
rect 6320 596 6360 684
rect 6320 564 6324 596
rect 6356 564 6360 596
rect 6320 516 6360 564
rect 6320 484 6324 516
rect 6356 484 6360 516
rect 6320 436 6360 484
rect 6320 404 6324 436
rect 6356 404 6360 436
rect 6320 356 6360 404
rect 6320 324 6324 356
rect 6356 324 6360 356
rect 6320 276 6360 324
rect 6320 244 6324 276
rect 6356 244 6360 276
rect 6320 196 6360 244
rect 6320 164 6324 196
rect 6356 164 6360 196
rect 6320 116 6360 164
rect 6320 84 6324 116
rect 6356 84 6360 116
rect 6320 36 6360 84
rect 6320 4 6324 36
rect 6356 4 6360 36
rect 6320 -40 6360 4
rect 6400 3995 6440 16640
rect 6400 3965 6405 3995
rect 6435 3965 6440 3995
rect 6400 -40 6440 3965
rect 6480 16596 6520 16644
rect 6640 16836 6680 16840
rect 6640 16644 6644 16836
rect 6676 16644 6680 16836
rect 6480 16564 6484 16596
rect 6516 16564 6520 16596
rect 6480 16516 6520 16564
rect 6480 16484 6484 16516
rect 6516 16484 6520 16516
rect 6480 16436 6520 16484
rect 6480 16404 6484 16436
rect 6516 16404 6520 16436
rect 6480 16356 6520 16404
rect 6480 16324 6484 16356
rect 6516 16324 6520 16356
rect 6480 16276 6520 16324
rect 6480 16244 6484 16276
rect 6516 16244 6520 16276
rect 6480 16196 6520 16244
rect 6480 16164 6484 16196
rect 6516 16164 6520 16196
rect 6480 16116 6520 16164
rect 6480 16084 6484 16116
rect 6516 16084 6520 16116
rect 6480 16036 6520 16084
rect 6480 16004 6484 16036
rect 6516 16004 6520 16036
rect 6480 15956 6520 16004
rect 6480 15924 6484 15956
rect 6516 15924 6520 15956
rect 6480 15436 6520 15924
rect 6480 15404 6484 15436
rect 6516 15404 6520 15436
rect 6480 15356 6520 15404
rect 6480 15324 6484 15356
rect 6516 15324 6520 15356
rect 6480 15276 6520 15324
rect 6480 15244 6484 15276
rect 6516 15244 6520 15276
rect 6480 15196 6520 15244
rect 6480 15164 6484 15196
rect 6516 15164 6520 15196
rect 6480 15116 6520 15164
rect 6480 15084 6484 15116
rect 6516 15084 6520 15116
rect 6480 15036 6520 15084
rect 6480 15004 6484 15036
rect 6516 15004 6520 15036
rect 6480 14956 6520 15004
rect 6480 14924 6484 14956
rect 6516 14924 6520 14956
rect 6480 14876 6520 14924
rect 6480 14844 6484 14876
rect 6516 14844 6520 14876
rect 6480 14796 6520 14844
rect 6480 14764 6484 14796
rect 6516 14764 6520 14796
rect 6480 14716 6520 14764
rect 6480 14684 6484 14716
rect 6516 14684 6520 14716
rect 6480 14636 6520 14684
rect 6480 14604 6484 14636
rect 6516 14604 6520 14636
rect 6480 14556 6520 14604
rect 6480 14524 6484 14556
rect 6516 14524 6520 14556
rect 6480 14476 6520 14524
rect 6480 14444 6484 14476
rect 6516 14444 6520 14476
rect 6480 13996 6520 14444
rect 6480 13964 6484 13996
rect 6516 13964 6520 13996
rect 6480 13876 6520 13964
rect 6480 13844 6484 13876
rect 6516 13844 6520 13876
rect 6480 13796 6520 13844
rect 6480 13764 6484 13796
rect 6516 13764 6520 13796
rect 6480 13716 6520 13764
rect 6480 13684 6484 13716
rect 6516 13684 6520 13716
rect 6480 13636 6520 13684
rect 6480 13604 6484 13636
rect 6516 13604 6520 13636
rect 6480 13556 6520 13604
rect 6480 13524 6484 13556
rect 6516 13524 6520 13556
rect 6480 13476 6520 13524
rect 6480 13444 6484 13476
rect 6516 13444 6520 13476
rect 6480 13396 6520 13444
rect 6480 13364 6484 13396
rect 6516 13364 6520 13396
rect 6480 13316 6520 13364
rect 6480 13284 6484 13316
rect 6516 13284 6520 13316
rect 6480 13236 6520 13284
rect 6480 13204 6484 13236
rect 6516 13204 6520 13236
rect 6480 13156 6520 13204
rect 6480 13124 6484 13156
rect 6516 13124 6520 13156
rect 6480 13076 6520 13124
rect 6480 13044 6484 13076
rect 6516 13044 6520 13076
rect 6480 12996 6520 13044
rect 6480 12964 6484 12996
rect 6516 12964 6520 12996
rect 6480 12516 6520 12964
rect 6480 12484 6484 12516
rect 6516 12484 6520 12516
rect 6480 12436 6520 12484
rect 6480 12404 6484 12436
rect 6516 12404 6520 12436
rect 6480 12316 6520 12404
rect 6480 12284 6484 12316
rect 6516 12284 6520 12316
rect 6480 12236 6520 12284
rect 6480 12204 6484 12236
rect 6516 12204 6520 12236
rect 6480 12156 6520 12204
rect 6480 12124 6484 12156
rect 6516 12124 6520 12156
rect 6480 12076 6520 12124
rect 6480 12044 6484 12076
rect 6516 12044 6520 12076
rect 6480 11996 6520 12044
rect 6480 11964 6484 11996
rect 6516 11964 6520 11996
rect 6480 11916 6520 11964
rect 6480 11884 6484 11916
rect 6516 11884 6520 11916
rect 6480 11836 6520 11884
rect 6480 11804 6484 11836
rect 6516 11804 6520 11836
rect 6480 11756 6520 11804
rect 6480 11724 6484 11756
rect 6516 11724 6520 11756
rect 6480 11676 6520 11724
rect 6480 11644 6484 11676
rect 6516 11644 6520 11676
rect 6480 11596 6520 11644
rect 6480 11564 6484 11596
rect 6516 11564 6520 11596
rect 6480 11516 6520 11564
rect 6480 11484 6484 11516
rect 6516 11484 6520 11516
rect 6480 11436 6520 11484
rect 6480 11404 6484 11436
rect 6516 11404 6520 11436
rect 6480 11356 6520 11404
rect 6480 11324 6484 11356
rect 6516 11324 6520 11356
rect 6480 11196 6520 11324
rect 6480 11164 6484 11196
rect 6516 11164 6520 11196
rect 6480 11116 6520 11164
rect 6480 11084 6484 11116
rect 6516 11084 6520 11116
rect 6480 11036 6520 11084
rect 6480 11004 6484 11036
rect 6516 11004 6520 11036
rect 6480 10876 6520 11004
rect 6480 10844 6484 10876
rect 6516 10844 6520 10876
rect 6480 10716 6520 10844
rect 6480 10684 6484 10716
rect 6516 10684 6520 10716
rect 6480 10636 6520 10684
rect 6480 10604 6484 10636
rect 6516 10604 6520 10636
rect 6480 10476 6520 10604
rect 6480 10444 6484 10476
rect 6516 10444 6520 10476
rect 6480 10316 6520 10444
rect 6480 10284 6484 10316
rect 6516 10284 6520 10316
rect 6480 10236 6520 10284
rect 6480 10204 6484 10236
rect 6516 10204 6520 10236
rect 6480 10156 6520 10204
rect 6480 10124 6484 10156
rect 6516 10124 6520 10156
rect 6480 10076 6520 10124
rect 6480 10044 6484 10076
rect 6516 10044 6520 10076
rect 6480 9996 6520 10044
rect 6480 9964 6484 9996
rect 6516 9964 6520 9996
rect 6480 9916 6520 9964
rect 6480 9884 6484 9916
rect 6516 9884 6520 9916
rect 6480 9836 6520 9884
rect 6480 9804 6484 9836
rect 6516 9804 6520 9836
rect 6480 9756 6520 9804
rect 6480 9724 6484 9756
rect 6516 9724 6520 9756
rect 6480 9676 6520 9724
rect 6480 9644 6484 9676
rect 6516 9644 6520 9676
rect 6480 9596 6520 9644
rect 6480 9564 6484 9596
rect 6516 9564 6520 9596
rect 6480 9516 6520 9564
rect 6480 9484 6484 9516
rect 6516 9484 6520 9516
rect 6480 9436 6520 9484
rect 6480 9404 6484 9436
rect 6516 9404 6520 9436
rect 6480 9356 6520 9404
rect 6480 9324 6484 9356
rect 6516 9324 6520 9356
rect 6480 9276 6520 9324
rect 6480 9244 6484 9276
rect 6516 9244 6520 9276
rect 6480 9116 6520 9244
rect 6480 9084 6484 9116
rect 6516 9084 6520 9116
rect 6480 9036 6520 9084
rect 6480 9004 6484 9036
rect 6516 9004 6520 9036
rect 6480 8956 6520 9004
rect 6480 8924 6484 8956
rect 6516 8924 6520 8956
rect 6480 8636 6520 8924
rect 6480 8604 6484 8636
rect 6516 8604 6520 8636
rect 6480 8556 6520 8604
rect 6480 8524 6484 8556
rect 6516 8524 6520 8556
rect 6480 8396 6520 8524
rect 6480 8364 6484 8396
rect 6516 8364 6520 8396
rect 6480 8236 6520 8364
rect 6480 8204 6484 8236
rect 6516 8204 6520 8236
rect 6480 8156 6520 8204
rect 6480 8124 6484 8156
rect 6516 8124 6520 8156
rect 6480 8076 6520 8124
rect 6480 8044 6484 8076
rect 6516 8044 6520 8076
rect 6480 7996 6520 8044
rect 6480 7964 6484 7996
rect 6516 7964 6520 7996
rect 6480 7916 6520 7964
rect 6480 7884 6484 7916
rect 6516 7884 6520 7916
rect 6480 7836 6520 7884
rect 6480 7804 6484 7836
rect 6516 7804 6520 7836
rect 6480 7756 6520 7804
rect 6480 7724 6484 7756
rect 6516 7724 6520 7756
rect 6480 7676 6520 7724
rect 6480 7644 6484 7676
rect 6516 7644 6520 7676
rect 6480 7596 6520 7644
rect 6480 7564 6484 7596
rect 6516 7564 6520 7596
rect 6480 7516 6520 7564
rect 6480 7484 6484 7516
rect 6516 7484 6520 7516
rect 6480 7436 6520 7484
rect 6480 7404 6484 7436
rect 6516 7404 6520 7436
rect 6480 7356 6520 7404
rect 6480 7324 6484 7356
rect 6516 7324 6520 7356
rect 6480 7276 6520 7324
rect 6480 7244 6484 7276
rect 6516 7244 6520 7276
rect 6480 7196 6520 7244
rect 6480 7164 6484 7196
rect 6516 7164 6520 7196
rect 6480 7116 6520 7164
rect 6480 7084 6484 7116
rect 6516 7084 6520 7116
rect 6480 7036 6520 7084
rect 6480 7004 6484 7036
rect 6516 7004 6520 7036
rect 6480 6956 6520 7004
rect 6480 6924 6484 6956
rect 6516 6924 6520 6956
rect 6480 6876 6520 6924
rect 6480 6844 6484 6876
rect 6516 6844 6520 6876
rect 6480 6796 6520 6844
rect 6480 6764 6484 6796
rect 6516 6764 6520 6796
rect 6480 6716 6520 6764
rect 6480 6684 6484 6716
rect 6516 6684 6520 6716
rect 6480 6636 6520 6684
rect 6480 6604 6484 6636
rect 6516 6604 6520 6636
rect 6480 6556 6520 6604
rect 6480 6524 6484 6556
rect 6516 6524 6520 6556
rect 6480 6476 6520 6524
rect 6480 6444 6484 6476
rect 6516 6444 6520 6476
rect 6480 6316 6520 6444
rect 6480 6284 6484 6316
rect 6516 6284 6520 6316
rect 6480 6236 6520 6284
rect 6480 6204 6484 6236
rect 6516 6204 6520 6236
rect 6480 6156 6520 6204
rect 6480 6124 6484 6156
rect 6516 6124 6520 6156
rect 6480 5996 6520 6124
rect 6480 5964 6484 5996
rect 6516 5964 6520 5996
rect 6480 5836 6520 5964
rect 6480 5804 6484 5836
rect 6516 5804 6520 5836
rect 6480 5756 6520 5804
rect 6480 5724 6484 5756
rect 6516 5724 6520 5756
rect 6480 5676 6520 5724
rect 6480 5644 6484 5676
rect 6516 5644 6520 5676
rect 6480 5596 6520 5644
rect 6480 5564 6484 5596
rect 6516 5564 6520 5596
rect 6480 5516 6520 5564
rect 6480 5484 6484 5516
rect 6516 5484 6520 5516
rect 6480 5436 6520 5484
rect 6480 5404 6484 5436
rect 6516 5404 6520 5436
rect 6480 5356 6520 5404
rect 6480 5324 6484 5356
rect 6516 5324 6520 5356
rect 6480 5276 6520 5324
rect 6480 5244 6484 5276
rect 6516 5244 6520 5276
rect 6480 5196 6520 5244
rect 6480 5164 6484 5196
rect 6516 5164 6520 5196
rect 6480 5116 6520 5164
rect 6480 5084 6484 5116
rect 6516 5084 6520 5116
rect 6480 5036 6520 5084
rect 6480 5004 6484 5036
rect 6516 5004 6520 5036
rect 6480 4956 6520 5004
rect 6480 4924 6484 4956
rect 6516 4924 6520 4956
rect 6480 4876 6520 4924
rect 6480 4844 6484 4876
rect 6516 4844 6520 4876
rect 6480 4796 6520 4844
rect 6480 4764 6484 4796
rect 6516 4764 6520 4796
rect 6480 4716 6520 4764
rect 6480 4684 6484 4716
rect 6516 4684 6520 4716
rect 6480 4636 6520 4684
rect 6480 4604 6484 4636
rect 6516 4604 6520 4636
rect 6480 4556 6520 4604
rect 6480 4524 6484 4556
rect 6516 4524 6520 4556
rect 6480 4476 6520 4524
rect 6480 4444 6484 4476
rect 6516 4444 6520 4476
rect 6480 4396 6520 4444
rect 6480 4364 6484 4396
rect 6516 4364 6520 4396
rect 6480 4316 6520 4364
rect 6480 4284 6484 4316
rect 6516 4284 6520 4316
rect 6480 4236 6520 4284
rect 6480 4204 6484 4236
rect 6516 4204 6520 4236
rect 6480 4156 6520 4204
rect 6480 4124 6484 4156
rect 6516 4124 6520 4156
rect 6480 4076 6520 4124
rect 6480 4044 6484 4076
rect 6516 4044 6520 4076
rect 6480 3996 6520 4044
rect 6480 3964 6484 3996
rect 6516 3964 6520 3996
rect 6480 3916 6520 3964
rect 6480 3884 6484 3916
rect 6516 3884 6520 3916
rect 6480 3836 6520 3884
rect 6480 3804 6484 3836
rect 6516 3804 6520 3836
rect 6480 3756 6520 3804
rect 6480 3724 6484 3756
rect 6516 3724 6520 3756
rect 6480 3596 6520 3724
rect 6480 3564 6484 3596
rect 6516 3564 6520 3596
rect 6480 3436 6520 3564
rect 6480 3404 6484 3436
rect 6516 3404 6520 3436
rect 6480 3356 6520 3404
rect 6480 3324 6484 3356
rect 6516 3324 6520 3356
rect 6480 3276 6520 3324
rect 6480 3244 6484 3276
rect 6516 3244 6520 3276
rect 6480 3196 6520 3244
rect 6480 3164 6484 3196
rect 6516 3164 6520 3196
rect 6480 3116 6520 3164
rect 6480 3084 6484 3116
rect 6516 3084 6520 3116
rect 6480 3036 6520 3084
rect 6480 3004 6484 3036
rect 6516 3004 6520 3036
rect 6480 2956 6520 3004
rect 6480 2924 6484 2956
rect 6516 2924 6520 2956
rect 6480 2876 6520 2924
rect 6480 2844 6484 2876
rect 6516 2844 6520 2876
rect 6480 2796 6520 2844
rect 6480 2764 6484 2796
rect 6516 2764 6520 2796
rect 6480 2716 6520 2764
rect 6480 2684 6484 2716
rect 6516 2684 6520 2716
rect 6480 2636 6520 2684
rect 6480 2604 6484 2636
rect 6516 2604 6520 2636
rect 6480 2556 6520 2604
rect 6480 2524 6484 2556
rect 6516 2524 6520 2556
rect 6480 2476 6520 2524
rect 6480 2444 6484 2476
rect 6516 2444 6520 2476
rect 6480 2396 6520 2444
rect 6480 2364 6484 2396
rect 6516 2364 6520 2396
rect 6480 2316 6520 2364
rect 6480 2284 6484 2316
rect 6516 2284 6520 2316
rect 6480 2236 6520 2284
rect 6480 2204 6484 2236
rect 6516 2204 6520 2236
rect 6480 2156 6520 2204
rect 6480 2124 6484 2156
rect 6516 2124 6520 2156
rect 6480 2076 6520 2124
rect 6480 2044 6484 2076
rect 6516 2044 6520 2076
rect 6480 1996 6520 2044
rect 6480 1964 6484 1996
rect 6516 1964 6520 1996
rect 6480 1916 6520 1964
rect 6480 1884 6484 1916
rect 6516 1884 6520 1916
rect 6480 1836 6520 1884
rect 6480 1804 6484 1836
rect 6516 1804 6520 1836
rect 6480 1756 6520 1804
rect 6480 1724 6484 1756
rect 6516 1724 6520 1756
rect 6480 1676 6520 1724
rect 6480 1644 6484 1676
rect 6516 1644 6520 1676
rect 6480 1596 6520 1644
rect 6480 1564 6484 1596
rect 6516 1564 6520 1596
rect 6480 1516 6520 1564
rect 6480 1484 6484 1516
rect 6516 1484 6520 1516
rect 6480 1436 6520 1484
rect 6480 1404 6484 1436
rect 6516 1404 6520 1436
rect 6480 1356 6520 1404
rect 6480 1324 6484 1356
rect 6516 1324 6520 1356
rect 6480 1276 6520 1324
rect 6480 1244 6484 1276
rect 6516 1244 6520 1276
rect 6480 1196 6520 1244
rect 6480 1164 6484 1196
rect 6516 1164 6520 1196
rect 6480 1116 6520 1164
rect 6480 1084 6484 1116
rect 6516 1084 6520 1116
rect 6480 1036 6520 1084
rect 6480 1004 6484 1036
rect 6516 1004 6520 1036
rect 6480 956 6520 1004
rect 6480 924 6484 956
rect 6516 924 6520 956
rect 6480 876 6520 924
rect 6480 844 6484 876
rect 6516 844 6520 876
rect 6480 796 6520 844
rect 6480 764 6484 796
rect 6516 764 6520 796
rect 6480 716 6520 764
rect 6480 684 6484 716
rect 6516 684 6520 716
rect 6480 596 6520 684
rect 6480 564 6484 596
rect 6516 564 6520 596
rect 6480 516 6520 564
rect 6480 484 6484 516
rect 6516 484 6520 516
rect 6480 436 6520 484
rect 6480 404 6484 436
rect 6516 404 6520 436
rect 6480 356 6520 404
rect 6480 324 6484 356
rect 6516 324 6520 356
rect 6480 276 6520 324
rect 6480 244 6484 276
rect 6516 244 6520 276
rect 6480 196 6520 244
rect 6480 164 6484 196
rect 6516 164 6520 196
rect 6480 116 6520 164
rect 6480 84 6484 116
rect 6516 84 6520 116
rect 6480 36 6520 84
rect 6480 4 6484 36
rect 6516 4 6520 36
rect 6480 -40 6520 4
rect 6560 6395 6600 16640
rect 6560 6365 6565 6395
rect 6595 6365 6600 6395
rect 6560 -40 6600 6365
rect 6640 16596 6680 16644
rect 6800 16836 6840 16840
rect 6800 16644 6804 16836
rect 6836 16644 6840 16836
rect 6640 16564 6644 16596
rect 6676 16564 6680 16596
rect 6640 16516 6680 16564
rect 6640 16484 6644 16516
rect 6676 16484 6680 16516
rect 6640 16436 6680 16484
rect 6640 16404 6644 16436
rect 6676 16404 6680 16436
rect 6640 16356 6680 16404
rect 6640 16324 6644 16356
rect 6676 16324 6680 16356
rect 6640 16276 6680 16324
rect 6640 16244 6644 16276
rect 6676 16244 6680 16276
rect 6640 16196 6680 16244
rect 6640 16164 6644 16196
rect 6676 16164 6680 16196
rect 6640 16116 6680 16164
rect 6640 16084 6644 16116
rect 6676 16084 6680 16116
rect 6640 16036 6680 16084
rect 6640 16004 6644 16036
rect 6676 16004 6680 16036
rect 6640 15956 6680 16004
rect 6640 15924 6644 15956
rect 6676 15924 6680 15956
rect 6640 15436 6680 15924
rect 6640 15404 6644 15436
rect 6676 15404 6680 15436
rect 6640 15356 6680 15404
rect 6640 15324 6644 15356
rect 6676 15324 6680 15356
rect 6640 15276 6680 15324
rect 6640 15244 6644 15276
rect 6676 15244 6680 15276
rect 6640 15196 6680 15244
rect 6640 15164 6644 15196
rect 6676 15164 6680 15196
rect 6640 15116 6680 15164
rect 6640 15084 6644 15116
rect 6676 15084 6680 15116
rect 6640 15036 6680 15084
rect 6640 15004 6644 15036
rect 6676 15004 6680 15036
rect 6640 14956 6680 15004
rect 6640 14924 6644 14956
rect 6676 14924 6680 14956
rect 6640 14876 6680 14924
rect 6640 14844 6644 14876
rect 6676 14844 6680 14876
rect 6640 14796 6680 14844
rect 6640 14764 6644 14796
rect 6676 14764 6680 14796
rect 6640 14716 6680 14764
rect 6640 14684 6644 14716
rect 6676 14684 6680 14716
rect 6640 14636 6680 14684
rect 6640 14604 6644 14636
rect 6676 14604 6680 14636
rect 6640 14556 6680 14604
rect 6640 14524 6644 14556
rect 6676 14524 6680 14556
rect 6640 14476 6680 14524
rect 6640 14444 6644 14476
rect 6676 14444 6680 14476
rect 6640 13996 6680 14444
rect 6640 13964 6644 13996
rect 6676 13964 6680 13996
rect 6640 13876 6680 13964
rect 6640 13844 6644 13876
rect 6676 13844 6680 13876
rect 6640 13796 6680 13844
rect 6640 13764 6644 13796
rect 6676 13764 6680 13796
rect 6640 13716 6680 13764
rect 6640 13684 6644 13716
rect 6676 13684 6680 13716
rect 6640 13636 6680 13684
rect 6640 13604 6644 13636
rect 6676 13604 6680 13636
rect 6640 13556 6680 13604
rect 6640 13524 6644 13556
rect 6676 13524 6680 13556
rect 6640 13476 6680 13524
rect 6640 13444 6644 13476
rect 6676 13444 6680 13476
rect 6640 13396 6680 13444
rect 6640 13364 6644 13396
rect 6676 13364 6680 13396
rect 6640 13316 6680 13364
rect 6640 13284 6644 13316
rect 6676 13284 6680 13316
rect 6640 13236 6680 13284
rect 6640 13204 6644 13236
rect 6676 13204 6680 13236
rect 6640 13156 6680 13204
rect 6640 13124 6644 13156
rect 6676 13124 6680 13156
rect 6640 13076 6680 13124
rect 6640 13044 6644 13076
rect 6676 13044 6680 13076
rect 6640 12996 6680 13044
rect 6640 12964 6644 12996
rect 6676 12964 6680 12996
rect 6640 12516 6680 12964
rect 6640 12484 6644 12516
rect 6676 12484 6680 12516
rect 6640 12436 6680 12484
rect 6640 12404 6644 12436
rect 6676 12404 6680 12436
rect 6640 12316 6680 12404
rect 6640 12284 6644 12316
rect 6676 12284 6680 12316
rect 6640 12236 6680 12284
rect 6640 12204 6644 12236
rect 6676 12204 6680 12236
rect 6640 12156 6680 12204
rect 6640 12124 6644 12156
rect 6676 12124 6680 12156
rect 6640 12076 6680 12124
rect 6640 12044 6644 12076
rect 6676 12044 6680 12076
rect 6640 11996 6680 12044
rect 6640 11964 6644 11996
rect 6676 11964 6680 11996
rect 6640 11916 6680 11964
rect 6640 11884 6644 11916
rect 6676 11884 6680 11916
rect 6640 11836 6680 11884
rect 6640 11804 6644 11836
rect 6676 11804 6680 11836
rect 6640 11756 6680 11804
rect 6640 11724 6644 11756
rect 6676 11724 6680 11756
rect 6640 11676 6680 11724
rect 6640 11644 6644 11676
rect 6676 11644 6680 11676
rect 6640 11596 6680 11644
rect 6640 11564 6644 11596
rect 6676 11564 6680 11596
rect 6640 11516 6680 11564
rect 6640 11484 6644 11516
rect 6676 11484 6680 11516
rect 6640 11436 6680 11484
rect 6640 11404 6644 11436
rect 6676 11404 6680 11436
rect 6640 11356 6680 11404
rect 6640 11324 6644 11356
rect 6676 11324 6680 11356
rect 6640 11196 6680 11324
rect 6640 11164 6644 11196
rect 6676 11164 6680 11196
rect 6640 11116 6680 11164
rect 6640 11084 6644 11116
rect 6676 11084 6680 11116
rect 6640 11036 6680 11084
rect 6640 11004 6644 11036
rect 6676 11004 6680 11036
rect 6640 10876 6680 11004
rect 6640 10844 6644 10876
rect 6676 10844 6680 10876
rect 6640 10716 6680 10844
rect 6640 10684 6644 10716
rect 6676 10684 6680 10716
rect 6640 10636 6680 10684
rect 6640 10604 6644 10636
rect 6676 10604 6680 10636
rect 6640 10476 6680 10604
rect 6640 10444 6644 10476
rect 6676 10444 6680 10476
rect 6640 10316 6680 10444
rect 6640 10284 6644 10316
rect 6676 10284 6680 10316
rect 6640 10236 6680 10284
rect 6640 10204 6644 10236
rect 6676 10204 6680 10236
rect 6640 10156 6680 10204
rect 6640 10124 6644 10156
rect 6676 10124 6680 10156
rect 6640 10076 6680 10124
rect 6640 10044 6644 10076
rect 6676 10044 6680 10076
rect 6640 9996 6680 10044
rect 6640 9964 6644 9996
rect 6676 9964 6680 9996
rect 6640 9916 6680 9964
rect 6640 9884 6644 9916
rect 6676 9884 6680 9916
rect 6640 9836 6680 9884
rect 6640 9804 6644 9836
rect 6676 9804 6680 9836
rect 6640 9756 6680 9804
rect 6640 9724 6644 9756
rect 6676 9724 6680 9756
rect 6640 9676 6680 9724
rect 6640 9644 6644 9676
rect 6676 9644 6680 9676
rect 6640 9596 6680 9644
rect 6640 9564 6644 9596
rect 6676 9564 6680 9596
rect 6640 9516 6680 9564
rect 6640 9484 6644 9516
rect 6676 9484 6680 9516
rect 6640 9436 6680 9484
rect 6640 9404 6644 9436
rect 6676 9404 6680 9436
rect 6640 9356 6680 9404
rect 6640 9324 6644 9356
rect 6676 9324 6680 9356
rect 6640 9276 6680 9324
rect 6640 9244 6644 9276
rect 6676 9244 6680 9276
rect 6640 9116 6680 9244
rect 6640 9084 6644 9116
rect 6676 9084 6680 9116
rect 6640 9036 6680 9084
rect 6640 9004 6644 9036
rect 6676 9004 6680 9036
rect 6640 8956 6680 9004
rect 6640 8924 6644 8956
rect 6676 8924 6680 8956
rect 6640 8636 6680 8924
rect 6640 8604 6644 8636
rect 6676 8604 6680 8636
rect 6640 8556 6680 8604
rect 6640 8524 6644 8556
rect 6676 8524 6680 8556
rect 6640 8396 6680 8524
rect 6640 8364 6644 8396
rect 6676 8364 6680 8396
rect 6640 8236 6680 8364
rect 6640 8204 6644 8236
rect 6676 8204 6680 8236
rect 6640 8156 6680 8204
rect 6640 8124 6644 8156
rect 6676 8124 6680 8156
rect 6640 8076 6680 8124
rect 6640 8044 6644 8076
rect 6676 8044 6680 8076
rect 6640 7996 6680 8044
rect 6640 7964 6644 7996
rect 6676 7964 6680 7996
rect 6640 7916 6680 7964
rect 6640 7884 6644 7916
rect 6676 7884 6680 7916
rect 6640 7836 6680 7884
rect 6640 7804 6644 7836
rect 6676 7804 6680 7836
rect 6640 7756 6680 7804
rect 6640 7724 6644 7756
rect 6676 7724 6680 7756
rect 6640 7676 6680 7724
rect 6640 7644 6644 7676
rect 6676 7644 6680 7676
rect 6640 7596 6680 7644
rect 6640 7564 6644 7596
rect 6676 7564 6680 7596
rect 6640 7516 6680 7564
rect 6640 7484 6644 7516
rect 6676 7484 6680 7516
rect 6640 7436 6680 7484
rect 6640 7404 6644 7436
rect 6676 7404 6680 7436
rect 6640 7356 6680 7404
rect 6640 7324 6644 7356
rect 6676 7324 6680 7356
rect 6640 7276 6680 7324
rect 6640 7244 6644 7276
rect 6676 7244 6680 7276
rect 6640 7196 6680 7244
rect 6640 7164 6644 7196
rect 6676 7164 6680 7196
rect 6640 7116 6680 7164
rect 6640 7084 6644 7116
rect 6676 7084 6680 7116
rect 6640 7036 6680 7084
rect 6640 7004 6644 7036
rect 6676 7004 6680 7036
rect 6640 6956 6680 7004
rect 6640 6924 6644 6956
rect 6676 6924 6680 6956
rect 6640 6876 6680 6924
rect 6640 6844 6644 6876
rect 6676 6844 6680 6876
rect 6640 6796 6680 6844
rect 6640 6764 6644 6796
rect 6676 6764 6680 6796
rect 6640 6716 6680 6764
rect 6640 6684 6644 6716
rect 6676 6684 6680 6716
rect 6640 6636 6680 6684
rect 6640 6604 6644 6636
rect 6676 6604 6680 6636
rect 6640 6556 6680 6604
rect 6640 6524 6644 6556
rect 6676 6524 6680 6556
rect 6640 6476 6680 6524
rect 6640 6444 6644 6476
rect 6676 6444 6680 6476
rect 6640 6396 6680 6444
rect 6640 6364 6644 6396
rect 6676 6364 6680 6396
rect 6640 6316 6680 6364
rect 6640 6284 6644 6316
rect 6676 6284 6680 6316
rect 6640 6236 6680 6284
rect 6640 6204 6644 6236
rect 6676 6204 6680 6236
rect 6640 6156 6680 6204
rect 6640 6124 6644 6156
rect 6676 6124 6680 6156
rect 6640 5996 6680 6124
rect 6640 5964 6644 5996
rect 6676 5964 6680 5996
rect 6640 5836 6680 5964
rect 6640 5804 6644 5836
rect 6676 5804 6680 5836
rect 6640 5756 6680 5804
rect 6640 5724 6644 5756
rect 6676 5724 6680 5756
rect 6640 5676 6680 5724
rect 6640 5644 6644 5676
rect 6676 5644 6680 5676
rect 6640 5596 6680 5644
rect 6640 5564 6644 5596
rect 6676 5564 6680 5596
rect 6640 5516 6680 5564
rect 6640 5484 6644 5516
rect 6676 5484 6680 5516
rect 6640 5436 6680 5484
rect 6640 5404 6644 5436
rect 6676 5404 6680 5436
rect 6640 5356 6680 5404
rect 6640 5324 6644 5356
rect 6676 5324 6680 5356
rect 6640 5276 6680 5324
rect 6640 5244 6644 5276
rect 6676 5244 6680 5276
rect 6640 5196 6680 5244
rect 6640 5164 6644 5196
rect 6676 5164 6680 5196
rect 6640 5116 6680 5164
rect 6640 5084 6644 5116
rect 6676 5084 6680 5116
rect 6640 5036 6680 5084
rect 6640 5004 6644 5036
rect 6676 5004 6680 5036
rect 6640 4956 6680 5004
rect 6640 4924 6644 4956
rect 6676 4924 6680 4956
rect 6640 4876 6680 4924
rect 6640 4844 6644 4876
rect 6676 4844 6680 4876
rect 6640 4796 6680 4844
rect 6640 4764 6644 4796
rect 6676 4764 6680 4796
rect 6640 4716 6680 4764
rect 6640 4684 6644 4716
rect 6676 4684 6680 4716
rect 6640 4636 6680 4684
rect 6640 4604 6644 4636
rect 6676 4604 6680 4636
rect 6640 4556 6680 4604
rect 6640 4524 6644 4556
rect 6676 4524 6680 4556
rect 6640 4476 6680 4524
rect 6640 4444 6644 4476
rect 6676 4444 6680 4476
rect 6640 4396 6680 4444
rect 6640 4364 6644 4396
rect 6676 4364 6680 4396
rect 6640 4316 6680 4364
rect 6640 4284 6644 4316
rect 6676 4284 6680 4316
rect 6640 4236 6680 4284
rect 6640 4204 6644 4236
rect 6676 4204 6680 4236
rect 6640 4156 6680 4204
rect 6640 4124 6644 4156
rect 6676 4124 6680 4156
rect 6640 4076 6680 4124
rect 6640 4044 6644 4076
rect 6676 4044 6680 4076
rect 6640 3996 6680 4044
rect 6640 3964 6644 3996
rect 6676 3964 6680 3996
rect 6640 3916 6680 3964
rect 6640 3884 6644 3916
rect 6676 3884 6680 3916
rect 6640 3836 6680 3884
rect 6640 3804 6644 3836
rect 6676 3804 6680 3836
rect 6640 3756 6680 3804
rect 6640 3724 6644 3756
rect 6676 3724 6680 3756
rect 6640 3596 6680 3724
rect 6640 3564 6644 3596
rect 6676 3564 6680 3596
rect 6640 3436 6680 3564
rect 6640 3404 6644 3436
rect 6676 3404 6680 3436
rect 6640 3356 6680 3404
rect 6640 3324 6644 3356
rect 6676 3324 6680 3356
rect 6640 3276 6680 3324
rect 6640 3244 6644 3276
rect 6676 3244 6680 3276
rect 6640 3196 6680 3244
rect 6640 3164 6644 3196
rect 6676 3164 6680 3196
rect 6640 3116 6680 3164
rect 6640 3084 6644 3116
rect 6676 3084 6680 3116
rect 6640 3036 6680 3084
rect 6640 3004 6644 3036
rect 6676 3004 6680 3036
rect 6640 2956 6680 3004
rect 6640 2924 6644 2956
rect 6676 2924 6680 2956
rect 6640 2876 6680 2924
rect 6640 2844 6644 2876
rect 6676 2844 6680 2876
rect 6640 2796 6680 2844
rect 6640 2764 6644 2796
rect 6676 2764 6680 2796
rect 6640 2716 6680 2764
rect 6640 2684 6644 2716
rect 6676 2684 6680 2716
rect 6640 2636 6680 2684
rect 6640 2604 6644 2636
rect 6676 2604 6680 2636
rect 6640 2556 6680 2604
rect 6640 2524 6644 2556
rect 6676 2524 6680 2556
rect 6640 2476 6680 2524
rect 6640 2444 6644 2476
rect 6676 2444 6680 2476
rect 6640 2396 6680 2444
rect 6640 2364 6644 2396
rect 6676 2364 6680 2396
rect 6640 2316 6680 2364
rect 6640 2284 6644 2316
rect 6676 2284 6680 2316
rect 6640 2236 6680 2284
rect 6640 2204 6644 2236
rect 6676 2204 6680 2236
rect 6640 2156 6680 2204
rect 6640 2124 6644 2156
rect 6676 2124 6680 2156
rect 6640 2076 6680 2124
rect 6640 2044 6644 2076
rect 6676 2044 6680 2076
rect 6640 1996 6680 2044
rect 6640 1964 6644 1996
rect 6676 1964 6680 1996
rect 6640 1916 6680 1964
rect 6640 1884 6644 1916
rect 6676 1884 6680 1916
rect 6640 1836 6680 1884
rect 6640 1804 6644 1836
rect 6676 1804 6680 1836
rect 6640 1756 6680 1804
rect 6640 1724 6644 1756
rect 6676 1724 6680 1756
rect 6640 1676 6680 1724
rect 6640 1644 6644 1676
rect 6676 1644 6680 1676
rect 6640 1596 6680 1644
rect 6640 1564 6644 1596
rect 6676 1564 6680 1596
rect 6640 1516 6680 1564
rect 6640 1484 6644 1516
rect 6676 1484 6680 1516
rect 6640 1436 6680 1484
rect 6640 1404 6644 1436
rect 6676 1404 6680 1436
rect 6640 1356 6680 1404
rect 6640 1324 6644 1356
rect 6676 1324 6680 1356
rect 6640 1276 6680 1324
rect 6640 1244 6644 1276
rect 6676 1244 6680 1276
rect 6640 1196 6680 1244
rect 6640 1164 6644 1196
rect 6676 1164 6680 1196
rect 6640 1116 6680 1164
rect 6640 1084 6644 1116
rect 6676 1084 6680 1116
rect 6640 1036 6680 1084
rect 6640 1004 6644 1036
rect 6676 1004 6680 1036
rect 6640 956 6680 1004
rect 6640 924 6644 956
rect 6676 924 6680 956
rect 6640 876 6680 924
rect 6640 844 6644 876
rect 6676 844 6680 876
rect 6640 796 6680 844
rect 6640 764 6644 796
rect 6676 764 6680 796
rect 6640 716 6680 764
rect 6640 684 6644 716
rect 6676 684 6680 716
rect 6640 596 6680 684
rect 6640 564 6644 596
rect 6676 564 6680 596
rect 6640 516 6680 564
rect 6640 484 6644 516
rect 6676 484 6680 516
rect 6640 436 6680 484
rect 6640 404 6644 436
rect 6676 404 6680 436
rect 6640 356 6680 404
rect 6640 324 6644 356
rect 6676 324 6680 356
rect 6640 276 6680 324
rect 6640 244 6644 276
rect 6676 244 6680 276
rect 6640 196 6680 244
rect 6640 164 6644 196
rect 6676 164 6680 196
rect 6640 116 6680 164
rect 6640 84 6644 116
rect 6676 84 6680 116
rect 6640 36 6680 84
rect 6640 4 6644 36
rect 6676 4 6680 36
rect 6640 -40 6680 4
rect 6720 8315 6760 16640
rect 6720 8285 6725 8315
rect 6755 8285 6760 8315
rect 6720 3515 6760 8285
rect 6720 3485 6725 3515
rect 6755 3485 6760 3515
rect 6720 -40 6760 3485
rect 6800 16596 6840 16644
rect 6960 16836 7000 16840
rect 6960 16644 6964 16836
rect 6996 16644 7000 16836
rect 6800 16564 6804 16596
rect 6836 16564 6840 16596
rect 6800 16516 6840 16564
rect 6800 16484 6804 16516
rect 6836 16484 6840 16516
rect 6800 16436 6840 16484
rect 6800 16404 6804 16436
rect 6836 16404 6840 16436
rect 6800 16356 6840 16404
rect 6800 16324 6804 16356
rect 6836 16324 6840 16356
rect 6800 16276 6840 16324
rect 6800 16244 6804 16276
rect 6836 16244 6840 16276
rect 6800 16196 6840 16244
rect 6800 16164 6804 16196
rect 6836 16164 6840 16196
rect 6800 16116 6840 16164
rect 6800 16084 6804 16116
rect 6836 16084 6840 16116
rect 6800 16036 6840 16084
rect 6800 16004 6804 16036
rect 6836 16004 6840 16036
rect 6800 15956 6840 16004
rect 6800 15924 6804 15956
rect 6836 15924 6840 15956
rect 6800 15436 6840 15924
rect 6800 15404 6804 15436
rect 6836 15404 6840 15436
rect 6800 15356 6840 15404
rect 6800 15324 6804 15356
rect 6836 15324 6840 15356
rect 6800 15276 6840 15324
rect 6800 15244 6804 15276
rect 6836 15244 6840 15276
rect 6800 15196 6840 15244
rect 6800 15164 6804 15196
rect 6836 15164 6840 15196
rect 6800 15116 6840 15164
rect 6800 15084 6804 15116
rect 6836 15084 6840 15116
rect 6800 15036 6840 15084
rect 6800 15004 6804 15036
rect 6836 15004 6840 15036
rect 6800 14956 6840 15004
rect 6800 14924 6804 14956
rect 6836 14924 6840 14956
rect 6800 14876 6840 14924
rect 6800 14844 6804 14876
rect 6836 14844 6840 14876
rect 6800 14796 6840 14844
rect 6800 14764 6804 14796
rect 6836 14764 6840 14796
rect 6800 14716 6840 14764
rect 6800 14684 6804 14716
rect 6836 14684 6840 14716
rect 6800 14636 6840 14684
rect 6800 14604 6804 14636
rect 6836 14604 6840 14636
rect 6800 14556 6840 14604
rect 6800 14524 6804 14556
rect 6836 14524 6840 14556
rect 6800 14476 6840 14524
rect 6800 14444 6804 14476
rect 6836 14444 6840 14476
rect 6800 13996 6840 14444
rect 6800 13964 6804 13996
rect 6836 13964 6840 13996
rect 6800 13876 6840 13964
rect 6800 13844 6804 13876
rect 6836 13844 6840 13876
rect 6800 13796 6840 13844
rect 6800 13764 6804 13796
rect 6836 13764 6840 13796
rect 6800 13716 6840 13764
rect 6800 13684 6804 13716
rect 6836 13684 6840 13716
rect 6800 13636 6840 13684
rect 6800 13604 6804 13636
rect 6836 13604 6840 13636
rect 6800 13556 6840 13604
rect 6800 13524 6804 13556
rect 6836 13524 6840 13556
rect 6800 13476 6840 13524
rect 6800 13444 6804 13476
rect 6836 13444 6840 13476
rect 6800 13396 6840 13444
rect 6800 13364 6804 13396
rect 6836 13364 6840 13396
rect 6800 13316 6840 13364
rect 6800 13284 6804 13316
rect 6836 13284 6840 13316
rect 6800 13236 6840 13284
rect 6800 13204 6804 13236
rect 6836 13204 6840 13236
rect 6800 13156 6840 13204
rect 6800 13124 6804 13156
rect 6836 13124 6840 13156
rect 6800 13076 6840 13124
rect 6800 13044 6804 13076
rect 6836 13044 6840 13076
rect 6800 12996 6840 13044
rect 6800 12964 6804 12996
rect 6836 12964 6840 12996
rect 6800 12516 6840 12964
rect 6800 12484 6804 12516
rect 6836 12484 6840 12516
rect 6800 12436 6840 12484
rect 6800 12404 6804 12436
rect 6836 12404 6840 12436
rect 6800 12316 6840 12404
rect 6800 12284 6804 12316
rect 6836 12284 6840 12316
rect 6800 12236 6840 12284
rect 6800 12204 6804 12236
rect 6836 12204 6840 12236
rect 6800 12156 6840 12204
rect 6800 12124 6804 12156
rect 6836 12124 6840 12156
rect 6800 12076 6840 12124
rect 6800 12044 6804 12076
rect 6836 12044 6840 12076
rect 6800 11996 6840 12044
rect 6800 11964 6804 11996
rect 6836 11964 6840 11996
rect 6800 11916 6840 11964
rect 6800 11884 6804 11916
rect 6836 11884 6840 11916
rect 6800 11836 6840 11884
rect 6800 11804 6804 11836
rect 6836 11804 6840 11836
rect 6800 11756 6840 11804
rect 6800 11724 6804 11756
rect 6836 11724 6840 11756
rect 6800 11676 6840 11724
rect 6800 11644 6804 11676
rect 6836 11644 6840 11676
rect 6800 11596 6840 11644
rect 6800 11564 6804 11596
rect 6836 11564 6840 11596
rect 6800 11516 6840 11564
rect 6800 11484 6804 11516
rect 6836 11484 6840 11516
rect 6800 11436 6840 11484
rect 6800 11404 6804 11436
rect 6836 11404 6840 11436
rect 6800 11356 6840 11404
rect 6800 11324 6804 11356
rect 6836 11324 6840 11356
rect 6800 11196 6840 11324
rect 6800 11164 6804 11196
rect 6836 11164 6840 11196
rect 6800 11116 6840 11164
rect 6800 11084 6804 11116
rect 6836 11084 6840 11116
rect 6800 11036 6840 11084
rect 6800 11004 6804 11036
rect 6836 11004 6840 11036
rect 6800 10876 6840 11004
rect 6800 10844 6804 10876
rect 6836 10844 6840 10876
rect 6800 10716 6840 10844
rect 6800 10684 6804 10716
rect 6836 10684 6840 10716
rect 6800 10636 6840 10684
rect 6800 10604 6804 10636
rect 6836 10604 6840 10636
rect 6800 10476 6840 10604
rect 6800 10444 6804 10476
rect 6836 10444 6840 10476
rect 6800 10316 6840 10444
rect 6800 10284 6804 10316
rect 6836 10284 6840 10316
rect 6800 10236 6840 10284
rect 6800 10204 6804 10236
rect 6836 10204 6840 10236
rect 6800 10156 6840 10204
rect 6800 10124 6804 10156
rect 6836 10124 6840 10156
rect 6800 10076 6840 10124
rect 6800 10044 6804 10076
rect 6836 10044 6840 10076
rect 6800 9996 6840 10044
rect 6800 9964 6804 9996
rect 6836 9964 6840 9996
rect 6800 9916 6840 9964
rect 6800 9884 6804 9916
rect 6836 9884 6840 9916
rect 6800 9836 6840 9884
rect 6800 9804 6804 9836
rect 6836 9804 6840 9836
rect 6800 9756 6840 9804
rect 6800 9724 6804 9756
rect 6836 9724 6840 9756
rect 6800 9676 6840 9724
rect 6800 9644 6804 9676
rect 6836 9644 6840 9676
rect 6800 9596 6840 9644
rect 6800 9564 6804 9596
rect 6836 9564 6840 9596
rect 6800 9516 6840 9564
rect 6800 9484 6804 9516
rect 6836 9484 6840 9516
rect 6800 9436 6840 9484
rect 6800 9404 6804 9436
rect 6836 9404 6840 9436
rect 6800 9356 6840 9404
rect 6800 9324 6804 9356
rect 6836 9324 6840 9356
rect 6800 9276 6840 9324
rect 6800 9244 6804 9276
rect 6836 9244 6840 9276
rect 6800 9116 6840 9244
rect 6800 9084 6804 9116
rect 6836 9084 6840 9116
rect 6800 9036 6840 9084
rect 6800 9004 6804 9036
rect 6836 9004 6840 9036
rect 6800 8956 6840 9004
rect 6800 8924 6804 8956
rect 6836 8924 6840 8956
rect 6800 8636 6840 8924
rect 6800 8604 6804 8636
rect 6836 8604 6840 8636
rect 6800 8556 6840 8604
rect 6800 8524 6804 8556
rect 6836 8524 6840 8556
rect 6800 8396 6840 8524
rect 6800 8364 6804 8396
rect 6836 8364 6840 8396
rect 6800 8316 6840 8364
rect 6800 8284 6804 8316
rect 6836 8284 6840 8316
rect 6800 8236 6840 8284
rect 6800 8204 6804 8236
rect 6836 8204 6840 8236
rect 6800 8156 6840 8204
rect 6800 8124 6804 8156
rect 6836 8124 6840 8156
rect 6800 8076 6840 8124
rect 6800 8044 6804 8076
rect 6836 8044 6840 8076
rect 6800 7996 6840 8044
rect 6800 7964 6804 7996
rect 6836 7964 6840 7996
rect 6800 7916 6840 7964
rect 6800 7884 6804 7916
rect 6836 7884 6840 7916
rect 6800 7836 6840 7884
rect 6800 7804 6804 7836
rect 6836 7804 6840 7836
rect 6800 7756 6840 7804
rect 6800 7724 6804 7756
rect 6836 7724 6840 7756
rect 6800 7676 6840 7724
rect 6800 7644 6804 7676
rect 6836 7644 6840 7676
rect 6800 7596 6840 7644
rect 6800 7564 6804 7596
rect 6836 7564 6840 7596
rect 6800 7516 6840 7564
rect 6800 7484 6804 7516
rect 6836 7484 6840 7516
rect 6800 7436 6840 7484
rect 6800 7404 6804 7436
rect 6836 7404 6840 7436
rect 6800 7356 6840 7404
rect 6800 7324 6804 7356
rect 6836 7324 6840 7356
rect 6800 7276 6840 7324
rect 6800 7244 6804 7276
rect 6836 7244 6840 7276
rect 6800 7196 6840 7244
rect 6800 7164 6804 7196
rect 6836 7164 6840 7196
rect 6800 7116 6840 7164
rect 6800 7084 6804 7116
rect 6836 7084 6840 7116
rect 6800 7036 6840 7084
rect 6800 7004 6804 7036
rect 6836 7004 6840 7036
rect 6800 6956 6840 7004
rect 6800 6924 6804 6956
rect 6836 6924 6840 6956
rect 6800 6876 6840 6924
rect 6800 6844 6804 6876
rect 6836 6844 6840 6876
rect 6800 6796 6840 6844
rect 6800 6764 6804 6796
rect 6836 6764 6840 6796
rect 6800 6716 6840 6764
rect 6800 6684 6804 6716
rect 6836 6684 6840 6716
rect 6800 6636 6840 6684
rect 6800 6604 6804 6636
rect 6836 6604 6840 6636
rect 6800 6556 6840 6604
rect 6800 6524 6804 6556
rect 6836 6524 6840 6556
rect 6800 6476 6840 6524
rect 6800 6444 6804 6476
rect 6836 6444 6840 6476
rect 6800 6396 6840 6444
rect 6800 6364 6804 6396
rect 6836 6364 6840 6396
rect 6800 6316 6840 6364
rect 6800 6284 6804 6316
rect 6836 6284 6840 6316
rect 6800 6236 6840 6284
rect 6800 6204 6804 6236
rect 6836 6204 6840 6236
rect 6800 6156 6840 6204
rect 6800 6124 6804 6156
rect 6836 6124 6840 6156
rect 6800 5996 6840 6124
rect 6800 5964 6804 5996
rect 6836 5964 6840 5996
rect 6800 5836 6840 5964
rect 6800 5804 6804 5836
rect 6836 5804 6840 5836
rect 6800 5756 6840 5804
rect 6800 5724 6804 5756
rect 6836 5724 6840 5756
rect 6800 5676 6840 5724
rect 6800 5644 6804 5676
rect 6836 5644 6840 5676
rect 6800 5596 6840 5644
rect 6800 5564 6804 5596
rect 6836 5564 6840 5596
rect 6800 5516 6840 5564
rect 6800 5484 6804 5516
rect 6836 5484 6840 5516
rect 6800 5436 6840 5484
rect 6800 5404 6804 5436
rect 6836 5404 6840 5436
rect 6800 5356 6840 5404
rect 6800 5324 6804 5356
rect 6836 5324 6840 5356
rect 6800 5276 6840 5324
rect 6800 5244 6804 5276
rect 6836 5244 6840 5276
rect 6800 5196 6840 5244
rect 6800 5164 6804 5196
rect 6836 5164 6840 5196
rect 6800 5116 6840 5164
rect 6800 5084 6804 5116
rect 6836 5084 6840 5116
rect 6800 5036 6840 5084
rect 6800 5004 6804 5036
rect 6836 5004 6840 5036
rect 6800 4956 6840 5004
rect 6800 4924 6804 4956
rect 6836 4924 6840 4956
rect 6800 4876 6840 4924
rect 6800 4844 6804 4876
rect 6836 4844 6840 4876
rect 6800 4796 6840 4844
rect 6800 4764 6804 4796
rect 6836 4764 6840 4796
rect 6800 4716 6840 4764
rect 6800 4684 6804 4716
rect 6836 4684 6840 4716
rect 6800 4636 6840 4684
rect 6800 4604 6804 4636
rect 6836 4604 6840 4636
rect 6800 4556 6840 4604
rect 6800 4524 6804 4556
rect 6836 4524 6840 4556
rect 6800 4476 6840 4524
rect 6800 4444 6804 4476
rect 6836 4444 6840 4476
rect 6800 4396 6840 4444
rect 6800 4364 6804 4396
rect 6836 4364 6840 4396
rect 6800 4316 6840 4364
rect 6800 4284 6804 4316
rect 6836 4284 6840 4316
rect 6800 4236 6840 4284
rect 6800 4204 6804 4236
rect 6836 4204 6840 4236
rect 6800 4156 6840 4204
rect 6800 4124 6804 4156
rect 6836 4124 6840 4156
rect 6800 4076 6840 4124
rect 6800 4044 6804 4076
rect 6836 4044 6840 4076
rect 6800 3996 6840 4044
rect 6800 3964 6804 3996
rect 6836 3964 6840 3996
rect 6800 3916 6840 3964
rect 6800 3884 6804 3916
rect 6836 3884 6840 3916
rect 6800 3836 6840 3884
rect 6800 3804 6804 3836
rect 6836 3804 6840 3836
rect 6800 3756 6840 3804
rect 6800 3724 6804 3756
rect 6836 3724 6840 3756
rect 6800 3596 6840 3724
rect 6800 3564 6804 3596
rect 6836 3564 6840 3596
rect 6800 3516 6840 3564
rect 6800 3484 6804 3516
rect 6836 3484 6840 3516
rect 6800 3436 6840 3484
rect 6800 3404 6804 3436
rect 6836 3404 6840 3436
rect 6800 3356 6840 3404
rect 6800 3324 6804 3356
rect 6836 3324 6840 3356
rect 6800 3276 6840 3324
rect 6800 3244 6804 3276
rect 6836 3244 6840 3276
rect 6800 3196 6840 3244
rect 6800 3164 6804 3196
rect 6836 3164 6840 3196
rect 6800 3116 6840 3164
rect 6800 3084 6804 3116
rect 6836 3084 6840 3116
rect 6800 3036 6840 3084
rect 6800 3004 6804 3036
rect 6836 3004 6840 3036
rect 6800 2956 6840 3004
rect 6800 2924 6804 2956
rect 6836 2924 6840 2956
rect 6800 2876 6840 2924
rect 6800 2844 6804 2876
rect 6836 2844 6840 2876
rect 6800 2796 6840 2844
rect 6800 2764 6804 2796
rect 6836 2764 6840 2796
rect 6800 2716 6840 2764
rect 6800 2684 6804 2716
rect 6836 2684 6840 2716
rect 6800 2636 6840 2684
rect 6800 2604 6804 2636
rect 6836 2604 6840 2636
rect 6800 2556 6840 2604
rect 6800 2524 6804 2556
rect 6836 2524 6840 2556
rect 6800 2476 6840 2524
rect 6800 2444 6804 2476
rect 6836 2444 6840 2476
rect 6800 2396 6840 2444
rect 6800 2364 6804 2396
rect 6836 2364 6840 2396
rect 6800 2316 6840 2364
rect 6800 2284 6804 2316
rect 6836 2284 6840 2316
rect 6800 2236 6840 2284
rect 6800 2204 6804 2236
rect 6836 2204 6840 2236
rect 6800 2156 6840 2204
rect 6800 2124 6804 2156
rect 6836 2124 6840 2156
rect 6800 2076 6840 2124
rect 6800 2044 6804 2076
rect 6836 2044 6840 2076
rect 6800 1996 6840 2044
rect 6800 1964 6804 1996
rect 6836 1964 6840 1996
rect 6800 1916 6840 1964
rect 6800 1884 6804 1916
rect 6836 1884 6840 1916
rect 6800 1836 6840 1884
rect 6800 1804 6804 1836
rect 6836 1804 6840 1836
rect 6800 1756 6840 1804
rect 6800 1724 6804 1756
rect 6836 1724 6840 1756
rect 6800 1676 6840 1724
rect 6800 1644 6804 1676
rect 6836 1644 6840 1676
rect 6800 1596 6840 1644
rect 6800 1564 6804 1596
rect 6836 1564 6840 1596
rect 6800 1516 6840 1564
rect 6800 1484 6804 1516
rect 6836 1484 6840 1516
rect 6800 1436 6840 1484
rect 6800 1404 6804 1436
rect 6836 1404 6840 1436
rect 6800 1356 6840 1404
rect 6800 1324 6804 1356
rect 6836 1324 6840 1356
rect 6800 1276 6840 1324
rect 6800 1244 6804 1276
rect 6836 1244 6840 1276
rect 6800 1196 6840 1244
rect 6800 1164 6804 1196
rect 6836 1164 6840 1196
rect 6800 1116 6840 1164
rect 6800 1084 6804 1116
rect 6836 1084 6840 1116
rect 6800 1036 6840 1084
rect 6800 1004 6804 1036
rect 6836 1004 6840 1036
rect 6800 956 6840 1004
rect 6800 924 6804 956
rect 6836 924 6840 956
rect 6800 876 6840 924
rect 6800 844 6804 876
rect 6836 844 6840 876
rect 6800 796 6840 844
rect 6800 764 6804 796
rect 6836 764 6840 796
rect 6800 716 6840 764
rect 6800 684 6804 716
rect 6836 684 6840 716
rect 6800 596 6840 684
rect 6800 564 6804 596
rect 6836 564 6840 596
rect 6800 516 6840 564
rect 6800 484 6804 516
rect 6836 484 6840 516
rect 6800 436 6840 484
rect 6800 404 6804 436
rect 6836 404 6840 436
rect 6800 356 6840 404
rect 6800 324 6804 356
rect 6836 324 6840 356
rect 6800 276 6840 324
rect 6800 244 6804 276
rect 6836 244 6840 276
rect 6800 196 6840 244
rect 6800 164 6804 196
rect 6836 164 6840 196
rect 6800 116 6840 164
rect 6800 84 6804 116
rect 6836 84 6840 116
rect 6800 36 6840 84
rect 6800 4 6804 36
rect 6836 4 6840 36
rect 6800 -40 6840 4
rect 6880 10395 6920 16640
rect 6880 10365 6885 10395
rect 6915 10365 6920 10395
rect 6880 5915 6920 10365
rect 6880 5885 6885 5915
rect 6915 5885 6920 5915
rect 6880 -40 6920 5885
rect 6960 16596 7000 16644
rect 7120 16836 7160 16840
rect 7120 16644 7124 16836
rect 7156 16644 7160 16836
rect 6960 16564 6964 16596
rect 6996 16564 7000 16596
rect 6960 16516 7000 16564
rect 6960 16484 6964 16516
rect 6996 16484 7000 16516
rect 6960 16436 7000 16484
rect 6960 16404 6964 16436
rect 6996 16404 7000 16436
rect 6960 16356 7000 16404
rect 6960 16324 6964 16356
rect 6996 16324 7000 16356
rect 6960 16276 7000 16324
rect 6960 16244 6964 16276
rect 6996 16244 7000 16276
rect 6960 16196 7000 16244
rect 6960 16164 6964 16196
rect 6996 16164 7000 16196
rect 6960 16116 7000 16164
rect 6960 16084 6964 16116
rect 6996 16084 7000 16116
rect 6960 16036 7000 16084
rect 6960 16004 6964 16036
rect 6996 16004 7000 16036
rect 6960 15956 7000 16004
rect 6960 15924 6964 15956
rect 6996 15924 7000 15956
rect 6960 15436 7000 15924
rect 6960 15404 6964 15436
rect 6996 15404 7000 15436
rect 6960 15356 7000 15404
rect 6960 15324 6964 15356
rect 6996 15324 7000 15356
rect 6960 15276 7000 15324
rect 6960 15244 6964 15276
rect 6996 15244 7000 15276
rect 6960 15196 7000 15244
rect 6960 15164 6964 15196
rect 6996 15164 7000 15196
rect 6960 15116 7000 15164
rect 6960 15084 6964 15116
rect 6996 15084 7000 15116
rect 6960 15036 7000 15084
rect 6960 15004 6964 15036
rect 6996 15004 7000 15036
rect 6960 14956 7000 15004
rect 6960 14924 6964 14956
rect 6996 14924 7000 14956
rect 6960 14876 7000 14924
rect 6960 14844 6964 14876
rect 6996 14844 7000 14876
rect 6960 14796 7000 14844
rect 6960 14764 6964 14796
rect 6996 14764 7000 14796
rect 6960 14716 7000 14764
rect 6960 14684 6964 14716
rect 6996 14684 7000 14716
rect 6960 14636 7000 14684
rect 6960 14604 6964 14636
rect 6996 14604 7000 14636
rect 6960 14556 7000 14604
rect 6960 14524 6964 14556
rect 6996 14524 7000 14556
rect 6960 14476 7000 14524
rect 6960 14444 6964 14476
rect 6996 14444 7000 14476
rect 6960 14395 7000 14444
rect 6960 14365 6965 14395
rect 6995 14365 7000 14395
rect 6960 14235 7000 14365
rect 6960 14205 6965 14235
rect 6995 14205 7000 14235
rect 6960 14075 7000 14205
rect 6960 14045 6965 14075
rect 6995 14045 7000 14075
rect 6960 13996 7000 14045
rect 6960 13964 6964 13996
rect 6996 13964 7000 13996
rect 6960 13876 7000 13964
rect 6960 13844 6964 13876
rect 6996 13844 7000 13876
rect 6960 13796 7000 13844
rect 6960 13764 6964 13796
rect 6996 13764 7000 13796
rect 6960 13716 7000 13764
rect 6960 13684 6964 13716
rect 6996 13684 7000 13716
rect 6960 13636 7000 13684
rect 6960 13604 6964 13636
rect 6996 13604 7000 13636
rect 6960 13556 7000 13604
rect 6960 13524 6964 13556
rect 6996 13524 7000 13556
rect 6960 13476 7000 13524
rect 6960 13444 6964 13476
rect 6996 13444 7000 13476
rect 6960 13396 7000 13444
rect 6960 13364 6964 13396
rect 6996 13364 7000 13396
rect 6960 13316 7000 13364
rect 6960 13284 6964 13316
rect 6996 13284 7000 13316
rect 6960 13236 7000 13284
rect 6960 13204 6964 13236
rect 6996 13204 7000 13236
rect 6960 13156 7000 13204
rect 6960 13124 6964 13156
rect 6996 13124 7000 13156
rect 6960 13076 7000 13124
rect 6960 13044 6964 13076
rect 6996 13044 7000 13076
rect 6960 12996 7000 13044
rect 6960 12964 6964 12996
rect 6996 12964 7000 12996
rect 6960 12516 7000 12964
rect 6960 12484 6964 12516
rect 6996 12484 7000 12516
rect 6960 12436 7000 12484
rect 6960 12404 6964 12436
rect 6996 12404 7000 12436
rect 6960 12316 7000 12404
rect 6960 12284 6964 12316
rect 6996 12284 7000 12316
rect 6960 12236 7000 12284
rect 6960 12204 6964 12236
rect 6996 12204 7000 12236
rect 6960 12156 7000 12204
rect 6960 12124 6964 12156
rect 6996 12124 7000 12156
rect 6960 12076 7000 12124
rect 6960 12044 6964 12076
rect 6996 12044 7000 12076
rect 6960 11996 7000 12044
rect 6960 11964 6964 11996
rect 6996 11964 7000 11996
rect 6960 11916 7000 11964
rect 6960 11884 6964 11916
rect 6996 11884 7000 11916
rect 6960 11836 7000 11884
rect 6960 11804 6964 11836
rect 6996 11804 7000 11836
rect 6960 11756 7000 11804
rect 6960 11724 6964 11756
rect 6996 11724 7000 11756
rect 6960 11676 7000 11724
rect 6960 11644 6964 11676
rect 6996 11644 7000 11676
rect 6960 11596 7000 11644
rect 6960 11564 6964 11596
rect 6996 11564 7000 11596
rect 6960 11516 7000 11564
rect 6960 11484 6964 11516
rect 6996 11484 7000 11516
rect 6960 11436 7000 11484
rect 6960 11404 6964 11436
rect 6996 11404 7000 11436
rect 6960 11356 7000 11404
rect 6960 11324 6964 11356
rect 6996 11324 7000 11356
rect 6960 11196 7000 11324
rect 6960 11164 6964 11196
rect 6996 11164 7000 11196
rect 6960 11116 7000 11164
rect 6960 11084 6964 11116
rect 6996 11084 7000 11116
rect 6960 11036 7000 11084
rect 6960 11004 6964 11036
rect 6996 11004 7000 11036
rect 6960 10876 7000 11004
rect 6960 10844 6964 10876
rect 6996 10844 7000 10876
rect 6960 10716 7000 10844
rect 6960 10684 6964 10716
rect 6996 10684 7000 10716
rect 6960 10636 7000 10684
rect 6960 10604 6964 10636
rect 6996 10604 7000 10636
rect 6960 10476 7000 10604
rect 6960 10444 6964 10476
rect 6996 10444 7000 10476
rect 6960 10396 7000 10444
rect 6960 10364 6964 10396
rect 6996 10364 7000 10396
rect 6960 10316 7000 10364
rect 6960 10284 6964 10316
rect 6996 10284 7000 10316
rect 6960 10236 7000 10284
rect 6960 10204 6964 10236
rect 6996 10204 7000 10236
rect 6960 10156 7000 10204
rect 6960 10124 6964 10156
rect 6996 10124 7000 10156
rect 6960 10076 7000 10124
rect 6960 10044 6964 10076
rect 6996 10044 7000 10076
rect 6960 9996 7000 10044
rect 6960 9964 6964 9996
rect 6996 9964 7000 9996
rect 6960 9916 7000 9964
rect 6960 9884 6964 9916
rect 6996 9884 7000 9916
rect 6960 9836 7000 9884
rect 6960 9804 6964 9836
rect 6996 9804 7000 9836
rect 6960 9756 7000 9804
rect 6960 9724 6964 9756
rect 6996 9724 7000 9756
rect 6960 9676 7000 9724
rect 6960 9644 6964 9676
rect 6996 9644 7000 9676
rect 6960 9596 7000 9644
rect 6960 9564 6964 9596
rect 6996 9564 7000 9596
rect 6960 9516 7000 9564
rect 6960 9484 6964 9516
rect 6996 9484 7000 9516
rect 6960 9436 7000 9484
rect 6960 9404 6964 9436
rect 6996 9404 7000 9436
rect 6960 9356 7000 9404
rect 6960 9324 6964 9356
rect 6996 9324 7000 9356
rect 6960 9276 7000 9324
rect 6960 9244 6964 9276
rect 6996 9244 7000 9276
rect 6960 9116 7000 9244
rect 6960 9084 6964 9116
rect 6996 9084 7000 9116
rect 6960 9036 7000 9084
rect 6960 9004 6964 9036
rect 6996 9004 7000 9036
rect 6960 8956 7000 9004
rect 6960 8924 6964 8956
rect 6996 8924 7000 8956
rect 6960 8636 7000 8924
rect 6960 8604 6964 8636
rect 6996 8604 7000 8636
rect 6960 8556 7000 8604
rect 6960 8524 6964 8556
rect 6996 8524 7000 8556
rect 6960 8396 7000 8524
rect 6960 8364 6964 8396
rect 6996 8364 7000 8396
rect 6960 8316 7000 8364
rect 6960 8284 6964 8316
rect 6996 8284 7000 8316
rect 6960 8236 7000 8284
rect 6960 8204 6964 8236
rect 6996 8204 7000 8236
rect 6960 8156 7000 8204
rect 6960 8124 6964 8156
rect 6996 8124 7000 8156
rect 6960 8076 7000 8124
rect 6960 8044 6964 8076
rect 6996 8044 7000 8076
rect 6960 7996 7000 8044
rect 6960 7964 6964 7996
rect 6996 7964 7000 7996
rect 6960 7916 7000 7964
rect 6960 7884 6964 7916
rect 6996 7884 7000 7916
rect 6960 7836 7000 7884
rect 6960 7804 6964 7836
rect 6996 7804 7000 7836
rect 6960 7756 7000 7804
rect 6960 7724 6964 7756
rect 6996 7724 7000 7756
rect 6960 7676 7000 7724
rect 6960 7644 6964 7676
rect 6996 7644 7000 7676
rect 6960 7596 7000 7644
rect 6960 7564 6964 7596
rect 6996 7564 7000 7596
rect 6960 7516 7000 7564
rect 6960 7484 6964 7516
rect 6996 7484 7000 7516
rect 6960 7436 7000 7484
rect 6960 7404 6964 7436
rect 6996 7404 7000 7436
rect 6960 7356 7000 7404
rect 6960 7324 6964 7356
rect 6996 7324 7000 7356
rect 6960 7276 7000 7324
rect 6960 7244 6964 7276
rect 6996 7244 7000 7276
rect 6960 7196 7000 7244
rect 6960 7164 6964 7196
rect 6996 7164 7000 7196
rect 6960 7116 7000 7164
rect 6960 7084 6964 7116
rect 6996 7084 7000 7116
rect 6960 7036 7000 7084
rect 6960 7004 6964 7036
rect 6996 7004 7000 7036
rect 6960 6956 7000 7004
rect 6960 6924 6964 6956
rect 6996 6924 7000 6956
rect 6960 6876 7000 6924
rect 6960 6844 6964 6876
rect 6996 6844 7000 6876
rect 6960 6796 7000 6844
rect 6960 6764 6964 6796
rect 6996 6764 7000 6796
rect 6960 6716 7000 6764
rect 6960 6684 6964 6716
rect 6996 6684 7000 6716
rect 6960 6636 7000 6684
rect 6960 6604 6964 6636
rect 6996 6604 7000 6636
rect 6960 6556 7000 6604
rect 6960 6524 6964 6556
rect 6996 6524 7000 6556
rect 6960 6476 7000 6524
rect 6960 6444 6964 6476
rect 6996 6444 7000 6476
rect 6960 6396 7000 6444
rect 6960 6364 6964 6396
rect 6996 6364 7000 6396
rect 6960 6316 7000 6364
rect 6960 6284 6964 6316
rect 6996 6284 7000 6316
rect 6960 6236 7000 6284
rect 6960 6204 6964 6236
rect 6996 6204 7000 6236
rect 6960 6156 7000 6204
rect 6960 6124 6964 6156
rect 6996 6124 7000 6156
rect 6960 5996 7000 6124
rect 6960 5964 6964 5996
rect 6996 5964 7000 5996
rect 6960 5916 7000 5964
rect 6960 5884 6964 5916
rect 6996 5884 7000 5916
rect 6960 5836 7000 5884
rect 6960 5804 6964 5836
rect 6996 5804 7000 5836
rect 6960 5756 7000 5804
rect 6960 5724 6964 5756
rect 6996 5724 7000 5756
rect 6960 5676 7000 5724
rect 6960 5644 6964 5676
rect 6996 5644 7000 5676
rect 6960 5596 7000 5644
rect 6960 5564 6964 5596
rect 6996 5564 7000 5596
rect 6960 5516 7000 5564
rect 6960 5484 6964 5516
rect 6996 5484 7000 5516
rect 6960 5436 7000 5484
rect 6960 5404 6964 5436
rect 6996 5404 7000 5436
rect 6960 5356 7000 5404
rect 6960 5324 6964 5356
rect 6996 5324 7000 5356
rect 6960 5276 7000 5324
rect 6960 5244 6964 5276
rect 6996 5244 7000 5276
rect 6960 5196 7000 5244
rect 6960 5164 6964 5196
rect 6996 5164 7000 5196
rect 6960 5116 7000 5164
rect 6960 5084 6964 5116
rect 6996 5084 7000 5116
rect 6960 5036 7000 5084
rect 6960 5004 6964 5036
rect 6996 5004 7000 5036
rect 6960 4956 7000 5004
rect 6960 4924 6964 4956
rect 6996 4924 7000 4956
rect 6960 4876 7000 4924
rect 6960 4844 6964 4876
rect 6996 4844 7000 4876
rect 6960 4796 7000 4844
rect 6960 4764 6964 4796
rect 6996 4764 7000 4796
rect 6960 4716 7000 4764
rect 6960 4684 6964 4716
rect 6996 4684 7000 4716
rect 6960 4636 7000 4684
rect 6960 4604 6964 4636
rect 6996 4604 7000 4636
rect 6960 4556 7000 4604
rect 6960 4524 6964 4556
rect 6996 4524 7000 4556
rect 6960 4476 7000 4524
rect 6960 4444 6964 4476
rect 6996 4444 7000 4476
rect 6960 4396 7000 4444
rect 6960 4364 6964 4396
rect 6996 4364 7000 4396
rect 6960 4316 7000 4364
rect 6960 4284 6964 4316
rect 6996 4284 7000 4316
rect 6960 4236 7000 4284
rect 6960 4204 6964 4236
rect 6996 4204 7000 4236
rect 6960 4156 7000 4204
rect 6960 4124 6964 4156
rect 6996 4124 7000 4156
rect 6960 4076 7000 4124
rect 6960 4044 6964 4076
rect 6996 4044 7000 4076
rect 6960 3996 7000 4044
rect 6960 3964 6964 3996
rect 6996 3964 7000 3996
rect 6960 3916 7000 3964
rect 6960 3884 6964 3916
rect 6996 3884 7000 3916
rect 6960 3836 7000 3884
rect 6960 3804 6964 3836
rect 6996 3804 7000 3836
rect 6960 3756 7000 3804
rect 6960 3724 6964 3756
rect 6996 3724 7000 3756
rect 6960 3596 7000 3724
rect 6960 3564 6964 3596
rect 6996 3564 7000 3596
rect 6960 3516 7000 3564
rect 6960 3484 6964 3516
rect 6996 3484 7000 3516
rect 6960 3436 7000 3484
rect 6960 3404 6964 3436
rect 6996 3404 7000 3436
rect 6960 3356 7000 3404
rect 6960 3324 6964 3356
rect 6996 3324 7000 3356
rect 6960 3276 7000 3324
rect 6960 3244 6964 3276
rect 6996 3244 7000 3276
rect 6960 3196 7000 3244
rect 6960 3164 6964 3196
rect 6996 3164 7000 3196
rect 6960 3116 7000 3164
rect 6960 3084 6964 3116
rect 6996 3084 7000 3116
rect 6960 3036 7000 3084
rect 6960 3004 6964 3036
rect 6996 3004 7000 3036
rect 6960 2956 7000 3004
rect 6960 2924 6964 2956
rect 6996 2924 7000 2956
rect 6960 2876 7000 2924
rect 6960 2844 6964 2876
rect 6996 2844 7000 2876
rect 6960 2796 7000 2844
rect 6960 2764 6964 2796
rect 6996 2764 7000 2796
rect 6960 2716 7000 2764
rect 6960 2684 6964 2716
rect 6996 2684 7000 2716
rect 6960 2636 7000 2684
rect 6960 2604 6964 2636
rect 6996 2604 7000 2636
rect 6960 2556 7000 2604
rect 6960 2524 6964 2556
rect 6996 2524 7000 2556
rect 6960 2476 7000 2524
rect 6960 2444 6964 2476
rect 6996 2444 7000 2476
rect 6960 2396 7000 2444
rect 6960 2364 6964 2396
rect 6996 2364 7000 2396
rect 6960 2316 7000 2364
rect 6960 2284 6964 2316
rect 6996 2284 7000 2316
rect 6960 2236 7000 2284
rect 6960 2204 6964 2236
rect 6996 2204 7000 2236
rect 6960 2156 7000 2204
rect 6960 2124 6964 2156
rect 6996 2124 7000 2156
rect 6960 2076 7000 2124
rect 6960 2044 6964 2076
rect 6996 2044 7000 2076
rect 6960 1996 7000 2044
rect 6960 1964 6964 1996
rect 6996 1964 7000 1996
rect 6960 1916 7000 1964
rect 6960 1884 6964 1916
rect 6996 1884 7000 1916
rect 6960 1836 7000 1884
rect 6960 1804 6964 1836
rect 6996 1804 7000 1836
rect 6960 1756 7000 1804
rect 6960 1724 6964 1756
rect 6996 1724 7000 1756
rect 6960 1676 7000 1724
rect 6960 1644 6964 1676
rect 6996 1644 7000 1676
rect 6960 1596 7000 1644
rect 6960 1564 6964 1596
rect 6996 1564 7000 1596
rect 6960 1516 7000 1564
rect 6960 1484 6964 1516
rect 6996 1484 7000 1516
rect 6960 1436 7000 1484
rect 6960 1404 6964 1436
rect 6996 1404 7000 1436
rect 6960 1356 7000 1404
rect 6960 1324 6964 1356
rect 6996 1324 7000 1356
rect 6960 1276 7000 1324
rect 6960 1244 6964 1276
rect 6996 1244 7000 1276
rect 6960 1196 7000 1244
rect 6960 1164 6964 1196
rect 6996 1164 7000 1196
rect 6960 1116 7000 1164
rect 6960 1084 6964 1116
rect 6996 1084 7000 1116
rect 6960 1036 7000 1084
rect 6960 1004 6964 1036
rect 6996 1004 7000 1036
rect 6960 956 7000 1004
rect 6960 924 6964 956
rect 6996 924 7000 956
rect 6960 876 7000 924
rect 6960 844 6964 876
rect 6996 844 7000 876
rect 6960 796 7000 844
rect 6960 764 6964 796
rect 6996 764 7000 796
rect 6960 716 7000 764
rect 6960 684 6964 716
rect 6996 684 7000 716
rect 6960 596 7000 684
rect 6960 564 6964 596
rect 6996 564 7000 596
rect 6960 516 7000 564
rect 6960 484 6964 516
rect 6996 484 7000 516
rect 6960 436 7000 484
rect 6960 404 6964 436
rect 6996 404 7000 436
rect 6960 356 7000 404
rect 6960 324 6964 356
rect 6996 324 7000 356
rect 6960 276 7000 324
rect 6960 244 6964 276
rect 6996 244 7000 276
rect 6960 196 7000 244
rect 6960 164 6964 196
rect 6996 164 7000 196
rect 6960 116 7000 164
rect 6960 84 6964 116
rect 6996 84 7000 116
rect 6960 36 7000 84
rect 6960 4 6964 36
rect 6996 4 7000 36
rect 6960 -40 7000 4
rect 7040 14155 7080 16640
rect 7040 14125 7045 14155
rect 7075 14125 7080 14155
rect 7040 10795 7080 14125
rect 7040 10765 7045 10795
rect 7075 10765 7080 10795
rect 7040 10555 7080 10765
rect 7040 10525 7045 10555
rect 7075 10525 7080 10555
rect 7040 8475 7080 10525
rect 7040 8445 7045 8475
rect 7075 8445 7080 8475
rect 7040 6075 7080 8445
rect 7040 6045 7045 6075
rect 7075 6045 7080 6075
rect 7040 3675 7080 6045
rect 7040 3645 7045 3675
rect 7075 3645 7080 3675
rect 7040 -40 7080 3645
rect 7120 16596 7160 16644
rect 7280 16836 7320 17124
rect 7280 16644 7284 16836
rect 7316 16644 7320 16836
rect 7120 16564 7124 16596
rect 7156 16564 7160 16596
rect 7120 16516 7160 16564
rect 7120 16484 7124 16516
rect 7156 16484 7160 16516
rect 7120 16436 7160 16484
rect 7120 16404 7124 16436
rect 7156 16404 7160 16436
rect 7120 16356 7160 16404
rect 7120 16324 7124 16356
rect 7156 16324 7160 16356
rect 7120 16276 7160 16324
rect 7120 16244 7124 16276
rect 7156 16244 7160 16276
rect 7120 16196 7160 16244
rect 7120 16164 7124 16196
rect 7156 16164 7160 16196
rect 7120 16116 7160 16164
rect 7120 16084 7124 16116
rect 7156 16084 7160 16116
rect 7120 16036 7160 16084
rect 7120 16004 7124 16036
rect 7156 16004 7160 16036
rect 7120 15956 7160 16004
rect 7120 15924 7124 15956
rect 7156 15924 7160 15956
rect 7120 15436 7160 15924
rect 7120 15404 7124 15436
rect 7156 15404 7160 15436
rect 7120 15356 7160 15404
rect 7120 15324 7124 15356
rect 7156 15324 7160 15356
rect 7120 15276 7160 15324
rect 7120 15244 7124 15276
rect 7156 15244 7160 15276
rect 7120 15196 7160 15244
rect 7120 15164 7124 15196
rect 7156 15164 7160 15196
rect 7120 15116 7160 15164
rect 7120 15084 7124 15116
rect 7156 15084 7160 15116
rect 7120 15036 7160 15084
rect 7120 15004 7124 15036
rect 7156 15004 7160 15036
rect 7120 14956 7160 15004
rect 7120 14924 7124 14956
rect 7156 14924 7160 14956
rect 7120 14876 7160 14924
rect 7120 14844 7124 14876
rect 7156 14844 7160 14876
rect 7120 14796 7160 14844
rect 7120 14764 7124 14796
rect 7156 14764 7160 14796
rect 7120 14716 7160 14764
rect 7120 14684 7124 14716
rect 7156 14684 7160 14716
rect 7120 14636 7160 14684
rect 7120 14604 7124 14636
rect 7156 14604 7160 14636
rect 7120 14556 7160 14604
rect 7120 14524 7124 14556
rect 7156 14524 7160 14556
rect 7120 14476 7160 14524
rect 7120 14444 7124 14476
rect 7156 14444 7160 14476
rect 7120 14395 7160 14444
rect 7120 14365 7125 14395
rect 7155 14365 7160 14395
rect 7120 14235 7160 14365
rect 7120 14205 7125 14235
rect 7155 14205 7160 14235
rect 7120 14075 7160 14205
rect 7120 14045 7125 14075
rect 7155 14045 7160 14075
rect 7120 13996 7160 14045
rect 7120 13964 7124 13996
rect 7156 13964 7160 13996
rect 7120 13876 7160 13964
rect 7120 13844 7124 13876
rect 7156 13844 7160 13876
rect 7120 13796 7160 13844
rect 7120 13764 7124 13796
rect 7156 13764 7160 13796
rect 7120 13716 7160 13764
rect 7120 13684 7124 13716
rect 7156 13684 7160 13716
rect 7120 13636 7160 13684
rect 7120 13604 7124 13636
rect 7156 13604 7160 13636
rect 7120 13556 7160 13604
rect 7120 13524 7124 13556
rect 7156 13524 7160 13556
rect 7120 13476 7160 13524
rect 7120 13444 7124 13476
rect 7156 13444 7160 13476
rect 7120 13396 7160 13444
rect 7120 13364 7124 13396
rect 7156 13364 7160 13396
rect 7120 13316 7160 13364
rect 7120 13284 7124 13316
rect 7156 13284 7160 13316
rect 7120 13236 7160 13284
rect 7120 13204 7124 13236
rect 7156 13204 7160 13236
rect 7120 13156 7160 13204
rect 7120 13124 7124 13156
rect 7156 13124 7160 13156
rect 7120 13076 7160 13124
rect 7120 13044 7124 13076
rect 7156 13044 7160 13076
rect 7120 12996 7160 13044
rect 7120 12964 7124 12996
rect 7156 12964 7160 12996
rect 7120 12516 7160 12964
rect 7120 12484 7124 12516
rect 7156 12484 7160 12516
rect 7120 12436 7160 12484
rect 7120 12404 7124 12436
rect 7156 12404 7160 12436
rect 7120 12316 7160 12404
rect 7120 12284 7124 12316
rect 7156 12284 7160 12316
rect 7120 12236 7160 12284
rect 7120 12204 7124 12236
rect 7156 12204 7160 12236
rect 7120 12156 7160 12204
rect 7120 12124 7124 12156
rect 7156 12124 7160 12156
rect 7120 12076 7160 12124
rect 7120 12044 7124 12076
rect 7156 12044 7160 12076
rect 7120 11996 7160 12044
rect 7120 11964 7124 11996
rect 7156 11964 7160 11996
rect 7120 11916 7160 11964
rect 7120 11884 7124 11916
rect 7156 11884 7160 11916
rect 7120 11836 7160 11884
rect 7120 11804 7124 11836
rect 7156 11804 7160 11836
rect 7120 11756 7160 11804
rect 7120 11724 7124 11756
rect 7156 11724 7160 11756
rect 7120 11676 7160 11724
rect 7120 11644 7124 11676
rect 7156 11644 7160 11676
rect 7120 11596 7160 11644
rect 7120 11564 7124 11596
rect 7156 11564 7160 11596
rect 7120 11516 7160 11564
rect 7120 11484 7124 11516
rect 7156 11484 7160 11516
rect 7120 11436 7160 11484
rect 7120 11404 7124 11436
rect 7156 11404 7160 11436
rect 7120 11356 7160 11404
rect 7120 11324 7124 11356
rect 7156 11324 7160 11356
rect 7120 11196 7160 11324
rect 7120 11164 7124 11196
rect 7156 11164 7160 11196
rect 7120 11116 7160 11164
rect 7120 11084 7124 11116
rect 7156 11084 7160 11116
rect 7120 11036 7160 11084
rect 7120 11004 7124 11036
rect 7156 11004 7160 11036
rect 7120 10876 7160 11004
rect 7120 10844 7124 10876
rect 7156 10844 7160 10876
rect 7120 10796 7160 10844
rect 7120 10764 7124 10796
rect 7156 10764 7160 10796
rect 7120 10716 7160 10764
rect 7120 10684 7124 10716
rect 7156 10684 7160 10716
rect 7120 10636 7160 10684
rect 7120 10604 7124 10636
rect 7156 10604 7160 10636
rect 7120 10556 7160 10604
rect 7120 10524 7124 10556
rect 7156 10524 7160 10556
rect 7120 10476 7160 10524
rect 7120 10444 7124 10476
rect 7156 10444 7160 10476
rect 7120 10396 7160 10444
rect 7120 10364 7124 10396
rect 7156 10364 7160 10396
rect 7120 10316 7160 10364
rect 7120 10284 7124 10316
rect 7156 10284 7160 10316
rect 7120 10236 7160 10284
rect 7120 10204 7124 10236
rect 7156 10204 7160 10236
rect 7120 10156 7160 10204
rect 7120 10124 7124 10156
rect 7156 10124 7160 10156
rect 7120 10076 7160 10124
rect 7120 10044 7124 10076
rect 7156 10044 7160 10076
rect 7120 9996 7160 10044
rect 7120 9964 7124 9996
rect 7156 9964 7160 9996
rect 7120 9916 7160 9964
rect 7120 9884 7124 9916
rect 7156 9884 7160 9916
rect 7120 9836 7160 9884
rect 7120 9804 7124 9836
rect 7156 9804 7160 9836
rect 7120 9756 7160 9804
rect 7120 9724 7124 9756
rect 7156 9724 7160 9756
rect 7120 9676 7160 9724
rect 7120 9644 7124 9676
rect 7156 9644 7160 9676
rect 7120 9596 7160 9644
rect 7120 9564 7124 9596
rect 7156 9564 7160 9596
rect 7120 9516 7160 9564
rect 7120 9484 7124 9516
rect 7156 9484 7160 9516
rect 7120 9436 7160 9484
rect 7120 9404 7124 9436
rect 7156 9404 7160 9436
rect 7120 9356 7160 9404
rect 7120 9324 7124 9356
rect 7156 9324 7160 9356
rect 7120 9276 7160 9324
rect 7120 9244 7124 9276
rect 7156 9244 7160 9276
rect 7120 9116 7160 9244
rect 7120 9084 7124 9116
rect 7156 9084 7160 9116
rect 7120 9036 7160 9084
rect 7120 9004 7124 9036
rect 7156 9004 7160 9036
rect 7120 8956 7160 9004
rect 7120 8924 7124 8956
rect 7156 8924 7160 8956
rect 7120 8636 7160 8924
rect 7120 8604 7124 8636
rect 7156 8604 7160 8636
rect 7120 8556 7160 8604
rect 7120 8524 7124 8556
rect 7156 8524 7160 8556
rect 7120 8476 7160 8524
rect 7120 8444 7124 8476
rect 7156 8444 7160 8476
rect 7120 8396 7160 8444
rect 7120 8364 7124 8396
rect 7156 8364 7160 8396
rect 7120 8316 7160 8364
rect 7120 8284 7124 8316
rect 7156 8284 7160 8316
rect 7120 8236 7160 8284
rect 7120 8204 7124 8236
rect 7156 8204 7160 8236
rect 7120 8156 7160 8204
rect 7120 8124 7124 8156
rect 7156 8124 7160 8156
rect 7120 8076 7160 8124
rect 7120 8044 7124 8076
rect 7156 8044 7160 8076
rect 7120 7996 7160 8044
rect 7120 7964 7124 7996
rect 7156 7964 7160 7996
rect 7120 7916 7160 7964
rect 7120 7884 7124 7916
rect 7156 7884 7160 7916
rect 7120 7836 7160 7884
rect 7120 7804 7124 7836
rect 7156 7804 7160 7836
rect 7120 7756 7160 7804
rect 7120 7724 7124 7756
rect 7156 7724 7160 7756
rect 7120 7676 7160 7724
rect 7120 7644 7124 7676
rect 7156 7644 7160 7676
rect 7120 7596 7160 7644
rect 7120 7564 7124 7596
rect 7156 7564 7160 7596
rect 7120 7516 7160 7564
rect 7120 7484 7124 7516
rect 7156 7484 7160 7516
rect 7120 7436 7160 7484
rect 7120 7404 7124 7436
rect 7156 7404 7160 7436
rect 7120 7356 7160 7404
rect 7120 7324 7124 7356
rect 7156 7324 7160 7356
rect 7120 7276 7160 7324
rect 7120 7244 7124 7276
rect 7156 7244 7160 7276
rect 7120 7196 7160 7244
rect 7120 7164 7124 7196
rect 7156 7164 7160 7196
rect 7120 7116 7160 7164
rect 7120 7084 7124 7116
rect 7156 7084 7160 7116
rect 7120 7036 7160 7084
rect 7120 7004 7124 7036
rect 7156 7004 7160 7036
rect 7120 6956 7160 7004
rect 7120 6924 7124 6956
rect 7156 6924 7160 6956
rect 7120 6876 7160 6924
rect 7120 6844 7124 6876
rect 7156 6844 7160 6876
rect 7120 6796 7160 6844
rect 7120 6764 7124 6796
rect 7156 6764 7160 6796
rect 7120 6716 7160 6764
rect 7120 6684 7124 6716
rect 7156 6684 7160 6716
rect 7120 6636 7160 6684
rect 7120 6604 7124 6636
rect 7156 6604 7160 6636
rect 7120 6556 7160 6604
rect 7120 6524 7124 6556
rect 7156 6524 7160 6556
rect 7120 6476 7160 6524
rect 7120 6444 7124 6476
rect 7156 6444 7160 6476
rect 7120 6396 7160 6444
rect 7120 6364 7124 6396
rect 7156 6364 7160 6396
rect 7120 6316 7160 6364
rect 7120 6284 7124 6316
rect 7156 6284 7160 6316
rect 7120 6236 7160 6284
rect 7120 6204 7124 6236
rect 7156 6204 7160 6236
rect 7120 6156 7160 6204
rect 7120 6124 7124 6156
rect 7156 6124 7160 6156
rect 7120 6076 7160 6124
rect 7120 6044 7124 6076
rect 7156 6044 7160 6076
rect 7120 5996 7160 6044
rect 7120 5964 7124 5996
rect 7156 5964 7160 5996
rect 7120 5916 7160 5964
rect 7120 5884 7124 5916
rect 7156 5884 7160 5916
rect 7120 5836 7160 5884
rect 7120 5804 7124 5836
rect 7156 5804 7160 5836
rect 7120 5756 7160 5804
rect 7120 5724 7124 5756
rect 7156 5724 7160 5756
rect 7120 5676 7160 5724
rect 7120 5644 7124 5676
rect 7156 5644 7160 5676
rect 7120 5596 7160 5644
rect 7120 5564 7124 5596
rect 7156 5564 7160 5596
rect 7120 5516 7160 5564
rect 7120 5484 7124 5516
rect 7156 5484 7160 5516
rect 7120 5436 7160 5484
rect 7120 5404 7124 5436
rect 7156 5404 7160 5436
rect 7120 5356 7160 5404
rect 7120 5324 7124 5356
rect 7156 5324 7160 5356
rect 7120 5276 7160 5324
rect 7120 5244 7124 5276
rect 7156 5244 7160 5276
rect 7120 5196 7160 5244
rect 7120 5164 7124 5196
rect 7156 5164 7160 5196
rect 7120 5116 7160 5164
rect 7120 5084 7124 5116
rect 7156 5084 7160 5116
rect 7120 5036 7160 5084
rect 7120 5004 7124 5036
rect 7156 5004 7160 5036
rect 7120 4956 7160 5004
rect 7120 4924 7124 4956
rect 7156 4924 7160 4956
rect 7120 4876 7160 4924
rect 7120 4844 7124 4876
rect 7156 4844 7160 4876
rect 7120 4796 7160 4844
rect 7120 4764 7124 4796
rect 7156 4764 7160 4796
rect 7120 4716 7160 4764
rect 7120 4684 7124 4716
rect 7156 4684 7160 4716
rect 7120 4636 7160 4684
rect 7120 4604 7124 4636
rect 7156 4604 7160 4636
rect 7120 4556 7160 4604
rect 7120 4524 7124 4556
rect 7156 4524 7160 4556
rect 7120 4476 7160 4524
rect 7120 4444 7124 4476
rect 7156 4444 7160 4476
rect 7120 4396 7160 4444
rect 7120 4364 7124 4396
rect 7156 4364 7160 4396
rect 7120 4316 7160 4364
rect 7120 4284 7124 4316
rect 7156 4284 7160 4316
rect 7120 4236 7160 4284
rect 7120 4204 7124 4236
rect 7156 4204 7160 4236
rect 7120 4156 7160 4204
rect 7120 4124 7124 4156
rect 7156 4124 7160 4156
rect 7120 4076 7160 4124
rect 7120 4044 7124 4076
rect 7156 4044 7160 4076
rect 7120 3996 7160 4044
rect 7120 3964 7124 3996
rect 7156 3964 7160 3996
rect 7120 3916 7160 3964
rect 7120 3884 7124 3916
rect 7156 3884 7160 3916
rect 7120 3836 7160 3884
rect 7120 3804 7124 3836
rect 7156 3804 7160 3836
rect 7120 3756 7160 3804
rect 7120 3724 7124 3756
rect 7156 3724 7160 3756
rect 7120 3676 7160 3724
rect 7120 3644 7124 3676
rect 7156 3644 7160 3676
rect 7120 3596 7160 3644
rect 7120 3564 7124 3596
rect 7156 3564 7160 3596
rect 7120 3516 7160 3564
rect 7120 3484 7124 3516
rect 7156 3484 7160 3516
rect 7120 3436 7160 3484
rect 7120 3404 7124 3436
rect 7156 3404 7160 3436
rect 7120 3356 7160 3404
rect 7120 3324 7124 3356
rect 7156 3324 7160 3356
rect 7120 3276 7160 3324
rect 7120 3244 7124 3276
rect 7156 3244 7160 3276
rect 7120 3196 7160 3244
rect 7120 3164 7124 3196
rect 7156 3164 7160 3196
rect 7120 3116 7160 3164
rect 7120 3084 7124 3116
rect 7156 3084 7160 3116
rect 7120 3036 7160 3084
rect 7120 3004 7124 3036
rect 7156 3004 7160 3036
rect 7120 2956 7160 3004
rect 7120 2924 7124 2956
rect 7156 2924 7160 2956
rect 7120 2876 7160 2924
rect 7120 2844 7124 2876
rect 7156 2844 7160 2876
rect 7120 2796 7160 2844
rect 7120 2764 7124 2796
rect 7156 2764 7160 2796
rect 7120 2716 7160 2764
rect 7120 2684 7124 2716
rect 7156 2684 7160 2716
rect 7120 2636 7160 2684
rect 7120 2604 7124 2636
rect 7156 2604 7160 2636
rect 7120 2556 7160 2604
rect 7120 2524 7124 2556
rect 7156 2524 7160 2556
rect 7120 2476 7160 2524
rect 7120 2444 7124 2476
rect 7156 2444 7160 2476
rect 7120 2396 7160 2444
rect 7120 2364 7124 2396
rect 7156 2364 7160 2396
rect 7120 2316 7160 2364
rect 7120 2284 7124 2316
rect 7156 2284 7160 2316
rect 7120 2236 7160 2284
rect 7120 2204 7124 2236
rect 7156 2204 7160 2236
rect 7120 2156 7160 2204
rect 7120 2124 7124 2156
rect 7156 2124 7160 2156
rect 7120 2076 7160 2124
rect 7120 2044 7124 2076
rect 7156 2044 7160 2076
rect 7120 1996 7160 2044
rect 7120 1964 7124 1996
rect 7156 1964 7160 1996
rect 7120 1916 7160 1964
rect 7120 1884 7124 1916
rect 7156 1884 7160 1916
rect 7120 1836 7160 1884
rect 7120 1804 7124 1836
rect 7156 1804 7160 1836
rect 7120 1756 7160 1804
rect 7120 1724 7124 1756
rect 7156 1724 7160 1756
rect 7120 1676 7160 1724
rect 7120 1644 7124 1676
rect 7156 1644 7160 1676
rect 7120 1596 7160 1644
rect 7120 1564 7124 1596
rect 7156 1564 7160 1596
rect 7120 1516 7160 1564
rect 7120 1484 7124 1516
rect 7156 1484 7160 1516
rect 7120 1436 7160 1484
rect 7120 1404 7124 1436
rect 7156 1404 7160 1436
rect 7120 1356 7160 1404
rect 7120 1324 7124 1356
rect 7156 1324 7160 1356
rect 7120 1276 7160 1324
rect 7120 1244 7124 1276
rect 7156 1244 7160 1276
rect 7120 1196 7160 1244
rect 7120 1164 7124 1196
rect 7156 1164 7160 1196
rect 7120 1116 7160 1164
rect 7120 1084 7124 1116
rect 7156 1084 7160 1116
rect 7120 1036 7160 1084
rect 7120 1004 7124 1036
rect 7156 1004 7160 1036
rect 7120 956 7160 1004
rect 7120 924 7124 956
rect 7156 924 7160 956
rect 7120 876 7160 924
rect 7120 844 7124 876
rect 7156 844 7160 876
rect 7120 796 7160 844
rect 7120 764 7124 796
rect 7156 764 7160 796
rect 7120 716 7160 764
rect 7120 684 7124 716
rect 7156 684 7160 716
rect 7120 596 7160 684
rect 7120 564 7124 596
rect 7156 564 7160 596
rect 7120 516 7160 564
rect 7120 484 7124 516
rect 7156 484 7160 516
rect 7120 436 7160 484
rect 7120 404 7124 436
rect 7156 404 7160 436
rect 7120 356 7160 404
rect 7120 324 7124 356
rect 7156 324 7160 356
rect 7120 276 7160 324
rect 7120 244 7124 276
rect 7156 244 7160 276
rect 7120 196 7160 244
rect 7120 164 7124 196
rect 7156 164 7160 196
rect 7120 116 7160 164
rect 7120 84 7124 116
rect 7156 84 7160 116
rect 7120 36 7160 84
rect 7120 4 7124 36
rect 7156 4 7160 36
rect 7120 -40 7160 4
rect 7200 14315 7240 16640
rect 7200 14285 7205 14315
rect 7235 14285 7240 14315
rect 7200 11275 7240 14285
rect 7200 11245 7205 11275
rect 7235 11245 7240 11275
rect 7200 10955 7240 11245
rect 7200 10925 7205 10955
rect 7235 10925 7240 10955
rect 7200 9195 7240 10925
rect 7200 9165 7205 9195
rect 7235 9165 7240 9195
rect 7200 -40 7240 9165
rect 7280 16596 7320 16644
rect 7280 16564 7284 16596
rect 7316 16564 7320 16596
rect 7280 16516 7320 16564
rect 7280 16484 7284 16516
rect 7316 16484 7320 16516
rect 7280 16436 7320 16484
rect 7280 16404 7284 16436
rect 7316 16404 7320 16436
rect 7280 16356 7320 16404
rect 7280 16324 7284 16356
rect 7316 16324 7320 16356
rect 7280 16276 7320 16324
rect 7280 16244 7284 16276
rect 7316 16244 7320 16276
rect 7280 16196 7320 16244
rect 7280 16164 7284 16196
rect 7316 16164 7320 16196
rect 7280 16116 7320 16164
rect 7280 16084 7284 16116
rect 7316 16084 7320 16116
rect 7280 16036 7320 16084
rect 7280 16004 7284 16036
rect 7316 16004 7320 16036
rect 7280 15956 7320 16004
rect 7280 15924 7284 15956
rect 7316 15924 7320 15956
rect 7280 15436 7320 15924
rect 7280 15404 7284 15436
rect 7316 15404 7320 15436
rect 7280 15356 7320 15404
rect 7280 15324 7284 15356
rect 7316 15324 7320 15356
rect 7280 15276 7320 15324
rect 7280 15244 7284 15276
rect 7316 15244 7320 15276
rect 7280 15196 7320 15244
rect 7280 15164 7284 15196
rect 7316 15164 7320 15196
rect 7280 15116 7320 15164
rect 7280 15084 7284 15116
rect 7316 15084 7320 15116
rect 7280 15036 7320 15084
rect 7280 15004 7284 15036
rect 7316 15004 7320 15036
rect 7280 14956 7320 15004
rect 7280 14924 7284 14956
rect 7316 14924 7320 14956
rect 7280 14876 7320 14924
rect 7280 14844 7284 14876
rect 7316 14844 7320 14876
rect 7280 14796 7320 14844
rect 7280 14764 7284 14796
rect 7316 14764 7320 14796
rect 7280 14716 7320 14764
rect 7280 14684 7284 14716
rect 7316 14684 7320 14716
rect 7280 14636 7320 14684
rect 7280 14604 7284 14636
rect 7316 14604 7320 14636
rect 7280 14556 7320 14604
rect 7280 14524 7284 14556
rect 7316 14524 7320 14556
rect 7280 14476 7320 14524
rect 7280 14444 7284 14476
rect 7316 14444 7320 14476
rect 7280 14395 7320 14444
rect 7280 14365 7285 14395
rect 7315 14365 7320 14395
rect 7280 14235 7320 14365
rect 7280 14205 7285 14235
rect 7315 14205 7320 14235
rect 7280 14075 7320 14205
rect 7280 14045 7285 14075
rect 7315 14045 7320 14075
rect 7280 13996 7320 14045
rect 7280 13964 7284 13996
rect 7316 13964 7320 13996
rect 7280 13876 7320 13964
rect 7280 13844 7284 13876
rect 7316 13844 7320 13876
rect 7280 13796 7320 13844
rect 7280 13764 7284 13796
rect 7316 13764 7320 13796
rect 7280 13716 7320 13764
rect 7280 13684 7284 13716
rect 7316 13684 7320 13716
rect 7280 13636 7320 13684
rect 7280 13604 7284 13636
rect 7316 13604 7320 13636
rect 7280 13556 7320 13604
rect 7280 13524 7284 13556
rect 7316 13524 7320 13556
rect 7280 13476 7320 13524
rect 7280 13444 7284 13476
rect 7316 13444 7320 13476
rect 7280 13396 7320 13444
rect 7280 13364 7284 13396
rect 7316 13364 7320 13396
rect 7280 13316 7320 13364
rect 7280 13284 7284 13316
rect 7316 13284 7320 13316
rect 7280 13236 7320 13284
rect 7280 13204 7284 13236
rect 7316 13204 7320 13236
rect 7280 13156 7320 13204
rect 7280 13124 7284 13156
rect 7316 13124 7320 13156
rect 7280 13076 7320 13124
rect 7280 13044 7284 13076
rect 7316 13044 7320 13076
rect 7280 12996 7320 13044
rect 7280 12964 7284 12996
rect 7316 12964 7320 12996
rect 7280 12516 7320 12964
rect 7280 12484 7284 12516
rect 7316 12484 7320 12516
rect 7280 12436 7320 12484
rect 7280 12404 7284 12436
rect 7316 12404 7320 12436
rect 7280 12316 7320 12404
rect 7280 12284 7284 12316
rect 7316 12284 7320 12316
rect 7280 12236 7320 12284
rect 7280 12204 7284 12236
rect 7316 12204 7320 12236
rect 7280 12156 7320 12204
rect 7280 12124 7284 12156
rect 7316 12124 7320 12156
rect 7280 12076 7320 12124
rect 7280 12044 7284 12076
rect 7316 12044 7320 12076
rect 7280 11996 7320 12044
rect 7280 11964 7284 11996
rect 7316 11964 7320 11996
rect 7280 11916 7320 11964
rect 7280 11884 7284 11916
rect 7316 11884 7320 11916
rect 7280 11836 7320 11884
rect 7280 11804 7284 11836
rect 7316 11804 7320 11836
rect 7280 11756 7320 11804
rect 7280 11724 7284 11756
rect 7316 11724 7320 11756
rect 7280 11676 7320 11724
rect 7280 11644 7284 11676
rect 7316 11644 7320 11676
rect 7280 11596 7320 11644
rect 7280 11564 7284 11596
rect 7316 11564 7320 11596
rect 7280 11516 7320 11564
rect 7280 11484 7284 11516
rect 7316 11484 7320 11516
rect 7280 11436 7320 11484
rect 7280 11404 7284 11436
rect 7316 11404 7320 11436
rect 7280 11356 7320 11404
rect 7280 11324 7284 11356
rect 7316 11324 7320 11356
rect 7280 11196 7320 11324
rect 7280 11164 7284 11196
rect 7316 11164 7320 11196
rect 7280 11116 7320 11164
rect 7280 11084 7284 11116
rect 7316 11084 7320 11116
rect 7280 11036 7320 11084
rect 7280 11004 7284 11036
rect 7316 11004 7320 11036
rect 7280 10876 7320 11004
rect 7280 10844 7284 10876
rect 7316 10844 7320 10876
rect 7280 10796 7320 10844
rect 7280 10764 7284 10796
rect 7316 10764 7320 10796
rect 7280 10716 7320 10764
rect 7280 10684 7284 10716
rect 7316 10684 7320 10716
rect 7280 10636 7320 10684
rect 7280 10604 7284 10636
rect 7316 10604 7320 10636
rect 7280 10556 7320 10604
rect 7280 10524 7284 10556
rect 7316 10524 7320 10556
rect 7280 10476 7320 10524
rect 7280 10444 7284 10476
rect 7316 10444 7320 10476
rect 7280 10396 7320 10444
rect 7280 10364 7284 10396
rect 7316 10364 7320 10396
rect 7280 10316 7320 10364
rect 7280 10284 7284 10316
rect 7316 10284 7320 10316
rect 7280 10236 7320 10284
rect 7280 10204 7284 10236
rect 7316 10204 7320 10236
rect 7280 10156 7320 10204
rect 7280 10124 7284 10156
rect 7316 10124 7320 10156
rect 7280 10076 7320 10124
rect 7280 10044 7284 10076
rect 7316 10044 7320 10076
rect 7280 9996 7320 10044
rect 7280 9964 7284 9996
rect 7316 9964 7320 9996
rect 7280 9916 7320 9964
rect 7280 9884 7284 9916
rect 7316 9884 7320 9916
rect 7280 9836 7320 9884
rect 7280 9804 7284 9836
rect 7316 9804 7320 9836
rect 7280 9756 7320 9804
rect 7280 9724 7284 9756
rect 7316 9724 7320 9756
rect 7280 9676 7320 9724
rect 7280 9644 7284 9676
rect 7316 9644 7320 9676
rect 7280 9596 7320 9644
rect 7280 9564 7284 9596
rect 7316 9564 7320 9596
rect 7280 9516 7320 9564
rect 7280 9484 7284 9516
rect 7316 9484 7320 9516
rect 7280 9436 7320 9484
rect 7280 9404 7284 9436
rect 7316 9404 7320 9436
rect 7280 9356 7320 9404
rect 7280 9324 7284 9356
rect 7316 9324 7320 9356
rect 7280 9276 7320 9324
rect 7280 9244 7284 9276
rect 7316 9244 7320 9276
rect 7280 9116 7320 9244
rect 7280 9084 7284 9116
rect 7316 9084 7320 9116
rect 7280 9036 7320 9084
rect 7280 9004 7284 9036
rect 7316 9004 7320 9036
rect 7280 8956 7320 9004
rect 7280 8924 7284 8956
rect 7316 8924 7320 8956
rect 7280 8636 7320 8924
rect 7280 8604 7284 8636
rect 7316 8604 7320 8636
rect 7280 8556 7320 8604
rect 7280 8524 7284 8556
rect 7316 8524 7320 8556
rect 7280 8476 7320 8524
rect 7280 8444 7284 8476
rect 7316 8444 7320 8476
rect 7280 8396 7320 8444
rect 7280 8364 7284 8396
rect 7316 8364 7320 8396
rect 7280 8316 7320 8364
rect 7280 8284 7284 8316
rect 7316 8284 7320 8316
rect 7280 8236 7320 8284
rect 7280 8204 7284 8236
rect 7316 8204 7320 8236
rect 7280 8156 7320 8204
rect 7280 8124 7284 8156
rect 7316 8124 7320 8156
rect 7280 8076 7320 8124
rect 7280 8044 7284 8076
rect 7316 8044 7320 8076
rect 7280 7996 7320 8044
rect 7280 7964 7284 7996
rect 7316 7964 7320 7996
rect 7280 7916 7320 7964
rect 7280 7884 7284 7916
rect 7316 7884 7320 7916
rect 7280 7836 7320 7884
rect 7280 7804 7284 7836
rect 7316 7804 7320 7836
rect 7280 7756 7320 7804
rect 7280 7724 7284 7756
rect 7316 7724 7320 7756
rect 7280 7676 7320 7724
rect 7280 7644 7284 7676
rect 7316 7644 7320 7676
rect 7280 7596 7320 7644
rect 7280 7564 7284 7596
rect 7316 7564 7320 7596
rect 7280 7516 7320 7564
rect 7280 7484 7284 7516
rect 7316 7484 7320 7516
rect 7280 7436 7320 7484
rect 7280 7404 7284 7436
rect 7316 7404 7320 7436
rect 7280 7356 7320 7404
rect 7280 7324 7284 7356
rect 7316 7324 7320 7356
rect 7280 7276 7320 7324
rect 7280 7244 7284 7276
rect 7316 7244 7320 7276
rect 7280 7196 7320 7244
rect 7280 7164 7284 7196
rect 7316 7164 7320 7196
rect 7280 7116 7320 7164
rect 7280 7084 7284 7116
rect 7316 7084 7320 7116
rect 7280 7036 7320 7084
rect 7280 7004 7284 7036
rect 7316 7004 7320 7036
rect 7280 6956 7320 7004
rect 7280 6924 7284 6956
rect 7316 6924 7320 6956
rect 7280 6876 7320 6924
rect 7280 6844 7284 6876
rect 7316 6844 7320 6876
rect 7280 6796 7320 6844
rect 7280 6764 7284 6796
rect 7316 6764 7320 6796
rect 7280 6716 7320 6764
rect 7280 6684 7284 6716
rect 7316 6684 7320 6716
rect 7280 6636 7320 6684
rect 7280 6604 7284 6636
rect 7316 6604 7320 6636
rect 7280 6556 7320 6604
rect 7280 6524 7284 6556
rect 7316 6524 7320 6556
rect 7280 6476 7320 6524
rect 7280 6444 7284 6476
rect 7316 6444 7320 6476
rect 7280 6396 7320 6444
rect 7280 6364 7284 6396
rect 7316 6364 7320 6396
rect 7280 6316 7320 6364
rect 7280 6284 7284 6316
rect 7316 6284 7320 6316
rect 7280 6236 7320 6284
rect 7280 6204 7284 6236
rect 7316 6204 7320 6236
rect 7280 6156 7320 6204
rect 7280 6124 7284 6156
rect 7316 6124 7320 6156
rect 7280 6076 7320 6124
rect 7280 6044 7284 6076
rect 7316 6044 7320 6076
rect 7280 5996 7320 6044
rect 7280 5964 7284 5996
rect 7316 5964 7320 5996
rect 7280 5916 7320 5964
rect 7280 5884 7284 5916
rect 7316 5884 7320 5916
rect 7280 5836 7320 5884
rect 7280 5804 7284 5836
rect 7316 5804 7320 5836
rect 7280 5756 7320 5804
rect 7280 5724 7284 5756
rect 7316 5724 7320 5756
rect 7280 5676 7320 5724
rect 7280 5644 7284 5676
rect 7316 5644 7320 5676
rect 7280 5596 7320 5644
rect 7280 5564 7284 5596
rect 7316 5564 7320 5596
rect 7280 5516 7320 5564
rect 7280 5484 7284 5516
rect 7316 5484 7320 5516
rect 7280 5436 7320 5484
rect 7280 5404 7284 5436
rect 7316 5404 7320 5436
rect 7280 5356 7320 5404
rect 7280 5324 7284 5356
rect 7316 5324 7320 5356
rect 7280 5276 7320 5324
rect 7280 5244 7284 5276
rect 7316 5244 7320 5276
rect 7280 5196 7320 5244
rect 7280 5164 7284 5196
rect 7316 5164 7320 5196
rect 7280 5116 7320 5164
rect 7280 5084 7284 5116
rect 7316 5084 7320 5116
rect 7280 5036 7320 5084
rect 7280 5004 7284 5036
rect 7316 5004 7320 5036
rect 7280 4956 7320 5004
rect 7280 4924 7284 4956
rect 7316 4924 7320 4956
rect 7280 4876 7320 4924
rect 7280 4844 7284 4876
rect 7316 4844 7320 4876
rect 7280 4796 7320 4844
rect 7280 4764 7284 4796
rect 7316 4764 7320 4796
rect 7280 4716 7320 4764
rect 7280 4684 7284 4716
rect 7316 4684 7320 4716
rect 7280 4636 7320 4684
rect 7280 4604 7284 4636
rect 7316 4604 7320 4636
rect 7280 4556 7320 4604
rect 7280 4524 7284 4556
rect 7316 4524 7320 4556
rect 7280 4476 7320 4524
rect 7280 4444 7284 4476
rect 7316 4444 7320 4476
rect 7280 4396 7320 4444
rect 7280 4364 7284 4396
rect 7316 4364 7320 4396
rect 7280 4316 7320 4364
rect 7280 4284 7284 4316
rect 7316 4284 7320 4316
rect 7280 4236 7320 4284
rect 7280 4204 7284 4236
rect 7316 4204 7320 4236
rect 7280 4156 7320 4204
rect 7280 4124 7284 4156
rect 7316 4124 7320 4156
rect 7280 4076 7320 4124
rect 7280 4044 7284 4076
rect 7316 4044 7320 4076
rect 7280 3996 7320 4044
rect 7280 3964 7284 3996
rect 7316 3964 7320 3996
rect 7280 3916 7320 3964
rect 7280 3884 7284 3916
rect 7316 3884 7320 3916
rect 7280 3836 7320 3884
rect 7280 3804 7284 3836
rect 7316 3804 7320 3836
rect 7280 3756 7320 3804
rect 7280 3724 7284 3756
rect 7316 3724 7320 3756
rect 7280 3676 7320 3724
rect 7280 3644 7284 3676
rect 7316 3644 7320 3676
rect 7280 3596 7320 3644
rect 7280 3564 7284 3596
rect 7316 3564 7320 3596
rect 7280 3516 7320 3564
rect 7280 3484 7284 3516
rect 7316 3484 7320 3516
rect 7280 3436 7320 3484
rect 7280 3404 7284 3436
rect 7316 3404 7320 3436
rect 7280 3356 7320 3404
rect 7280 3324 7284 3356
rect 7316 3324 7320 3356
rect 7280 3276 7320 3324
rect 7280 3244 7284 3276
rect 7316 3244 7320 3276
rect 7280 3196 7320 3244
rect 7280 3164 7284 3196
rect 7316 3164 7320 3196
rect 7280 3116 7320 3164
rect 7280 3084 7284 3116
rect 7316 3084 7320 3116
rect 7280 3036 7320 3084
rect 7280 3004 7284 3036
rect 7316 3004 7320 3036
rect 7280 2956 7320 3004
rect 7280 2924 7284 2956
rect 7316 2924 7320 2956
rect 7280 2876 7320 2924
rect 7280 2844 7284 2876
rect 7316 2844 7320 2876
rect 7280 2796 7320 2844
rect 7280 2764 7284 2796
rect 7316 2764 7320 2796
rect 7280 2716 7320 2764
rect 7280 2684 7284 2716
rect 7316 2684 7320 2716
rect 7280 2636 7320 2684
rect 7280 2604 7284 2636
rect 7316 2604 7320 2636
rect 7280 2556 7320 2604
rect 7280 2524 7284 2556
rect 7316 2524 7320 2556
rect 7280 2476 7320 2524
rect 7280 2444 7284 2476
rect 7316 2444 7320 2476
rect 7280 2396 7320 2444
rect 7280 2364 7284 2396
rect 7316 2364 7320 2396
rect 7280 2316 7320 2364
rect 7280 2284 7284 2316
rect 7316 2284 7320 2316
rect 7280 2236 7320 2284
rect 7280 2204 7284 2236
rect 7316 2204 7320 2236
rect 7280 2156 7320 2204
rect 7280 2124 7284 2156
rect 7316 2124 7320 2156
rect 7280 2076 7320 2124
rect 7280 2044 7284 2076
rect 7316 2044 7320 2076
rect 7280 1996 7320 2044
rect 7280 1964 7284 1996
rect 7316 1964 7320 1996
rect 7280 1916 7320 1964
rect 7280 1884 7284 1916
rect 7316 1884 7320 1916
rect 7280 1836 7320 1884
rect 7280 1804 7284 1836
rect 7316 1804 7320 1836
rect 7280 1756 7320 1804
rect 7280 1724 7284 1756
rect 7316 1724 7320 1756
rect 7280 1676 7320 1724
rect 7280 1644 7284 1676
rect 7316 1644 7320 1676
rect 7280 1596 7320 1644
rect 7280 1564 7284 1596
rect 7316 1564 7320 1596
rect 7280 1516 7320 1564
rect 7280 1484 7284 1516
rect 7316 1484 7320 1516
rect 7280 1436 7320 1484
rect 7280 1404 7284 1436
rect 7316 1404 7320 1436
rect 7280 1356 7320 1404
rect 7280 1324 7284 1356
rect 7316 1324 7320 1356
rect 7280 1276 7320 1324
rect 7280 1244 7284 1276
rect 7316 1244 7320 1276
rect 7280 1196 7320 1244
rect 7280 1164 7284 1196
rect 7316 1164 7320 1196
rect 7280 1116 7320 1164
rect 7280 1084 7284 1116
rect 7316 1084 7320 1116
rect 7280 1036 7320 1084
rect 7280 1004 7284 1036
rect 7316 1004 7320 1036
rect 7280 956 7320 1004
rect 7280 924 7284 956
rect 7316 924 7320 956
rect 7280 876 7320 924
rect 7280 844 7284 876
rect 7316 844 7320 876
rect 7280 796 7320 844
rect 7280 764 7284 796
rect 7316 764 7320 796
rect 7280 716 7320 764
rect 7280 684 7284 716
rect 7316 684 7320 716
rect 7280 596 7320 684
rect 7280 564 7284 596
rect 7316 564 7320 596
rect 7280 516 7320 564
rect 7280 484 7284 516
rect 7316 484 7320 516
rect 7280 436 7320 484
rect 7280 404 7284 436
rect 7316 404 7320 436
rect 7280 356 7320 404
rect 7280 324 7284 356
rect 7316 324 7320 356
rect 7280 276 7320 324
rect 7280 244 7284 276
rect 7316 244 7320 276
rect 7280 196 7320 244
rect 7280 164 7284 196
rect 7316 164 7320 196
rect 7280 116 7320 164
rect 7280 84 7284 116
rect 7316 84 7320 116
rect 7280 36 7320 84
rect 7280 4 7284 36
rect 7316 4 7320 36
rect 7280 -40 7320 4
rect 7360 18516 7400 19684
rect 7520 19716 7560 19720
rect 7520 19684 7524 19716
rect 7556 19684 7560 19716
rect 7360 18484 7364 18516
rect 7396 18484 7400 18516
rect 7360 18436 7400 18484
rect 7360 18404 7364 18436
rect 7396 18404 7400 18436
rect 7360 16596 7400 18404
rect 7360 16564 7364 16596
rect 7396 16564 7400 16596
rect 7360 16516 7400 16564
rect 7360 16484 7364 16516
rect 7396 16484 7400 16516
rect 7360 16436 7400 16484
rect 7360 16404 7364 16436
rect 7396 16404 7400 16436
rect 7360 16356 7400 16404
rect 7360 16324 7364 16356
rect 7396 16324 7400 16356
rect 7360 16276 7400 16324
rect 7360 16244 7364 16276
rect 7396 16244 7400 16276
rect 7360 16196 7400 16244
rect 7360 16164 7364 16196
rect 7396 16164 7400 16196
rect 7360 16116 7400 16164
rect 7360 16084 7364 16116
rect 7396 16084 7400 16116
rect 7360 16036 7400 16084
rect 7360 16004 7364 16036
rect 7396 16004 7400 16036
rect 7360 15956 7400 16004
rect 7360 15924 7364 15956
rect 7396 15924 7400 15956
rect 7360 15875 7400 15924
rect 7360 15845 7365 15875
rect 7395 15845 7400 15875
rect 7360 15715 7400 15845
rect 7360 15685 7365 15715
rect 7395 15685 7400 15715
rect 7360 15555 7400 15685
rect 7360 15525 7365 15555
rect 7395 15525 7400 15555
rect 7360 15436 7400 15525
rect 7360 15404 7364 15436
rect 7396 15404 7400 15436
rect 7360 15356 7400 15404
rect 7360 15324 7364 15356
rect 7396 15324 7400 15356
rect 7360 15276 7400 15324
rect 7360 15244 7364 15276
rect 7396 15244 7400 15276
rect 7360 15196 7400 15244
rect 7360 15164 7364 15196
rect 7396 15164 7400 15196
rect 7360 15116 7400 15164
rect 7360 15084 7364 15116
rect 7396 15084 7400 15116
rect 7360 15036 7400 15084
rect 7360 15004 7364 15036
rect 7396 15004 7400 15036
rect 7360 14956 7400 15004
rect 7360 14924 7364 14956
rect 7396 14924 7400 14956
rect 7360 14876 7400 14924
rect 7360 14844 7364 14876
rect 7396 14844 7400 14876
rect 7360 14796 7400 14844
rect 7360 14764 7364 14796
rect 7396 14764 7400 14796
rect 7360 14716 7400 14764
rect 7360 14684 7364 14716
rect 7396 14684 7400 14716
rect 7360 14636 7400 14684
rect 7360 14604 7364 14636
rect 7396 14604 7400 14636
rect 7360 14556 7400 14604
rect 7360 14524 7364 14556
rect 7396 14524 7400 14556
rect 7360 14476 7400 14524
rect 7360 14444 7364 14476
rect 7396 14444 7400 14476
rect 7360 14396 7400 14444
rect 7360 14364 7364 14396
rect 7396 14364 7400 14396
rect 7360 14316 7400 14364
rect 7360 14284 7364 14316
rect 7396 14284 7400 14316
rect 7360 14236 7400 14284
rect 7360 14204 7364 14236
rect 7396 14204 7400 14236
rect 7360 14156 7400 14204
rect 7360 14124 7364 14156
rect 7396 14124 7400 14156
rect 7360 14076 7400 14124
rect 7360 14044 7364 14076
rect 7396 14044 7400 14076
rect 7360 13996 7400 14044
rect 7360 13964 7364 13996
rect 7396 13964 7400 13996
rect 7360 13876 7400 13964
rect 7360 13844 7364 13876
rect 7396 13844 7400 13876
rect 7360 13796 7400 13844
rect 7360 13764 7364 13796
rect 7396 13764 7400 13796
rect 7360 13716 7400 13764
rect 7360 13684 7364 13716
rect 7396 13684 7400 13716
rect 7360 13636 7400 13684
rect 7360 13604 7364 13636
rect 7396 13604 7400 13636
rect 7360 13556 7400 13604
rect 7360 13524 7364 13556
rect 7396 13524 7400 13556
rect 7360 13476 7400 13524
rect 7360 13444 7364 13476
rect 7396 13444 7400 13476
rect 7360 13396 7400 13444
rect 7360 13364 7364 13396
rect 7396 13364 7400 13396
rect 7360 13316 7400 13364
rect 7360 13284 7364 13316
rect 7396 13284 7400 13316
rect 7360 13236 7400 13284
rect 7360 13204 7364 13236
rect 7396 13204 7400 13236
rect 7360 13156 7400 13204
rect 7360 13124 7364 13156
rect 7396 13124 7400 13156
rect 7360 13076 7400 13124
rect 7360 13044 7364 13076
rect 7396 13044 7400 13076
rect 7360 12996 7400 13044
rect 7360 12964 7364 12996
rect 7396 12964 7400 12996
rect 7360 12915 7400 12964
rect 7360 12885 7365 12915
rect 7395 12885 7400 12915
rect 7360 12755 7400 12885
rect 7360 12725 7365 12755
rect 7395 12725 7400 12755
rect 7360 12595 7400 12725
rect 7360 12565 7365 12595
rect 7395 12565 7400 12595
rect 7360 12476 7400 12565
rect 7360 12444 7364 12476
rect 7396 12444 7400 12476
rect 7360 12396 7400 12444
rect 7360 12364 7364 12396
rect 7396 12364 7400 12396
rect 7360 12316 7400 12364
rect 7360 12284 7364 12316
rect 7396 12284 7400 12316
rect 7360 12236 7400 12284
rect 7360 12204 7364 12236
rect 7396 12204 7400 12236
rect 7360 12156 7400 12204
rect 7360 12124 7364 12156
rect 7396 12124 7400 12156
rect 7360 12076 7400 12124
rect 7360 12044 7364 12076
rect 7396 12044 7400 12076
rect 7360 11996 7400 12044
rect 7360 11964 7364 11996
rect 7396 11964 7400 11996
rect 7360 11916 7400 11964
rect 7360 11884 7364 11916
rect 7396 11884 7400 11916
rect 7360 11836 7400 11884
rect 7360 11804 7364 11836
rect 7396 11804 7400 11836
rect 7360 11756 7400 11804
rect 7360 11724 7364 11756
rect 7396 11724 7400 11756
rect 7360 11676 7400 11724
rect 7360 11644 7364 11676
rect 7396 11644 7400 11676
rect 7360 11596 7400 11644
rect 7360 11564 7364 11596
rect 7396 11564 7400 11596
rect 7360 11516 7400 11564
rect 7360 11484 7364 11516
rect 7396 11484 7400 11516
rect 7360 11436 7400 11484
rect 7360 11404 7364 11436
rect 7396 11404 7400 11436
rect 7360 11356 7400 11404
rect 7360 11324 7364 11356
rect 7396 11324 7400 11356
rect 7360 11276 7400 11324
rect 7360 11244 7364 11276
rect 7396 11244 7400 11276
rect 7360 11196 7400 11244
rect 7360 11164 7364 11196
rect 7396 11164 7400 11196
rect 7360 11116 7400 11164
rect 7360 11084 7364 11116
rect 7396 11084 7400 11116
rect 7360 11036 7400 11084
rect 7360 11004 7364 11036
rect 7396 11004 7400 11036
rect 7360 10956 7400 11004
rect 7360 10924 7364 10956
rect 7396 10924 7400 10956
rect 7360 10876 7400 10924
rect 7360 10844 7364 10876
rect 7396 10844 7400 10876
rect 7360 10796 7400 10844
rect 7360 10764 7364 10796
rect 7396 10764 7400 10796
rect 7360 10716 7400 10764
rect 7360 10684 7364 10716
rect 7396 10684 7400 10716
rect 7360 10636 7400 10684
rect 7360 10604 7364 10636
rect 7396 10604 7400 10636
rect 7360 10556 7400 10604
rect 7360 10524 7364 10556
rect 7396 10524 7400 10556
rect 7360 10476 7400 10524
rect 7360 10444 7364 10476
rect 7396 10444 7400 10476
rect 7360 10396 7400 10444
rect 7360 10364 7364 10396
rect 7396 10364 7400 10396
rect 7360 10316 7400 10364
rect 7360 10284 7364 10316
rect 7396 10284 7400 10316
rect 7360 10236 7400 10284
rect 7360 10204 7364 10236
rect 7396 10204 7400 10236
rect 7360 10156 7400 10204
rect 7360 10124 7364 10156
rect 7396 10124 7400 10156
rect 7360 10076 7400 10124
rect 7360 10044 7364 10076
rect 7396 10044 7400 10076
rect 7360 9996 7400 10044
rect 7360 9964 7364 9996
rect 7396 9964 7400 9996
rect 7360 9916 7400 9964
rect 7360 9884 7364 9916
rect 7396 9884 7400 9916
rect 7360 9836 7400 9884
rect 7360 9804 7364 9836
rect 7396 9804 7400 9836
rect 7360 9756 7400 9804
rect 7360 9724 7364 9756
rect 7396 9724 7400 9756
rect 7360 9676 7400 9724
rect 7360 9644 7364 9676
rect 7396 9644 7400 9676
rect 7360 9596 7400 9644
rect 7360 9564 7364 9596
rect 7396 9564 7400 9596
rect 7360 9516 7400 9564
rect 7360 9484 7364 9516
rect 7396 9484 7400 9516
rect 7360 9436 7400 9484
rect 7360 9404 7364 9436
rect 7396 9404 7400 9436
rect 7360 9356 7400 9404
rect 7360 9324 7364 9356
rect 7396 9324 7400 9356
rect 7360 9276 7400 9324
rect 7360 9244 7364 9276
rect 7396 9244 7400 9276
rect 7360 9196 7400 9244
rect 7360 9164 7364 9196
rect 7396 9164 7400 9196
rect 7360 9116 7400 9164
rect 7360 9084 7364 9116
rect 7396 9084 7400 9116
rect 7360 9036 7400 9084
rect 7360 9004 7364 9036
rect 7396 9004 7400 9036
rect 7360 8956 7400 9004
rect 7360 8924 7364 8956
rect 7396 8924 7400 8956
rect 7360 8795 7400 8924
rect 7360 8765 7365 8795
rect 7395 8765 7400 8795
rect 7360 8636 7400 8765
rect 7360 8604 7364 8636
rect 7396 8604 7400 8636
rect 7360 8556 7400 8604
rect 7360 8524 7364 8556
rect 7396 8524 7400 8556
rect 7360 8476 7400 8524
rect 7360 8444 7364 8476
rect 7396 8444 7400 8476
rect 7360 8396 7400 8444
rect 7360 8364 7364 8396
rect 7396 8364 7400 8396
rect 7360 8316 7400 8364
rect 7360 8284 7364 8316
rect 7396 8284 7400 8316
rect 7360 8236 7400 8284
rect 7360 8204 7364 8236
rect 7396 8204 7400 8236
rect 7360 8156 7400 8204
rect 7360 8124 7364 8156
rect 7396 8124 7400 8156
rect 7360 8076 7400 8124
rect 7360 8044 7364 8076
rect 7396 8044 7400 8076
rect 7360 7996 7400 8044
rect 7360 7964 7364 7996
rect 7396 7964 7400 7996
rect 7360 7916 7400 7964
rect 7360 7884 7364 7916
rect 7396 7884 7400 7916
rect 7360 7836 7400 7884
rect 7360 7804 7364 7836
rect 7396 7804 7400 7836
rect 7360 7756 7400 7804
rect 7360 7724 7364 7756
rect 7396 7724 7400 7756
rect 7360 7676 7400 7724
rect 7360 7644 7364 7676
rect 7396 7644 7400 7676
rect 7360 7596 7400 7644
rect 7360 7564 7364 7596
rect 7396 7564 7400 7596
rect 7360 7516 7400 7564
rect 7360 7484 7364 7516
rect 7396 7484 7400 7516
rect 7360 7436 7400 7484
rect 7360 7404 7364 7436
rect 7396 7404 7400 7436
rect 7360 7356 7400 7404
rect 7360 7324 7364 7356
rect 7396 7324 7400 7356
rect 7360 7276 7400 7324
rect 7360 7244 7364 7276
rect 7396 7244 7400 7276
rect 7360 7196 7400 7244
rect 7360 7164 7364 7196
rect 7396 7164 7400 7196
rect 7360 7116 7400 7164
rect 7360 7084 7364 7116
rect 7396 7084 7400 7116
rect 7360 7036 7400 7084
rect 7360 7004 7364 7036
rect 7396 7004 7400 7036
rect 7360 6956 7400 7004
rect 7360 6924 7364 6956
rect 7396 6924 7400 6956
rect 7360 6876 7400 6924
rect 7360 6844 7364 6876
rect 7396 6844 7400 6876
rect 7360 6796 7400 6844
rect 7360 6764 7364 6796
rect 7396 6764 7400 6796
rect 7360 6716 7400 6764
rect 7360 6684 7364 6716
rect 7396 6684 7400 6716
rect 7360 6636 7400 6684
rect 7360 6604 7364 6636
rect 7396 6604 7400 6636
rect 7360 6556 7400 6604
rect 7360 6524 7364 6556
rect 7396 6524 7400 6556
rect 7360 6476 7400 6524
rect 7360 6444 7364 6476
rect 7396 6444 7400 6476
rect 7360 6396 7400 6444
rect 7360 6364 7364 6396
rect 7396 6364 7400 6396
rect 7360 6316 7400 6364
rect 7360 6284 7364 6316
rect 7396 6284 7400 6316
rect 7360 6236 7400 6284
rect 7360 6204 7364 6236
rect 7396 6204 7400 6236
rect 7360 6156 7400 6204
rect 7360 6124 7364 6156
rect 7396 6124 7400 6156
rect 7360 6076 7400 6124
rect 7360 6044 7364 6076
rect 7396 6044 7400 6076
rect 7360 5996 7400 6044
rect 7360 5964 7364 5996
rect 7396 5964 7400 5996
rect 7360 5916 7400 5964
rect 7360 5884 7364 5916
rect 7396 5884 7400 5916
rect 7360 5836 7400 5884
rect 7360 5804 7364 5836
rect 7396 5804 7400 5836
rect 7360 5756 7400 5804
rect 7360 5724 7364 5756
rect 7396 5724 7400 5756
rect 7360 5676 7400 5724
rect 7360 5644 7364 5676
rect 7396 5644 7400 5676
rect 7360 5596 7400 5644
rect 7360 5564 7364 5596
rect 7396 5564 7400 5596
rect 7360 5516 7400 5564
rect 7360 5484 7364 5516
rect 7396 5484 7400 5516
rect 7360 5436 7400 5484
rect 7360 5404 7364 5436
rect 7396 5404 7400 5436
rect 7360 5356 7400 5404
rect 7360 5324 7364 5356
rect 7396 5324 7400 5356
rect 7360 5276 7400 5324
rect 7360 5244 7364 5276
rect 7396 5244 7400 5276
rect 7360 5196 7400 5244
rect 7360 5164 7364 5196
rect 7396 5164 7400 5196
rect 7360 5116 7400 5164
rect 7360 5084 7364 5116
rect 7396 5084 7400 5116
rect 7360 5036 7400 5084
rect 7360 5004 7364 5036
rect 7396 5004 7400 5036
rect 7360 4956 7400 5004
rect 7360 4924 7364 4956
rect 7396 4924 7400 4956
rect 7360 4876 7400 4924
rect 7360 4844 7364 4876
rect 7396 4844 7400 4876
rect 7360 4796 7400 4844
rect 7360 4764 7364 4796
rect 7396 4764 7400 4796
rect 7360 4716 7400 4764
rect 7360 4684 7364 4716
rect 7396 4684 7400 4716
rect 7360 4636 7400 4684
rect 7360 4604 7364 4636
rect 7396 4604 7400 4636
rect 7360 4556 7400 4604
rect 7360 4524 7364 4556
rect 7396 4524 7400 4556
rect 7360 4476 7400 4524
rect 7360 4444 7364 4476
rect 7396 4444 7400 4476
rect 7360 4396 7400 4444
rect 7360 4364 7364 4396
rect 7396 4364 7400 4396
rect 7360 4316 7400 4364
rect 7360 4284 7364 4316
rect 7396 4284 7400 4316
rect 7360 4236 7400 4284
rect 7360 4204 7364 4236
rect 7396 4204 7400 4236
rect 7360 4156 7400 4204
rect 7360 4124 7364 4156
rect 7396 4124 7400 4156
rect 7360 4076 7400 4124
rect 7360 4044 7364 4076
rect 7396 4044 7400 4076
rect 7360 3996 7400 4044
rect 7360 3964 7364 3996
rect 7396 3964 7400 3996
rect 7360 3916 7400 3964
rect 7360 3884 7364 3916
rect 7396 3884 7400 3916
rect 7360 3836 7400 3884
rect 7360 3804 7364 3836
rect 7396 3804 7400 3836
rect 7360 3756 7400 3804
rect 7360 3724 7364 3756
rect 7396 3724 7400 3756
rect 7360 3676 7400 3724
rect 7360 3644 7364 3676
rect 7396 3644 7400 3676
rect 7360 3596 7400 3644
rect 7360 3564 7364 3596
rect 7396 3564 7400 3596
rect 7360 3516 7400 3564
rect 7360 3484 7364 3516
rect 7396 3484 7400 3516
rect 7360 3436 7400 3484
rect 7360 3404 7364 3436
rect 7396 3404 7400 3436
rect 7360 3356 7400 3404
rect 7360 3324 7364 3356
rect 7396 3324 7400 3356
rect 7360 3276 7400 3324
rect 7360 3244 7364 3276
rect 7396 3244 7400 3276
rect 7360 3196 7400 3244
rect 7360 3164 7364 3196
rect 7396 3164 7400 3196
rect 7360 3116 7400 3164
rect 7360 3084 7364 3116
rect 7396 3084 7400 3116
rect 7360 3036 7400 3084
rect 7360 3004 7364 3036
rect 7396 3004 7400 3036
rect 7360 2956 7400 3004
rect 7360 2924 7364 2956
rect 7396 2924 7400 2956
rect 7360 2876 7400 2924
rect 7360 2844 7364 2876
rect 7396 2844 7400 2876
rect 7360 2796 7400 2844
rect 7360 2764 7364 2796
rect 7396 2764 7400 2796
rect 7360 2716 7400 2764
rect 7360 2684 7364 2716
rect 7396 2684 7400 2716
rect 7360 2636 7400 2684
rect 7360 2604 7364 2636
rect 7396 2604 7400 2636
rect 7360 2556 7400 2604
rect 7360 2524 7364 2556
rect 7396 2524 7400 2556
rect 7360 2476 7400 2524
rect 7360 2444 7364 2476
rect 7396 2444 7400 2476
rect 7360 2396 7400 2444
rect 7360 2364 7364 2396
rect 7396 2364 7400 2396
rect 7360 2316 7400 2364
rect 7360 2284 7364 2316
rect 7396 2284 7400 2316
rect 7360 2236 7400 2284
rect 7360 2204 7364 2236
rect 7396 2204 7400 2236
rect 7360 2156 7400 2204
rect 7360 2124 7364 2156
rect 7396 2124 7400 2156
rect 7360 2076 7400 2124
rect 7360 2044 7364 2076
rect 7396 2044 7400 2076
rect 7360 1996 7400 2044
rect 7360 1964 7364 1996
rect 7396 1964 7400 1996
rect 7360 1916 7400 1964
rect 7360 1884 7364 1916
rect 7396 1884 7400 1916
rect 7360 1836 7400 1884
rect 7360 1804 7364 1836
rect 7396 1804 7400 1836
rect 7360 1756 7400 1804
rect 7360 1724 7364 1756
rect 7396 1724 7400 1756
rect 7360 1676 7400 1724
rect 7360 1644 7364 1676
rect 7396 1644 7400 1676
rect 7360 1596 7400 1644
rect 7360 1564 7364 1596
rect 7396 1564 7400 1596
rect 7360 1516 7400 1564
rect 7360 1484 7364 1516
rect 7396 1484 7400 1516
rect 7360 1436 7400 1484
rect 7360 1404 7364 1436
rect 7396 1404 7400 1436
rect 7360 1356 7400 1404
rect 7360 1324 7364 1356
rect 7396 1324 7400 1356
rect 7360 1276 7400 1324
rect 7360 1244 7364 1276
rect 7396 1244 7400 1276
rect 7360 1196 7400 1244
rect 7360 1164 7364 1196
rect 7396 1164 7400 1196
rect 7360 1116 7400 1164
rect 7360 1084 7364 1116
rect 7396 1084 7400 1116
rect 7360 1036 7400 1084
rect 7360 1004 7364 1036
rect 7396 1004 7400 1036
rect 7360 956 7400 1004
rect 7360 924 7364 956
rect 7396 924 7400 956
rect 7360 876 7400 924
rect 7360 844 7364 876
rect 7396 844 7400 876
rect 7360 796 7400 844
rect 7360 764 7364 796
rect 7396 764 7400 796
rect 7360 716 7400 764
rect 7360 684 7364 716
rect 7396 684 7400 716
rect 7360 596 7400 684
rect 7360 564 7364 596
rect 7396 564 7400 596
rect 7360 516 7400 564
rect 7360 484 7364 516
rect 7396 484 7400 516
rect 7360 436 7400 484
rect 7360 404 7364 436
rect 7396 404 7400 436
rect 7360 356 7400 404
rect 7360 324 7364 356
rect 7396 324 7400 356
rect 7360 276 7400 324
rect 7360 244 7364 276
rect 7396 244 7400 276
rect 7360 196 7400 244
rect 7360 164 7364 196
rect 7396 164 7400 196
rect 7360 116 7400 164
rect 7360 84 7364 116
rect 7396 84 7400 116
rect 7360 36 7400 84
rect 7360 4 7364 36
rect 7396 4 7400 36
rect 7360 -40 7400 4
rect 7440 19636 7480 19640
rect 7440 19604 7444 19636
rect 7476 19604 7480 19636
rect 7440 15635 7480 19604
rect 7520 18516 7560 19684
rect 7520 18484 7524 18516
rect 7556 18484 7560 18516
rect 7520 18480 7560 18484
rect 7520 18436 7560 18440
rect 7520 18404 7524 18436
rect 7556 18404 7560 18436
rect 7520 17200 7560 18404
rect 7600 17400 7640 19720
rect 7680 19716 7720 19720
rect 7680 19684 7684 19716
rect 7716 19684 7720 19716
rect 7680 18516 7720 19684
rect 7680 18484 7684 18516
rect 7716 18484 7720 18516
rect 7680 18480 7720 18484
rect 7760 18480 7800 19680
rect 7680 18436 7720 18440
rect 7680 18404 7684 18436
rect 7716 18404 7720 18436
rect 7600 17316 7640 17320
rect 7600 17284 7604 17316
rect 7636 17284 7640 17316
rect 7520 16640 7560 17080
rect 7440 15605 7445 15635
rect 7475 15605 7480 15635
rect 7440 12675 7480 15605
rect 7440 12645 7445 12675
rect 7475 12645 7480 12675
rect 7440 8715 7480 12645
rect 7440 8685 7445 8715
rect 7475 8685 7480 8715
rect 7440 -40 7480 8685
rect 7520 16596 7560 16600
rect 7520 16564 7524 16596
rect 7556 16564 7560 16596
rect 7520 16516 7560 16564
rect 7520 16484 7524 16516
rect 7556 16484 7560 16516
rect 7520 16436 7560 16484
rect 7520 16404 7524 16436
rect 7556 16404 7560 16436
rect 7520 16356 7560 16404
rect 7520 16324 7524 16356
rect 7556 16324 7560 16356
rect 7520 16276 7560 16324
rect 7520 16244 7524 16276
rect 7556 16244 7560 16276
rect 7520 16196 7560 16244
rect 7520 16164 7524 16196
rect 7556 16164 7560 16196
rect 7520 16116 7560 16164
rect 7520 16084 7524 16116
rect 7556 16084 7560 16116
rect 7520 16036 7560 16084
rect 7520 16004 7524 16036
rect 7556 16004 7560 16036
rect 7520 15956 7560 16004
rect 7520 15924 7524 15956
rect 7556 15924 7560 15956
rect 7520 15875 7560 15924
rect 7520 15845 7525 15875
rect 7555 15845 7560 15875
rect 7520 15715 7560 15845
rect 7520 15685 7525 15715
rect 7555 15685 7560 15715
rect 7520 15555 7560 15685
rect 7520 15525 7525 15555
rect 7555 15525 7560 15555
rect 7520 15436 7560 15525
rect 7520 15404 7524 15436
rect 7556 15404 7560 15436
rect 7520 15356 7560 15404
rect 7520 15324 7524 15356
rect 7556 15324 7560 15356
rect 7520 15276 7560 15324
rect 7520 15244 7524 15276
rect 7556 15244 7560 15276
rect 7520 15196 7560 15244
rect 7520 15164 7524 15196
rect 7556 15164 7560 15196
rect 7520 15116 7560 15164
rect 7520 15084 7524 15116
rect 7556 15084 7560 15116
rect 7520 15036 7560 15084
rect 7520 15004 7524 15036
rect 7556 15004 7560 15036
rect 7520 14956 7560 15004
rect 7520 14924 7524 14956
rect 7556 14924 7560 14956
rect 7520 14876 7560 14924
rect 7520 14844 7524 14876
rect 7556 14844 7560 14876
rect 7520 14796 7560 14844
rect 7520 14764 7524 14796
rect 7556 14764 7560 14796
rect 7520 14716 7560 14764
rect 7520 14684 7524 14716
rect 7556 14684 7560 14716
rect 7520 14636 7560 14684
rect 7520 14604 7524 14636
rect 7556 14604 7560 14636
rect 7520 14556 7560 14604
rect 7520 14524 7524 14556
rect 7556 14524 7560 14556
rect 7520 14476 7560 14524
rect 7520 14444 7524 14476
rect 7556 14444 7560 14476
rect 7520 14396 7560 14444
rect 7520 14364 7524 14396
rect 7556 14364 7560 14396
rect 7520 14316 7560 14364
rect 7520 14284 7524 14316
rect 7556 14284 7560 14316
rect 7520 14236 7560 14284
rect 7520 14204 7524 14236
rect 7556 14204 7560 14236
rect 7520 14156 7560 14204
rect 7520 14124 7524 14156
rect 7556 14124 7560 14156
rect 7520 14076 7560 14124
rect 7520 14044 7524 14076
rect 7556 14044 7560 14076
rect 7520 13996 7560 14044
rect 7520 13964 7524 13996
rect 7556 13964 7560 13996
rect 7520 13876 7560 13964
rect 7520 13844 7524 13876
rect 7556 13844 7560 13876
rect 7520 13796 7560 13844
rect 7520 13764 7524 13796
rect 7556 13764 7560 13796
rect 7520 13716 7560 13764
rect 7520 13684 7524 13716
rect 7556 13684 7560 13716
rect 7520 13636 7560 13684
rect 7520 13604 7524 13636
rect 7556 13604 7560 13636
rect 7520 13556 7560 13604
rect 7520 13524 7524 13556
rect 7556 13524 7560 13556
rect 7520 13476 7560 13524
rect 7520 13444 7524 13476
rect 7556 13444 7560 13476
rect 7520 13396 7560 13444
rect 7520 13364 7524 13396
rect 7556 13364 7560 13396
rect 7520 13316 7560 13364
rect 7520 13284 7524 13316
rect 7556 13284 7560 13316
rect 7520 13236 7560 13284
rect 7520 13204 7524 13236
rect 7556 13204 7560 13236
rect 7520 13156 7560 13204
rect 7520 13124 7524 13156
rect 7556 13124 7560 13156
rect 7520 13076 7560 13124
rect 7520 13044 7524 13076
rect 7556 13044 7560 13076
rect 7520 12996 7560 13044
rect 7520 12964 7524 12996
rect 7556 12964 7560 12996
rect 7520 12915 7560 12964
rect 7520 12885 7525 12915
rect 7555 12885 7560 12915
rect 7520 12755 7560 12885
rect 7520 12725 7525 12755
rect 7555 12725 7560 12755
rect 7520 12595 7560 12725
rect 7520 12565 7525 12595
rect 7555 12565 7560 12595
rect 7520 12476 7560 12565
rect 7520 12444 7524 12476
rect 7556 12444 7560 12476
rect 7520 12396 7560 12444
rect 7520 12364 7524 12396
rect 7556 12364 7560 12396
rect 7520 12316 7560 12364
rect 7520 12284 7524 12316
rect 7556 12284 7560 12316
rect 7520 12236 7560 12284
rect 7520 12204 7524 12236
rect 7556 12204 7560 12236
rect 7520 12156 7560 12204
rect 7520 12124 7524 12156
rect 7556 12124 7560 12156
rect 7520 12076 7560 12124
rect 7520 12044 7524 12076
rect 7556 12044 7560 12076
rect 7520 11996 7560 12044
rect 7520 11964 7524 11996
rect 7556 11964 7560 11996
rect 7520 11916 7560 11964
rect 7520 11884 7524 11916
rect 7556 11884 7560 11916
rect 7520 11836 7560 11884
rect 7520 11804 7524 11836
rect 7556 11804 7560 11836
rect 7520 11756 7560 11804
rect 7520 11724 7524 11756
rect 7556 11724 7560 11756
rect 7520 11676 7560 11724
rect 7520 11644 7524 11676
rect 7556 11644 7560 11676
rect 7520 11596 7560 11644
rect 7520 11564 7524 11596
rect 7556 11564 7560 11596
rect 7520 11516 7560 11564
rect 7520 11484 7524 11516
rect 7556 11484 7560 11516
rect 7520 11436 7560 11484
rect 7520 11404 7524 11436
rect 7556 11404 7560 11436
rect 7520 11356 7560 11404
rect 7520 11324 7524 11356
rect 7556 11324 7560 11356
rect 7520 11276 7560 11324
rect 7520 11244 7524 11276
rect 7556 11244 7560 11276
rect 7520 11196 7560 11244
rect 7520 11164 7524 11196
rect 7556 11164 7560 11196
rect 7520 11116 7560 11164
rect 7520 11084 7524 11116
rect 7556 11084 7560 11116
rect 7520 11036 7560 11084
rect 7520 11004 7524 11036
rect 7556 11004 7560 11036
rect 7520 10956 7560 11004
rect 7520 10924 7524 10956
rect 7556 10924 7560 10956
rect 7520 10876 7560 10924
rect 7520 10844 7524 10876
rect 7556 10844 7560 10876
rect 7520 10796 7560 10844
rect 7520 10764 7524 10796
rect 7556 10764 7560 10796
rect 7520 10716 7560 10764
rect 7520 10684 7524 10716
rect 7556 10684 7560 10716
rect 7520 10636 7560 10684
rect 7520 10604 7524 10636
rect 7556 10604 7560 10636
rect 7520 10556 7560 10604
rect 7520 10524 7524 10556
rect 7556 10524 7560 10556
rect 7520 10476 7560 10524
rect 7520 10444 7524 10476
rect 7556 10444 7560 10476
rect 7520 10396 7560 10444
rect 7520 10364 7524 10396
rect 7556 10364 7560 10396
rect 7520 10316 7560 10364
rect 7520 10284 7524 10316
rect 7556 10284 7560 10316
rect 7520 10236 7560 10284
rect 7520 10204 7524 10236
rect 7556 10204 7560 10236
rect 7520 10156 7560 10204
rect 7520 10124 7524 10156
rect 7556 10124 7560 10156
rect 7520 10076 7560 10124
rect 7520 10044 7524 10076
rect 7556 10044 7560 10076
rect 7520 9996 7560 10044
rect 7520 9964 7524 9996
rect 7556 9964 7560 9996
rect 7520 9916 7560 9964
rect 7520 9884 7524 9916
rect 7556 9884 7560 9916
rect 7520 9836 7560 9884
rect 7520 9804 7524 9836
rect 7556 9804 7560 9836
rect 7520 9756 7560 9804
rect 7520 9724 7524 9756
rect 7556 9724 7560 9756
rect 7520 9676 7560 9724
rect 7520 9644 7524 9676
rect 7556 9644 7560 9676
rect 7520 9596 7560 9644
rect 7520 9564 7524 9596
rect 7556 9564 7560 9596
rect 7520 9516 7560 9564
rect 7520 9484 7524 9516
rect 7556 9484 7560 9516
rect 7520 9436 7560 9484
rect 7520 9404 7524 9436
rect 7556 9404 7560 9436
rect 7520 9356 7560 9404
rect 7520 9324 7524 9356
rect 7556 9324 7560 9356
rect 7520 9276 7560 9324
rect 7520 9244 7524 9276
rect 7556 9244 7560 9276
rect 7520 9196 7560 9244
rect 7520 9164 7524 9196
rect 7556 9164 7560 9196
rect 7520 9116 7560 9164
rect 7520 9084 7524 9116
rect 7556 9084 7560 9116
rect 7520 9036 7560 9084
rect 7520 9004 7524 9036
rect 7556 9004 7560 9036
rect 7520 8956 7560 9004
rect 7520 8924 7524 8956
rect 7556 8924 7560 8956
rect 7520 8795 7560 8924
rect 7520 8765 7525 8795
rect 7555 8765 7560 8795
rect 7520 8636 7560 8765
rect 7520 8604 7524 8636
rect 7556 8604 7560 8636
rect 7520 8556 7560 8604
rect 7520 8524 7524 8556
rect 7556 8524 7560 8556
rect 7520 8476 7560 8524
rect 7520 8444 7524 8476
rect 7556 8444 7560 8476
rect 7520 8396 7560 8444
rect 7520 8364 7524 8396
rect 7556 8364 7560 8396
rect 7520 8316 7560 8364
rect 7520 8284 7524 8316
rect 7556 8284 7560 8316
rect 7520 8236 7560 8284
rect 7520 8204 7524 8236
rect 7556 8204 7560 8236
rect 7520 8156 7560 8204
rect 7520 8124 7524 8156
rect 7556 8124 7560 8156
rect 7520 8076 7560 8124
rect 7520 8044 7524 8076
rect 7556 8044 7560 8076
rect 7520 7996 7560 8044
rect 7520 7964 7524 7996
rect 7556 7964 7560 7996
rect 7520 7916 7560 7964
rect 7520 7884 7524 7916
rect 7556 7884 7560 7916
rect 7520 7836 7560 7884
rect 7520 7804 7524 7836
rect 7556 7804 7560 7836
rect 7520 7756 7560 7804
rect 7520 7724 7524 7756
rect 7556 7724 7560 7756
rect 7520 7676 7560 7724
rect 7520 7644 7524 7676
rect 7556 7644 7560 7676
rect 7520 7596 7560 7644
rect 7520 7564 7524 7596
rect 7556 7564 7560 7596
rect 7520 7516 7560 7564
rect 7520 7484 7524 7516
rect 7556 7484 7560 7516
rect 7520 7436 7560 7484
rect 7520 7404 7524 7436
rect 7556 7404 7560 7436
rect 7520 7356 7560 7404
rect 7520 7324 7524 7356
rect 7556 7324 7560 7356
rect 7520 7276 7560 7324
rect 7520 7244 7524 7276
rect 7556 7244 7560 7276
rect 7520 7196 7560 7244
rect 7520 7164 7524 7196
rect 7556 7164 7560 7196
rect 7520 7116 7560 7164
rect 7520 7084 7524 7116
rect 7556 7084 7560 7116
rect 7520 7036 7560 7084
rect 7520 7004 7524 7036
rect 7556 7004 7560 7036
rect 7520 6956 7560 7004
rect 7520 6924 7524 6956
rect 7556 6924 7560 6956
rect 7520 6876 7560 6924
rect 7520 6844 7524 6876
rect 7556 6844 7560 6876
rect 7520 6796 7560 6844
rect 7520 6764 7524 6796
rect 7556 6764 7560 6796
rect 7520 6716 7560 6764
rect 7520 6684 7524 6716
rect 7556 6684 7560 6716
rect 7520 6636 7560 6684
rect 7520 6604 7524 6636
rect 7556 6604 7560 6636
rect 7520 6556 7560 6604
rect 7520 6524 7524 6556
rect 7556 6524 7560 6556
rect 7520 6476 7560 6524
rect 7520 6444 7524 6476
rect 7556 6444 7560 6476
rect 7520 6396 7560 6444
rect 7520 6364 7524 6396
rect 7556 6364 7560 6396
rect 7520 6316 7560 6364
rect 7520 6284 7524 6316
rect 7556 6284 7560 6316
rect 7520 6236 7560 6284
rect 7520 6204 7524 6236
rect 7556 6204 7560 6236
rect 7520 6156 7560 6204
rect 7520 6124 7524 6156
rect 7556 6124 7560 6156
rect 7520 6076 7560 6124
rect 7520 6044 7524 6076
rect 7556 6044 7560 6076
rect 7520 5996 7560 6044
rect 7520 5964 7524 5996
rect 7556 5964 7560 5996
rect 7520 5916 7560 5964
rect 7520 5884 7524 5916
rect 7556 5884 7560 5916
rect 7520 5836 7560 5884
rect 7520 5804 7524 5836
rect 7556 5804 7560 5836
rect 7520 5756 7560 5804
rect 7520 5724 7524 5756
rect 7556 5724 7560 5756
rect 7520 5676 7560 5724
rect 7520 5644 7524 5676
rect 7556 5644 7560 5676
rect 7520 5596 7560 5644
rect 7520 5564 7524 5596
rect 7556 5564 7560 5596
rect 7520 5516 7560 5564
rect 7520 5484 7524 5516
rect 7556 5484 7560 5516
rect 7520 5436 7560 5484
rect 7520 5404 7524 5436
rect 7556 5404 7560 5436
rect 7520 5356 7560 5404
rect 7520 5324 7524 5356
rect 7556 5324 7560 5356
rect 7520 5276 7560 5324
rect 7520 5244 7524 5276
rect 7556 5244 7560 5276
rect 7520 5196 7560 5244
rect 7520 5164 7524 5196
rect 7556 5164 7560 5196
rect 7520 5116 7560 5164
rect 7520 5084 7524 5116
rect 7556 5084 7560 5116
rect 7520 5036 7560 5084
rect 7520 5004 7524 5036
rect 7556 5004 7560 5036
rect 7520 4956 7560 5004
rect 7520 4924 7524 4956
rect 7556 4924 7560 4956
rect 7520 4876 7560 4924
rect 7520 4844 7524 4876
rect 7556 4844 7560 4876
rect 7520 4796 7560 4844
rect 7520 4764 7524 4796
rect 7556 4764 7560 4796
rect 7520 4716 7560 4764
rect 7520 4684 7524 4716
rect 7556 4684 7560 4716
rect 7520 4636 7560 4684
rect 7520 4604 7524 4636
rect 7556 4604 7560 4636
rect 7520 4556 7560 4604
rect 7520 4524 7524 4556
rect 7556 4524 7560 4556
rect 7520 4476 7560 4524
rect 7520 4444 7524 4476
rect 7556 4444 7560 4476
rect 7520 4396 7560 4444
rect 7520 4364 7524 4396
rect 7556 4364 7560 4396
rect 7520 4316 7560 4364
rect 7520 4284 7524 4316
rect 7556 4284 7560 4316
rect 7520 4236 7560 4284
rect 7520 4204 7524 4236
rect 7556 4204 7560 4236
rect 7520 4156 7560 4204
rect 7520 4124 7524 4156
rect 7556 4124 7560 4156
rect 7520 4076 7560 4124
rect 7520 4044 7524 4076
rect 7556 4044 7560 4076
rect 7520 3996 7560 4044
rect 7520 3964 7524 3996
rect 7556 3964 7560 3996
rect 7520 3916 7560 3964
rect 7520 3884 7524 3916
rect 7556 3884 7560 3916
rect 7520 3836 7560 3884
rect 7520 3804 7524 3836
rect 7556 3804 7560 3836
rect 7520 3756 7560 3804
rect 7520 3724 7524 3756
rect 7556 3724 7560 3756
rect 7520 3676 7560 3724
rect 7520 3644 7524 3676
rect 7556 3644 7560 3676
rect 7520 3596 7560 3644
rect 7520 3564 7524 3596
rect 7556 3564 7560 3596
rect 7520 3516 7560 3564
rect 7520 3484 7524 3516
rect 7556 3484 7560 3516
rect 7520 3436 7560 3484
rect 7520 3404 7524 3436
rect 7556 3404 7560 3436
rect 7520 3356 7560 3404
rect 7520 3324 7524 3356
rect 7556 3324 7560 3356
rect 7520 3276 7560 3324
rect 7520 3244 7524 3276
rect 7556 3244 7560 3276
rect 7520 3196 7560 3244
rect 7520 3164 7524 3196
rect 7556 3164 7560 3196
rect 7520 3116 7560 3164
rect 7520 3084 7524 3116
rect 7556 3084 7560 3116
rect 7520 3036 7560 3084
rect 7520 3004 7524 3036
rect 7556 3004 7560 3036
rect 7520 2956 7560 3004
rect 7520 2924 7524 2956
rect 7556 2924 7560 2956
rect 7520 2876 7560 2924
rect 7520 2844 7524 2876
rect 7556 2844 7560 2876
rect 7520 2796 7560 2844
rect 7520 2764 7524 2796
rect 7556 2764 7560 2796
rect 7520 2716 7560 2764
rect 7520 2684 7524 2716
rect 7556 2684 7560 2716
rect 7520 2636 7560 2684
rect 7520 2604 7524 2636
rect 7556 2604 7560 2636
rect 7520 2556 7560 2604
rect 7520 2524 7524 2556
rect 7556 2524 7560 2556
rect 7520 2476 7560 2524
rect 7520 2444 7524 2476
rect 7556 2444 7560 2476
rect 7520 2396 7560 2444
rect 7520 2364 7524 2396
rect 7556 2364 7560 2396
rect 7520 2316 7560 2364
rect 7520 2284 7524 2316
rect 7556 2284 7560 2316
rect 7520 2236 7560 2284
rect 7520 2204 7524 2236
rect 7556 2204 7560 2236
rect 7520 2156 7560 2204
rect 7520 2124 7524 2156
rect 7556 2124 7560 2156
rect 7520 2076 7560 2124
rect 7520 2044 7524 2076
rect 7556 2044 7560 2076
rect 7520 1996 7560 2044
rect 7520 1964 7524 1996
rect 7556 1964 7560 1996
rect 7520 1916 7560 1964
rect 7520 1884 7524 1916
rect 7556 1884 7560 1916
rect 7520 1836 7560 1884
rect 7520 1804 7524 1836
rect 7556 1804 7560 1836
rect 7520 1756 7560 1804
rect 7520 1724 7524 1756
rect 7556 1724 7560 1756
rect 7520 1676 7560 1724
rect 7520 1644 7524 1676
rect 7556 1644 7560 1676
rect 7520 1596 7560 1644
rect 7520 1564 7524 1596
rect 7556 1564 7560 1596
rect 7520 1516 7560 1564
rect 7520 1484 7524 1516
rect 7556 1484 7560 1516
rect 7520 1436 7560 1484
rect 7520 1404 7524 1436
rect 7556 1404 7560 1436
rect 7520 1356 7560 1404
rect 7520 1324 7524 1356
rect 7556 1324 7560 1356
rect 7520 1276 7560 1324
rect 7520 1244 7524 1276
rect 7556 1244 7560 1276
rect 7520 1196 7560 1244
rect 7520 1164 7524 1196
rect 7556 1164 7560 1196
rect 7520 1116 7560 1164
rect 7520 1084 7524 1116
rect 7556 1084 7560 1116
rect 7520 1036 7560 1084
rect 7520 1004 7524 1036
rect 7556 1004 7560 1036
rect 7520 956 7560 1004
rect 7520 924 7524 956
rect 7556 924 7560 956
rect 7520 876 7560 924
rect 7520 844 7524 876
rect 7556 844 7560 876
rect 7520 796 7560 844
rect 7520 764 7524 796
rect 7556 764 7560 796
rect 7520 716 7560 764
rect 7520 684 7524 716
rect 7556 684 7560 716
rect 7520 596 7560 684
rect 7520 564 7524 596
rect 7556 564 7560 596
rect 7520 516 7560 564
rect 7520 484 7524 516
rect 7556 484 7560 516
rect 7520 436 7560 484
rect 7520 404 7524 436
rect 7556 404 7560 436
rect 7520 356 7560 404
rect 7520 324 7524 356
rect 7556 324 7560 356
rect 7520 276 7560 324
rect 7520 244 7524 276
rect 7556 244 7560 276
rect 7520 196 7560 244
rect 7520 164 7524 196
rect 7556 164 7560 196
rect 7520 116 7560 164
rect 7520 84 7524 116
rect 7556 84 7560 116
rect 7520 36 7560 84
rect 7520 4 7524 36
rect 7556 4 7560 36
rect 7520 -40 7560 4
rect 7600 15795 7640 17284
rect 7680 17200 7720 18404
rect 7760 17200 7800 18440
rect 7760 16836 7800 17080
rect 7760 16644 7764 16836
rect 7796 16644 7800 16836
rect 7600 15765 7605 15795
rect 7635 15765 7640 15795
rect 7600 12835 7640 15765
rect 7600 12805 7605 12835
rect 7635 12805 7640 12835
rect 7600 8875 7640 12805
rect 7600 8845 7605 8875
rect 7635 8845 7640 8875
rect 7600 -40 7640 8845
rect 7680 16596 7720 16600
rect 7680 16564 7684 16596
rect 7716 16564 7720 16596
rect 7680 16516 7720 16564
rect 7680 16484 7684 16516
rect 7716 16484 7720 16516
rect 7680 16436 7720 16484
rect 7680 16404 7684 16436
rect 7716 16404 7720 16436
rect 7680 16356 7720 16404
rect 7680 16324 7684 16356
rect 7716 16324 7720 16356
rect 7680 16276 7720 16324
rect 7680 16244 7684 16276
rect 7716 16244 7720 16276
rect 7680 16196 7720 16244
rect 7680 16164 7684 16196
rect 7716 16164 7720 16196
rect 7680 16116 7720 16164
rect 7680 16084 7684 16116
rect 7716 16084 7720 16116
rect 7680 16036 7720 16084
rect 7680 16004 7684 16036
rect 7716 16004 7720 16036
rect 7680 15956 7720 16004
rect 7680 15924 7684 15956
rect 7716 15924 7720 15956
rect 7680 15875 7720 15924
rect 7680 15845 7685 15875
rect 7715 15845 7720 15875
rect 7680 15715 7720 15845
rect 7680 15685 7685 15715
rect 7715 15685 7720 15715
rect 7680 15555 7720 15685
rect 7680 15525 7685 15555
rect 7715 15525 7720 15555
rect 7680 15436 7720 15525
rect 7680 15404 7684 15436
rect 7716 15404 7720 15436
rect 7680 15356 7720 15404
rect 7680 15324 7684 15356
rect 7716 15324 7720 15356
rect 7680 15276 7720 15324
rect 7680 15244 7684 15276
rect 7716 15244 7720 15276
rect 7680 15196 7720 15244
rect 7680 15164 7684 15196
rect 7716 15164 7720 15196
rect 7680 15116 7720 15164
rect 7680 15084 7684 15116
rect 7716 15084 7720 15116
rect 7680 15036 7720 15084
rect 7680 15004 7684 15036
rect 7716 15004 7720 15036
rect 7680 14956 7720 15004
rect 7680 14924 7684 14956
rect 7716 14924 7720 14956
rect 7680 14876 7720 14924
rect 7680 14844 7684 14876
rect 7716 14844 7720 14876
rect 7680 14796 7720 14844
rect 7680 14764 7684 14796
rect 7716 14764 7720 14796
rect 7680 14716 7720 14764
rect 7680 14684 7684 14716
rect 7716 14684 7720 14716
rect 7680 14636 7720 14684
rect 7680 14604 7684 14636
rect 7716 14604 7720 14636
rect 7680 14556 7720 14604
rect 7680 14524 7684 14556
rect 7716 14524 7720 14556
rect 7680 14476 7720 14524
rect 7680 14444 7684 14476
rect 7716 14444 7720 14476
rect 7680 14396 7720 14444
rect 7680 14364 7684 14396
rect 7716 14364 7720 14396
rect 7680 14316 7720 14364
rect 7680 14284 7684 14316
rect 7716 14284 7720 14316
rect 7680 14236 7720 14284
rect 7680 14204 7684 14236
rect 7716 14204 7720 14236
rect 7680 14156 7720 14204
rect 7680 14124 7684 14156
rect 7716 14124 7720 14156
rect 7680 14076 7720 14124
rect 7680 14044 7684 14076
rect 7716 14044 7720 14076
rect 7680 13996 7720 14044
rect 7680 13964 7684 13996
rect 7716 13964 7720 13996
rect 7680 13876 7720 13964
rect 7680 13844 7684 13876
rect 7716 13844 7720 13876
rect 7680 13796 7720 13844
rect 7680 13764 7684 13796
rect 7716 13764 7720 13796
rect 7680 13716 7720 13764
rect 7680 13684 7684 13716
rect 7716 13684 7720 13716
rect 7680 13636 7720 13684
rect 7680 13604 7684 13636
rect 7716 13604 7720 13636
rect 7680 13556 7720 13604
rect 7680 13524 7684 13556
rect 7716 13524 7720 13556
rect 7680 13476 7720 13524
rect 7680 13444 7684 13476
rect 7716 13444 7720 13476
rect 7680 13396 7720 13444
rect 7680 13364 7684 13396
rect 7716 13364 7720 13396
rect 7680 13316 7720 13364
rect 7680 13284 7684 13316
rect 7716 13284 7720 13316
rect 7680 13236 7720 13284
rect 7680 13204 7684 13236
rect 7716 13204 7720 13236
rect 7680 13156 7720 13204
rect 7680 13124 7684 13156
rect 7716 13124 7720 13156
rect 7680 13076 7720 13124
rect 7680 13044 7684 13076
rect 7716 13044 7720 13076
rect 7680 12996 7720 13044
rect 7680 12964 7684 12996
rect 7716 12964 7720 12996
rect 7680 12915 7720 12964
rect 7680 12885 7685 12915
rect 7715 12885 7720 12915
rect 7680 12755 7720 12885
rect 7680 12725 7685 12755
rect 7715 12725 7720 12755
rect 7680 12595 7720 12725
rect 7680 12565 7685 12595
rect 7715 12565 7720 12595
rect 7680 12476 7720 12565
rect 7680 12444 7684 12476
rect 7716 12444 7720 12476
rect 7680 12396 7720 12444
rect 7680 12364 7684 12396
rect 7716 12364 7720 12396
rect 7680 12316 7720 12364
rect 7680 12284 7684 12316
rect 7716 12284 7720 12316
rect 7680 12236 7720 12284
rect 7680 12204 7684 12236
rect 7716 12204 7720 12236
rect 7680 12156 7720 12204
rect 7680 12124 7684 12156
rect 7716 12124 7720 12156
rect 7680 12076 7720 12124
rect 7680 12044 7684 12076
rect 7716 12044 7720 12076
rect 7680 11996 7720 12044
rect 7680 11964 7684 11996
rect 7716 11964 7720 11996
rect 7680 11916 7720 11964
rect 7680 11884 7684 11916
rect 7716 11884 7720 11916
rect 7680 11836 7720 11884
rect 7680 11804 7684 11836
rect 7716 11804 7720 11836
rect 7680 11756 7720 11804
rect 7680 11724 7684 11756
rect 7716 11724 7720 11756
rect 7680 11676 7720 11724
rect 7680 11644 7684 11676
rect 7716 11644 7720 11676
rect 7680 11596 7720 11644
rect 7680 11564 7684 11596
rect 7716 11564 7720 11596
rect 7680 11516 7720 11564
rect 7680 11484 7684 11516
rect 7716 11484 7720 11516
rect 7680 11436 7720 11484
rect 7680 11404 7684 11436
rect 7716 11404 7720 11436
rect 7680 11356 7720 11404
rect 7680 11324 7684 11356
rect 7716 11324 7720 11356
rect 7680 11276 7720 11324
rect 7680 11244 7684 11276
rect 7716 11244 7720 11276
rect 7680 11196 7720 11244
rect 7680 11164 7684 11196
rect 7716 11164 7720 11196
rect 7680 11116 7720 11164
rect 7680 11084 7684 11116
rect 7716 11084 7720 11116
rect 7680 11036 7720 11084
rect 7680 11004 7684 11036
rect 7716 11004 7720 11036
rect 7680 10956 7720 11004
rect 7680 10924 7684 10956
rect 7716 10924 7720 10956
rect 7680 10876 7720 10924
rect 7680 10844 7684 10876
rect 7716 10844 7720 10876
rect 7680 10796 7720 10844
rect 7680 10764 7684 10796
rect 7716 10764 7720 10796
rect 7680 10716 7720 10764
rect 7680 10684 7684 10716
rect 7716 10684 7720 10716
rect 7680 10636 7720 10684
rect 7680 10604 7684 10636
rect 7716 10604 7720 10636
rect 7680 10556 7720 10604
rect 7680 10524 7684 10556
rect 7716 10524 7720 10556
rect 7680 10476 7720 10524
rect 7680 10444 7684 10476
rect 7716 10444 7720 10476
rect 7680 10396 7720 10444
rect 7680 10364 7684 10396
rect 7716 10364 7720 10396
rect 7680 10316 7720 10364
rect 7680 10284 7684 10316
rect 7716 10284 7720 10316
rect 7680 10236 7720 10284
rect 7680 10204 7684 10236
rect 7716 10204 7720 10236
rect 7680 10156 7720 10204
rect 7680 10124 7684 10156
rect 7716 10124 7720 10156
rect 7680 10076 7720 10124
rect 7680 10044 7684 10076
rect 7716 10044 7720 10076
rect 7680 9996 7720 10044
rect 7680 9964 7684 9996
rect 7716 9964 7720 9996
rect 7680 9916 7720 9964
rect 7680 9884 7684 9916
rect 7716 9884 7720 9916
rect 7680 9836 7720 9884
rect 7680 9804 7684 9836
rect 7716 9804 7720 9836
rect 7680 9756 7720 9804
rect 7680 9724 7684 9756
rect 7716 9724 7720 9756
rect 7680 9676 7720 9724
rect 7680 9644 7684 9676
rect 7716 9644 7720 9676
rect 7680 9596 7720 9644
rect 7680 9564 7684 9596
rect 7716 9564 7720 9596
rect 7680 9516 7720 9564
rect 7680 9484 7684 9516
rect 7716 9484 7720 9516
rect 7680 9436 7720 9484
rect 7680 9404 7684 9436
rect 7716 9404 7720 9436
rect 7680 9356 7720 9404
rect 7680 9324 7684 9356
rect 7716 9324 7720 9356
rect 7680 9276 7720 9324
rect 7680 9244 7684 9276
rect 7716 9244 7720 9276
rect 7680 9196 7720 9244
rect 7680 9164 7684 9196
rect 7716 9164 7720 9196
rect 7680 9116 7720 9164
rect 7680 9084 7684 9116
rect 7716 9084 7720 9116
rect 7680 9036 7720 9084
rect 7680 9004 7684 9036
rect 7716 9004 7720 9036
rect 7680 8956 7720 9004
rect 7680 8924 7684 8956
rect 7716 8924 7720 8956
rect 7680 8795 7720 8924
rect 7680 8765 7685 8795
rect 7715 8765 7720 8795
rect 7680 8636 7720 8765
rect 7680 8604 7684 8636
rect 7716 8604 7720 8636
rect 7680 8556 7720 8604
rect 7680 8524 7684 8556
rect 7716 8524 7720 8556
rect 7680 8476 7720 8524
rect 7680 8444 7684 8476
rect 7716 8444 7720 8476
rect 7680 8396 7720 8444
rect 7680 8364 7684 8396
rect 7716 8364 7720 8396
rect 7680 8316 7720 8364
rect 7680 8284 7684 8316
rect 7716 8284 7720 8316
rect 7680 8236 7720 8284
rect 7680 8204 7684 8236
rect 7716 8204 7720 8236
rect 7680 8156 7720 8204
rect 7680 8124 7684 8156
rect 7716 8124 7720 8156
rect 7680 8076 7720 8124
rect 7680 8044 7684 8076
rect 7716 8044 7720 8076
rect 7680 7996 7720 8044
rect 7680 7964 7684 7996
rect 7716 7964 7720 7996
rect 7680 7916 7720 7964
rect 7680 7884 7684 7916
rect 7716 7884 7720 7916
rect 7680 7836 7720 7884
rect 7680 7804 7684 7836
rect 7716 7804 7720 7836
rect 7680 7756 7720 7804
rect 7680 7724 7684 7756
rect 7716 7724 7720 7756
rect 7680 7676 7720 7724
rect 7680 7644 7684 7676
rect 7716 7644 7720 7676
rect 7680 7596 7720 7644
rect 7680 7564 7684 7596
rect 7716 7564 7720 7596
rect 7680 7516 7720 7564
rect 7680 7484 7684 7516
rect 7716 7484 7720 7516
rect 7680 7436 7720 7484
rect 7680 7404 7684 7436
rect 7716 7404 7720 7436
rect 7680 7356 7720 7404
rect 7680 7324 7684 7356
rect 7716 7324 7720 7356
rect 7680 7276 7720 7324
rect 7680 7244 7684 7276
rect 7716 7244 7720 7276
rect 7680 7196 7720 7244
rect 7680 7164 7684 7196
rect 7716 7164 7720 7196
rect 7680 7116 7720 7164
rect 7680 7084 7684 7116
rect 7716 7084 7720 7116
rect 7680 7036 7720 7084
rect 7680 7004 7684 7036
rect 7716 7004 7720 7036
rect 7680 6956 7720 7004
rect 7680 6924 7684 6956
rect 7716 6924 7720 6956
rect 7680 6876 7720 6924
rect 7680 6844 7684 6876
rect 7716 6844 7720 6876
rect 7680 6796 7720 6844
rect 7680 6764 7684 6796
rect 7716 6764 7720 6796
rect 7680 6716 7720 6764
rect 7680 6684 7684 6716
rect 7716 6684 7720 6716
rect 7680 6636 7720 6684
rect 7680 6604 7684 6636
rect 7716 6604 7720 6636
rect 7680 6556 7720 6604
rect 7680 6524 7684 6556
rect 7716 6524 7720 6556
rect 7680 6476 7720 6524
rect 7680 6444 7684 6476
rect 7716 6444 7720 6476
rect 7680 6396 7720 6444
rect 7680 6364 7684 6396
rect 7716 6364 7720 6396
rect 7680 6316 7720 6364
rect 7680 6284 7684 6316
rect 7716 6284 7720 6316
rect 7680 6236 7720 6284
rect 7680 6204 7684 6236
rect 7716 6204 7720 6236
rect 7680 6156 7720 6204
rect 7680 6124 7684 6156
rect 7716 6124 7720 6156
rect 7680 6076 7720 6124
rect 7680 6044 7684 6076
rect 7716 6044 7720 6076
rect 7680 5996 7720 6044
rect 7680 5964 7684 5996
rect 7716 5964 7720 5996
rect 7680 5916 7720 5964
rect 7680 5884 7684 5916
rect 7716 5884 7720 5916
rect 7680 5836 7720 5884
rect 7680 5804 7684 5836
rect 7716 5804 7720 5836
rect 7680 5756 7720 5804
rect 7680 5724 7684 5756
rect 7716 5724 7720 5756
rect 7680 5676 7720 5724
rect 7680 5644 7684 5676
rect 7716 5644 7720 5676
rect 7680 5596 7720 5644
rect 7680 5564 7684 5596
rect 7716 5564 7720 5596
rect 7680 5516 7720 5564
rect 7680 5484 7684 5516
rect 7716 5484 7720 5516
rect 7680 5436 7720 5484
rect 7680 5404 7684 5436
rect 7716 5404 7720 5436
rect 7680 5356 7720 5404
rect 7680 5324 7684 5356
rect 7716 5324 7720 5356
rect 7680 5276 7720 5324
rect 7680 5244 7684 5276
rect 7716 5244 7720 5276
rect 7680 5196 7720 5244
rect 7680 5164 7684 5196
rect 7716 5164 7720 5196
rect 7680 5116 7720 5164
rect 7680 5084 7684 5116
rect 7716 5084 7720 5116
rect 7680 5036 7720 5084
rect 7680 5004 7684 5036
rect 7716 5004 7720 5036
rect 7680 4956 7720 5004
rect 7680 4924 7684 4956
rect 7716 4924 7720 4956
rect 7680 4876 7720 4924
rect 7680 4844 7684 4876
rect 7716 4844 7720 4876
rect 7680 4796 7720 4844
rect 7680 4764 7684 4796
rect 7716 4764 7720 4796
rect 7680 4716 7720 4764
rect 7680 4684 7684 4716
rect 7716 4684 7720 4716
rect 7680 4636 7720 4684
rect 7680 4604 7684 4636
rect 7716 4604 7720 4636
rect 7680 4556 7720 4604
rect 7680 4524 7684 4556
rect 7716 4524 7720 4556
rect 7680 4476 7720 4524
rect 7680 4444 7684 4476
rect 7716 4444 7720 4476
rect 7680 4396 7720 4444
rect 7680 4364 7684 4396
rect 7716 4364 7720 4396
rect 7680 4316 7720 4364
rect 7680 4284 7684 4316
rect 7716 4284 7720 4316
rect 7680 4236 7720 4284
rect 7680 4204 7684 4236
rect 7716 4204 7720 4236
rect 7680 4156 7720 4204
rect 7680 4124 7684 4156
rect 7716 4124 7720 4156
rect 7680 4076 7720 4124
rect 7680 4044 7684 4076
rect 7716 4044 7720 4076
rect 7680 3996 7720 4044
rect 7680 3964 7684 3996
rect 7716 3964 7720 3996
rect 7680 3916 7720 3964
rect 7680 3884 7684 3916
rect 7716 3884 7720 3916
rect 7680 3836 7720 3884
rect 7680 3804 7684 3836
rect 7716 3804 7720 3836
rect 7680 3756 7720 3804
rect 7680 3724 7684 3756
rect 7716 3724 7720 3756
rect 7680 3676 7720 3724
rect 7680 3644 7684 3676
rect 7716 3644 7720 3676
rect 7680 3596 7720 3644
rect 7680 3564 7684 3596
rect 7716 3564 7720 3596
rect 7680 3516 7720 3564
rect 7680 3484 7684 3516
rect 7716 3484 7720 3516
rect 7680 3436 7720 3484
rect 7680 3404 7684 3436
rect 7716 3404 7720 3436
rect 7680 3356 7720 3404
rect 7680 3324 7684 3356
rect 7716 3324 7720 3356
rect 7680 3276 7720 3324
rect 7680 3244 7684 3276
rect 7716 3244 7720 3276
rect 7680 3196 7720 3244
rect 7680 3164 7684 3196
rect 7716 3164 7720 3196
rect 7680 3116 7720 3164
rect 7680 3084 7684 3116
rect 7716 3084 7720 3116
rect 7680 3036 7720 3084
rect 7680 3004 7684 3036
rect 7716 3004 7720 3036
rect 7680 2956 7720 3004
rect 7680 2924 7684 2956
rect 7716 2924 7720 2956
rect 7680 2876 7720 2924
rect 7680 2844 7684 2876
rect 7716 2844 7720 2876
rect 7680 2796 7720 2844
rect 7680 2764 7684 2796
rect 7716 2764 7720 2796
rect 7680 2716 7720 2764
rect 7680 2684 7684 2716
rect 7716 2684 7720 2716
rect 7680 2636 7720 2684
rect 7680 2604 7684 2636
rect 7716 2604 7720 2636
rect 7680 2556 7720 2604
rect 7680 2524 7684 2556
rect 7716 2524 7720 2556
rect 7680 2476 7720 2524
rect 7680 2444 7684 2476
rect 7716 2444 7720 2476
rect 7680 2396 7720 2444
rect 7680 2364 7684 2396
rect 7716 2364 7720 2396
rect 7680 2316 7720 2364
rect 7680 2284 7684 2316
rect 7716 2284 7720 2316
rect 7680 2236 7720 2284
rect 7680 2204 7684 2236
rect 7716 2204 7720 2236
rect 7680 2156 7720 2204
rect 7680 2124 7684 2156
rect 7716 2124 7720 2156
rect 7680 2076 7720 2124
rect 7680 2044 7684 2076
rect 7716 2044 7720 2076
rect 7680 1996 7720 2044
rect 7680 1964 7684 1996
rect 7716 1964 7720 1996
rect 7680 1916 7720 1964
rect 7680 1884 7684 1916
rect 7716 1884 7720 1916
rect 7680 1836 7720 1884
rect 7680 1804 7684 1836
rect 7716 1804 7720 1836
rect 7680 1756 7720 1804
rect 7680 1724 7684 1756
rect 7716 1724 7720 1756
rect 7680 1676 7720 1724
rect 7680 1644 7684 1676
rect 7716 1644 7720 1676
rect 7680 1596 7720 1644
rect 7680 1564 7684 1596
rect 7716 1564 7720 1596
rect 7680 1516 7720 1564
rect 7680 1484 7684 1516
rect 7716 1484 7720 1516
rect 7680 1436 7720 1484
rect 7680 1404 7684 1436
rect 7716 1404 7720 1436
rect 7680 1356 7720 1404
rect 7680 1324 7684 1356
rect 7716 1324 7720 1356
rect 7680 1276 7720 1324
rect 7680 1244 7684 1276
rect 7716 1244 7720 1276
rect 7680 1196 7720 1244
rect 7680 1164 7684 1196
rect 7716 1164 7720 1196
rect 7680 1116 7720 1164
rect 7680 1084 7684 1116
rect 7716 1084 7720 1116
rect 7680 1036 7720 1084
rect 7680 1004 7684 1036
rect 7716 1004 7720 1036
rect 7680 956 7720 1004
rect 7680 924 7684 956
rect 7716 924 7720 956
rect 7680 876 7720 924
rect 7680 844 7684 876
rect 7716 844 7720 876
rect 7680 796 7720 844
rect 7680 764 7684 796
rect 7716 764 7720 796
rect 7680 716 7720 764
rect 7680 684 7684 716
rect 7716 684 7720 716
rect 7680 596 7720 684
rect 7680 564 7684 596
rect 7716 564 7720 596
rect 7680 516 7720 564
rect 7680 484 7684 516
rect 7716 484 7720 516
rect 7680 436 7720 484
rect 7680 404 7684 436
rect 7716 404 7720 436
rect 7680 356 7720 404
rect 7680 324 7684 356
rect 7716 324 7720 356
rect 7680 276 7720 324
rect 7680 244 7684 276
rect 7716 244 7720 276
rect 7680 196 7720 244
rect 7680 164 7684 196
rect 7716 164 7720 196
rect 7680 116 7720 164
rect 7680 84 7684 116
rect 7716 84 7720 116
rect 7680 36 7720 84
rect 7680 4 7684 36
rect 7716 4 7720 36
rect 7680 -40 7720 4
rect 7760 -40 7800 16644
<< via3 >>
rect 7364 19684 7396 19716
rect 564 19604 1636 19636
rect 1684 19604 2756 19636
rect 2804 19604 3876 19636
rect 3924 19604 4996 19636
rect 5044 19604 6116 19636
rect 6164 19604 7236 19636
rect 564 17284 1636 17316
rect 1684 17284 2756 17316
rect 2804 17284 3876 17316
rect 3924 17284 4996 17316
rect 5044 17284 6116 17316
rect 6164 17284 7236 17316
rect 7284 17124 7316 17156
rect 5524 16644 5556 16836
rect 5684 16644 5716 16836
rect 5524 16595 5556 16596
rect 5524 16565 5525 16595
rect 5525 16565 5555 16595
rect 5555 16565 5556 16595
rect 5524 16564 5556 16565
rect 5524 16515 5556 16516
rect 5524 16485 5525 16515
rect 5525 16485 5555 16515
rect 5555 16485 5556 16515
rect 5524 16484 5556 16485
rect 5524 16435 5556 16436
rect 5524 16405 5525 16435
rect 5525 16405 5555 16435
rect 5555 16405 5556 16435
rect 5524 16404 5556 16405
rect 5524 16355 5556 16356
rect 5524 16325 5525 16355
rect 5525 16325 5555 16355
rect 5555 16325 5556 16355
rect 5524 16324 5556 16325
rect 5524 16275 5556 16276
rect 5524 16245 5525 16275
rect 5525 16245 5555 16275
rect 5555 16245 5556 16275
rect 5524 16244 5556 16245
rect 5524 16195 5556 16196
rect 5524 16165 5525 16195
rect 5525 16165 5555 16195
rect 5555 16165 5556 16195
rect 5524 16164 5556 16165
rect 5524 16115 5556 16116
rect 5524 16085 5525 16115
rect 5525 16085 5555 16115
rect 5555 16085 5556 16115
rect 5524 16084 5556 16085
rect 5524 16035 5556 16036
rect 5524 16005 5525 16035
rect 5525 16005 5555 16035
rect 5555 16005 5556 16035
rect 5524 16004 5556 16005
rect 5524 15955 5556 15956
rect 5524 15925 5525 15955
rect 5525 15925 5555 15955
rect 5555 15925 5556 15955
rect 5524 15924 5556 15925
rect 5524 15435 5556 15436
rect 5524 15405 5525 15435
rect 5525 15405 5555 15435
rect 5555 15405 5556 15435
rect 5524 15404 5556 15405
rect 5524 15355 5556 15356
rect 5524 15325 5525 15355
rect 5525 15325 5555 15355
rect 5555 15325 5556 15355
rect 5524 15324 5556 15325
rect 5524 15275 5556 15276
rect 5524 15245 5525 15275
rect 5525 15245 5555 15275
rect 5555 15245 5556 15275
rect 5524 15244 5556 15245
rect 5524 15195 5556 15196
rect 5524 15165 5525 15195
rect 5525 15165 5555 15195
rect 5555 15165 5556 15195
rect 5524 15164 5556 15165
rect 5524 15115 5556 15116
rect 5524 15085 5525 15115
rect 5525 15085 5555 15115
rect 5555 15085 5556 15115
rect 5524 15084 5556 15085
rect 5524 14955 5556 14956
rect 5524 14925 5525 14955
rect 5525 14925 5555 14955
rect 5555 14925 5556 14955
rect 5524 14924 5556 14925
rect 5524 14875 5556 14876
rect 5524 14845 5525 14875
rect 5525 14845 5555 14875
rect 5555 14845 5556 14875
rect 5524 14844 5556 14845
rect 5524 14795 5556 14796
rect 5524 14765 5525 14795
rect 5525 14765 5555 14795
rect 5555 14765 5556 14795
rect 5524 14764 5556 14765
rect 5524 14715 5556 14716
rect 5524 14685 5525 14715
rect 5525 14685 5555 14715
rect 5555 14685 5556 14715
rect 5524 14684 5556 14685
rect 5524 14555 5556 14556
rect 5524 14525 5525 14555
rect 5525 14525 5555 14555
rect 5555 14525 5556 14555
rect 5524 14524 5556 14525
rect 5524 14475 5556 14476
rect 5524 14445 5525 14475
rect 5525 14445 5555 14475
rect 5555 14445 5556 14475
rect 5524 14444 5556 14445
rect 5524 13995 5556 13996
rect 5524 13965 5525 13995
rect 5525 13965 5555 13995
rect 5555 13965 5556 13995
rect 5524 13964 5556 13965
rect 5524 13795 5556 13796
rect 5524 13765 5525 13795
rect 5525 13765 5555 13795
rect 5555 13765 5556 13795
rect 5524 13764 5556 13765
rect 5524 13715 5556 13716
rect 5524 13685 5525 13715
rect 5525 13685 5555 13715
rect 5555 13685 5556 13715
rect 5524 13684 5556 13685
rect 5524 13635 5556 13636
rect 5524 13605 5525 13635
rect 5525 13605 5555 13635
rect 5555 13605 5556 13635
rect 5524 13604 5556 13605
rect 5524 13475 5556 13476
rect 5524 13445 5525 13475
rect 5525 13445 5555 13475
rect 5555 13445 5556 13475
rect 5524 13444 5556 13445
rect 5524 13395 5556 13396
rect 5524 13365 5525 13395
rect 5525 13365 5555 13395
rect 5555 13365 5556 13395
rect 5524 13364 5556 13365
rect 5524 13315 5556 13316
rect 5524 13285 5525 13315
rect 5525 13285 5555 13315
rect 5555 13285 5556 13315
rect 5524 13284 5556 13285
rect 5524 13235 5556 13236
rect 5524 13205 5525 13235
rect 5525 13205 5555 13235
rect 5555 13205 5556 13235
rect 5524 13204 5556 13205
rect 5524 13075 5556 13076
rect 5524 13045 5525 13075
rect 5525 13045 5555 13075
rect 5555 13045 5556 13075
rect 5524 13044 5556 13045
rect 5524 12995 5556 12996
rect 5524 12965 5525 12995
rect 5525 12965 5555 12995
rect 5555 12965 5556 12995
rect 5524 12964 5556 12965
rect 5524 12515 5556 12516
rect 5524 12485 5525 12515
rect 5525 12485 5555 12515
rect 5555 12485 5556 12515
rect 5524 12484 5556 12485
rect 5524 12315 5556 12316
rect 5524 12285 5525 12315
rect 5525 12285 5555 12315
rect 5555 12285 5556 12315
rect 5524 12284 5556 12285
rect 5524 12235 5556 12236
rect 5524 12205 5525 12235
rect 5525 12205 5555 12235
rect 5555 12205 5556 12235
rect 5524 12204 5556 12205
rect 5524 12155 5556 12156
rect 5524 12125 5525 12155
rect 5525 12125 5555 12155
rect 5555 12125 5556 12155
rect 5524 12124 5556 12125
rect 5524 12075 5556 12076
rect 5524 12045 5525 12075
rect 5525 12045 5555 12075
rect 5555 12045 5556 12075
rect 5524 12044 5556 12045
rect 5524 11995 5556 11996
rect 5524 11965 5525 11995
rect 5525 11965 5555 11995
rect 5555 11965 5556 11995
rect 5524 11964 5556 11965
rect 5524 11915 5556 11916
rect 5524 11885 5525 11915
rect 5525 11885 5555 11915
rect 5555 11885 5556 11915
rect 5524 11884 5556 11885
rect 5524 11835 5556 11836
rect 5524 11805 5525 11835
rect 5525 11805 5555 11835
rect 5555 11805 5556 11835
rect 5524 11804 5556 11805
rect 5524 11755 5556 11756
rect 5524 11725 5525 11755
rect 5525 11725 5555 11755
rect 5555 11725 5556 11755
rect 5524 11724 5556 11725
rect 5524 11675 5556 11676
rect 5524 11645 5525 11675
rect 5525 11645 5555 11675
rect 5555 11645 5556 11675
rect 5524 11644 5556 11645
rect 5524 11595 5556 11596
rect 5524 11565 5525 11595
rect 5525 11565 5555 11595
rect 5555 11565 5556 11595
rect 5524 11564 5556 11565
rect 5524 11515 5556 11516
rect 5524 11485 5525 11515
rect 5525 11485 5555 11515
rect 5555 11485 5556 11515
rect 5524 11484 5556 11485
rect 5524 11435 5556 11436
rect 5524 11405 5525 11435
rect 5525 11405 5555 11435
rect 5555 11405 5556 11435
rect 5524 11404 5556 11405
rect 5524 11355 5556 11356
rect 5524 11325 5525 11355
rect 5525 11325 5555 11355
rect 5555 11325 5556 11355
rect 5524 11324 5556 11325
rect 5524 11195 5556 11196
rect 5524 11165 5525 11195
rect 5525 11165 5555 11195
rect 5555 11165 5556 11195
rect 5524 11164 5556 11165
rect 5524 11115 5556 11116
rect 5524 11085 5525 11115
rect 5525 11085 5555 11115
rect 5555 11085 5556 11115
rect 5524 11084 5556 11085
rect 5524 11035 5556 11036
rect 5524 11005 5525 11035
rect 5525 11005 5555 11035
rect 5555 11005 5556 11035
rect 5524 11004 5556 11005
rect 5524 10875 5556 10876
rect 5524 10845 5525 10875
rect 5525 10845 5555 10875
rect 5555 10845 5556 10875
rect 5524 10844 5556 10845
rect 5524 10715 5556 10716
rect 5524 10685 5525 10715
rect 5525 10685 5555 10715
rect 5555 10685 5556 10715
rect 5524 10684 5556 10685
rect 5524 10635 5556 10636
rect 5524 10605 5525 10635
rect 5525 10605 5555 10635
rect 5555 10605 5556 10635
rect 5524 10604 5556 10605
rect 5524 10475 5556 10476
rect 5524 10445 5525 10475
rect 5525 10445 5555 10475
rect 5555 10445 5556 10475
rect 5524 10444 5556 10445
rect 5524 10315 5556 10316
rect 5524 10285 5525 10315
rect 5525 10285 5555 10315
rect 5555 10285 5556 10315
rect 5524 10284 5556 10285
rect 5524 10235 5556 10236
rect 5524 10205 5525 10235
rect 5525 10205 5555 10235
rect 5555 10205 5556 10235
rect 5524 10204 5556 10205
rect 5524 10155 5556 10156
rect 5524 10125 5525 10155
rect 5525 10125 5555 10155
rect 5555 10125 5556 10155
rect 5524 10124 5556 10125
rect 5524 10075 5556 10076
rect 5524 10045 5525 10075
rect 5525 10045 5555 10075
rect 5555 10045 5556 10075
rect 5524 10044 5556 10045
rect 5524 9995 5556 9996
rect 5524 9965 5525 9995
rect 5525 9965 5555 9995
rect 5555 9965 5556 9995
rect 5524 9964 5556 9965
rect 5524 9915 5556 9916
rect 5524 9885 5525 9915
rect 5525 9885 5555 9915
rect 5555 9885 5556 9915
rect 5524 9884 5556 9885
rect 5524 9835 5556 9836
rect 5524 9805 5525 9835
rect 5525 9805 5555 9835
rect 5555 9805 5556 9835
rect 5524 9804 5556 9805
rect 5524 9755 5556 9756
rect 5524 9725 5525 9755
rect 5525 9725 5555 9755
rect 5555 9725 5556 9755
rect 5524 9724 5556 9725
rect 5524 9675 5556 9676
rect 5524 9645 5525 9675
rect 5525 9645 5555 9675
rect 5555 9645 5556 9675
rect 5524 9644 5556 9645
rect 5524 9595 5556 9596
rect 5524 9565 5525 9595
rect 5525 9565 5555 9595
rect 5555 9565 5556 9595
rect 5524 9564 5556 9565
rect 5524 9515 5556 9516
rect 5524 9485 5525 9515
rect 5525 9485 5555 9515
rect 5555 9485 5556 9515
rect 5524 9484 5556 9485
rect 5524 9435 5556 9436
rect 5524 9405 5525 9435
rect 5525 9405 5555 9435
rect 5555 9405 5556 9435
rect 5524 9404 5556 9405
rect 5524 9355 5556 9356
rect 5524 9325 5525 9355
rect 5525 9325 5555 9355
rect 5555 9325 5556 9355
rect 5524 9324 5556 9325
rect 5524 9275 5556 9276
rect 5524 9245 5525 9275
rect 5525 9245 5555 9275
rect 5555 9245 5556 9275
rect 5524 9244 5556 9245
rect 5524 9115 5556 9116
rect 5524 9085 5525 9115
rect 5525 9085 5555 9115
rect 5555 9085 5556 9115
rect 5524 9084 5556 9085
rect 5524 9035 5556 9036
rect 5524 9005 5525 9035
rect 5525 9005 5555 9035
rect 5555 9005 5556 9035
rect 5524 9004 5556 9005
rect 5524 8955 5556 8956
rect 5524 8925 5525 8955
rect 5525 8925 5555 8955
rect 5555 8925 5556 8955
rect 5524 8924 5556 8925
rect 5524 8635 5556 8636
rect 5524 8605 5525 8635
rect 5525 8605 5555 8635
rect 5555 8605 5556 8635
rect 5524 8604 5556 8605
rect 5524 8555 5556 8556
rect 5524 8525 5525 8555
rect 5525 8525 5555 8555
rect 5555 8525 5556 8555
rect 5524 8524 5556 8525
rect 5524 8395 5556 8396
rect 5524 8365 5525 8395
rect 5525 8365 5555 8395
rect 5555 8365 5556 8395
rect 5524 8364 5556 8365
rect 5524 8235 5556 8236
rect 5524 8205 5525 8235
rect 5525 8205 5555 8235
rect 5555 8205 5556 8235
rect 5524 8204 5556 8205
rect 5524 8155 5556 8156
rect 5524 8125 5525 8155
rect 5525 8125 5555 8155
rect 5555 8125 5556 8155
rect 5524 8124 5556 8125
rect 5524 8075 5556 8076
rect 5524 8045 5525 8075
rect 5525 8045 5555 8075
rect 5555 8045 5556 8075
rect 5524 8044 5556 8045
rect 5524 7995 5556 7996
rect 5524 7965 5525 7995
rect 5525 7965 5555 7995
rect 5555 7965 5556 7995
rect 5524 7964 5556 7965
rect 5524 7915 5556 7916
rect 5524 7885 5525 7915
rect 5525 7885 5555 7915
rect 5555 7885 5556 7915
rect 5524 7884 5556 7885
rect 5524 7835 5556 7836
rect 5524 7805 5525 7835
rect 5525 7805 5555 7835
rect 5555 7805 5556 7835
rect 5524 7804 5556 7805
rect 5524 7755 5556 7756
rect 5524 7725 5525 7755
rect 5525 7725 5555 7755
rect 5555 7725 5556 7755
rect 5524 7724 5556 7725
rect 5524 7675 5556 7676
rect 5524 7645 5525 7675
rect 5525 7645 5555 7675
rect 5555 7645 5556 7675
rect 5524 7644 5556 7645
rect 5524 7595 5556 7596
rect 5524 7565 5525 7595
rect 5525 7565 5555 7595
rect 5555 7565 5556 7595
rect 5524 7564 5556 7565
rect 5524 7515 5556 7516
rect 5524 7485 5525 7515
rect 5525 7485 5555 7515
rect 5555 7485 5556 7515
rect 5524 7484 5556 7485
rect 5524 7435 5556 7436
rect 5524 7405 5525 7435
rect 5525 7405 5555 7435
rect 5555 7405 5556 7435
rect 5524 7404 5556 7405
rect 5524 7355 5556 7356
rect 5524 7325 5525 7355
rect 5525 7325 5555 7355
rect 5555 7325 5556 7355
rect 5524 7324 5556 7325
rect 5524 7275 5556 7276
rect 5524 7245 5525 7275
rect 5525 7245 5555 7275
rect 5555 7245 5556 7275
rect 5524 7244 5556 7245
rect 5524 7195 5556 7196
rect 5524 7165 5525 7195
rect 5525 7165 5555 7195
rect 5555 7165 5556 7195
rect 5524 7164 5556 7165
rect 5524 7035 5556 7036
rect 5524 7005 5525 7035
rect 5525 7005 5555 7035
rect 5555 7005 5556 7035
rect 5524 7004 5556 7005
rect 5524 6955 5556 6956
rect 5524 6925 5525 6955
rect 5525 6925 5555 6955
rect 5555 6925 5556 6955
rect 5524 6924 5556 6925
rect 5524 6795 5556 6796
rect 5524 6765 5525 6795
rect 5525 6765 5555 6795
rect 5555 6765 5556 6795
rect 5524 6764 5556 6765
rect 5524 6715 5556 6716
rect 5524 6685 5525 6715
rect 5525 6685 5555 6715
rect 5555 6685 5556 6715
rect 5524 6684 5556 6685
rect 5524 6635 5556 6636
rect 5524 6605 5525 6635
rect 5525 6605 5555 6635
rect 5555 6605 5556 6635
rect 5524 6604 5556 6605
rect 5524 6555 5556 6556
rect 5524 6525 5525 6555
rect 5525 6525 5555 6555
rect 5555 6525 5556 6555
rect 5524 6524 5556 6525
rect 5524 6475 5556 6476
rect 5524 6445 5525 6475
rect 5525 6445 5555 6475
rect 5555 6445 5556 6475
rect 5524 6444 5556 6445
rect 5524 6315 5556 6316
rect 5524 6285 5525 6315
rect 5525 6285 5555 6315
rect 5555 6285 5556 6315
rect 5524 6284 5556 6285
rect 5524 6235 5556 6236
rect 5524 6205 5525 6235
rect 5525 6205 5555 6235
rect 5555 6205 5556 6235
rect 5524 6204 5556 6205
rect 5524 6155 5556 6156
rect 5524 6125 5525 6155
rect 5525 6125 5555 6155
rect 5555 6125 5556 6155
rect 5524 6124 5556 6125
rect 5524 5995 5556 5996
rect 5524 5965 5525 5995
rect 5525 5965 5555 5995
rect 5555 5965 5556 5995
rect 5524 5964 5556 5965
rect 5524 5835 5556 5836
rect 5524 5805 5525 5835
rect 5525 5805 5555 5835
rect 5555 5805 5556 5835
rect 5524 5804 5556 5805
rect 5524 5755 5556 5756
rect 5524 5725 5525 5755
rect 5525 5725 5555 5755
rect 5555 5725 5556 5755
rect 5524 5724 5556 5725
rect 5524 5675 5556 5676
rect 5524 5645 5525 5675
rect 5525 5645 5555 5675
rect 5555 5645 5556 5675
rect 5524 5644 5556 5645
rect 5524 5595 5556 5596
rect 5524 5565 5525 5595
rect 5525 5565 5555 5595
rect 5555 5565 5556 5595
rect 5524 5564 5556 5565
rect 5524 5515 5556 5516
rect 5524 5485 5525 5515
rect 5525 5485 5555 5515
rect 5555 5485 5556 5515
rect 5524 5484 5556 5485
rect 5524 5435 5556 5436
rect 5524 5405 5525 5435
rect 5525 5405 5555 5435
rect 5555 5405 5556 5435
rect 5524 5404 5556 5405
rect 5524 5355 5556 5356
rect 5524 5325 5525 5355
rect 5525 5325 5555 5355
rect 5555 5325 5556 5355
rect 5524 5324 5556 5325
rect 5524 5275 5556 5276
rect 5524 5245 5525 5275
rect 5525 5245 5555 5275
rect 5555 5245 5556 5275
rect 5524 5244 5556 5245
rect 5524 5195 5556 5196
rect 5524 5165 5525 5195
rect 5525 5165 5555 5195
rect 5555 5165 5556 5195
rect 5524 5164 5556 5165
rect 5524 5115 5556 5116
rect 5524 5085 5525 5115
rect 5525 5085 5555 5115
rect 5555 5085 5556 5115
rect 5524 5084 5556 5085
rect 5524 5035 5556 5036
rect 5524 5005 5525 5035
rect 5525 5005 5555 5035
rect 5555 5005 5556 5035
rect 5524 5004 5556 5005
rect 5524 4955 5556 4956
rect 5524 4925 5525 4955
rect 5525 4925 5555 4955
rect 5555 4925 5556 4955
rect 5524 4924 5556 4925
rect 5524 4875 5556 4876
rect 5524 4845 5525 4875
rect 5525 4845 5555 4875
rect 5555 4845 5556 4875
rect 5524 4844 5556 4845
rect 5524 4795 5556 4796
rect 5524 4765 5525 4795
rect 5525 4765 5555 4795
rect 5555 4765 5556 4795
rect 5524 4764 5556 4765
rect 5524 4635 5556 4636
rect 5524 4605 5525 4635
rect 5525 4605 5555 4635
rect 5555 4605 5556 4635
rect 5524 4604 5556 4605
rect 5524 4555 5556 4556
rect 5524 4525 5525 4555
rect 5525 4525 5555 4555
rect 5555 4525 5556 4555
rect 5524 4524 5556 4525
rect 5524 4395 5556 4396
rect 5524 4365 5525 4395
rect 5525 4365 5555 4395
rect 5555 4365 5556 4395
rect 5524 4364 5556 4365
rect 5524 4315 5556 4316
rect 5524 4285 5525 4315
rect 5525 4285 5555 4315
rect 5555 4285 5556 4315
rect 5524 4284 5556 4285
rect 5524 4235 5556 4236
rect 5524 4205 5525 4235
rect 5525 4205 5555 4235
rect 5555 4205 5556 4235
rect 5524 4204 5556 4205
rect 5524 4155 5556 4156
rect 5524 4125 5525 4155
rect 5525 4125 5555 4155
rect 5555 4125 5556 4155
rect 5524 4124 5556 4125
rect 5524 4075 5556 4076
rect 5524 4045 5525 4075
rect 5525 4045 5555 4075
rect 5555 4045 5556 4075
rect 5524 4044 5556 4045
rect 5524 3915 5556 3916
rect 5524 3885 5525 3915
rect 5525 3885 5555 3915
rect 5555 3885 5556 3915
rect 5524 3884 5556 3885
rect 5524 3835 5556 3836
rect 5524 3805 5525 3835
rect 5525 3805 5555 3835
rect 5555 3805 5556 3835
rect 5524 3804 5556 3805
rect 5524 3755 5556 3756
rect 5524 3725 5525 3755
rect 5525 3725 5555 3755
rect 5555 3725 5556 3755
rect 5524 3724 5556 3725
rect 5524 3595 5556 3596
rect 5524 3565 5525 3595
rect 5525 3565 5555 3595
rect 5555 3565 5556 3595
rect 5524 3564 5556 3565
rect 5524 3435 5556 3436
rect 5524 3405 5525 3435
rect 5525 3405 5555 3435
rect 5555 3405 5556 3435
rect 5524 3404 5556 3405
rect 5524 3355 5556 3356
rect 5524 3325 5525 3355
rect 5525 3325 5555 3355
rect 5555 3325 5556 3355
rect 5524 3324 5556 3325
rect 5524 3275 5556 3276
rect 5524 3245 5525 3275
rect 5525 3245 5555 3275
rect 5555 3245 5556 3275
rect 5524 3244 5556 3245
rect 5524 3195 5556 3196
rect 5524 3165 5525 3195
rect 5525 3165 5555 3195
rect 5555 3165 5556 3195
rect 5524 3164 5556 3165
rect 5524 3115 5556 3116
rect 5524 3085 5525 3115
rect 5525 3085 5555 3115
rect 5555 3085 5556 3115
rect 5524 3084 5556 3085
rect 5524 3035 5556 3036
rect 5524 3005 5525 3035
rect 5525 3005 5555 3035
rect 5555 3005 5556 3035
rect 5524 3004 5556 3005
rect 5524 2955 5556 2956
rect 5524 2925 5525 2955
rect 5525 2925 5555 2955
rect 5555 2925 5556 2955
rect 5524 2924 5556 2925
rect 5524 2875 5556 2876
rect 5524 2845 5525 2875
rect 5525 2845 5555 2875
rect 5555 2845 5556 2875
rect 5524 2844 5556 2845
rect 5524 2795 5556 2796
rect 5524 2765 5525 2795
rect 5525 2765 5555 2795
rect 5555 2765 5556 2795
rect 5524 2764 5556 2765
rect 5524 2715 5556 2716
rect 5524 2685 5525 2715
rect 5525 2685 5555 2715
rect 5555 2685 5556 2715
rect 5524 2684 5556 2685
rect 5524 2635 5556 2636
rect 5524 2605 5525 2635
rect 5525 2605 5555 2635
rect 5555 2605 5556 2635
rect 5524 2604 5556 2605
rect 5524 2555 5556 2556
rect 5524 2525 5525 2555
rect 5525 2525 5555 2555
rect 5555 2525 5556 2555
rect 5524 2524 5556 2525
rect 5524 2475 5556 2476
rect 5524 2445 5525 2475
rect 5525 2445 5555 2475
rect 5555 2445 5556 2475
rect 5524 2444 5556 2445
rect 5524 2395 5556 2396
rect 5524 2365 5525 2395
rect 5525 2365 5555 2395
rect 5555 2365 5556 2395
rect 5524 2364 5556 2365
rect 5524 2235 5556 2236
rect 5524 2205 5525 2235
rect 5525 2205 5555 2235
rect 5555 2205 5556 2235
rect 5524 2204 5556 2205
rect 5524 2155 5556 2156
rect 5524 2125 5525 2155
rect 5525 2125 5555 2155
rect 5555 2125 5556 2155
rect 5524 2124 5556 2125
rect 5524 2075 5556 2076
rect 5524 2045 5525 2075
rect 5525 2045 5555 2075
rect 5555 2045 5556 2075
rect 5524 2044 5556 2045
rect 5524 1995 5556 1996
rect 5524 1965 5525 1995
rect 5525 1965 5555 1995
rect 5555 1965 5556 1995
rect 5524 1964 5556 1965
rect 5524 1915 5556 1916
rect 5524 1885 5525 1915
rect 5525 1885 5555 1915
rect 5555 1885 5556 1915
rect 5524 1884 5556 1885
rect 5524 1835 5556 1836
rect 5524 1805 5525 1835
rect 5525 1805 5555 1835
rect 5555 1805 5556 1835
rect 5524 1804 5556 1805
rect 5524 1755 5556 1756
rect 5524 1725 5525 1755
rect 5525 1725 5555 1755
rect 5555 1725 5556 1755
rect 5524 1724 5556 1725
rect 5524 1675 5556 1676
rect 5524 1645 5525 1675
rect 5525 1645 5555 1675
rect 5555 1645 5556 1675
rect 5524 1644 5556 1645
rect 5524 1515 5556 1516
rect 5524 1485 5525 1515
rect 5525 1485 5555 1515
rect 5555 1485 5556 1515
rect 5524 1484 5556 1485
rect 5524 1435 5556 1436
rect 5524 1405 5525 1435
rect 5525 1405 5555 1435
rect 5555 1405 5556 1435
rect 5524 1404 5556 1405
rect 5524 1355 5556 1356
rect 5524 1325 5525 1355
rect 5525 1325 5555 1355
rect 5555 1325 5556 1355
rect 5524 1324 5556 1325
rect 5524 1195 5556 1196
rect 5524 1165 5525 1195
rect 5525 1165 5555 1195
rect 5555 1165 5556 1195
rect 5524 1164 5556 1165
rect 5524 1115 5556 1116
rect 5524 1085 5525 1115
rect 5525 1085 5555 1115
rect 5555 1085 5556 1115
rect 5524 1084 5556 1085
rect 5524 1035 5556 1036
rect 5524 1005 5525 1035
rect 5525 1005 5555 1035
rect 5555 1005 5556 1035
rect 5524 1004 5556 1005
rect 5524 955 5556 956
rect 5524 925 5525 955
rect 5525 925 5555 955
rect 5555 925 5556 955
rect 5524 924 5556 925
rect 5524 875 5556 876
rect 5524 845 5525 875
rect 5525 845 5555 875
rect 5555 845 5556 875
rect 5524 844 5556 845
rect 5524 795 5556 796
rect 5524 765 5525 795
rect 5525 765 5555 795
rect 5555 765 5556 795
rect 5524 764 5556 765
rect 5524 595 5556 596
rect 5524 565 5525 595
rect 5525 565 5555 595
rect 5555 565 5556 595
rect 5524 564 5556 565
rect 5524 515 5556 516
rect 5524 485 5525 515
rect 5525 485 5555 515
rect 5555 485 5556 515
rect 5524 484 5556 485
rect 5524 355 5556 356
rect 5524 325 5525 355
rect 5525 325 5555 355
rect 5555 325 5556 355
rect 5524 324 5556 325
rect 5524 275 5556 276
rect 5524 245 5525 275
rect 5525 245 5555 275
rect 5555 245 5556 275
rect 5524 244 5556 245
rect 5524 195 5556 196
rect 5524 165 5525 195
rect 5525 165 5555 195
rect 5555 165 5556 195
rect 5524 164 5556 165
rect 5524 115 5556 116
rect 5524 85 5525 115
rect 5525 85 5555 115
rect 5555 85 5556 115
rect 5524 84 5556 85
rect 5524 35 5556 36
rect 5524 5 5525 35
rect 5525 5 5555 35
rect 5555 5 5556 35
rect 5524 4 5556 5
rect 5844 16644 5876 16836
rect 5684 16595 5716 16596
rect 5684 16565 5685 16595
rect 5685 16565 5715 16595
rect 5715 16565 5716 16595
rect 5684 16564 5716 16565
rect 5684 16515 5716 16516
rect 5684 16485 5685 16515
rect 5685 16485 5715 16515
rect 5715 16485 5716 16515
rect 5684 16484 5716 16485
rect 5684 16435 5716 16436
rect 5684 16405 5685 16435
rect 5685 16405 5715 16435
rect 5715 16405 5716 16435
rect 5684 16404 5716 16405
rect 5684 16355 5716 16356
rect 5684 16325 5685 16355
rect 5685 16325 5715 16355
rect 5715 16325 5716 16355
rect 5684 16324 5716 16325
rect 5684 16275 5716 16276
rect 5684 16245 5685 16275
rect 5685 16245 5715 16275
rect 5715 16245 5716 16275
rect 5684 16244 5716 16245
rect 5684 16195 5716 16196
rect 5684 16165 5685 16195
rect 5685 16165 5715 16195
rect 5715 16165 5716 16195
rect 5684 16164 5716 16165
rect 5684 16115 5716 16116
rect 5684 16085 5685 16115
rect 5685 16085 5715 16115
rect 5715 16085 5716 16115
rect 5684 16084 5716 16085
rect 5684 16035 5716 16036
rect 5684 16005 5685 16035
rect 5685 16005 5715 16035
rect 5715 16005 5716 16035
rect 5684 16004 5716 16005
rect 5684 15955 5716 15956
rect 5684 15925 5685 15955
rect 5685 15925 5715 15955
rect 5715 15925 5716 15955
rect 5684 15924 5716 15925
rect 5684 15435 5716 15436
rect 5684 15405 5685 15435
rect 5685 15405 5715 15435
rect 5715 15405 5716 15435
rect 5684 15404 5716 15405
rect 5684 15355 5716 15356
rect 5684 15325 5685 15355
rect 5685 15325 5715 15355
rect 5715 15325 5716 15355
rect 5684 15324 5716 15325
rect 5684 15275 5716 15276
rect 5684 15245 5685 15275
rect 5685 15245 5715 15275
rect 5715 15245 5716 15275
rect 5684 15244 5716 15245
rect 5684 15195 5716 15196
rect 5684 15165 5685 15195
rect 5685 15165 5715 15195
rect 5715 15165 5716 15195
rect 5684 15164 5716 15165
rect 5684 15115 5716 15116
rect 5684 15085 5685 15115
rect 5685 15085 5715 15115
rect 5715 15085 5716 15115
rect 5684 15084 5716 15085
rect 5684 14955 5716 14956
rect 5684 14925 5685 14955
rect 5685 14925 5715 14955
rect 5715 14925 5716 14955
rect 5684 14924 5716 14925
rect 5684 14875 5716 14876
rect 5684 14845 5685 14875
rect 5685 14845 5715 14875
rect 5715 14845 5716 14875
rect 5684 14844 5716 14845
rect 5684 14795 5716 14796
rect 5684 14765 5685 14795
rect 5685 14765 5715 14795
rect 5715 14765 5716 14795
rect 5684 14764 5716 14765
rect 5684 14715 5716 14716
rect 5684 14685 5685 14715
rect 5685 14685 5715 14715
rect 5715 14685 5716 14715
rect 5684 14684 5716 14685
rect 5684 14555 5716 14556
rect 5684 14525 5685 14555
rect 5685 14525 5715 14555
rect 5715 14525 5716 14555
rect 5684 14524 5716 14525
rect 5684 14475 5716 14476
rect 5684 14445 5685 14475
rect 5685 14445 5715 14475
rect 5715 14445 5716 14475
rect 5684 14444 5716 14445
rect 5684 13995 5716 13996
rect 5684 13965 5685 13995
rect 5685 13965 5715 13995
rect 5715 13965 5716 13995
rect 5684 13964 5716 13965
rect 5684 13795 5716 13796
rect 5684 13765 5685 13795
rect 5685 13765 5715 13795
rect 5715 13765 5716 13795
rect 5684 13764 5716 13765
rect 5684 13715 5716 13716
rect 5684 13685 5685 13715
rect 5685 13685 5715 13715
rect 5715 13685 5716 13715
rect 5684 13684 5716 13685
rect 5684 13635 5716 13636
rect 5684 13605 5685 13635
rect 5685 13605 5715 13635
rect 5715 13605 5716 13635
rect 5684 13604 5716 13605
rect 5684 13475 5716 13476
rect 5684 13445 5685 13475
rect 5685 13445 5715 13475
rect 5715 13445 5716 13475
rect 5684 13444 5716 13445
rect 5684 13395 5716 13396
rect 5684 13365 5685 13395
rect 5685 13365 5715 13395
rect 5715 13365 5716 13395
rect 5684 13364 5716 13365
rect 5684 13315 5716 13316
rect 5684 13285 5685 13315
rect 5685 13285 5715 13315
rect 5715 13285 5716 13315
rect 5684 13284 5716 13285
rect 5684 13235 5716 13236
rect 5684 13205 5685 13235
rect 5685 13205 5715 13235
rect 5715 13205 5716 13235
rect 5684 13204 5716 13205
rect 5684 13075 5716 13076
rect 5684 13045 5685 13075
rect 5685 13045 5715 13075
rect 5715 13045 5716 13075
rect 5684 13044 5716 13045
rect 5684 12995 5716 12996
rect 5684 12965 5685 12995
rect 5685 12965 5715 12995
rect 5715 12965 5716 12995
rect 5684 12964 5716 12965
rect 5684 12515 5716 12516
rect 5684 12485 5685 12515
rect 5685 12485 5715 12515
rect 5715 12485 5716 12515
rect 5684 12484 5716 12485
rect 5684 12315 5716 12316
rect 5684 12285 5685 12315
rect 5685 12285 5715 12315
rect 5715 12285 5716 12315
rect 5684 12284 5716 12285
rect 5684 12235 5716 12236
rect 5684 12205 5685 12235
rect 5685 12205 5715 12235
rect 5715 12205 5716 12235
rect 5684 12204 5716 12205
rect 5684 12155 5716 12156
rect 5684 12125 5685 12155
rect 5685 12125 5715 12155
rect 5715 12125 5716 12155
rect 5684 12124 5716 12125
rect 5684 12075 5716 12076
rect 5684 12045 5685 12075
rect 5685 12045 5715 12075
rect 5715 12045 5716 12075
rect 5684 12044 5716 12045
rect 5684 11995 5716 11996
rect 5684 11965 5685 11995
rect 5685 11965 5715 11995
rect 5715 11965 5716 11995
rect 5684 11964 5716 11965
rect 5684 11915 5716 11916
rect 5684 11885 5685 11915
rect 5685 11885 5715 11915
rect 5715 11885 5716 11915
rect 5684 11884 5716 11885
rect 5684 11835 5716 11836
rect 5684 11805 5685 11835
rect 5685 11805 5715 11835
rect 5715 11805 5716 11835
rect 5684 11804 5716 11805
rect 5684 11755 5716 11756
rect 5684 11725 5685 11755
rect 5685 11725 5715 11755
rect 5715 11725 5716 11755
rect 5684 11724 5716 11725
rect 5684 11675 5716 11676
rect 5684 11645 5685 11675
rect 5685 11645 5715 11675
rect 5715 11645 5716 11675
rect 5684 11644 5716 11645
rect 5684 11595 5716 11596
rect 5684 11565 5685 11595
rect 5685 11565 5715 11595
rect 5715 11565 5716 11595
rect 5684 11564 5716 11565
rect 5684 11515 5716 11516
rect 5684 11485 5685 11515
rect 5685 11485 5715 11515
rect 5715 11485 5716 11515
rect 5684 11484 5716 11485
rect 5684 11435 5716 11436
rect 5684 11405 5685 11435
rect 5685 11405 5715 11435
rect 5715 11405 5716 11435
rect 5684 11404 5716 11405
rect 5684 11355 5716 11356
rect 5684 11325 5685 11355
rect 5685 11325 5715 11355
rect 5715 11325 5716 11355
rect 5684 11324 5716 11325
rect 5684 11195 5716 11196
rect 5684 11165 5685 11195
rect 5685 11165 5715 11195
rect 5715 11165 5716 11195
rect 5684 11164 5716 11165
rect 5684 11115 5716 11116
rect 5684 11085 5685 11115
rect 5685 11085 5715 11115
rect 5715 11085 5716 11115
rect 5684 11084 5716 11085
rect 5684 11035 5716 11036
rect 5684 11005 5685 11035
rect 5685 11005 5715 11035
rect 5715 11005 5716 11035
rect 5684 11004 5716 11005
rect 5684 10875 5716 10876
rect 5684 10845 5685 10875
rect 5685 10845 5715 10875
rect 5715 10845 5716 10875
rect 5684 10844 5716 10845
rect 5684 10715 5716 10716
rect 5684 10685 5685 10715
rect 5685 10685 5715 10715
rect 5715 10685 5716 10715
rect 5684 10684 5716 10685
rect 5684 10635 5716 10636
rect 5684 10605 5685 10635
rect 5685 10605 5715 10635
rect 5715 10605 5716 10635
rect 5684 10604 5716 10605
rect 5684 10475 5716 10476
rect 5684 10445 5685 10475
rect 5685 10445 5715 10475
rect 5715 10445 5716 10475
rect 5684 10444 5716 10445
rect 5684 10315 5716 10316
rect 5684 10285 5685 10315
rect 5685 10285 5715 10315
rect 5715 10285 5716 10315
rect 5684 10284 5716 10285
rect 5684 10235 5716 10236
rect 5684 10205 5685 10235
rect 5685 10205 5715 10235
rect 5715 10205 5716 10235
rect 5684 10204 5716 10205
rect 5684 10155 5716 10156
rect 5684 10125 5685 10155
rect 5685 10125 5715 10155
rect 5715 10125 5716 10155
rect 5684 10124 5716 10125
rect 5684 10075 5716 10076
rect 5684 10045 5685 10075
rect 5685 10045 5715 10075
rect 5715 10045 5716 10075
rect 5684 10044 5716 10045
rect 5684 9995 5716 9996
rect 5684 9965 5685 9995
rect 5685 9965 5715 9995
rect 5715 9965 5716 9995
rect 5684 9964 5716 9965
rect 5684 9915 5716 9916
rect 5684 9885 5685 9915
rect 5685 9885 5715 9915
rect 5715 9885 5716 9915
rect 5684 9884 5716 9885
rect 5684 9835 5716 9836
rect 5684 9805 5685 9835
rect 5685 9805 5715 9835
rect 5715 9805 5716 9835
rect 5684 9804 5716 9805
rect 5684 9755 5716 9756
rect 5684 9725 5685 9755
rect 5685 9725 5715 9755
rect 5715 9725 5716 9755
rect 5684 9724 5716 9725
rect 5684 9675 5716 9676
rect 5684 9645 5685 9675
rect 5685 9645 5715 9675
rect 5715 9645 5716 9675
rect 5684 9644 5716 9645
rect 5684 9595 5716 9596
rect 5684 9565 5685 9595
rect 5685 9565 5715 9595
rect 5715 9565 5716 9595
rect 5684 9564 5716 9565
rect 5684 9515 5716 9516
rect 5684 9485 5685 9515
rect 5685 9485 5715 9515
rect 5715 9485 5716 9515
rect 5684 9484 5716 9485
rect 5684 9435 5716 9436
rect 5684 9405 5685 9435
rect 5685 9405 5715 9435
rect 5715 9405 5716 9435
rect 5684 9404 5716 9405
rect 5684 9355 5716 9356
rect 5684 9325 5685 9355
rect 5685 9325 5715 9355
rect 5715 9325 5716 9355
rect 5684 9324 5716 9325
rect 5684 9275 5716 9276
rect 5684 9245 5685 9275
rect 5685 9245 5715 9275
rect 5715 9245 5716 9275
rect 5684 9244 5716 9245
rect 5684 9115 5716 9116
rect 5684 9085 5685 9115
rect 5685 9085 5715 9115
rect 5715 9085 5716 9115
rect 5684 9084 5716 9085
rect 5684 9035 5716 9036
rect 5684 9005 5685 9035
rect 5685 9005 5715 9035
rect 5715 9005 5716 9035
rect 5684 9004 5716 9005
rect 5684 8955 5716 8956
rect 5684 8925 5685 8955
rect 5685 8925 5715 8955
rect 5715 8925 5716 8955
rect 5684 8924 5716 8925
rect 5684 8635 5716 8636
rect 5684 8605 5685 8635
rect 5685 8605 5715 8635
rect 5715 8605 5716 8635
rect 5684 8604 5716 8605
rect 5684 8555 5716 8556
rect 5684 8525 5685 8555
rect 5685 8525 5715 8555
rect 5715 8525 5716 8555
rect 5684 8524 5716 8525
rect 5684 8395 5716 8396
rect 5684 8365 5685 8395
rect 5685 8365 5715 8395
rect 5715 8365 5716 8395
rect 5684 8364 5716 8365
rect 5684 8235 5716 8236
rect 5684 8205 5685 8235
rect 5685 8205 5715 8235
rect 5715 8205 5716 8235
rect 5684 8204 5716 8205
rect 5684 8155 5716 8156
rect 5684 8125 5685 8155
rect 5685 8125 5715 8155
rect 5715 8125 5716 8155
rect 5684 8124 5716 8125
rect 5684 8075 5716 8076
rect 5684 8045 5685 8075
rect 5685 8045 5715 8075
rect 5715 8045 5716 8075
rect 5684 8044 5716 8045
rect 5684 7995 5716 7996
rect 5684 7965 5685 7995
rect 5685 7965 5715 7995
rect 5715 7965 5716 7995
rect 5684 7964 5716 7965
rect 5684 7915 5716 7916
rect 5684 7885 5685 7915
rect 5685 7885 5715 7915
rect 5715 7885 5716 7915
rect 5684 7884 5716 7885
rect 5684 7835 5716 7836
rect 5684 7805 5685 7835
rect 5685 7805 5715 7835
rect 5715 7805 5716 7835
rect 5684 7804 5716 7805
rect 5684 7755 5716 7756
rect 5684 7725 5685 7755
rect 5685 7725 5715 7755
rect 5715 7725 5716 7755
rect 5684 7724 5716 7725
rect 5684 7675 5716 7676
rect 5684 7645 5685 7675
rect 5685 7645 5715 7675
rect 5715 7645 5716 7675
rect 5684 7644 5716 7645
rect 5684 7595 5716 7596
rect 5684 7565 5685 7595
rect 5685 7565 5715 7595
rect 5715 7565 5716 7595
rect 5684 7564 5716 7565
rect 5684 7515 5716 7516
rect 5684 7485 5685 7515
rect 5685 7485 5715 7515
rect 5715 7485 5716 7515
rect 5684 7484 5716 7485
rect 5684 7435 5716 7436
rect 5684 7405 5685 7435
rect 5685 7405 5715 7435
rect 5715 7405 5716 7435
rect 5684 7404 5716 7405
rect 5684 7355 5716 7356
rect 5684 7325 5685 7355
rect 5685 7325 5715 7355
rect 5715 7325 5716 7355
rect 5684 7324 5716 7325
rect 5684 7275 5716 7276
rect 5684 7245 5685 7275
rect 5685 7245 5715 7275
rect 5715 7245 5716 7275
rect 5684 7244 5716 7245
rect 5684 7195 5716 7196
rect 5684 7165 5685 7195
rect 5685 7165 5715 7195
rect 5715 7165 5716 7195
rect 5684 7164 5716 7165
rect 5684 7035 5716 7036
rect 5684 7005 5685 7035
rect 5685 7005 5715 7035
rect 5715 7005 5716 7035
rect 5684 7004 5716 7005
rect 5684 6955 5716 6956
rect 5684 6925 5685 6955
rect 5685 6925 5715 6955
rect 5715 6925 5716 6955
rect 5684 6924 5716 6925
rect 5684 6795 5716 6796
rect 5684 6765 5685 6795
rect 5685 6765 5715 6795
rect 5715 6765 5716 6795
rect 5684 6764 5716 6765
rect 5684 6715 5716 6716
rect 5684 6685 5685 6715
rect 5685 6685 5715 6715
rect 5715 6685 5716 6715
rect 5684 6684 5716 6685
rect 5684 6635 5716 6636
rect 5684 6605 5685 6635
rect 5685 6605 5715 6635
rect 5715 6605 5716 6635
rect 5684 6604 5716 6605
rect 5684 6555 5716 6556
rect 5684 6525 5685 6555
rect 5685 6525 5715 6555
rect 5715 6525 5716 6555
rect 5684 6524 5716 6525
rect 5684 6475 5716 6476
rect 5684 6445 5685 6475
rect 5685 6445 5715 6475
rect 5715 6445 5716 6475
rect 5684 6444 5716 6445
rect 5684 6315 5716 6316
rect 5684 6285 5685 6315
rect 5685 6285 5715 6315
rect 5715 6285 5716 6315
rect 5684 6284 5716 6285
rect 5684 6235 5716 6236
rect 5684 6205 5685 6235
rect 5685 6205 5715 6235
rect 5715 6205 5716 6235
rect 5684 6204 5716 6205
rect 5684 6155 5716 6156
rect 5684 6125 5685 6155
rect 5685 6125 5715 6155
rect 5715 6125 5716 6155
rect 5684 6124 5716 6125
rect 5684 5995 5716 5996
rect 5684 5965 5685 5995
rect 5685 5965 5715 5995
rect 5715 5965 5716 5995
rect 5684 5964 5716 5965
rect 5684 5835 5716 5836
rect 5684 5805 5685 5835
rect 5685 5805 5715 5835
rect 5715 5805 5716 5835
rect 5684 5804 5716 5805
rect 5684 5755 5716 5756
rect 5684 5725 5685 5755
rect 5685 5725 5715 5755
rect 5715 5725 5716 5755
rect 5684 5724 5716 5725
rect 5684 5675 5716 5676
rect 5684 5645 5685 5675
rect 5685 5645 5715 5675
rect 5715 5645 5716 5675
rect 5684 5644 5716 5645
rect 5684 5595 5716 5596
rect 5684 5565 5685 5595
rect 5685 5565 5715 5595
rect 5715 5565 5716 5595
rect 5684 5564 5716 5565
rect 5684 5515 5716 5516
rect 5684 5485 5685 5515
rect 5685 5485 5715 5515
rect 5715 5485 5716 5515
rect 5684 5484 5716 5485
rect 5684 5435 5716 5436
rect 5684 5405 5685 5435
rect 5685 5405 5715 5435
rect 5715 5405 5716 5435
rect 5684 5404 5716 5405
rect 5684 5355 5716 5356
rect 5684 5325 5685 5355
rect 5685 5325 5715 5355
rect 5715 5325 5716 5355
rect 5684 5324 5716 5325
rect 5684 5275 5716 5276
rect 5684 5245 5685 5275
rect 5685 5245 5715 5275
rect 5715 5245 5716 5275
rect 5684 5244 5716 5245
rect 5684 5195 5716 5196
rect 5684 5165 5685 5195
rect 5685 5165 5715 5195
rect 5715 5165 5716 5195
rect 5684 5164 5716 5165
rect 5684 5115 5716 5116
rect 5684 5085 5685 5115
rect 5685 5085 5715 5115
rect 5715 5085 5716 5115
rect 5684 5084 5716 5085
rect 5684 5035 5716 5036
rect 5684 5005 5685 5035
rect 5685 5005 5715 5035
rect 5715 5005 5716 5035
rect 5684 5004 5716 5005
rect 5684 4955 5716 4956
rect 5684 4925 5685 4955
rect 5685 4925 5715 4955
rect 5715 4925 5716 4955
rect 5684 4924 5716 4925
rect 5684 4875 5716 4876
rect 5684 4845 5685 4875
rect 5685 4845 5715 4875
rect 5715 4845 5716 4875
rect 5684 4844 5716 4845
rect 5684 4795 5716 4796
rect 5684 4765 5685 4795
rect 5685 4765 5715 4795
rect 5715 4765 5716 4795
rect 5684 4764 5716 4765
rect 5684 4635 5716 4636
rect 5684 4605 5685 4635
rect 5685 4605 5715 4635
rect 5715 4605 5716 4635
rect 5684 4604 5716 4605
rect 5684 4555 5716 4556
rect 5684 4525 5685 4555
rect 5685 4525 5715 4555
rect 5715 4525 5716 4555
rect 5684 4524 5716 4525
rect 5684 4395 5716 4396
rect 5684 4365 5685 4395
rect 5685 4365 5715 4395
rect 5715 4365 5716 4395
rect 5684 4364 5716 4365
rect 5684 4315 5716 4316
rect 5684 4285 5685 4315
rect 5685 4285 5715 4315
rect 5715 4285 5716 4315
rect 5684 4284 5716 4285
rect 5684 4235 5716 4236
rect 5684 4205 5685 4235
rect 5685 4205 5715 4235
rect 5715 4205 5716 4235
rect 5684 4204 5716 4205
rect 5684 4155 5716 4156
rect 5684 4125 5685 4155
rect 5685 4125 5715 4155
rect 5715 4125 5716 4155
rect 5684 4124 5716 4125
rect 5684 4075 5716 4076
rect 5684 4045 5685 4075
rect 5685 4045 5715 4075
rect 5715 4045 5716 4075
rect 5684 4044 5716 4045
rect 5684 3915 5716 3916
rect 5684 3885 5685 3915
rect 5685 3885 5715 3915
rect 5715 3885 5716 3915
rect 5684 3884 5716 3885
rect 5684 3835 5716 3836
rect 5684 3805 5685 3835
rect 5685 3805 5715 3835
rect 5715 3805 5716 3835
rect 5684 3804 5716 3805
rect 5684 3755 5716 3756
rect 5684 3725 5685 3755
rect 5685 3725 5715 3755
rect 5715 3725 5716 3755
rect 5684 3724 5716 3725
rect 5684 3595 5716 3596
rect 5684 3565 5685 3595
rect 5685 3565 5715 3595
rect 5715 3565 5716 3595
rect 5684 3564 5716 3565
rect 5684 3435 5716 3436
rect 5684 3405 5685 3435
rect 5685 3405 5715 3435
rect 5715 3405 5716 3435
rect 5684 3404 5716 3405
rect 5684 3355 5716 3356
rect 5684 3325 5685 3355
rect 5685 3325 5715 3355
rect 5715 3325 5716 3355
rect 5684 3324 5716 3325
rect 5684 3275 5716 3276
rect 5684 3245 5685 3275
rect 5685 3245 5715 3275
rect 5715 3245 5716 3275
rect 5684 3244 5716 3245
rect 5684 3195 5716 3196
rect 5684 3165 5685 3195
rect 5685 3165 5715 3195
rect 5715 3165 5716 3195
rect 5684 3164 5716 3165
rect 5684 3115 5716 3116
rect 5684 3085 5685 3115
rect 5685 3085 5715 3115
rect 5715 3085 5716 3115
rect 5684 3084 5716 3085
rect 5684 3035 5716 3036
rect 5684 3005 5685 3035
rect 5685 3005 5715 3035
rect 5715 3005 5716 3035
rect 5684 3004 5716 3005
rect 5684 2955 5716 2956
rect 5684 2925 5685 2955
rect 5685 2925 5715 2955
rect 5715 2925 5716 2955
rect 5684 2924 5716 2925
rect 5684 2875 5716 2876
rect 5684 2845 5685 2875
rect 5685 2845 5715 2875
rect 5715 2845 5716 2875
rect 5684 2844 5716 2845
rect 5684 2795 5716 2796
rect 5684 2765 5685 2795
rect 5685 2765 5715 2795
rect 5715 2765 5716 2795
rect 5684 2764 5716 2765
rect 5684 2715 5716 2716
rect 5684 2685 5685 2715
rect 5685 2685 5715 2715
rect 5715 2685 5716 2715
rect 5684 2684 5716 2685
rect 5684 2635 5716 2636
rect 5684 2605 5685 2635
rect 5685 2605 5715 2635
rect 5715 2605 5716 2635
rect 5684 2604 5716 2605
rect 5684 2555 5716 2556
rect 5684 2525 5685 2555
rect 5685 2525 5715 2555
rect 5715 2525 5716 2555
rect 5684 2524 5716 2525
rect 5684 2475 5716 2476
rect 5684 2445 5685 2475
rect 5685 2445 5715 2475
rect 5715 2445 5716 2475
rect 5684 2444 5716 2445
rect 5684 2395 5716 2396
rect 5684 2365 5685 2395
rect 5685 2365 5715 2395
rect 5715 2365 5716 2395
rect 5684 2364 5716 2365
rect 5684 2235 5716 2236
rect 5684 2205 5685 2235
rect 5685 2205 5715 2235
rect 5715 2205 5716 2235
rect 5684 2204 5716 2205
rect 5684 2155 5716 2156
rect 5684 2125 5685 2155
rect 5685 2125 5715 2155
rect 5715 2125 5716 2155
rect 5684 2124 5716 2125
rect 5684 2075 5716 2076
rect 5684 2045 5685 2075
rect 5685 2045 5715 2075
rect 5715 2045 5716 2075
rect 5684 2044 5716 2045
rect 5684 1995 5716 1996
rect 5684 1965 5685 1995
rect 5685 1965 5715 1995
rect 5715 1965 5716 1995
rect 5684 1964 5716 1965
rect 5684 1915 5716 1916
rect 5684 1885 5685 1915
rect 5685 1885 5715 1915
rect 5715 1885 5716 1915
rect 5684 1884 5716 1885
rect 5684 1835 5716 1836
rect 5684 1805 5685 1835
rect 5685 1805 5715 1835
rect 5715 1805 5716 1835
rect 5684 1804 5716 1805
rect 5684 1755 5716 1756
rect 5684 1725 5685 1755
rect 5685 1725 5715 1755
rect 5715 1725 5716 1755
rect 5684 1724 5716 1725
rect 5684 1675 5716 1676
rect 5684 1645 5685 1675
rect 5685 1645 5715 1675
rect 5715 1645 5716 1675
rect 5684 1644 5716 1645
rect 5684 1515 5716 1516
rect 5684 1485 5685 1515
rect 5685 1485 5715 1515
rect 5715 1485 5716 1515
rect 5684 1484 5716 1485
rect 5684 1435 5716 1436
rect 5684 1405 5685 1435
rect 5685 1405 5715 1435
rect 5715 1405 5716 1435
rect 5684 1404 5716 1405
rect 5684 1355 5716 1356
rect 5684 1325 5685 1355
rect 5685 1325 5715 1355
rect 5715 1325 5716 1355
rect 5684 1324 5716 1325
rect 5684 1275 5716 1276
rect 5684 1245 5685 1275
rect 5685 1245 5715 1275
rect 5715 1245 5716 1275
rect 5684 1244 5716 1245
rect 5684 1195 5716 1196
rect 5684 1165 5685 1195
rect 5685 1165 5715 1195
rect 5715 1165 5716 1195
rect 5684 1164 5716 1165
rect 5684 1115 5716 1116
rect 5684 1085 5685 1115
rect 5685 1085 5715 1115
rect 5715 1085 5716 1115
rect 5684 1084 5716 1085
rect 5684 1035 5716 1036
rect 5684 1005 5685 1035
rect 5685 1005 5715 1035
rect 5715 1005 5716 1035
rect 5684 1004 5716 1005
rect 5684 955 5716 956
rect 5684 925 5685 955
rect 5685 925 5715 955
rect 5715 925 5716 955
rect 5684 924 5716 925
rect 5684 875 5716 876
rect 5684 845 5685 875
rect 5685 845 5715 875
rect 5715 845 5716 875
rect 5684 844 5716 845
rect 5684 795 5716 796
rect 5684 765 5685 795
rect 5685 765 5715 795
rect 5715 765 5716 795
rect 5684 764 5716 765
rect 5684 595 5716 596
rect 5684 565 5685 595
rect 5685 565 5715 595
rect 5715 565 5716 595
rect 5684 564 5716 565
rect 5684 515 5716 516
rect 5684 485 5685 515
rect 5685 485 5715 515
rect 5715 485 5716 515
rect 5684 484 5716 485
rect 5684 435 5716 436
rect 5684 405 5685 435
rect 5685 405 5715 435
rect 5715 405 5716 435
rect 5684 404 5716 405
rect 5684 355 5716 356
rect 5684 325 5685 355
rect 5685 325 5715 355
rect 5715 325 5716 355
rect 5684 324 5716 325
rect 5684 275 5716 276
rect 5684 245 5685 275
rect 5685 245 5715 275
rect 5715 245 5716 275
rect 5684 244 5716 245
rect 5684 195 5716 196
rect 5684 165 5685 195
rect 5685 165 5715 195
rect 5715 165 5716 195
rect 5684 164 5716 165
rect 5684 115 5716 116
rect 5684 85 5685 115
rect 5685 85 5715 115
rect 5715 85 5716 115
rect 5684 84 5716 85
rect 5684 35 5716 36
rect 5684 5 5685 35
rect 5685 5 5715 35
rect 5715 5 5716 35
rect 5684 4 5716 5
rect 6004 16644 6036 16836
rect 5844 16595 5876 16596
rect 5844 16565 5845 16595
rect 5845 16565 5875 16595
rect 5875 16565 5876 16595
rect 5844 16564 5876 16565
rect 5844 16515 5876 16516
rect 5844 16485 5845 16515
rect 5845 16485 5875 16515
rect 5875 16485 5876 16515
rect 5844 16484 5876 16485
rect 5844 16435 5876 16436
rect 5844 16405 5845 16435
rect 5845 16405 5875 16435
rect 5875 16405 5876 16435
rect 5844 16404 5876 16405
rect 5844 16355 5876 16356
rect 5844 16325 5845 16355
rect 5845 16325 5875 16355
rect 5875 16325 5876 16355
rect 5844 16324 5876 16325
rect 5844 16275 5876 16276
rect 5844 16245 5845 16275
rect 5845 16245 5875 16275
rect 5875 16245 5876 16275
rect 5844 16244 5876 16245
rect 5844 16195 5876 16196
rect 5844 16165 5845 16195
rect 5845 16165 5875 16195
rect 5875 16165 5876 16195
rect 5844 16164 5876 16165
rect 5844 16115 5876 16116
rect 5844 16085 5845 16115
rect 5845 16085 5875 16115
rect 5875 16085 5876 16115
rect 5844 16084 5876 16085
rect 5844 16035 5876 16036
rect 5844 16005 5845 16035
rect 5845 16005 5875 16035
rect 5875 16005 5876 16035
rect 5844 16004 5876 16005
rect 5844 15955 5876 15956
rect 5844 15925 5845 15955
rect 5845 15925 5875 15955
rect 5875 15925 5876 15955
rect 5844 15924 5876 15925
rect 5844 15435 5876 15436
rect 5844 15405 5845 15435
rect 5845 15405 5875 15435
rect 5875 15405 5876 15435
rect 5844 15404 5876 15405
rect 5844 15355 5876 15356
rect 5844 15325 5845 15355
rect 5845 15325 5875 15355
rect 5875 15325 5876 15355
rect 5844 15324 5876 15325
rect 5844 15275 5876 15276
rect 5844 15245 5845 15275
rect 5845 15245 5875 15275
rect 5875 15245 5876 15275
rect 5844 15244 5876 15245
rect 5844 15195 5876 15196
rect 5844 15165 5845 15195
rect 5845 15165 5875 15195
rect 5875 15165 5876 15195
rect 5844 15164 5876 15165
rect 5844 15115 5876 15116
rect 5844 15085 5845 15115
rect 5845 15085 5875 15115
rect 5875 15085 5876 15115
rect 5844 15084 5876 15085
rect 5844 14955 5876 14956
rect 5844 14925 5845 14955
rect 5845 14925 5875 14955
rect 5875 14925 5876 14955
rect 5844 14924 5876 14925
rect 5844 14875 5876 14876
rect 5844 14845 5845 14875
rect 5845 14845 5875 14875
rect 5875 14845 5876 14875
rect 5844 14844 5876 14845
rect 5844 14795 5876 14796
rect 5844 14765 5845 14795
rect 5845 14765 5875 14795
rect 5875 14765 5876 14795
rect 5844 14764 5876 14765
rect 5844 14715 5876 14716
rect 5844 14685 5845 14715
rect 5845 14685 5875 14715
rect 5875 14685 5876 14715
rect 5844 14684 5876 14685
rect 5844 14555 5876 14556
rect 5844 14525 5845 14555
rect 5845 14525 5875 14555
rect 5875 14525 5876 14555
rect 5844 14524 5876 14525
rect 5844 14475 5876 14476
rect 5844 14445 5845 14475
rect 5845 14445 5875 14475
rect 5875 14445 5876 14475
rect 5844 14444 5876 14445
rect 5844 13995 5876 13996
rect 5844 13965 5845 13995
rect 5845 13965 5875 13995
rect 5875 13965 5876 13995
rect 5844 13964 5876 13965
rect 5844 13875 5876 13876
rect 5844 13845 5845 13875
rect 5845 13845 5875 13875
rect 5875 13845 5876 13875
rect 5844 13844 5876 13845
rect 5844 13795 5876 13796
rect 5844 13765 5845 13795
rect 5845 13765 5875 13795
rect 5875 13765 5876 13795
rect 5844 13764 5876 13765
rect 5844 13715 5876 13716
rect 5844 13685 5845 13715
rect 5845 13685 5875 13715
rect 5875 13685 5876 13715
rect 5844 13684 5876 13685
rect 5844 13635 5876 13636
rect 5844 13605 5845 13635
rect 5845 13605 5875 13635
rect 5875 13605 5876 13635
rect 5844 13604 5876 13605
rect 5844 13475 5876 13476
rect 5844 13445 5845 13475
rect 5845 13445 5875 13475
rect 5875 13445 5876 13475
rect 5844 13444 5876 13445
rect 5844 13395 5876 13396
rect 5844 13365 5845 13395
rect 5845 13365 5875 13395
rect 5875 13365 5876 13395
rect 5844 13364 5876 13365
rect 5844 13315 5876 13316
rect 5844 13285 5845 13315
rect 5845 13285 5875 13315
rect 5875 13285 5876 13315
rect 5844 13284 5876 13285
rect 5844 13235 5876 13236
rect 5844 13205 5845 13235
rect 5845 13205 5875 13235
rect 5875 13205 5876 13235
rect 5844 13204 5876 13205
rect 5844 13075 5876 13076
rect 5844 13045 5845 13075
rect 5845 13045 5875 13075
rect 5875 13045 5876 13075
rect 5844 13044 5876 13045
rect 5844 12995 5876 12996
rect 5844 12965 5845 12995
rect 5845 12965 5875 12995
rect 5875 12965 5876 12995
rect 5844 12964 5876 12965
rect 5844 12515 5876 12516
rect 5844 12485 5845 12515
rect 5845 12485 5875 12515
rect 5875 12485 5876 12515
rect 5844 12484 5876 12485
rect 5844 12435 5876 12436
rect 5844 12405 5845 12435
rect 5845 12405 5875 12435
rect 5875 12405 5876 12435
rect 5844 12404 5876 12405
rect 5844 12315 5876 12316
rect 5844 12285 5845 12315
rect 5845 12285 5875 12315
rect 5875 12285 5876 12315
rect 5844 12284 5876 12285
rect 5844 12235 5876 12236
rect 5844 12205 5845 12235
rect 5845 12205 5875 12235
rect 5875 12205 5876 12235
rect 5844 12204 5876 12205
rect 5844 12155 5876 12156
rect 5844 12125 5845 12155
rect 5845 12125 5875 12155
rect 5875 12125 5876 12155
rect 5844 12124 5876 12125
rect 5844 12075 5876 12076
rect 5844 12045 5845 12075
rect 5845 12045 5875 12075
rect 5875 12045 5876 12075
rect 5844 12044 5876 12045
rect 5844 11995 5876 11996
rect 5844 11965 5845 11995
rect 5845 11965 5875 11995
rect 5875 11965 5876 11995
rect 5844 11964 5876 11965
rect 5844 11915 5876 11916
rect 5844 11885 5845 11915
rect 5845 11885 5875 11915
rect 5875 11885 5876 11915
rect 5844 11884 5876 11885
rect 5844 11835 5876 11836
rect 5844 11805 5845 11835
rect 5845 11805 5875 11835
rect 5875 11805 5876 11835
rect 5844 11804 5876 11805
rect 5844 11755 5876 11756
rect 5844 11725 5845 11755
rect 5845 11725 5875 11755
rect 5875 11725 5876 11755
rect 5844 11724 5876 11725
rect 5844 11675 5876 11676
rect 5844 11645 5845 11675
rect 5845 11645 5875 11675
rect 5875 11645 5876 11675
rect 5844 11644 5876 11645
rect 5844 11595 5876 11596
rect 5844 11565 5845 11595
rect 5845 11565 5875 11595
rect 5875 11565 5876 11595
rect 5844 11564 5876 11565
rect 5844 11515 5876 11516
rect 5844 11485 5845 11515
rect 5845 11485 5875 11515
rect 5875 11485 5876 11515
rect 5844 11484 5876 11485
rect 5844 11435 5876 11436
rect 5844 11405 5845 11435
rect 5845 11405 5875 11435
rect 5875 11405 5876 11435
rect 5844 11404 5876 11405
rect 5844 11355 5876 11356
rect 5844 11325 5845 11355
rect 5845 11325 5875 11355
rect 5875 11325 5876 11355
rect 5844 11324 5876 11325
rect 5844 11195 5876 11196
rect 5844 11165 5845 11195
rect 5845 11165 5875 11195
rect 5875 11165 5876 11195
rect 5844 11164 5876 11165
rect 5844 11115 5876 11116
rect 5844 11085 5845 11115
rect 5845 11085 5875 11115
rect 5875 11085 5876 11115
rect 5844 11084 5876 11085
rect 5844 11035 5876 11036
rect 5844 11005 5845 11035
rect 5845 11005 5875 11035
rect 5875 11005 5876 11035
rect 5844 11004 5876 11005
rect 5844 10875 5876 10876
rect 5844 10845 5845 10875
rect 5845 10845 5875 10875
rect 5875 10845 5876 10875
rect 5844 10844 5876 10845
rect 5844 10715 5876 10716
rect 5844 10685 5845 10715
rect 5845 10685 5875 10715
rect 5875 10685 5876 10715
rect 5844 10684 5876 10685
rect 5844 10635 5876 10636
rect 5844 10605 5845 10635
rect 5845 10605 5875 10635
rect 5875 10605 5876 10635
rect 5844 10604 5876 10605
rect 5844 10475 5876 10476
rect 5844 10445 5845 10475
rect 5845 10445 5875 10475
rect 5875 10445 5876 10475
rect 5844 10444 5876 10445
rect 5844 10315 5876 10316
rect 5844 10285 5845 10315
rect 5845 10285 5875 10315
rect 5875 10285 5876 10315
rect 5844 10284 5876 10285
rect 5844 10235 5876 10236
rect 5844 10205 5845 10235
rect 5845 10205 5875 10235
rect 5875 10205 5876 10235
rect 5844 10204 5876 10205
rect 5844 10155 5876 10156
rect 5844 10125 5845 10155
rect 5845 10125 5875 10155
rect 5875 10125 5876 10155
rect 5844 10124 5876 10125
rect 5844 10075 5876 10076
rect 5844 10045 5845 10075
rect 5845 10045 5875 10075
rect 5875 10045 5876 10075
rect 5844 10044 5876 10045
rect 5844 9995 5876 9996
rect 5844 9965 5845 9995
rect 5845 9965 5875 9995
rect 5875 9965 5876 9995
rect 5844 9964 5876 9965
rect 5844 9915 5876 9916
rect 5844 9885 5845 9915
rect 5845 9885 5875 9915
rect 5875 9885 5876 9915
rect 5844 9884 5876 9885
rect 5844 9835 5876 9836
rect 5844 9805 5845 9835
rect 5845 9805 5875 9835
rect 5875 9805 5876 9835
rect 5844 9804 5876 9805
rect 5844 9755 5876 9756
rect 5844 9725 5845 9755
rect 5845 9725 5875 9755
rect 5875 9725 5876 9755
rect 5844 9724 5876 9725
rect 5844 9675 5876 9676
rect 5844 9645 5845 9675
rect 5845 9645 5875 9675
rect 5875 9645 5876 9675
rect 5844 9644 5876 9645
rect 5844 9595 5876 9596
rect 5844 9565 5845 9595
rect 5845 9565 5875 9595
rect 5875 9565 5876 9595
rect 5844 9564 5876 9565
rect 5844 9515 5876 9516
rect 5844 9485 5845 9515
rect 5845 9485 5875 9515
rect 5875 9485 5876 9515
rect 5844 9484 5876 9485
rect 5844 9435 5876 9436
rect 5844 9405 5845 9435
rect 5845 9405 5875 9435
rect 5875 9405 5876 9435
rect 5844 9404 5876 9405
rect 5844 9355 5876 9356
rect 5844 9325 5845 9355
rect 5845 9325 5875 9355
rect 5875 9325 5876 9355
rect 5844 9324 5876 9325
rect 5844 9275 5876 9276
rect 5844 9245 5845 9275
rect 5845 9245 5875 9275
rect 5875 9245 5876 9275
rect 5844 9244 5876 9245
rect 5844 9115 5876 9116
rect 5844 9085 5845 9115
rect 5845 9085 5875 9115
rect 5875 9085 5876 9115
rect 5844 9084 5876 9085
rect 5844 9035 5876 9036
rect 5844 9005 5845 9035
rect 5845 9005 5875 9035
rect 5875 9005 5876 9035
rect 5844 9004 5876 9005
rect 5844 8955 5876 8956
rect 5844 8925 5845 8955
rect 5845 8925 5875 8955
rect 5875 8925 5876 8955
rect 5844 8924 5876 8925
rect 5844 8635 5876 8636
rect 5844 8605 5845 8635
rect 5845 8605 5875 8635
rect 5875 8605 5876 8635
rect 5844 8604 5876 8605
rect 5844 8555 5876 8556
rect 5844 8525 5845 8555
rect 5845 8525 5875 8555
rect 5875 8525 5876 8555
rect 5844 8524 5876 8525
rect 5844 8395 5876 8396
rect 5844 8365 5845 8395
rect 5845 8365 5875 8395
rect 5875 8365 5876 8395
rect 5844 8364 5876 8365
rect 5844 8235 5876 8236
rect 5844 8205 5845 8235
rect 5845 8205 5875 8235
rect 5875 8205 5876 8235
rect 5844 8204 5876 8205
rect 5844 8155 5876 8156
rect 5844 8125 5845 8155
rect 5845 8125 5875 8155
rect 5875 8125 5876 8155
rect 5844 8124 5876 8125
rect 5844 8075 5876 8076
rect 5844 8045 5845 8075
rect 5845 8045 5875 8075
rect 5875 8045 5876 8075
rect 5844 8044 5876 8045
rect 5844 7995 5876 7996
rect 5844 7965 5845 7995
rect 5845 7965 5875 7995
rect 5875 7965 5876 7995
rect 5844 7964 5876 7965
rect 5844 7915 5876 7916
rect 5844 7885 5845 7915
rect 5845 7885 5875 7915
rect 5875 7885 5876 7915
rect 5844 7884 5876 7885
rect 5844 7835 5876 7836
rect 5844 7805 5845 7835
rect 5845 7805 5875 7835
rect 5875 7805 5876 7835
rect 5844 7804 5876 7805
rect 5844 7755 5876 7756
rect 5844 7725 5845 7755
rect 5845 7725 5875 7755
rect 5875 7725 5876 7755
rect 5844 7724 5876 7725
rect 5844 7675 5876 7676
rect 5844 7645 5845 7675
rect 5845 7645 5875 7675
rect 5875 7645 5876 7675
rect 5844 7644 5876 7645
rect 5844 7595 5876 7596
rect 5844 7565 5845 7595
rect 5845 7565 5875 7595
rect 5875 7565 5876 7595
rect 5844 7564 5876 7565
rect 5844 7515 5876 7516
rect 5844 7485 5845 7515
rect 5845 7485 5875 7515
rect 5875 7485 5876 7515
rect 5844 7484 5876 7485
rect 5844 7435 5876 7436
rect 5844 7405 5845 7435
rect 5845 7405 5875 7435
rect 5875 7405 5876 7435
rect 5844 7404 5876 7405
rect 5844 7355 5876 7356
rect 5844 7325 5845 7355
rect 5845 7325 5875 7355
rect 5875 7325 5876 7355
rect 5844 7324 5876 7325
rect 5844 7275 5876 7276
rect 5844 7245 5845 7275
rect 5845 7245 5875 7275
rect 5875 7245 5876 7275
rect 5844 7244 5876 7245
rect 5844 7195 5876 7196
rect 5844 7165 5845 7195
rect 5845 7165 5875 7195
rect 5875 7165 5876 7195
rect 5844 7164 5876 7165
rect 5844 7035 5876 7036
rect 5844 7005 5845 7035
rect 5845 7005 5875 7035
rect 5875 7005 5876 7035
rect 5844 7004 5876 7005
rect 5844 6955 5876 6956
rect 5844 6925 5845 6955
rect 5845 6925 5875 6955
rect 5875 6925 5876 6955
rect 5844 6924 5876 6925
rect 5844 6795 5876 6796
rect 5844 6765 5845 6795
rect 5845 6765 5875 6795
rect 5875 6765 5876 6795
rect 5844 6764 5876 6765
rect 5844 6715 5876 6716
rect 5844 6685 5845 6715
rect 5845 6685 5875 6715
rect 5875 6685 5876 6715
rect 5844 6684 5876 6685
rect 5844 6635 5876 6636
rect 5844 6605 5845 6635
rect 5845 6605 5875 6635
rect 5875 6605 5876 6635
rect 5844 6604 5876 6605
rect 5844 6555 5876 6556
rect 5844 6525 5845 6555
rect 5845 6525 5875 6555
rect 5875 6525 5876 6555
rect 5844 6524 5876 6525
rect 5844 6475 5876 6476
rect 5844 6445 5845 6475
rect 5845 6445 5875 6475
rect 5875 6445 5876 6475
rect 5844 6444 5876 6445
rect 5844 6315 5876 6316
rect 5844 6285 5845 6315
rect 5845 6285 5875 6315
rect 5875 6285 5876 6315
rect 5844 6284 5876 6285
rect 5844 6235 5876 6236
rect 5844 6205 5845 6235
rect 5845 6205 5875 6235
rect 5875 6205 5876 6235
rect 5844 6204 5876 6205
rect 5844 6155 5876 6156
rect 5844 6125 5845 6155
rect 5845 6125 5875 6155
rect 5875 6125 5876 6155
rect 5844 6124 5876 6125
rect 5844 5995 5876 5996
rect 5844 5965 5845 5995
rect 5845 5965 5875 5995
rect 5875 5965 5876 5995
rect 5844 5964 5876 5965
rect 5844 5835 5876 5836
rect 5844 5805 5845 5835
rect 5845 5805 5875 5835
rect 5875 5805 5876 5835
rect 5844 5804 5876 5805
rect 5844 5755 5876 5756
rect 5844 5725 5845 5755
rect 5845 5725 5875 5755
rect 5875 5725 5876 5755
rect 5844 5724 5876 5725
rect 5844 5675 5876 5676
rect 5844 5645 5845 5675
rect 5845 5645 5875 5675
rect 5875 5645 5876 5675
rect 5844 5644 5876 5645
rect 5844 5595 5876 5596
rect 5844 5565 5845 5595
rect 5845 5565 5875 5595
rect 5875 5565 5876 5595
rect 5844 5564 5876 5565
rect 5844 5515 5876 5516
rect 5844 5485 5845 5515
rect 5845 5485 5875 5515
rect 5875 5485 5876 5515
rect 5844 5484 5876 5485
rect 5844 5435 5876 5436
rect 5844 5405 5845 5435
rect 5845 5405 5875 5435
rect 5875 5405 5876 5435
rect 5844 5404 5876 5405
rect 5844 5355 5876 5356
rect 5844 5325 5845 5355
rect 5845 5325 5875 5355
rect 5875 5325 5876 5355
rect 5844 5324 5876 5325
rect 5844 5275 5876 5276
rect 5844 5245 5845 5275
rect 5845 5245 5875 5275
rect 5875 5245 5876 5275
rect 5844 5244 5876 5245
rect 5844 5195 5876 5196
rect 5844 5165 5845 5195
rect 5845 5165 5875 5195
rect 5875 5165 5876 5195
rect 5844 5164 5876 5165
rect 5844 5115 5876 5116
rect 5844 5085 5845 5115
rect 5845 5085 5875 5115
rect 5875 5085 5876 5115
rect 5844 5084 5876 5085
rect 5844 5035 5876 5036
rect 5844 5005 5845 5035
rect 5845 5005 5875 5035
rect 5875 5005 5876 5035
rect 5844 5004 5876 5005
rect 5844 4955 5876 4956
rect 5844 4925 5845 4955
rect 5845 4925 5875 4955
rect 5875 4925 5876 4955
rect 5844 4924 5876 4925
rect 5844 4875 5876 4876
rect 5844 4845 5845 4875
rect 5845 4845 5875 4875
rect 5875 4845 5876 4875
rect 5844 4844 5876 4845
rect 5844 4795 5876 4796
rect 5844 4765 5845 4795
rect 5845 4765 5875 4795
rect 5875 4765 5876 4795
rect 5844 4764 5876 4765
rect 5844 4635 5876 4636
rect 5844 4605 5845 4635
rect 5845 4605 5875 4635
rect 5875 4605 5876 4635
rect 5844 4604 5876 4605
rect 5844 4555 5876 4556
rect 5844 4525 5845 4555
rect 5845 4525 5875 4555
rect 5875 4525 5876 4555
rect 5844 4524 5876 4525
rect 5844 4395 5876 4396
rect 5844 4365 5845 4395
rect 5845 4365 5875 4395
rect 5875 4365 5876 4395
rect 5844 4364 5876 4365
rect 5844 4315 5876 4316
rect 5844 4285 5845 4315
rect 5845 4285 5875 4315
rect 5875 4285 5876 4315
rect 5844 4284 5876 4285
rect 5844 4235 5876 4236
rect 5844 4205 5845 4235
rect 5845 4205 5875 4235
rect 5875 4205 5876 4235
rect 5844 4204 5876 4205
rect 5844 4155 5876 4156
rect 5844 4125 5845 4155
rect 5845 4125 5875 4155
rect 5875 4125 5876 4155
rect 5844 4124 5876 4125
rect 5844 4075 5876 4076
rect 5844 4045 5845 4075
rect 5845 4045 5875 4075
rect 5875 4045 5876 4075
rect 5844 4044 5876 4045
rect 5844 3915 5876 3916
rect 5844 3885 5845 3915
rect 5845 3885 5875 3915
rect 5875 3885 5876 3915
rect 5844 3884 5876 3885
rect 5844 3835 5876 3836
rect 5844 3805 5845 3835
rect 5845 3805 5875 3835
rect 5875 3805 5876 3835
rect 5844 3804 5876 3805
rect 5844 3755 5876 3756
rect 5844 3725 5845 3755
rect 5845 3725 5875 3755
rect 5875 3725 5876 3755
rect 5844 3724 5876 3725
rect 5844 3595 5876 3596
rect 5844 3565 5845 3595
rect 5845 3565 5875 3595
rect 5875 3565 5876 3595
rect 5844 3564 5876 3565
rect 5844 3435 5876 3436
rect 5844 3405 5845 3435
rect 5845 3405 5875 3435
rect 5875 3405 5876 3435
rect 5844 3404 5876 3405
rect 5844 3355 5876 3356
rect 5844 3325 5845 3355
rect 5845 3325 5875 3355
rect 5875 3325 5876 3355
rect 5844 3324 5876 3325
rect 5844 3275 5876 3276
rect 5844 3245 5845 3275
rect 5845 3245 5875 3275
rect 5875 3245 5876 3275
rect 5844 3244 5876 3245
rect 5844 3195 5876 3196
rect 5844 3165 5845 3195
rect 5845 3165 5875 3195
rect 5875 3165 5876 3195
rect 5844 3164 5876 3165
rect 5844 3115 5876 3116
rect 5844 3085 5845 3115
rect 5845 3085 5875 3115
rect 5875 3085 5876 3115
rect 5844 3084 5876 3085
rect 5844 3035 5876 3036
rect 5844 3005 5845 3035
rect 5845 3005 5875 3035
rect 5875 3005 5876 3035
rect 5844 3004 5876 3005
rect 5844 2955 5876 2956
rect 5844 2925 5845 2955
rect 5845 2925 5875 2955
rect 5875 2925 5876 2955
rect 5844 2924 5876 2925
rect 5844 2875 5876 2876
rect 5844 2845 5845 2875
rect 5845 2845 5875 2875
rect 5875 2845 5876 2875
rect 5844 2844 5876 2845
rect 5844 2795 5876 2796
rect 5844 2765 5845 2795
rect 5845 2765 5875 2795
rect 5875 2765 5876 2795
rect 5844 2764 5876 2765
rect 5844 2715 5876 2716
rect 5844 2685 5845 2715
rect 5845 2685 5875 2715
rect 5875 2685 5876 2715
rect 5844 2684 5876 2685
rect 5844 2635 5876 2636
rect 5844 2605 5845 2635
rect 5845 2605 5875 2635
rect 5875 2605 5876 2635
rect 5844 2604 5876 2605
rect 5844 2555 5876 2556
rect 5844 2525 5845 2555
rect 5845 2525 5875 2555
rect 5875 2525 5876 2555
rect 5844 2524 5876 2525
rect 5844 2475 5876 2476
rect 5844 2445 5845 2475
rect 5845 2445 5875 2475
rect 5875 2445 5876 2475
rect 5844 2444 5876 2445
rect 5844 2395 5876 2396
rect 5844 2365 5845 2395
rect 5845 2365 5875 2395
rect 5875 2365 5876 2395
rect 5844 2364 5876 2365
rect 5844 2235 5876 2236
rect 5844 2205 5845 2235
rect 5845 2205 5875 2235
rect 5875 2205 5876 2235
rect 5844 2204 5876 2205
rect 5844 2155 5876 2156
rect 5844 2125 5845 2155
rect 5845 2125 5875 2155
rect 5875 2125 5876 2155
rect 5844 2124 5876 2125
rect 5844 2075 5876 2076
rect 5844 2045 5845 2075
rect 5845 2045 5875 2075
rect 5875 2045 5876 2075
rect 5844 2044 5876 2045
rect 5844 1995 5876 1996
rect 5844 1965 5845 1995
rect 5845 1965 5875 1995
rect 5875 1965 5876 1995
rect 5844 1964 5876 1965
rect 5844 1915 5876 1916
rect 5844 1885 5845 1915
rect 5845 1885 5875 1915
rect 5875 1885 5876 1915
rect 5844 1884 5876 1885
rect 5844 1835 5876 1836
rect 5844 1805 5845 1835
rect 5845 1805 5875 1835
rect 5875 1805 5876 1835
rect 5844 1804 5876 1805
rect 5844 1755 5876 1756
rect 5844 1725 5845 1755
rect 5845 1725 5875 1755
rect 5875 1725 5876 1755
rect 5844 1724 5876 1725
rect 5844 1675 5876 1676
rect 5844 1645 5845 1675
rect 5845 1645 5875 1675
rect 5875 1645 5876 1675
rect 5844 1644 5876 1645
rect 5844 1515 5876 1516
rect 5844 1485 5845 1515
rect 5845 1485 5875 1515
rect 5875 1485 5876 1515
rect 5844 1484 5876 1485
rect 5844 1435 5876 1436
rect 5844 1405 5845 1435
rect 5845 1405 5875 1435
rect 5875 1405 5876 1435
rect 5844 1404 5876 1405
rect 5844 1355 5876 1356
rect 5844 1325 5845 1355
rect 5845 1325 5875 1355
rect 5875 1325 5876 1355
rect 5844 1324 5876 1325
rect 5844 1275 5876 1276
rect 5844 1245 5845 1275
rect 5845 1245 5875 1275
rect 5875 1245 5876 1275
rect 5844 1244 5876 1245
rect 5844 1195 5876 1196
rect 5844 1165 5845 1195
rect 5845 1165 5875 1195
rect 5875 1165 5876 1195
rect 5844 1164 5876 1165
rect 5844 1115 5876 1116
rect 5844 1085 5845 1115
rect 5845 1085 5875 1115
rect 5875 1085 5876 1115
rect 5844 1084 5876 1085
rect 5844 1035 5876 1036
rect 5844 1005 5845 1035
rect 5845 1005 5875 1035
rect 5875 1005 5876 1035
rect 5844 1004 5876 1005
rect 5844 955 5876 956
rect 5844 925 5845 955
rect 5845 925 5875 955
rect 5875 925 5876 955
rect 5844 924 5876 925
rect 5844 875 5876 876
rect 5844 845 5845 875
rect 5845 845 5875 875
rect 5875 845 5876 875
rect 5844 844 5876 845
rect 5844 795 5876 796
rect 5844 765 5845 795
rect 5845 765 5875 795
rect 5875 765 5876 795
rect 5844 764 5876 765
rect 5844 715 5876 716
rect 5844 685 5845 715
rect 5845 685 5875 715
rect 5875 685 5876 715
rect 5844 684 5876 685
rect 5844 595 5876 596
rect 5844 565 5845 595
rect 5845 565 5875 595
rect 5875 565 5876 595
rect 5844 564 5876 565
rect 5844 515 5876 516
rect 5844 485 5845 515
rect 5845 485 5875 515
rect 5875 485 5876 515
rect 5844 484 5876 485
rect 5844 435 5876 436
rect 5844 405 5845 435
rect 5845 405 5875 435
rect 5875 405 5876 435
rect 5844 404 5876 405
rect 5844 355 5876 356
rect 5844 325 5845 355
rect 5845 325 5875 355
rect 5875 325 5876 355
rect 5844 324 5876 325
rect 5844 275 5876 276
rect 5844 245 5845 275
rect 5845 245 5875 275
rect 5875 245 5876 275
rect 5844 244 5876 245
rect 5844 195 5876 196
rect 5844 165 5845 195
rect 5845 165 5875 195
rect 5875 165 5876 195
rect 5844 164 5876 165
rect 5844 115 5876 116
rect 5844 85 5845 115
rect 5845 85 5875 115
rect 5875 85 5876 115
rect 5844 84 5876 85
rect 5844 35 5876 36
rect 5844 5 5845 35
rect 5845 5 5875 35
rect 5875 5 5876 35
rect 5844 4 5876 5
rect 6164 16644 6196 16836
rect 6004 16595 6036 16596
rect 6004 16565 6005 16595
rect 6005 16565 6035 16595
rect 6035 16565 6036 16595
rect 6004 16564 6036 16565
rect 6004 16515 6036 16516
rect 6004 16485 6005 16515
rect 6005 16485 6035 16515
rect 6035 16485 6036 16515
rect 6004 16484 6036 16485
rect 6004 16435 6036 16436
rect 6004 16405 6005 16435
rect 6005 16405 6035 16435
rect 6035 16405 6036 16435
rect 6004 16404 6036 16405
rect 6004 16355 6036 16356
rect 6004 16325 6005 16355
rect 6005 16325 6035 16355
rect 6035 16325 6036 16355
rect 6004 16324 6036 16325
rect 6004 16275 6036 16276
rect 6004 16245 6005 16275
rect 6005 16245 6035 16275
rect 6035 16245 6036 16275
rect 6004 16244 6036 16245
rect 6004 16195 6036 16196
rect 6004 16165 6005 16195
rect 6005 16165 6035 16195
rect 6035 16165 6036 16195
rect 6004 16164 6036 16165
rect 6004 16115 6036 16116
rect 6004 16085 6005 16115
rect 6005 16085 6035 16115
rect 6035 16085 6036 16115
rect 6004 16084 6036 16085
rect 6004 16035 6036 16036
rect 6004 16005 6005 16035
rect 6005 16005 6035 16035
rect 6035 16005 6036 16035
rect 6004 16004 6036 16005
rect 6004 15955 6036 15956
rect 6004 15925 6005 15955
rect 6005 15925 6035 15955
rect 6035 15925 6036 15955
rect 6004 15924 6036 15925
rect 6004 15435 6036 15436
rect 6004 15405 6005 15435
rect 6005 15405 6035 15435
rect 6035 15405 6036 15435
rect 6004 15404 6036 15405
rect 6004 15355 6036 15356
rect 6004 15325 6005 15355
rect 6005 15325 6035 15355
rect 6035 15325 6036 15355
rect 6004 15324 6036 15325
rect 6004 15275 6036 15276
rect 6004 15245 6005 15275
rect 6005 15245 6035 15275
rect 6035 15245 6036 15275
rect 6004 15244 6036 15245
rect 6004 15195 6036 15196
rect 6004 15165 6005 15195
rect 6005 15165 6035 15195
rect 6035 15165 6036 15195
rect 6004 15164 6036 15165
rect 6004 15115 6036 15116
rect 6004 15085 6005 15115
rect 6005 15085 6035 15115
rect 6035 15085 6036 15115
rect 6004 15084 6036 15085
rect 6004 14955 6036 14956
rect 6004 14925 6005 14955
rect 6005 14925 6035 14955
rect 6035 14925 6036 14955
rect 6004 14924 6036 14925
rect 6004 14875 6036 14876
rect 6004 14845 6005 14875
rect 6005 14845 6035 14875
rect 6035 14845 6036 14875
rect 6004 14844 6036 14845
rect 6004 14795 6036 14796
rect 6004 14765 6005 14795
rect 6005 14765 6035 14795
rect 6035 14765 6036 14795
rect 6004 14764 6036 14765
rect 6004 14715 6036 14716
rect 6004 14685 6005 14715
rect 6005 14685 6035 14715
rect 6035 14685 6036 14715
rect 6004 14684 6036 14685
rect 6004 14635 6036 14636
rect 6004 14605 6005 14635
rect 6005 14605 6035 14635
rect 6035 14605 6036 14635
rect 6004 14604 6036 14605
rect 6004 14555 6036 14556
rect 6004 14525 6005 14555
rect 6005 14525 6035 14555
rect 6035 14525 6036 14555
rect 6004 14524 6036 14525
rect 6004 14475 6036 14476
rect 6004 14445 6005 14475
rect 6005 14445 6035 14475
rect 6035 14445 6036 14475
rect 6004 14444 6036 14445
rect 6004 13995 6036 13996
rect 6004 13965 6005 13995
rect 6005 13965 6035 13995
rect 6035 13965 6036 13995
rect 6004 13964 6036 13965
rect 6004 13875 6036 13876
rect 6004 13845 6005 13875
rect 6005 13845 6035 13875
rect 6035 13845 6036 13875
rect 6004 13844 6036 13845
rect 6004 13795 6036 13796
rect 6004 13765 6005 13795
rect 6005 13765 6035 13795
rect 6035 13765 6036 13795
rect 6004 13764 6036 13765
rect 6004 13715 6036 13716
rect 6004 13685 6005 13715
rect 6005 13685 6035 13715
rect 6035 13685 6036 13715
rect 6004 13684 6036 13685
rect 6004 13635 6036 13636
rect 6004 13605 6005 13635
rect 6005 13605 6035 13635
rect 6035 13605 6036 13635
rect 6004 13604 6036 13605
rect 6004 13475 6036 13476
rect 6004 13445 6005 13475
rect 6005 13445 6035 13475
rect 6035 13445 6036 13475
rect 6004 13444 6036 13445
rect 6004 13395 6036 13396
rect 6004 13365 6005 13395
rect 6005 13365 6035 13395
rect 6035 13365 6036 13395
rect 6004 13364 6036 13365
rect 6004 13315 6036 13316
rect 6004 13285 6005 13315
rect 6005 13285 6035 13315
rect 6035 13285 6036 13315
rect 6004 13284 6036 13285
rect 6004 13235 6036 13236
rect 6004 13205 6005 13235
rect 6005 13205 6035 13235
rect 6035 13205 6036 13235
rect 6004 13204 6036 13205
rect 6004 13155 6036 13156
rect 6004 13125 6005 13155
rect 6005 13125 6035 13155
rect 6035 13125 6036 13155
rect 6004 13124 6036 13125
rect 6004 13075 6036 13076
rect 6004 13045 6005 13075
rect 6005 13045 6035 13075
rect 6035 13045 6036 13075
rect 6004 13044 6036 13045
rect 6004 12995 6036 12996
rect 6004 12965 6005 12995
rect 6005 12965 6035 12995
rect 6035 12965 6036 12995
rect 6004 12964 6036 12965
rect 6004 12515 6036 12516
rect 6004 12485 6005 12515
rect 6005 12485 6035 12515
rect 6035 12485 6036 12515
rect 6004 12484 6036 12485
rect 6004 12435 6036 12436
rect 6004 12405 6005 12435
rect 6005 12405 6035 12435
rect 6035 12405 6036 12435
rect 6004 12404 6036 12405
rect 6004 12315 6036 12316
rect 6004 12285 6005 12315
rect 6005 12285 6035 12315
rect 6035 12285 6036 12315
rect 6004 12284 6036 12285
rect 6004 12235 6036 12236
rect 6004 12205 6005 12235
rect 6005 12205 6035 12235
rect 6035 12205 6036 12235
rect 6004 12204 6036 12205
rect 6004 12155 6036 12156
rect 6004 12125 6005 12155
rect 6005 12125 6035 12155
rect 6035 12125 6036 12155
rect 6004 12124 6036 12125
rect 6004 12075 6036 12076
rect 6004 12045 6005 12075
rect 6005 12045 6035 12075
rect 6035 12045 6036 12075
rect 6004 12044 6036 12045
rect 6004 11995 6036 11996
rect 6004 11965 6005 11995
rect 6005 11965 6035 11995
rect 6035 11965 6036 11995
rect 6004 11964 6036 11965
rect 6004 11915 6036 11916
rect 6004 11885 6005 11915
rect 6005 11885 6035 11915
rect 6035 11885 6036 11915
rect 6004 11884 6036 11885
rect 6004 11835 6036 11836
rect 6004 11805 6005 11835
rect 6005 11805 6035 11835
rect 6035 11805 6036 11835
rect 6004 11804 6036 11805
rect 6004 11755 6036 11756
rect 6004 11725 6005 11755
rect 6005 11725 6035 11755
rect 6035 11725 6036 11755
rect 6004 11724 6036 11725
rect 6004 11675 6036 11676
rect 6004 11645 6005 11675
rect 6005 11645 6035 11675
rect 6035 11645 6036 11675
rect 6004 11644 6036 11645
rect 6004 11595 6036 11596
rect 6004 11565 6005 11595
rect 6005 11565 6035 11595
rect 6035 11565 6036 11595
rect 6004 11564 6036 11565
rect 6004 11515 6036 11516
rect 6004 11485 6005 11515
rect 6005 11485 6035 11515
rect 6035 11485 6036 11515
rect 6004 11484 6036 11485
rect 6004 11435 6036 11436
rect 6004 11405 6005 11435
rect 6005 11405 6035 11435
rect 6035 11405 6036 11435
rect 6004 11404 6036 11405
rect 6004 11355 6036 11356
rect 6004 11325 6005 11355
rect 6005 11325 6035 11355
rect 6035 11325 6036 11355
rect 6004 11324 6036 11325
rect 6004 11195 6036 11196
rect 6004 11165 6005 11195
rect 6005 11165 6035 11195
rect 6035 11165 6036 11195
rect 6004 11164 6036 11165
rect 6004 11115 6036 11116
rect 6004 11085 6005 11115
rect 6005 11085 6035 11115
rect 6035 11085 6036 11115
rect 6004 11084 6036 11085
rect 6004 11035 6036 11036
rect 6004 11005 6005 11035
rect 6005 11005 6035 11035
rect 6035 11005 6036 11035
rect 6004 11004 6036 11005
rect 6004 10875 6036 10876
rect 6004 10845 6005 10875
rect 6005 10845 6035 10875
rect 6035 10845 6036 10875
rect 6004 10844 6036 10845
rect 6004 10715 6036 10716
rect 6004 10685 6005 10715
rect 6005 10685 6035 10715
rect 6035 10685 6036 10715
rect 6004 10684 6036 10685
rect 6004 10635 6036 10636
rect 6004 10605 6005 10635
rect 6005 10605 6035 10635
rect 6035 10605 6036 10635
rect 6004 10604 6036 10605
rect 6004 10475 6036 10476
rect 6004 10445 6005 10475
rect 6005 10445 6035 10475
rect 6035 10445 6036 10475
rect 6004 10444 6036 10445
rect 6004 10315 6036 10316
rect 6004 10285 6005 10315
rect 6005 10285 6035 10315
rect 6035 10285 6036 10315
rect 6004 10284 6036 10285
rect 6004 10235 6036 10236
rect 6004 10205 6005 10235
rect 6005 10205 6035 10235
rect 6035 10205 6036 10235
rect 6004 10204 6036 10205
rect 6004 10155 6036 10156
rect 6004 10125 6005 10155
rect 6005 10125 6035 10155
rect 6035 10125 6036 10155
rect 6004 10124 6036 10125
rect 6004 10075 6036 10076
rect 6004 10045 6005 10075
rect 6005 10045 6035 10075
rect 6035 10045 6036 10075
rect 6004 10044 6036 10045
rect 6004 9995 6036 9996
rect 6004 9965 6005 9995
rect 6005 9965 6035 9995
rect 6035 9965 6036 9995
rect 6004 9964 6036 9965
rect 6004 9915 6036 9916
rect 6004 9885 6005 9915
rect 6005 9885 6035 9915
rect 6035 9885 6036 9915
rect 6004 9884 6036 9885
rect 6004 9835 6036 9836
rect 6004 9805 6005 9835
rect 6005 9805 6035 9835
rect 6035 9805 6036 9835
rect 6004 9804 6036 9805
rect 6004 9755 6036 9756
rect 6004 9725 6005 9755
rect 6005 9725 6035 9755
rect 6035 9725 6036 9755
rect 6004 9724 6036 9725
rect 6004 9675 6036 9676
rect 6004 9645 6005 9675
rect 6005 9645 6035 9675
rect 6035 9645 6036 9675
rect 6004 9644 6036 9645
rect 6004 9595 6036 9596
rect 6004 9565 6005 9595
rect 6005 9565 6035 9595
rect 6035 9565 6036 9595
rect 6004 9564 6036 9565
rect 6004 9515 6036 9516
rect 6004 9485 6005 9515
rect 6005 9485 6035 9515
rect 6035 9485 6036 9515
rect 6004 9484 6036 9485
rect 6004 9435 6036 9436
rect 6004 9405 6005 9435
rect 6005 9405 6035 9435
rect 6035 9405 6036 9435
rect 6004 9404 6036 9405
rect 6004 9355 6036 9356
rect 6004 9325 6005 9355
rect 6005 9325 6035 9355
rect 6035 9325 6036 9355
rect 6004 9324 6036 9325
rect 6004 9275 6036 9276
rect 6004 9245 6005 9275
rect 6005 9245 6035 9275
rect 6035 9245 6036 9275
rect 6004 9244 6036 9245
rect 6004 9115 6036 9116
rect 6004 9085 6005 9115
rect 6005 9085 6035 9115
rect 6035 9085 6036 9115
rect 6004 9084 6036 9085
rect 6004 9035 6036 9036
rect 6004 9005 6005 9035
rect 6005 9005 6035 9035
rect 6035 9005 6036 9035
rect 6004 9004 6036 9005
rect 6004 8955 6036 8956
rect 6004 8925 6005 8955
rect 6005 8925 6035 8955
rect 6035 8925 6036 8955
rect 6004 8924 6036 8925
rect 6004 8635 6036 8636
rect 6004 8605 6005 8635
rect 6005 8605 6035 8635
rect 6035 8605 6036 8635
rect 6004 8604 6036 8605
rect 6004 8555 6036 8556
rect 6004 8525 6005 8555
rect 6005 8525 6035 8555
rect 6035 8525 6036 8555
rect 6004 8524 6036 8525
rect 6004 8395 6036 8396
rect 6004 8365 6005 8395
rect 6005 8365 6035 8395
rect 6035 8365 6036 8395
rect 6004 8364 6036 8365
rect 6004 8235 6036 8236
rect 6004 8205 6005 8235
rect 6005 8205 6035 8235
rect 6035 8205 6036 8235
rect 6004 8204 6036 8205
rect 6004 8155 6036 8156
rect 6004 8125 6005 8155
rect 6005 8125 6035 8155
rect 6035 8125 6036 8155
rect 6004 8124 6036 8125
rect 6004 8075 6036 8076
rect 6004 8045 6005 8075
rect 6005 8045 6035 8075
rect 6035 8045 6036 8075
rect 6004 8044 6036 8045
rect 6004 7995 6036 7996
rect 6004 7965 6005 7995
rect 6005 7965 6035 7995
rect 6035 7965 6036 7995
rect 6004 7964 6036 7965
rect 6004 7915 6036 7916
rect 6004 7885 6005 7915
rect 6005 7885 6035 7915
rect 6035 7885 6036 7915
rect 6004 7884 6036 7885
rect 6004 7835 6036 7836
rect 6004 7805 6005 7835
rect 6005 7805 6035 7835
rect 6035 7805 6036 7835
rect 6004 7804 6036 7805
rect 6004 7755 6036 7756
rect 6004 7725 6005 7755
rect 6005 7725 6035 7755
rect 6035 7725 6036 7755
rect 6004 7724 6036 7725
rect 6004 7675 6036 7676
rect 6004 7645 6005 7675
rect 6005 7645 6035 7675
rect 6035 7645 6036 7675
rect 6004 7644 6036 7645
rect 6004 7595 6036 7596
rect 6004 7565 6005 7595
rect 6005 7565 6035 7595
rect 6035 7565 6036 7595
rect 6004 7564 6036 7565
rect 6004 7515 6036 7516
rect 6004 7485 6005 7515
rect 6005 7485 6035 7515
rect 6035 7485 6036 7515
rect 6004 7484 6036 7485
rect 6004 7435 6036 7436
rect 6004 7405 6005 7435
rect 6005 7405 6035 7435
rect 6035 7405 6036 7435
rect 6004 7404 6036 7405
rect 6004 7355 6036 7356
rect 6004 7325 6005 7355
rect 6005 7325 6035 7355
rect 6035 7325 6036 7355
rect 6004 7324 6036 7325
rect 6004 7275 6036 7276
rect 6004 7245 6005 7275
rect 6005 7245 6035 7275
rect 6035 7245 6036 7275
rect 6004 7244 6036 7245
rect 6004 7195 6036 7196
rect 6004 7165 6005 7195
rect 6005 7165 6035 7195
rect 6035 7165 6036 7195
rect 6004 7164 6036 7165
rect 6004 7035 6036 7036
rect 6004 7005 6005 7035
rect 6005 7005 6035 7035
rect 6035 7005 6036 7035
rect 6004 7004 6036 7005
rect 6004 6955 6036 6956
rect 6004 6925 6005 6955
rect 6005 6925 6035 6955
rect 6035 6925 6036 6955
rect 6004 6924 6036 6925
rect 6004 6795 6036 6796
rect 6004 6765 6005 6795
rect 6005 6765 6035 6795
rect 6035 6765 6036 6795
rect 6004 6764 6036 6765
rect 6004 6715 6036 6716
rect 6004 6685 6005 6715
rect 6005 6685 6035 6715
rect 6035 6685 6036 6715
rect 6004 6684 6036 6685
rect 6004 6635 6036 6636
rect 6004 6605 6005 6635
rect 6005 6605 6035 6635
rect 6035 6605 6036 6635
rect 6004 6604 6036 6605
rect 6004 6555 6036 6556
rect 6004 6525 6005 6555
rect 6005 6525 6035 6555
rect 6035 6525 6036 6555
rect 6004 6524 6036 6525
rect 6004 6475 6036 6476
rect 6004 6445 6005 6475
rect 6005 6445 6035 6475
rect 6035 6445 6036 6475
rect 6004 6444 6036 6445
rect 6004 6315 6036 6316
rect 6004 6285 6005 6315
rect 6005 6285 6035 6315
rect 6035 6285 6036 6315
rect 6004 6284 6036 6285
rect 6004 6235 6036 6236
rect 6004 6205 6005 6235
rect 6005 6205 6035 6235
rect 6035 6205 6036 6235
rect 6004 6204 6036 6205
rect 6004 6155 6036 6156
rect 6004 6125 6005 6155
rect 6005 6125 6035 6155
rect 6035 6125 6036 6155
rect 6004 6124 6036 6125
rect 6004 5995 6036 5996
rect 6004 5965 6005 5995
rect 6005 5965 6035 5995
rect 6035 5965 6036 5995
rect 6004 5964 6036 5965
rect 6004 5835 6036 5836
rect 6004 5805 6005 5835
rect 6005 5805 6035 5835
rect 6035 5805 6036 5835
rect 6004 5804 6036 5805
rect 6004 5755 6036 5756
rect 6004 5725 6005 5755
rect 6005 5725 6035 5755
rect 6035 5725 6036 5755
rect 6004 5724 6036 5725
rect 6004 5675 6036 5676
rect 6004 5645 6005 5675
rect 6005 5645 6035 5675
rect 6035 5645 6036 5675
rect 6004 5644 6036 5645
rect 6004 5595 6036 5596
rect 6004 5565 6005 5595
rect 6005 5565 6035 5595
rect 6035 5565 6036 5595
rect 6004 5564 6036 5565
rect 6004 5515 6036 5516
rect 6004 5485 6005 5515
rect 6005 5485 6035 5515
rect 6035 5485 6036 5515
rect 6004 5484 6036 5485
rect 6004 5435 6036 5436
rect 6004 5405 6005 5435
rect 6005 5405 6035 5435
rect 6035 5405 6036 5435
rect 6004 5404 6036 5405
rect 6004 5355 6036 5356
rect 6004 5325 6005 5355
rect 6005 5325 6035 5355
rect 6035 5325 6036 5355
rect 6004 5324 6036 5325
rect 6004 5275 6036 5276
rect 6004 5245 6005 5275
rect 6005 5245 6035 5275
rect 6035 5245 6036 5275
rect 6004 5244 6036 5245
rect 6004 5195 6036 5196
rect 6004 5165 6005 5195
rect 6005 5165 6035 5195
rect 6035 5165 6036 5195
rect 6004 5164 6036 5165
rect 6004 5115 6036 5116
rect 6004 5085 6005 5115
rect 6005 5085 6035 5115
rect 6035 5085 6036 5115
rect 6004 5084 6036 5085
rect 6004 5035 6036 5036
rect 6004 5005 6005 5035
rect 6005 5005 6035 5035
rect 6035 5005 6036 5035
rect 6004 5004 6036 5005
rect 6004 4955 6036 4956
rect 6004 4925 6005 4955
rect 6005 4925 6035 4955
rect 6035 4925 6036 4955
rect 6004 4924 6036 4925
rect 6004 4875 6036 4876
rect 6004 4845 6005 4875
rect 6005 4845 6035 4875
rect 6035 4845 6036 4875
rect 6004 4844 6036 4845
rect 6004 4795 6036 4796
rect 6004 4765 6005 4795
rect 6005 4765 6035 4795
rect 6035 4765 6036 4795
rect 6004 4764 6036 4765
rect 6004 4635 6036 4636
rect 6004 4605 6005 4635
rect 6005 4605 6035 4635
rect 6035 4605 6036 4635
rect 6004 4604 6036 4605
rect 6004 4555 6036 4556
rect 6004 4525 6005 4555
rect 6005 4525 6035 4555
rect 6035 4525 6036 4555
rect 6004 4524 6036 4525
rect 6004 4395 6036 4396
rect 6004 4365 6005 4395
rect 6005 4365 6035 4395
rect 6035 4365 6036 4395
rect 6004 4364 6036 4365
rect 6004 4315 6036 4316
rect 6004 4285 6005 4315
rect 6005 4285 6035 4315
rect 6035 4285 6036 4315
rect 6004 4284 6036 4285
rect 6004 4235 6036 4236
rect 6004 4205 6005 4235
rect 6005 4205 6035 4235
rect 6035 4205 6036 4235
rect 6004 4204 6036 4205
rect 6004 4155 6036 4156
rect 6004 4125 6005 4155
rect 6005 4125 6035 4155
rect 6035 4125 6036 4155
rect 6004 4124 6036 4125
rect 6004 4075 6036 4076
rect 6004 4045 6005 4075
rect 6005 4045 6035 4075
rect 6035 4045 6036 4075
rect 6004 4044 6036 4045
rect 6004 3915 6036 3916
rect 6004 3885 6005 3915
rect 6005 3885 6035 3915
rect 6035 3885 6036 3915
rect 6004 3884 6036 3885
rect 6004 3835 6036 3836
rect 6004 3805 6005 3835
rect 6005 3805 6035 3835
rect 6035 3805 6036 3835
rect 6004 3804 6036 3805
rect 6004 3755 6036 3756
rect 6004 3725 6005 3755
rect 6005 3725 6035 3755
rect 6035 3725 6036 3755
rect 6004 3724 6036 3725
rect 6004 3595 6036 3596
rect 6004 3565 6005 3595
rect 6005 3565 6035 3595
rect 6035 3565 6036 3595
rect 6004 3564 6036 3565
rect 6004 3435 6036 3436
rect 6004 3405 6005 3435
rect 6005 3405 6035 3435
rect 6035 3405 6036 3435
rect 6004 3404 6036 3405
rect 6004 3355 6036 3356
rect 6004 3325 6005 3355
rect 6005 3325 6035 3355
rect 6035 3325 6036 3355
rect 6004 3324 6036 3325
rect 6004 3275 6036 3276
rect 6004 3245 6005 3275
rect 6005 3245 6035 3275
rect 6035 3245 6036 3275
rect 6004 3244 6036 3245
rect 6004 3195 6036 3196
rect 6004 3165 6005 3195
rect 6005 3165 6035 3195
rect 6035 3165 6036 3195
rect 6004 3164 6036 3165
rect 6004 3115 6036 3116
rect 6004 3085 6005 3115
rect 6005 3085 6035 3115
rect 6035 3085 6036 3115
rect 6004 3084 6036 3085
rect 6004 3035 6036 3036
rect 6004 3005 6005 3035
rect 6005 3005 6035 3035
rect 6035 3005 6036 3035
rect 6004 3004 6036 3005
rect 6004 2955 6036 2956
rect 6004 2925 6005 2955
rect 6005 2925 6035 2955
rect 6035 2925 6036 2955
rect 6004 2924 6036 2925
rect 6004 2875 6036 2876
rect 6004 2845 6005 2875
rect 6005 2845 6035 2875
rect 6035 2845 6036 2875
rect 6004 2844 6036 2845
rect 6004 2795 6036 2796
rect 6004 2765 6005 2795
rect 6005 2765 6035 2795
rect 6035 2765 6036 2795
rect 6004 2764 6036 2765
rect 6004 2715 6036 2716
rect 6004 2685 6005 2715
rect 6005 2685 6035 2715
rect 6035 2685 6036 2715
rect 6004 2684 6036 2685
rect 6004 2635 6036 2636
rect 6004 2605 6005 2635
rect 6005 2605 6035 2635
rect 6035 2605 6036 2635
rect 6004 2604 6036 2605
rect 6004 2555 6036 2556
rect 6004 2525 6005 2555
rect 6005 2525 6035 2555
rect 6035 2525 6036 2555
rect 6004 2524 6036 2525
rect 6004 2475 6036 2476
rect 6004 2445 6005 2475
rect 6005 2445 6035 2475
rect 6035 2445 6036 2475
rect 6004 2444 6036 2445
rect 6004 2395 6036 2396
rect 6004 2365 6005 2395
rect 6005 2365 6035 2395
rect 6035 2365 6036 2395
rect 6004 2364 6036 2365
rect 6004 2235 6036 2236
rect 6004 2205 6005 2235
rect 6005 2205 6035 2235
rect 6035 2205 6036 2235
rect 6004 2204 6036 2205
rect 6004 2155 6036 2156
rect 6004 2125 6005 2155
rect 6005 2125 6035 2155
rect 6035 2125 6036 2155
rect 6004 2124 6036 2125
rect 6004 2075 6036 2076
rect 6004 2045 6005 2075
rect 6005 2045 6035 2075
rect 6035 2045 6036 2075
rect 6004 2044 6036 2045
rect 6004 1995 6036 1996
rect 6004 1965 6005 1995
rect 6005 1965 6035 1995
rect 6035 1965 6036 1995
rect 6004 1964 6036 1965
rect 6004 1915 6036 1916
rect 6004 1885 6005 1915
rect 6005 1885 6035 1915
rect 6035 1885 6036 1915
rect 6004 1884 6036 1885
rect 6004 1835 6036 1836
rect 6004 1805 6005 1835
rect 6005 1805 6035 1835
rect 6035 1805 6036 1835
rect 6004 1804 6036 1805
rect 6004 1755 6036 1756
rect 6004 1725 6005 1755
rect 6005 1725 6035 1755
rect 6035 1725 6036 1755
rect 6004 1724 6036 1725
rect 6004 1675 6036 1676
rect 6004 1645 6005 1675
rect 6005 1645 6035 1675
rect 6035 1645 6036 1675
rect 6004 1644 6036 1645
rect 6004 1595 6036 1596
rect 6004 1565 6005 1595
rect 6005 1565 6035 1595
rect 6035 1565 6036 1595
rect 6004 1564 6036 1565
rect 6004 1515 6036 1516
rect 6004 1485 6005 1515
rect 6005 1485 6035 1515
rect 6035 1485 6036 1515
rect 6004 1484 6036 1485
rect 6004 1435 6036 1436
rect 6004 1405 6005 1435
rect 6005 1405 6035 1435
rect 6035 1405 6036 1435
rect 6004 1404 6036 1405
rect 6004 1355 6036 1356
rect 6004 1325 6005 1355
rect 6005 1325 6035 1355
rect 6035 1325 6036 1355
rect 6004 1324 6036 1325
rect 6004 1275 6036 1276
rect 6004 1245 6005 1275
rect 6005 1245 6035 1275
rect 6035 1245 6036 1275
rect 6004 1244 6036 1245
rect 6004 1195 6036 1196
rect 6004 1165 6005 1195
rect 6005 1165 6035 1195
rect 6035 1165 6036 1195
rect 6004 1164 6036 1165
rect 6004 1115 6036 1116
rect 6004 1085 6005 1115
rect 6005 1085 6035 1115
rect 6035 1085 6036 1115
rect 6004 1084 6036 1085
rect 6004 1035 6036 1036
rect 6004 1005 6005 1035
rect 6005 1005 6035 1035
rect 6035 1005 6036 1035
rect 6004 1004 6036 1005
rect 6004 955 6036 956
rect 6004 925 6005 955
rect 6005 925 6035 955
rect 6035 925 6036 955
rect 6004 924 6036 925
rect 6004 875 6036 876
rect 6004 845 6005 875
rect 6005 845 6035 875
rect 6035 845 6036 875
rect 6004 844 6036 845
rect 6004 795 6036 796
rect 6004 765 6005 795
rect 6005 765 6035 795
rect 6035 765 6036 795
rect 6004 764 6036 765
rect 6004 715 6036 716
rect 6004 685 6005 715
rect 6005 685 6035 715
rect 6035 685 6036 715
rect 6004 684 6036 685
rect 6004 595 6036 596
rect 6004 565 6005 595
rect 6005 565 6035 595
rect 6035 565 6036 595
rect 6004 564 6036 565
rect 6004 515 6036 516
rect 6004 485 6005 515
rect 6005 485 6035 515
rect 6035 485 6036 515
rect 6004 484 6036 485
rect 6004 435 6036 436
rect 6004 405 6005 435
rect 6005 405 6035 435
rect 6035 405 6036 435
rect 6004 404 6036 405
rect 6004 355 6036 356
rect 6004 325 6005 355
rect 6005 325 6035 355
rect 6035 325 6036 355
rect 6004 324 6036 325
rect 6004 275 6036 276
rect 6004 245 6005 275
rect 6005 245 6035 275
rect 6035 245 6036 275
rect 6004 244 6036 245
rect 6004 195 6036 196
rect 6004 165 6005 195
rect 6005 165 6035 195
rect 6035 165 6036 195
rect 6004 164 6036 165
rect 6004 115 6036 116
rect 6004 85 6005 115
rect 6005 85 6035 115
rect 6035 85 6036 115
rect 6004 84 6036 85
rect 6004 35 6036 36
rect 6004 5 6005 35
rect 6005 5 6035 35
rect 6035 5 6036 35
rect 6004 4 6036 5
rect 6324 16644 6356 16836
rect 6164 16595 6196 16596
rect 6164 16565 6165 16595
rect 6165 16565 6195 16595
rect 6195 16565 6196 16595
rect 6164 16564 6196 16565
rect 6164 16515 6196 16516
rect 6164 16485 6165 16515
rect 6165 16485 6195 16515
rect 6195 16485 6196 16515
rect 6164 16484 6196 16485
rect 6164 16435 6196 16436
rect 6164 16405 6165 16435
rect 6165 16405 6195 16435
rect 6195 16405 6196 16435
rect 6164 16404 6196 16405
rect 6164 16355 6196 16356
rect 6164 16325 6165 16355
rect 6165 16325 6195 16355
rect 6195 16325 6196 16355
rect 6164 16324 6196 16325
rect 6164 16275 6196 16276
rect 6164 16245 6165 16275
rect 6165 16245 6195 16275
rect 6195 16245 6196 16275
rect 6164 16244 6196 16245
rect 6164 16195 6196 16196
rect 6164 16165 6165 16195
rect 6165 16165 6195 16195
rect 6195 16165 6196 16195
rect 6164 16164 6196 16165
rect 6164 16115 6196 16116
rect 6164 16085 6165 16115
rect 6165 16085 6195 16115
rect 6195 16085 6196 16115
rect 6164 16084 6196 16085
rect 6164 16035 6196 16036
rect 6164 16005 6165 16035
rect 6165 16005 6195 16035
rect 6195 16005 6196 16035
rect 6164 16004 6196 16005
rect 6164 15955 6196 15956
rect 6164 15925 6165 15955
rect 6165 15925 6195 15955
rect 6195 15925 6196 15955
rect 6164 15924 6196 15925
rect 6164 15435 6196 15436
rect 6164 15405 6165 15435
rect 6165 15405 6195 15435
rect 6195 15405 6196 15435
rect 6164 15404 6196 15405
rect 6164 15355 6196 15356
rect 6164 15325 6165 15355
rect 6165 15325 6195 15355
rect 6195 15325 6196 15355
rect 6164 15324 6196 15325
rect 6164 15275 6196 15276
rect 6164 15245 6165 15275
rect 6165 15245 6195 15275
rect 6195 15245 6196 15275
rect 6164 15244 6196 15245
rect 6164 15195 6196 15196
rect 6164 15165 6165 15195
rect 6165 15165 6195 15195
rect 6195 15165 6196 15195
rect 6164 15164 6196 15165
rect 6164 15115 6196 15116
rect 6164 15085 6165 15115
rect 6165 15085 6195 15115
rect 6195 15085 6196 15115
rect 6164 15084 6196 15085
rect 6164 15035 6196 15036
rect 6164 15005 6165 15035
rect 6165 15005 6195 15035
rect 6195 15005 6196 15035
rect 6164 15004 6196 15005
rect 6164 14955 6196 14956
rect 6164 14925 6165 14955
rect 6165 14925 6195 14955
rect 6195 14925 6196 14955
rect 6164 14924 6196 14925
rect 6164 14875 6196 14876
rect 6164 14845 6165 14875
rect 6165 14845 6195 14875
rect 6195 14845 6196 14875
rect 6164 14844 6196 14845
rect 6164 14795 6196 14796
rect 6164 14765 6165 14795
rect 6165 14765 6195 14795
rect 6195 14765 6196 14795
rect 6164 14764 6196 14765
rect 6164 14715 6196 14716
rect 6164 14685 6165 14715
rect 6165 14685 6195 14715
rect 6195 14685 6196 14715
rect 6164 14684 6196 14685
rect 6164 14635 6196 14636
rect 6164 14605 6165 14635
rect 6165 14605 6195 14635
rect 6195 14605 6196 14635
rect 6164 14604 6196 14605
rect 6164 14555 6196 14556
rect 6164 14525 6165 14555
rect 6165 14525 6195 14555
rect 6195 14525 6196 14555
rect 6164 14524 6196 14525
rect 6164 14475 6196 14476
rect 6164 14445 6165 14475
rect 6165 14445 6195 14475
rect 6195 14445 6196 14475
rect 6164 14444 6196 14445
rect 6164 13995 6196 13996
rect 6164 13965 6165 13995
rect 6165 13965 6195 13995
rect 6195 13965 6196 13995
rect 6164 13964 6196 13965
rect 6164 13875 6196 13876
rect 6164 13845 6165 13875
rect 6165 13845 6195 13875
rect 6195 13845 6196 13875
rect 6164 13844 6196 13845
rect 6164 13795 6196 13796
rect 6164 13765 6165 13795
rect 6165 13765 6195 13795
rect 6195 13765 6196 13795
rect 6164 13764 6196 13765
rect 6164 13715 6196 13716
rect 6164 13685 6165 13715
rect 6165 13685 6195 13715
rect 6195 13685 6196 13715
rect 6164 13684 6196 13685
rect 6164 13635 6196 13636
rect 6164 13605 6165 13635
rect 6165 13605 6195 13635
rect 6195 13605 6196 13635
rect 6164 13604 6196 13605
rect 6164 13555 6196 13556
rect 6164 13525 6165 13555
rect 6165 13525 6195 13555
rect 6195 13525 6196 13555
rect 6164 13524 6196 13525
rect 6164 13475 6196 13476
rect 6164 13445 6165 13475
rect 6165 13445 6195 13475
rect 6195 13445 6196 13475
rect 6164 13444 6196 13445
rect 6164 13395 6196 13396
rect 6164 13365 6165 13395
rect 6165 13365 6195 13395
rect 6195 13365 6196 13395
rect 6164 13364 6196 13365
rect 6164 13315 6196 13316
rect 6164 13285 6165 13315
rect 6165 13285 6195 13315
rect 6195 13285 6196 13315
rect 6164 13284 6196 13285
rect 6164 13235 6196 13236
rect 6164 13205 6165 13235
rect 6165 13205 6195 13235
rect 6195 13205 6196 13235
rect 6164 13204 6196 13205
rect 6164 13155 6196 13156
rect 6164 13125 6165 13155
rect 6165 13125 6195 13155
rect 6195 13125 6196 13155
rect 6164 13124 6196 13125
rect 6164 13075 6196 13076
rect 6164 13045 6165 13075
rect 6165 13045 6195 13075
rect 6195 13045 6196 13075
rect 6164 13044 6196 13045
rect 6164 12995 6196 12996
rect 6164 12965 6165 12995
rect 6165 12965 6195 12995
rect 6195 12965 6196 12995
rect 6164 12964 6196 12965
rect 6164 12515 6196 12516
rect 6164 12485 6165 12515
rect 6165 12485 6195 12515
rect 6195 12485 6196 12515
rect 6164 12484 6196 12485
rect 6164 12435 6196 12436
rect 6164 12405 6165 12435
rect 6165 12405 6195 12435
rect 6195 12405 6196 12435
rect 6164 12404 6196 12405
rect 6164 12315 6196 12316
rect 6164 12285 6165 12315
rect 6165 12285 6195 12315
rect 6195 12285 6196 12315
rect 6164 12284 6196 12285
rect 6164 12235 6196 12236
rect 6164 12205 6165 12235
rect 6165 12205 6195 12235
rect 6195 12205 6196 12235
rect 6164 12204 6196 12205
rect 6164 12155 6196 12156
rect 6164 12125 6165 12155
rect 6165 12125 6195 12155
rect 6195 12125 6196 12155
rect 6164 12124 6196 12125
rect 6164 12075 6196 12076
rect 6164 12045 6165 12075
rect 6165 12045 6195 12075
rect 6195 12045 6196 12075
rect 6164 12044 6196 12045
rect 6164 11995 6196 11996
rect 6164 11965 6165 11995
rect 6165 11965 6195 11995
rect 6195 11965 6196 11995
rect 6164 11964 6196 11965
rect 6164 11915 6196 11916
rect 6164 11885 6165 11915
rect 6165 11885 6195 11915
rect 6195 11885 6196 11915
rect 6164 11884 6196 11885
rect 6164 11835 6196 11836
rect 6164 11805 6165 11835
rect 6165 11805 6195 11835
rect 6195 11805 6196 11835
rect 6164 11804 6196 11805
rect 6164 11755 6196 11756
rect 6164 11725 6165 11755
rect 6165 11725 6195 11755
rect 6195 11725 6196 11755
rect 6164 11724 6196 11725
rect 6164 11675 6196 11676
rect 6164 11645 6165 11675
rect 6165 11645 6195 11675
rect 6195 11645 6196 11675
rect 6164 11644 6196 11645
rect 6164 11595 6196 11596
rect 6164 11565 6165 11595
rect 6165 11565 6195 11595
rect 6195 11565 6196 11595
rect 6164 11564 6196 11565
rect 6164 11515 6196 11516
rect 6164 11485 6165 11515
rect 6165 11485 6195 11515
rect 6195 11485 6196 11515
rect 6164 11484 6196 11485
rect 6164 11435 6196 11436
rect 6164 11405 6165 11435
rect 6165 11405 6195 11435
rect 6195 11405 6196 11435
rect 6164 11404 6196 11405
rect 6164 11355 6196 11356
rect 6164 11325 6165 11355
rect 6165 11325 6195 11355
rect 6195 11325 6196 11355
rect 6164 11324 6196 11325
rect 6164 11195 6196 11196
rect 6164 11165 6165 11195
rect 6165 11165 6195 11195
rect 6195 11165 6196 11195
rect 6164 11164 6196 11165
rect 6164 11115 6196 11116
rect 6164 11085 6165 11115
rect 6165 11085 6195 11115
rect 6195 11085 6196 11115
rect 6164 11084 6196 11085
rect 6164 11035 6196 11036
rect 6164 11005 6165 11035
rect 6165 11005 6195 11035
rect 6195 11005 6196 11035
rect 6164 11004 6196 11005
rect 6164 10875 6196 10876
rect 6164 10845 6165 10875
rect 6165 10845 6195 10875
rect 6195 10845 6196 10875
rect 6164 10844 6196 10845
rect 6164 10715 6196 10716
rect 6164 10685 6165 10715
rect 6165 10685 6195 10715
rect 6195 10685 6196 10715
rect 6164 10684 6196 10685
rect 6164 10635 6196 10636
rect 6164 10605 6165 10635
rect 6165 10605 6195 10635
rect 6195 10605 6196 10635
rect 6164 10604 6196 10605
rect 6164 10475 6196 10476
rect 6164 10445 6165 10475
rect 6165 10445 6195 10475
rect 6195 10445 6196 10475
rect 6164 10444 6196 10445
rect 6164 10315 6196 10316
rect 6164 10285 6165 10315
rect 6165 10285 6195 10315
rect 6195 10285 6196 10315
rect 6164 10284 6196 10285
rect 6164 10235 6196 10236
rect 6164 10205 6165 10235
rect 6165 10205 6195 10235
rect 6195 10205 6196 10235
rect 6164 10204 6196 10205
rect 6164 10155 6196 10156
rect 6164 10125 6165 10155
rect 6165 10125 6195 10155
rect 6195 10125 6196 10155
rect 6164 10124 6196 10125
rect 6164 10075 6196 10076
rect 6164 10045 6165 10075
rect 6165 10045 6195 10075
rect 6195 10045 6196 10075
rect 6164 10044 6196 10045
rect 6164 9995 6196 9996
rect 6164 9965 6165 9995
rect 6165 9965 6195 9995
rect 6195 9965 6196 9995
rect 6164 9964 6196 9965
rect 6164 9915 6196 9916
rect 6164 9885 6165 9915
rect 6165 9885 6195 9915
rect 6195 9885 6196 9915
rect 6164 9884 6196 9885
rect 6164 9835 6196 9836
rect 6164 9805 6165 9835
rect 6165 9805 6195 9835
rect 6195 9805 6196 9835
rect 6164 9804 6196 9805
rect 6164 9755 6196 9756
rect 6164 9725 6165 9755
rect 6165 9725 6195 9755
rect 6195 9725 6196 9755
rect 6164 9724 6196 9725
rect 6164 9675 6196 9676
rect 6164 9645 6165 9675
rect 6165 9645 6195 9675
rect 6195 9645 6196 9675
rect 6164 9644 6196 9645
rect 6164 9595 6196 9596
rect 6164 9565 6165 9595
rect 6165 9565 6195 9595
rect 6195 9565 6196 9595
rect 6164 9564 6196 9565
rect 6164 9515 6196 9516
rect 6164 9485 6165 9515
rect 6165 9485 6195 9515
rect 6195 9485 6196 9515
rect 6164 9484 6196 9485
rect 6164 9435 6196 9436
rect 6164 9405 6165 9435
rect 6165 9405 6195 9435
rect 6195 9405 6196 9435
rect 6164 9404 6196 9405
rect 6164 9355 6196 9356
rect 6164 9325 6165 9355
rect 6165 9325 6195 9355
rect 6195 9325 6196 9355
rect 6164 9324 6196 9325
rect 6164 9275 6196 9276
rect 6164 9245 6165 9275
rect 6165 9245 6195 9275
rect 6195 9245 6196 9275
rect 6164 9244 6196 9245
rect 6164 9115 6196 9116
rect 6164 9085 6165 9115
rect 6165 9085 6195 9115
rect 6195 9085 6196 9115
rect 6164 9084 6196 9085
rect 6164 9035 6196 9036
rect 6164 9005 6165 9035
rect 6165 9005 6195 9035
rect 6195 9005 6196 9035
rect 6164 9004 6196 9005
rect 6164 8955 6196 8956
rect 6164 8925 6165 8955
rect 6165 8925 6195 8955
rect 6195 8925 6196 8955
rect 6164 8924 6196 8925
rect 6164 8635 6196 8636
rect 6164 8605 6165 8635
rect 6165 8605 6195 8635
rect 6195 8605 6196 8635
rect 6164 8604 6196 8605
rect 6164 8555 6196 8556
rect 6164 8525 6165 8555
rect 6165 8525 6195 8555
rect 6195 8525 6196 8555
rect 6164 8524 6196 8525
rect 6164 8395 6196 8396
rect 6164 8365 6165 8395
rect 6165 8365 6195 8395
rect 6195 8365 6196 8395
rect 6164 8364 6196 8365
rect 6164 8235 6196 8236
rect 6164 8205 6165 8235
rect 6165 8205 6195 8235
rect 6195 8205 6196 8235
rect 6164 8204 6196 8205
rect 6164 8155 6196 8156
rect 6164 8125 6165 8155
rect 6165 8125 6195 8155
rect 6195 8125 6196 8155
rect 6164 8124 6196 8125
rect 6164 8075 6196 8076
rect 6164 8045 6165 8075
rect 6165 8045 6195 8075
rect 6195 8045 6196 8075
rect 6164 8044 6196 8045
rect 6164 7995 6196 7996
rect 6164 7965 6165 7995
rect 6165 7965 6195 7995
rect 6195 7965 6196 7995
rect 6164 7964 6196 7965
rect 6164 7915 6196 7916
rect 6164 7885 6165 7915
rect 6165 7885 6195 7915
rect 6195 7885 6196 7915
rect 6164 7884 6196 7885
rect 6164 7835 6196 7836
rect 6164 7805 6165 7835
rect 6165 7805 6195 7835
rect 6195 7805 6196 7835
rect 6164 7804 6196 7805
rect 6164 7755 6196 7756
rect 6164 7725 6165 7755
rect 6165 7725 6195 7755
rect 6195 7725 6196 7755
rect 6164 7724 6196 7725
rect 6164 7675 6196 7676
rect 6164 7645 6165 7675
rect 6165 7645 6195 7675
rect 6195 7645 6196 7675
rect 6164 7644 6196 7645
rect 6164 7595 6196 7596
rect 6164 7565 6165 7595
rect 6165 7565 6195 7595
rect 6195 7565 6196 7595
rect 6164 7564 6196 7565
rect 6164 7515 6196 7516
rect 6164 7485 6165 7515
rect 6165 7485 6195 7515
rect 6195 7485 6196 7515
rect 6164 7484 6196 7485
rect 6164 7435 6196 7436
rect 6164 7405 6165 7435
rect 6165 7405 6195 7435
rect 6195 7405 6196 7435
rect 6164 7404 6196 7405
rect 6164 7355 6196 7356
rect 6164 7325 6165 7355
rect 6165 7325 6195 7355
rect 6195 7325 6196 7355
rect 6164 7324 6196 7325
rect 6164 7275 6196 7276
rect 6164 7245 6165 7275
rect 6165 7245 6195 7275
rect 6195 7245 6196 7275
rect 6164 7244 6196 7245
rect 6164 7195 6196 7196
rect 6164 7165 6165 7195
rect 6165 7165 6195 7195
rect 6195 7165 6196 7195
rect 6164 7164 6196 7165
rect 6164 7115 6196 7116
rect 6164 7085 6165 7115
rect 6165 7085 6195 7115
rect 6195 7085 6196 7115
rect 6164 7084 6196 7085
rect 6164 7035 6196 7036
rect 6164 7005 6165 7035
rect 6165 7005 6195 7035
rect 6195 7005 6196 7035
rect 6164 7004 6196 7005
rect 6164 6955 6196 6956
rect 6164 6925 6165 6955
rect 6165 6925 6195 6955
rect 6195 6925 6196 6955
rect 6164 6924 6196 6925
rect 6164 6795 6196 6796
rect 6164 6765 6165 6795
rect 6165 6765 6195 6795
rect 6195 6765 6196 6795
rect 6164 6764 6196 6765
rect 6164 6715 6196 6716
rect 6164 6685 6165 6715
rect 6165 6685 6195 6715
rect 6195 6685 6196 6715
rect 6164 6684 6196 6685
rect 6164 6635 6196 6636
rect 6164 6605 6165 6635
rect 6165 6605 6195 6635
rect 6195 6605 6196 6635
rect 6164 6604 6196 6605
rect 6164 6555 6196 6556
rect 6164 6525 6165 6555
rect 6165 6525 6195 6555
rect 6195 6525 6196 6555
rect 6164 6524 6196 6525
rect 6164 6475 6196 6476
rect 6164 6445 6165 6475
rect 6165 6445 6195 6475
rect 6195 6445 6196 6475
rect 6164 6444 6196 6445
rect 6164 6315 6196 6316
rect 6164 6285 6165 6315
rect 6165 6285 6195 6315
rect 6195 6285 6196 6315
rect 6164 6284 6196 6285
rect 6164 6235 6196 6236
rect 6164 6205 6165 6235
rect 6165 6205 6195 6235
rect 6195 6205 6196 6235
rect 6164 6204 6196 6205
rect 6164 6155 6196 6156
rect 6164 6125 6165 6155
rect 6165 6125 6195 6155
rect 6195 6125 6196 6155
rect 6164 6124 6196 6125
rect 6164 5995 6196 5996
rect 6164 5965 6165 5995
rect 6165 5965 6195 5995
rect 6195 5965 6196 5995
rect 6164 5964 6196 5965
rect 6164 5835 6196 5836
rect 6164 5805 6165 5835
rect 6165 5805 6195 5835
rect 6195 5805 6196 5835
rect 6164 5804 6196 5805
rect 6164 5755 6196 5756
rect 6164 5725 6165 5755
rect 6165 5725 6195 5755
rect 6195 5725 6196 5755
rect 6164 5724 6196 5725
rect 6164 5675 6196 5676
rect 6164 5645 6165 5675
rect 6165 5645 6195 5675
rect 6195 5645 6196 5675
rect 6164 5644 6196 5645
rect 6164 5595 6196 5596
rect 6164 5565 6165 5595
rect 6165 5565 6195 5595
rect 6195 5565 6196 5595
rect 6164 5564 6196 5565
rect 6164 5515 6196 5516
rect 6164 5485 6165 5515
rect 6165 5485 6195 5515
rect 6195 5485 6196 5515
rect 6164 5484 6196 5485
rect 6164 5435 6196 5436
rect 6164 5405 6165 5435
rect 6165 5405 6195 5435
rect 6195 5405 6196 5435
rect 6164 5404 6196 5405
rect 6164 5355 6196 5356
rect 6164 5325 6165 5355
rect 6165 5325 6195 5355
rect 6195 5325 6196 5355
rect 6164 5324 6196 5325
rect 6164 5275 6196 5276
rect 6164 5245 6165 5275
rect 6165 5245 6195 5275
rect 6195 5245 6196 5275
rect 6164 5244 6196 5245
rect 6164 5195 6196 5196
rect 6164 5165 6165 5195
rect 6165 5165 6195 5195
rect 6195 5165 6196 5195
rect 6164 5164 6196 5165
rect 6164 5115 6196 5116
rect 6164 5085 6165 5115
rect 6165 5085 6195 5115
rect 6195 5085 6196 5115
rect 6164 5084 6196 5085
rect 6164 5035 6196 5036
rect 6164 5005 6165 5035
rect 6165 5005 6195 5035
rect 6195 5005 6196 5035
rect 6164 5004 6196 5005
rect 6164 4955 6196 4956
rect 6164 4925 6165 4955
rect 6165 4925 6195 4955
rect 6195 4925 6196 4955
rect 6164 4924 6196 4925
rect 6164 4875 6196 4876
rect 6164 4845 6165 4875
rect 6165 4845 6195 4875
rect 6195 4845 6196 4875
rect 6164 4844 6196 4845
rect 6164 4795 6196 4796
rect 6164 4765 6165 4795
rect 6165 4765 6195 4795
rect 6195 4765 6196 4795
rect 6164 4764 6196 4765
rect 6164 4715 6196 4716
rect 6164 4685 6165 4715
rect 6165 4685 6195 4715
rect 6195 4685 6196 4715
rect 6164 4684 6196 4685
rect 6164 4635 6196 4636
rect 6164 4605 6165 4635
rect 6165 4605 6195 4635
rect 6195 4605 6196 4635
rect 6164 4604 6196 4605
rect 6164 4555 6196 4556
rect 6164 4525 6165 4555
rect 6165 4525 6195 4555
rect 6195 4525 6196 4555
rect 6164 4524 6196 4525
rect 6164 4395 6196 4396
rect 6164 4365 6165 4395
rect 6165 4365 6195 4395
rect 6195 4365 6196 4395
rect 6164 4364 6196 4365
rect 6164 4315 6196 4316
rect 6164 4285 6165 4315
rect 6165 4285 6195 4315
rect 6195 4285 6196 4315
rect 6164 4284 6196 4285
rect 6164 4235 6196 4236
rect 6164 4205 6165 4235
rect 6165 4205 6195 4235
rect 6195 4205 6196 4235
rect 6164 4204 6196 4205
rect 6164 4155 6196 4156
rect 6164 4125 6165 4155
rect 6165 4125 6195 4155
rect 6195 4125 6196 4155
rect 6164 4124 6196 4125
rect 6164 4075 6196 4076
rect 6164 4045 6165 4075
rect 6165 4045 6195 4075
rect 6195 4045 6196 4075
rect 6164 4044 6196 4045
rect 6164 3915 6196 3916
rect 6164 3885 6165 3915
rect 6165 3885 6195 3915
rect 6195 3885 6196 3915
rect 6164 3884 6196 3885
rect 6164 3835 6196 3836
rect 6164 3805 6165 3835
rect 6165 3805 6195 3835
rect 6195 3805 6196 3835
rect 6164 3804 6196 3805
rect 6164 3755 6196 3756
rect 6164 3725 6165 3755
rect 6165 3725 6195 3755
rect 6195 3725 6196 3755
rect 6164 3724 6196 3725
rect 6164 3595 6196 3596
rect 6164 3565 6165 3595
rect 6165 3565 6195 3595
rect 6195 3565 6196 3595
rect 6164 3564 6196 3565
rect 6164 3435 6196 3436
rect 6164 3405 6165 3435
rect 6165 3405 6195 3435
rect 6195 3405 6196 3435
rect 6164 3404 6196 3405
rect 6164 3355 6196 3356
rect 6164 3325 6165 3355
rect 6165 3325 6195 3355
rect 6195 3325 6196 3355
rect 6164 3324 6196 3325
rect 6164 3275 6196 3276
rect 6164 3245 6165 3275
rect 6165 3245 6195 3275
rect 6195 3245 6196 3275
rect 6164 3244 6196 3245
rect 6164 3195 6196 3196
rect 6164 3165 6165 3195
rect 6165 3165 6195 3195
rect 6195 3165 6196 3195
rect 6164 3164 6196 3165
rect 6164 3115 6196 3116
rect 6164 3085 6165 3115
rect 6165 3085 6195 3115
rect 6195 3085 6196 3115
rect 6164 3084 6196 3085
rect 6164 3035 6196 3036
rect 6164 3005 6165 3035
rect 6165 3005 6195 3035
rect 6195 3005 6196 3035
rect 6164 3004 6196 3005
rect 6164 2955 6196 2956
rect 6164 2925 6165 2955
rect 6165 2925 6195 2955
rect 6195 2925 6196 2955
rect 6164 2924 6196 2925
rect 6164 2875 6196 2876
rect 6164 2845 6165 2875
rect 6165 2845 6195 2875
rect 6195 2845 6196 2875
rect 6164 2844 6196 2845
rect 6164 2795 6196 2796
rect 6164 2765 6165 2795
rect 6165 2765 6195 2795
rect 6195 2765 6196 2795
rect 6164 2764 6196 2765
rect 6164 2715 6196 2716
rect 6164 2685 6165 2715
rect 6165 2685 6195 2715
rect 6195 2685 6196 2715
rect 6164 2684 6196 2685
rect 6164 2635 6196 2636
rect 6164 2605 6165 2635
rect 6165 2605 6195 2635
rect 6195 2605 6196 2635
rect 6164 2604 6196 2605
rect 6164 2555 6196 2556
rect 6164 2525 6165 2555
rect 6165 2525 6195 2555
rect 6195 2525 6196 2555
rect 6164 2524 6196 2525
rect 6164 2475 6196 2476
rect 6164 2445 6165 2475
rect 6165 2445 6195 2475
rect 6195 2445 6196 2475
rect 6164 2444 6196 2445
rect 6164 2395 6196 2396
rect 6164 2365 6165 2395
rect 6165 2365 6195 2395
rect 6195 2365 6196 2395
rect 6164 2364 6196 2365
rect 6164 2315 6196 2316
rect 6164 2285 6165 2315
rect 6165 2285 6195 2315
rect 6195 2285 6196 2315
rect 6164 2284 6196 2285
rect 6164 2235 6196 2236
rect 6164 2205 6165 2235
rect 6165 2205 6195 2235
rect 6195 2205 6196 2235
rect 6164 2204 6196 2205
rect 6164 2155 6196 2156
rect 6164 2125 6165 2155
rect 6165 2125 6195 2155
rect 6195 2125 6196 2155
rect 6164 2124 6196 2125
rect 6164 2075 6196 2076
rect 6164 2045 6165 2075
rect 6165 2045 6195 2075
rect 6195 2045 6196 2075
rect 6164 2044 6196 2045
rect 6164 1995 6196 1996
rect 6164 1965 6165 1995
rect 6165 1965 6195 1995
rect 6195 1965 6196 1995
rect 6164 1964 6196 1965
rect 6164 1915 6196 1916
rect 6164 1885 6165 1915
rect 6165 1885 6195 1915
rect 6195 1885 6196 1915
rect 6164 1884 6196 1885
rect 6164 1835 6196 1836
rect 6164 1805 6165 1835
rect 6165 1805 6195 1835
rect 6195 1805 6196 1835
rect 6164 1804 6196 1805
rect 6164 1755 6196 1756
rect 6164 1725 6165 1755
rect 6165 1725 6195 1755
rect 6195 1725 6196 1755
rect 6164 1724 6196 1725
rect 6164 1675 6196 1676
rect 6164 1645 6165 1675
rect 6165 1645 6195 1675
rect 6195 1645 6196 1675
rect 6164 1644 6196 1645
rect 6164 1595 6196 1596
rect 6164 1565 6165 1595
rect 6165 1565 6195 1595
rect 6195 1565 6196 1595
rect 6164 1564 6196 1565
rect 6164 1515 6196 1516
rect 6164 1485 6165 1515
rect 6165 1485 6195 1515
rect 6195 1485 6196 1515
rect 6164 1484 6196 1485
rect 6164 1435 6196 1436
rect 6164 1405 6165 1435
rect 6165 1405 6195 1435
rect 6195 1405 6196 1435
rect 6164 1404 6196 1405
rect 6164 1355 6196 1356
rect 6164 1325 6165 1355
rect 6165 1325 6195 1355
rect 6195 1325 6196 1355
rect 6164 1324 6196 1325
rect 6164 1275 6196 1276
rect 6164 1245 6165 1275
rect 6165 1245 6195 1275
rect 6195 1245 6196 1275
rect 6164 1244 6196 1245
rect 6164 1195 6196 1196
rect 6164 1165 6165 1195
rect 6165 1165 6195 1195
rect 6195 1165 6196 1195
rect 6164 1164 6196 1165
rect 6164 1115 6196 1116
rect 6164 1085 6165 1115
rect 6165 1085 6195 1115
rect 6195 1085 6196 1115
rect 6164 1084 6196 1085
rect 6164 1035 6196 1036
rect 6164 1005 6165 1035
rect 6165 1005 6195 1035
rect 6195 1005 6196 1035
rect 6164 1004 6196 1005
rect 6164 955 6196 956
rect 6164 925 6165 955
rect 6165 925 6195 955
rect 6195 925 6196 955
rect 6164 924 6196 925
rect 6164 875 6196 876
rect 6164 845 6165 875
rect 6165 845 6195 875
rect 6195 845 6196 875
rect 6164 844 6196 845
rect 6164 795 6196 796
rect 6164 765 6165 795
rect 6165 765 6195 795
rect 6195 765 6196 795
rect 6164 764 6196 765
rect 6164 715 6196 716
rect 6164 685 6165 715
rect 6165 685 6195 715
rect 6195 685 6196 715
rect 6164 684 6196 685
rect 6164 595 6196 596
rect 6164 565 6165 595
rect 6165 565 6195 595
rect 6195 565 6196 595
rect 6164 564 6196 565
rect 6164 515 6196 516
rect 6164 485 6165 515
rect 6165 485 6195 515
rect 6195 485 6196 515
rect 6164 484 6196 485
rect 6164 435 6196 436
rect 6164 405 6165 435
rect 6165 405 6195 435
rect 6195 405 6196 435
rect 6164 404 6196 405
rect 6164 355 6196 356
rect 6164 325 6165 355
rect 6165 325 6195 355
rect 6195 325 6196 355
rect 6164 324 6196 325
rect 6164 275 6196 276
rect 6164 245 6165 275
rect 6165 245 6195 275
rect 6195 245 6196 275
rect 6164 244 6196 245
rect 6164 195 6196 196
rect 6164 165 6165 195
rect 6165 165 6195 195
rect 6195 165 6196 195
rect 6164 164 6196 165
rect 6164 115 6196 116
rect 6164 85 6165 115
rect 6165 85 6195 115
rect 6195 85 6196 115
rect 6164 84 6196 85
rect 6164 35 6196 36
rect 6164 5 6165 35
rect 6165 5 6195 35
rect 6195 5 6196 35
rect 6164 4 6196 5
rect 6484 16644 6516 16836
rect 6324 16595 6356 16596
rect 6324 16565 6325 16595
rect 6325 16565 6355 16595
rect 6355 16565 6356 16595
rect 6324 16564 6356 16565
rect 6324 16515 6356 16516
rect 6324 16485 6325 16515
rect 6325 16485 6355 16515
rect 6355 16485 6356 16515
rect 6324 16484 6356 16485
rect 6324 16435 6356 16436
rect 6324 16405 6325 16435
rect 6325 16405 6355 16435
rect 6355 16405 6356 16435
rect 6324 16404 6356 16405
rect 6324 16355 6356 16356
rect 6324 16325 6325 16355
rect 6325 16325 6355 16355
rect 6355 16325 6356 16355
rect 6324 16324 6356 16325
rect 6324 16275 6356 16276
rect 6324 16245 6325 16275
rect 6325 16245 6355 16275
rect 6355 16245 6356 16275
rect 6324 16244 6356 16245
rect 6324 16195 6356 16196
rect 6324 16165 6325 16195
rect 6325 16165 6355 16195
rect 6355 16165 6356 16195
rect 6324 16164 6356 16165
rect 6324 16115 6356 16116
rect 6324 16085 6325 16115
rect 6325 16085 6355 16115
rect 6355 16085 6356 16115
rect 6324 16084 6356 16085
rect 6324 16035 6356 16036
rect 6324 16005 6325 16035
rect 6325 16005 6355 16035
rect 6355 16005 6356 16035
rect 6324 16004 6356 16005
rect 6324 15955 6356 15956
rect 6324 15925 6325 15955
rect 6325 15925 6355 15955
rect 6355 15925 6356 15955
rect 6324 15924 6356 15925
rect 6324 15435 6356 15436
rect 6324 15405 6325 15435
rect 6325 15405 6355 15435
rect 6355 15405 6356 15435
rect 6324 15404 6356 15405
rect 6324 15355 6356 15356
rect 6324 15325 6325 15355
rect 6325 15325 6355 15355
rect 6355 15325 6356 15355
rect 6324 15324 6356 15325
rect 6324 15275 6356 15276
rect 6324 15245 6325 15275
rect 6325 15245 6355 15275
rect 6355 15245 6356 15275
rect 6324 15244 6356 15245
rect 6324 15195 6356 15196
rect 6324 15165 6325 15195
rect 6325 15165 6355 15195
rect 6355 15165 6356 15195
rect 6324 15164 6356 15165
rect 6324 15115 6356 15116
rect 6324 15085 6325 15115
rect 6325 15085 6355 15115
rect 6355 15085 6356 15115
rect 6324 15084 6356 15085
rect 6324 15035 6356 15036
rect 6324 15005 6325 15035
rect 6325 15005 6355 15035
rect 6355 15005 6356 15035
rect 6324 15004 6356 15005
rect 6324 14955 6356 14956
rect 6324 14925 6325 14955
rect 6325 14925 6355 14955
rect 6355 14925 6356 14955
rect 6324 14924 6356 14925
rect 6324 14875 6356 14876
rect 6324 14845 6325 14875
rect 6325 14845 6355 14875
rect 6355 14845 6356 14875
rect 6324 14844 6356 14845
rect 6324 14795 6356 14796
rect 6324 14765 6325 14795
rect 6325 14765 6355 14795
rect 6355 14765 6356 14795
rect 6324 14764 6356 14765
rect 6324 14715 6356 14716
rect 6324 14685 6325 14715
rect 6325 14685 6355 14715
rect 6355 14685 6356 14715
rect 6324 14684 6356 14685
rect 6324 14635 6356 14636
rect 6324 14605 6325 14635
rect 6325 14605 6355 14635
rect 6355 14605 6356 14635
rect 6324 14604 6356 14605
rect 6324 14555 6356 14556
rect 6324 14525 6325 14555
rect 6325 14525 6355 14555
rect 6355 14525 6356 14555
rect 6324 14524 6356 14525
rect 6324 14475 6356 14476
rect 6324 14445 6325 14475
rect 6325 14445 6355 14475
rect 6355 14445 6356 14475
rect 6324 14444 6356 14445
rect 6324 13995 6356 13996
rect 6324 13965 6325 13995
rect 6325 13965 6355 13995
rect 6355 13965 6356 13995
rect 6324 13964 6356 13965
rect 6324 13875 6356 13876
rect 6324 13845 6325 13875
rect 6325 13845 6355 13875
rect 6355 13845 6356 13875
rect 6324 13844 6356 13845
rect 6324 13795 6356 13796
rect 6324 13765 6325 13795
rect 6325 13765 6355 13795
rect 6355 13765 6356 13795
rect 6324 13764 6356 13765
rect 6324 13715 6356 13716
rect 6324 13685 6325 13715
rect 6325 13685 6355 13715
rect 6355 13685 6356 13715
rect 6324 13684 6356 13685
rect 6324 13635 6356 13636
rect 6324 13605 6325 13635
rect 6325 13605 6355 13635
rect 6355 13605 6356 13635
rect 6324 13604 6356 13605
rect 6324 13555 6356 13556
rect 6324 13525 6325 13555
rect 6325 13525 6355 13555
rect 6355 13525 6356 13555
rect 6324 13524 6356 13525
rect 6324 13475 6356 13476
rect 6324 13445 6325 13475
rect 6325 13445 6355 13475
rect 6355 13445 6356 13475
rect 6324 13444 6356 13445
rect 6324 13395 6356 13396
rect 6324 13365 6325 13395
rect 6325 13365 6355 13395
rect 6355 13365 6356 13395
rect 6324 13364 6356 13365
rect 6324 13315 6356 13316
rect 6324 13285 6325 13315
rect 6325 13285 6355 13315
rect 6355 13285 6356 13315
rect 6324 13284 6356 13285
rect 6324 13235 6356 13236
rect 6324 13205 6325 13235
rect 6325 13205 6355 13235
rect 6355 13205 6356 13235
rect 6324 13204 6356 13205
rect 6324 13155 6356 13156
rect 6324 13125 6325 13155
rect 6325 13125 6355 13155
rect 6355 13125 6356 13155
rect 6324 13124 6356 13125
rect 6324 13075 6356 13076
rect 6324 13045 6325 13075
rect 6325 13045 6355 13075
rect 6355 13045 6356 13075
rect 6324 13044 6356 13045
rect 6324 12995 6356 12996
rect 6324 12965 6325 12995
rect 6325 12965 6355 12995
rect 6355 12965 6356 12995
rect 6324 12964 6356 12965
rect 6324 12515 6356 12516
rect 6324 12485 6325 12515
rect 6325 12485 6355 12515
rect 6355 12485 6356 12515
rect 6324 12484 6356 12485
rect 6324 12435 6356 12436
rect 6324 12405 6325 12435
rect 6325 12405 6355 12435
rect 6355 12405 6356 12435
rect 6324 12404 6356 12405
rect 6324 12315 6356 12316
rect 6324 12285 6325 12315
rect 6325 12285 6355 12315
rect 6355 12285 6356 12315
rect 6324 12284 6356 12285
rect 6324 12235 6356 12236
rect 6324 12205 6325 12235
rect 6325 12205 6355 12235
rect 6355 12205 6356 12235
rect 6324 12204 6356 12205
rect 6324 12155 6356 12156
rect 6324 12125 6325 12155
rect 6325 12125 6355 12155
rect 6355 12125 6356 12155
rect 6324 12124 6356 12125
rect 6324 12075 6356 12076
rect 6324 12045 6325 12075
rect 6325 12045 6355 12075
rect 6355 12045 6356 12075
rect 6324 12044 6356 12045
rect 6324 11995 6356 11996
rect 6324 11965 6325 11995
rect 6325 11965 6355 11995
rect 6355 11965 6356 11995
rect 6324 11964 6356 11965
rect 6324 11915 6356 11916
rect 6324 11885 6325 11915
rect 6325 11885 6355 11915
rect 6355 11885 6356 11915
rect 6324 11884 6356 11885
rect 6324 11835 6356 11836
rect 6324 11805 6325 11835
rect 6325 11805 6355 11835
rect 6355 11805 6356 11835
rect 6324 11804 6356 11805
rect 6324 11755 6356 11756
rect 6324 11725 6325 11755
rect 6325 11725 6355 11755
rect 6355 11725 6356 11755
rect 6324 11724 6356 11725
rect 6324 11675 6356 11676
rect 6324 11645 6325 11675
rect 6325 11645 6355 11675
rect 6355 11645 6356 11675
rect 6324 11644 6356 11645
rect 6324 11595 6356 11596
rect 6324 11565 6325 11595
rect 6325 11565 6355 11595
rect 6355 11565 6356 11595
rect 6324 11564 6356 11565
rect 6324 11515 6356 11516
rect 6324 11485 6325 11515
rect 6325 11485 6355 11515
rect 6355 11485 6356 11515
rect 6324 11484 6356 11485
rect 6324 11435 6356 11436
rect 6324 11405 6325 11435
rect 6325 11405 6355 11435
rect 6355 11405 6356 11435
rect 6324 11404 6356 11405
rect 6324 11355 6356 11356
rect 6324 11325 6325 11355
rect 6325 11325 6355 11355
rect 6355 11325 6356 11355
rect 6324 11324 6356 11325
rect 6324 11195 6356 11196
rect 6324 11165 6325 11195
rect 6325 11165 6355 11195
rect 6355 11165 6356 11195
rect 6324 11164 6356 11165
rect 6324 11115 6356 11116
rect 6324 11085 6325 11115
rect 6325 11085 6355 11115
rect 6355 11085 6356 11115
rect 6324 11084 6356 11085
rect 6324 11035 6356 11036
rect 6324 11005 6325 11035
rect 6325 11005 6355 11035
rect 6355 11005 6356 11035
rect 6324 11004 6356 11005
rect 6324 10875 6356 10876
rect 6324 10845 6325 10875
rect 6325 10845 6355 10875
rect 6355 10845 6356 10875
rect 6324 10844 6356 10845
rect 6324 10715 6356 10716
rect 6324 10685 6325 10715
rect 6325 10685 6355 10715
rect 6355 10685 6356 10715
rect 6324 10684 6356 10685
rect 6324 10635 6356 10636
rect 6324 10605 6325 10635
rect 6325 10605 6355 10635
rect 6355 10605 6356 10635
rect 6324 10604 6356 10605
rect 6324 10475 6356 10476
rect 6324 10445 6325 10475
rect 6325 10445 6355 10475
rect 6355 10445 6356 10475
rect 6324 10444 6356 10445
rect 6324 10315 6356 10316
rect 6324 10285 6325 10315
rect 6325 10285 6355 10315
rect 6355 10285 6356 10315
rect 6324 10284 6356 10285
rect 6324 10235 6356 10236
rect 6324 10205 6325 10235
rect 6325 10205 6355 10235
rect 6355 10205 6356 10235
rect 6324 10204 6356 10205
rect 6324 10155 6356 10156
rect 6324 10125 6325 10155
rect 6325 10125 6355 10155
rect 6355 10125 6356 10155
rect 6324 10124 6356 10125
rect 6324 10075 6356 10076
rect 6324 10045 6325 10075
rect 6325 10045 6355 10075
rect 6355 10045 6356 10075
rect 6324 10044 6356 10045
rect 6324 9995 6356 9996
rect 6324 9965 6325 9995
rect 6325 9965 6355 9995
rect 6355 9965 6356 9995
rect 6324 9964 6356 9965
rect 6324 9915 6356 9916
rect 6324 9885 6325 9915
rect 6325 9885 6355 9915
rect 6355 9885 6356 9915
rect 6324 9884 6356 9885
rect 6324 9835 6356 9836
rect 6324 9805 6325 9835
rect 6325 9805 6355 9835
rect 6355 9805 6356 9835
rect 6324 9804 6356 9805
rect 6324 9755 6356 9756
rect 6324 9725 6325 9755
rect 6325 9725 6355 9755
rect 6355 9725 6356 9755
rect 6324 9724 6356 9725
rect 6324 9675 6356 9676
rect 6324 9645 6325 9675
rect 6325 9645 6355 9675
rect 6355 9645 6356 9675
rect 6324 9644 6356 9645
rect 6324 9595 6356 9596
rect 6324 9565 6325 9595
rect 6325 9565 6355 9595
rect 6355 9565 6356 9595
rect 6324 9564 6356 9565
rect 6324 9515 6356 9516
rect 6324 9485 6325 9515
rect 6325 9485 6355 9515
rect 6355 9485 6356 9515
rect 6324 9484 6356 9485
rect 6324 9435 6356 9436
rect 6324 9405 6325 9435
rect 6325 9405 6355 9435
rect 6355 9405 6356 9435
rect 6324 9404 6356 9405
rect 6324 9355 6356 9356
rect 6324 9325 6325 9355
rect 6325 9325 6355 9355
rect 6355 9325 6356 9355
rect 6324 9324 6356 9325
rect 6324 9275 6356 9276
rect 6324 9245 6325 9275
rect 6325 9245 6355 9275
rect 6355 9245 6356 9275
rect 6324 9244 6356 9245
rect 6324 9115 6356 9116
rect 6324 9085 6325 9115
rect 6325 9085 6355 9115
rect 6355 9085 6356 9115
rect 6324 9084 6356 9085
rect 6324 9035 6356 9036
rect 6324 9005 6325 9035
rect 6325 9005 6355 9035
rect 6355 9005 6356 9035
rect 6324 9004 6356 9005
rect 6324 8955 6356 8956
rect 6324 8925 6325 8955
rect 6325 8925 6355 8955
rect 6355 8925 6356 8955
rect 6324 8924 6356 8925
rect 6324 8635 6356 8636
rect 6324 8605 6325 8635
rect 6325 8605 6355 8635
rect 6355 8605 6356 8635
rect 6324 8604 6356 8605
rect 6324 8555 6356 8556
rect 6324 8525 6325 8555
rect 6325 8525 6355 8555
rect 6355 8525 6356 8555
rect 6324 8524 6356 8525
rect 6324 8395 6356 8396
rect 6324 8365 6325 8395
rect 6325 8365 6355 8395
rect 6355 8365 6356 8395
rect 6324 8364 6356 8365
rect 6324 8235 6356 8236
rect 6324 8205 6325 8235
rect 6325 8205 6355 8235
rect 6355 8205 6356 8235
rect 6324 8204 6356 8205
rect 6324 8155 6356 8156
rect 6324 8125 6325 8155
rect 6325 8125 6355 8155
rect 6355 8125 6356 8155
rect 6324 8124 6356 8125
rect 6324 8075 6356 8076
rect 6324 8045 6325 8075
rect 6325 8045 6355 8075
rect 6355 8045 6356 8075
rect 6324 8044 6356 8045
rect 6324 7995 6356 7996
rect 6324 7965 6325 7995
rect 6325 7965 6355 7995
rect 6355 7965 6356 7995
rect 6324 7964 6356 7965
rect 6324 7915 6356 7916
rect 6324 7885 6325 7915
rect 6325 7885 6355 7915
rect 6355 7885 6356 7915
rect 6324 7884 6356 7885
rect 6324 7835 6356 7836
rect 6324 7805 6325 7835
rect 6325 7805 6355 7835
rect 6355 7805 6356 7835
rect 6324 7804 6356 7805
rect 6324 7755 6356 7756
rect 6324 7725 6325 7755
rect 6325 7725 6355 7755
rect 6355 7725 6356 7755
rect 6324 7724 6356 7725
rect 6324 7675 6356 7676
rect 6324 7645 6325 7675
rect 6325 7645 6355 7675
rect 6355 7645 6356 7675
rect 6324 7644 6356 7645
rect 6324 7595 6356 7596
rect 6324 7565 6325 7595
rect 6325 7565 6355 7595
rect 6355 7565 6356 7595
rect 6324 7564 6356 7565
rect 6324 7515 6356 7516
rect 6324 7485 6325 7515
rect 6325 7485 6355 7515
rect 6355 7485 6356 7515
rect 6324 7484 6356 7485
rect 6324 7435 6356 7436
rect 6324 7405 6325 7435
rect 6325 7405 6355 7435
rect 6355 7405 6356 7435
rect 6324 7404 6356 7405
rect 6324 7355 6356 7356
rect 6324 7325 6325 7355
rect 6325 7325 6355 7355
rect 6355 7325 6356 7355
rect 6324 7324 6356 7325
rect 6324 7275 6356 7276
rect 6324 7245 6325 7275
rect 6325 7245 6355 7275
rect 6355 7245 6356 7275
rect 6324 7244 6356 7245
rect 6324 7195 6356 7196
rect 6324 7165 6325 7195
rect 6325 7165 6355 7195
rect 6355 7165 6356 7195
rect 6324 7164 6356 7165
rect 6324 7115 6356 7116
rect 6324 7085 6325 7115
rect 6325 7085 6355 7115
rect 6355 7085 6356 7115
rect 6324 7084 6356 7085
rect 6324 7035 6356 7036
rect 6324 7005 6325 7035
rect 6325 7005 6355 7035
rect 6355 7005 6356 7035
rect 6324 7004 6356 7005
rect 6324 6955 6356 6956
rect 6324 6925 6325 6955
rect 6325 6925 6355 6955
rect 6355 6925 6356 6955
rect 6324 6924 6356 6925
rect 6324 6875 6356 6876
rect 6324 6845 6325 6875
rect 6325 6845 6355 6875
rect 6355 6845 6356 6875
rect 6324 6844 6356 6845
rect 6324 6795 6356 6796
rect 6324 6765 6325 6795
rect 6325 6765 6355 6795
rect 6355 6765 6356 6795
rect 6324 6764 6356 6765
rect 6324 6715 6356 6716
rect 6324 6685 6325 6715
rect 6325 6685 6355 6715
rect 6355 6685 6356 6715
rect 6324 6684 6356 6685
rect 6324 6635 6356 6636
rect 6324 6605 6325 6635
rect 6325 6605 6355 6635
rect 6355 6605 6356 6635
rect 6324 6604 6356 6605
rect 6324 6555 6356 6556
rect 6324 6525 6325 6555
rect 6325 6525 6355 6555
rect 6355 6525 6356 6555
rect 6324 6524 6356 6525
rect 6324 6475 6356 6476
rect 6324 6445 6325 6475
rect 6325 6445 6355 6475
rect 6355 6445 6356 6475
rect 6324 6444 6356 6445
rect 6324 6315 6356 6316
rect 6324 6285 6325 6315
rect 6325 6285 6355 6315
rect 6355 6285 6356 6315
rect 6324 6284 6356 6285
rect 6324 6235 6356 6236
rect 6324 6205 6325 6235
rect 6325 6205 6355 6235
rect 6355 6205 6356 6235
rect 6324 6204 6356 6205
rect 6324 6155 6356 6156
rect 6324 6125 6325 6155
rect 6325 6125 6355 6155
rect 6355 6125 6356 6155
rect 6324 6124 6356 6125
rect 6324 5995 6356 5996
rect 6324 5965 6325 5995
rect 6325 5965 6355 5995
rect 6355 5965 6356 5995
rect 6324 5964 6356 5965
rect 6324 5835 6356 5836
rect 6324 5805 6325 5835
rect 6325 5805 6355 5835
rect 6355 5805 6356 5835
rect 6324 5804 6356 5805
rect 6324 5755 6356 5756
rect 6324 5725 6325 5755
rect 6325 5725 6355 5755
rect 6355 5725 6356 5755
rect 6324 5724 6356 5725
rect 6324 5675 6356 5676
rect 6324 5645 6325 5675
rect 6325 5645 6355 5675
rect 6355 5645 6356 5675
rect 6324 5644 6356 5645
rect 6324 5595 6356 5596
rect 6324 5565 6325 5595
rect 6325 5565 6355 5595
rect 6355 5565 6356 5595
rect 6324 5564 6356 5565
rect 6324 5515 6356 5516
rect 6324 5485 6325 5515
rect 6325 5485 6355 5515
rect 6355 5485 6356 5515
rect 6324 5484 6356 5485
rect 6324 5435 6356 5436
rect 6324 5405 6325 5435
rect 6325 5405 6355 5435
rect 6355 5405 6356 5435
rect 6324 5404 6356 5405
rect 6324 5355 6356 5356
rect 6324 5325 6325 5355
rect 6325 5325 6355 5355
rect 6355 5325 6356 5355
rect 6324 5324 6356 5325
rect 6324 5275 6356 5276
rect 6324 5245 6325 5275
rect 6325 5245 6355 5275
rect 6355 5245 6356 5275
rect 6324 5244 6356 5245
rect 6324 5195 6356 5196
rect 6324 5165 6325 5195
rect 6325 5165 6355 5195
rect 6355 5165 6356 5195
rect 6324 5164 6356 5165
rect 6324 5115 6356 5116
rect 6324 5085 6325 5115
rect 6325 5085 6355 5115
rect 6355 5085 6356 5115
rect 6324 5084 6356 5085
rect 6324 5035 6356 5036
rect 6324 5005 6325 5035
rect 6325 5005 6355 5035
rect 6355 5005 6356 5035
rect 6324 5004 6356 5005
rect 6324 4955 6356 4956
rect 6324 4925 6325 4955
rect 6325 4925 6355 4955
rect 6355 4925 6356 4955
rect 6324 4924 6356 4925
rect 6324 4875 6356 4876
rect 6324 4845 6325 4875
rect 6325 4845 6355 4875
rect 6355 4845 6356 4875
rect 6324 4844 6356 4845
rect 6324 4795 6356 4796
rect 6324 4765 6325 4795
rect 6325 4765 6355 4795
rect 6355 4765 6356 4795
rect 6324 4764 6356 4765
rect 6324 4715 6356 4716
rect 6324 4685 6325 4715
rect 6325 4685 6355 4715
rect 6355 4685 6356 4715
rect 6324 4684 6356 4685
rect 6324 4635 6356 4636
rect 6324 4605 6325 4635
rect 6325 4605 6355 4635
rect 6355 4605 6356 4635
rect 6324 4604 6356 4605
rect 6324 4555 6356 4556
rect 6324 4525 6325 4555
rect 6325 4525 6355 4555
rect 6355 4525 6356 4555
rect 6324 4524 6356 4525
rect 6324 4475 6356 4476
rect 6324 4445 6325 4475
rect 6325 4445 6355 4475
rect 6355 4445 6356 4475
rect 6324 4444 6356 4445
rect 6324 4395 6356 4396
rect 6324 4365 6325 4395
rect 6325 4365 6355 4395
rect 6355 4365 6356 4395
rect 6324 4364 6356 4365
rect 6324 4315 6356 4316
rect 6324 4285 6325 4315
rect 6325 4285 6355 4315
rect 6355 4285 6356 4315
rect 6324 4284 6356 4285
rect 6324 4235 6356 4236
rect 6324 4205 6325 4235
rect 6325 4205 6355 4235
rect 6355 4205 6356 4235
rect 6324 4204 6356 4205
rect 6324 4155 6356 4156
rect 6324 4125 6325 4155
rect 6325 4125 6355 4155
rect 6355 4125 6356 4155
rect 6324 4124 6356 4125
rect 6324 4075 6356 4076
rect 6324 4045 6325 4075
rect 6325 4045 6355 4075
rect 6355 4045 6356 4075
rect 6324 4044 6356 4045
rect 6324 3915 6356 3916
rect 6324 3885 6325 3915
rect 6325 3885 6355 3915
rect 6355 3885 6356 3915
rect 6324 3884 6356 3885
rect 6324 3835 6356 3836
rect 6324 3805 6325 3835
rect 6325 3805 6355 3835
rect 6355 3805 6356 3835
rect 6324 3804 6356 3805
rect 6324 3755 6356 3756
rect 6324 3725 6325 3755
rect 6325 3725 6355 3755
rect 6355 3725 6356 3755
rect 6324 3724 6356 3725
rect 6324 3595 6356 3596
rect 6324 3565 6325 3595
rect 6325 3565 6355 3595
rect 6355 3565 6356 3595
rect 6324 3564 6356 3565
rect 6324 3435 6356 3436
rect 6324 3405 6325 3435
rect 6325 3405 6355 3435
rect 6355 3405 6356 3435
rect 6324 3404 6356 3405
rect 6324 3355 6356 3356
rect 6324 3325 6325 3355
rect 6325 3325 6355 3355
rect 6355 3325 6356 3355
rect 6324 3324 6356 3325
rect 6324 3275 6356 3276
rect 6324 3245 6325 3275
rect 6325 3245 6355 3275
rect 6355 3245 6356 3275
rect 6324 3244 6356 3245
rect 6324 3195 6356 3196
rect 6324 3165 6325 3195
rect 6325 3165 6355 3195
rect 6355 3165 6356 3195
rect 6324 3164 6356 3165
rect 6324 3115 6356 3116
rect 6324 3085 6325 3115
rect 6325 3085 6355 3115
rect 6355 3085 6356 3115
rect 6324 3084 6356 3085
rect 6324 3035 6356 3036
rect 6324 3005 6325 3035
rect 6325 3005 6355 3035
rect 6355 3005 6356 3035
rect 6324 3004 6356 3005
rect 6324 2955 6356 2956
rect 6324 2925 6325 2955
rect 6325 2925 6355 2955
rect 6355 2925 6356 2955
rect 6324 2924 6356 2925
rect 6324 2875 6356 2876
rect 6324 2845 6325 2875
rect 6325 2845 6355 2875
rect 6355 2845 6356 2875
rect 6324 2844 6356 2845
rect 6324 2795 6356 2796
rect 6324 2765 6325 2795
rect 6325 2765 6355 2795
rect 6355 2765 6356 2795
rect 6324 2764 6356 2765
rect 6324 2715 6356 2716
rect 6324 2685 6325 2715
rect 6325 2685 6355 2715
rect 6355 2685 6356 2715
rect 6324 2684 6356 2685
rect 6324 2635 6356 2636
rect 6324 2605 6325 2635
rect 6325 2605 6355 2635
rect 6355 2605 6356 2635
rect 6324 2604 6356 2605
rect 6324 2555 6356 2556
rect 6324 2525 6325 2555
rect 6325 2525 6355 2555
rect 6355 2525 6356 2555
rect 6324 2524 6356 2525
rect 6324 2475 6356 2476
rect 6324 2445 6325 2475
rect 6325 2445 6355 2475
rect 6355 2445 6356 2475
rect 6324 2444 6356 2445
rect 6324 2395 6356 2396
rect 6324 2365 6325 2395
rect 6325 2365 6355 2395
rect 6355 2365 6356 2395
rect 6324 2364 6356 2365
rect 6324 2315 6356 2316
rect 6324 2285 6325 2315
rect 6325 2285 6355 2315
rect 6355 2285 6356 2315
rect 6324 2284 6356 2285
rect 6324 2235 6356 2236
rect 6324 2205 6325 2235
rect 6325 2205 6355 2235
rect 6355 2205 6356 2235
rect 6324 2204 6356 2205
rect 6324 2155 6356 2156
rect 6324 2125 6325 2155
rect 6325 2125 6355 2155
rect 6355 2125 6356 2155
rect 6324 2124 6356 2125
rect 6324 2075 6356 2076
rect 6324 2045 6325 2075
rect 6325 2045 6355 2075
rect 6355 2045 6356 2075
rect 6324 2044 6356 2045
rect 6324 1995 6356 1996
rect 6324 1965 6325 1995
rect 6325 1965 6355 1995
rect 6355 1965 6356 1995
rect 6324 1964 6356 1965
rect 6324 1915 6356 1916
rect 6324 1885 6325 1915
rect 6325 1885 6355 1915
rect 6355 1885 6356 1915
rect 6324 1884 6356 1885
rect 6324 1835 6356 1836
rect 6324 1805 6325 1835
rect 6325 1805 6355 1835
rect 6355 1805 6356 1835
rect 6324 1804 6356 1805
rect 6324 1755 6356 1756
rect 6324 1725 6325 1755
rect 6325 1725 6355 1755
rect 6355 1725 6356 1755
rect 6324 1724 6356 1725
rect 6324 1675 6356 1676
rect 6324 1645 6325 1675
rect 6325 1645 6355 1675
rect 6355 1645 6356 1675
rect 6324 1644 6356 1645
rect 6324 1595 6356 1596
rect 6324 1565 6325 1595
rect 6325 1565 6355 1595
rect 6355 1565 6356 1595
rect 6324 1564 6356 1565
rect 6324 1515 6356 1516
rect 6324 1485 6325 1515
rect 6325 1485 6355 1515
rect 6355 1485 6356 1515
rect 6324 1484 6356 1485
rect 6324 1435 6356 1436
rect 6324 1405 6325 1435
rect 6325 1405 6355 1435
rect 6355 1405 6356 1435
rect 6324 1404 6356 1405
rect 6324 1355 6356 1356
rect 6324 1325 6325 1355
rect 6325 1325 6355 1355
rect 6355 1325 6356 1355
rect 6324 1324 6356 1325
rect 6324 1275 6356 1276
rect 6324 1245 6325 1275
rect 6325 1245 6355 1275
rect 6355 1245 6356 1275
rect 6324 1244 6356 1245
rect 6324 1195 6356 1196
rect 6324 1165 6325 1195
rect 6325 1165 6355 1195
rect 6355 1165 6356 1195
rect 6324 1164 6356 1165
rect 6324 1115 6356 1116
rect 6324 1085 6325 1115
rect 6325 1085 6355 1115
rect 6355 1085 6356 1115
rect 6324 1084 6356 1085
rect 6324 1035 6356 1036
rect 6324 1005 6325 1035
rect 6325 1005 6355 1035
rect 6355 1005 6356 1035
rect 6324 1004 6356 1005
rect 6324 955 6356 956
rect 6324 925 6325 955
rect 6325 925 6355 955
rect 6355 925 6356 955
rect 6324 924 6356 925
rect 6324 875 6356 876
rect 6324 845 6325 875
rect 6325 845 6355 875
rect 6355 845 6356 875
rect 6324 844 6356 845
rect 6324 795 6356 796
rect 6324 765 6325 795
rect 6325 765 6355 795
rect 6355 765 6356 795
rect 6324 764 6356 765
rect 6324 715 6356 716
rect 6324 685 6325 715
rect 6325 685 6355 715
rect 6355 685 6356 715
rect 6324 684 6356 685
rect 6324 595 6356 596
rect 6324 565 6325 595
rect 6325 565 6355 595
rect 6355 565 6356 595
rect 6324 564 6356 565
rect 6324 515 6356 516
rect 6324 485 6325 515
rect 6325 485 6355 515
rect 6355 485 6356 515
rect 6324 484 6356 485
rect 6324 435 6356 436
rect 6324 405 6325 435
rect 6325 405 6355 435
rect 6355 405 6356 435
rect 6324 404 6356 405
rect 6324 355 6356 356
rect 6324 325 6325 355
rect 6325 325 6355 355
rect 6355 325 6356 355
rect 6324 324 6356 325
rect 6324 275 6356 276
rect 6324 245 6325 275
rect 6325 245 6355 275
rect 6355 245 6356 275
rect 6324 244 6356 245
rect 6324 195 6356 196
rect 6324 165 6325 195
rect 6325 165 6355 195
rect 6355 165 6356 195
rect 6324 164 6356 165
rect 6324 115 6356 116
rect 6324 85 6325 115
rect 6325 85 6355 115
rect 6355 85 6356 115
rect 6324 84 6356 85
rect 6324 35 6356 36
rect 6324 5 6325 35
rect 6325 5 6355 35
rect 6355 5 6356 35
rect 6324 4 6356 5
rect 6644 16644 6676 16836
rect 6484 16595 6516 16596
rect 6484 16565 6485 16595
rect 6485 16565 6515 16595
rect 6515 16565 6516 16595
rect 6484 16564 6516 16565
rect 6484 16515 6516 16516
rect 6484 16485 6485 16515
rect 6485 16485 6515 16515
rect 6515 16485 6516 16515
rect 6484 16484 6516 16485
rect 6484 16435 6516 16436
rect 6484 16405 6485 16435
rect 6485 16405 6515 16435
rect 6515 16405 6516 16435
rect 6484 16404 6516 16405
rect 6484 16355 6516 16356
rect 6484 16325 6485 16355
rect 6485 16325 6515 16355
rect 6515 16325 6516 16355
rect 6484 16324 6516 16325
rect 6484 16275 6516 16276
rect 6484 16245 6485 16275
rect 6485 16245 6515 16275
rect 6515 16245 6516 16275
rect 6484 16244 6516 16245
rect 6484 16195 6516 16196
rect 6484 16165 6485 16195
rect 6485 16165 6515 16195
rect 6515 16165 6516 16195
rect 6484 16164 6516 16165
rect 6484 16115 6516 16116
rect 6484 16085 6485 16115
rect 6485 16085 6515 16115
rect 6515 16085 6516 16115
rect 6484 16084 6516 16085
rect 6484 16035 6516 16036
rect 6484 16005 6485 16035
rect 6485 16005 6515 16035
rect 6515 16005 6516 16035
rect 6484 16004 6516 16005
rect 6484 15955 6516 15956
rect 6484 15925 6485 15955
rect 6485 15925 6515 15955
rect 6515 15925 6516 15955
rect 6484 15924 6516 15925
rect 6484 15435 6516 15436
rect 6484 15405 6485 15435
rect 6485 15405 6515 15435
rect 6515 15405 6516 15435
rect 6484 15404 6516 15405
rect 6484 15355 6516 15356
rect 6484 15325 6485 15355
rect 6485 15325 6515 15355
rect 6515 15325 6516 15355
rect 6484 15324 6516 15325
rect 6484 15275 6516 15276
rect 6484 15245 6485 15275
rect 6485 15245 6515 15275
rect 6515 15245 6516 15275
rect 6484 15244 6516 15245
rect 6484 15195 6516 15196
rect 6484 15165 6485 15195
rect 6485 15165 6515 15195
rect 6515 15165 6516 15195
rect 6484 15164 6516 15165
rect 6484 15115 6516 15116
rect 6484 15085 6485 15115
rect 6485 15085 6515 15115
rect 6515 15085 6516 15115
rect 6484 15084 6516 15085
rect 6484 15035 6516 15036
rect 6484 15005 6485 15035
rect 6485 15005 6515 15035
rect 6515 15005 6516 15035
rect 6484 15004 6516 15005
rect 6484 14955 6516 14956
rect 6484 14925 6485 14955
rect 6485 14925 6515 14955
rect 6515 14925 6516 14955
rect 6484 14924 6516 14925
rect 6484 14875 6516 14876
rect 6484 14845 6485 14875
rect 6485 14845 6515 14875
rect 6515 14845 6516 14875
rect 6484 14844 6516 14845
rect 6484 14795 6516 14796
rect 6484 14765 6485 14795
rect 6485 14765 6515 14795
rect 6515 14765 6516 14795
rect 6484 14764 6516 14765
rect 6484 14715 6516 14716
rect 6484 14685 6485 14715
rect 6485 14685 6515 14715
rect 6515 14685 6516 14715
rect 6484 14684 6516 14685
rect 6484 14635 6516 14636
rect 6484 14605 6485 14635
rect 6485 14605 6515 14635
rect 6515 14605 6516 14635
rect 6484 14604 6516 14605
rect 6484 14555 6516 14556
rect 6484 14525 6485 14555
rect 6485 14525 6515 14555
rect 6515 14525 6516 14555
rect 6484 14524 6516 14525
rect 6484 14475 6516 14476
rect 6484 14445 6485 14475
rect 6485 14445 6515 14475
rect 6515 14445 6516 14475
rect 6484 14444 6516 14445
rect 6484 13995 6516 13996
rect 6484 13965 6485 13995
rect 6485 13965 6515 13995
rect 6515 13965 6516 13995
rect 6484 13964 6516 13965
rect 6484 13875 6516 13876
rect 6484 13845 6485 13875
rect 6485 13845 6515 13875
rect 6515 13845 6516 13875
rect 6484 13844 6516 13845
rect 6484 13795 6516 13796
rect 6484 13765 6485 13795
rect 6485 13765 6515 13795
rect 6515 13765 6516 13795
rect 6484 13764 6516 13765
rect 6484 13715 6516 13716
rect 6484 13685 6485 13715
rect 6485 13685 6515 13715
rect 6515 13685 6516 13715
rect 6484 13684 6516 13685
rect 6484 13635 6516 13636
rect 6484 13605 6485 13635
rect 6485 13605 6515 13635
rect 6515 13605 6516 13635
rect 6484 13604 6516 13605
rect 6484 13555 6516 13556
rect 6484 13525 6485 13555
rect 6485 13525 6515 13555
rect 6515 13525 6516 13555
rect 6484 13524 6516 13525
rect 6484 13475 6516 13476
rect 6484 13445 6485 13475
rect 6485 13445 6515 13475
rect 6515 13445 6516 13475
rect 6484 13444 6516 13445
rect 6484 13395 6516 13396
rect 6484 13365 6485 13395
rect 6485 13365 6515 13395
rect 6515 13365 6516 13395
rect 6484 13364 6516 13365
rect 6484 13315 6516 13316
rect 6484 13285 6485 13315
rect 6485 13285 6515 13315
rect 6515 13285 6516 13315
rect 6484 13284 6516 13285
rect 6484 13235 6516 13236
rect 6484 13205 6485 13235
rect 6485 13205 6515 13235
rect 6515 13205 6516 13235
rect 6484 13204 6516 13205
rect 6484 13155 6516 13156
rect 6484 13125 6485 13155
rect 6485 13125 6515 13155
rect 6515 13125 6516 13155
rect 6484 13124 6516 13125
rect 6484 13075 6516 13076
rect 6484 13045 6485 13075
rect 6485 13045 6515 13075
rect 6515 13045 6516 13075
rect 6484 13044 6516 13045
rect 6484 12995 6516 12996
rect 6484 12965 6485 12995
rect 6485 12965 6515 12995
rect 6515 12965 6516 12995
rect 6484 12964 6516 12965
rect 6484 12515 6516 12516
rect 6484 12485 6485 12515
rect 6485 12485 6515 12515
rect 6515 12485 6516 12515
rect 6484 12484 6516 12485
rect 6484 12435 6516 12436
rect 6484 12405 6485 12435
rect 6485 12405 6515 12435
rect 6515 12405 6516 12435
rect 6484 12404 6516 12405
rect 6484 12315 6516 12316
rect 6484 12285 6485 12315
rect 6485 12285 6515 12315
rect 6515 12285 6516 12315
rect 6484 12284 6516 12285
rect 6484 12235 6516 12236
rect 6484 12205 6485 12235
rect 6485 12205 6515 12235
rect 6515 12205 6516 12235
rect 6484 12204 6516 12205
rect 6484 12155 6516 12156
rect 6484 12125 6485 12155
rect 6485 12125 6515 12155
rect 6515 12125 6516 12155
rect 6484 12124 6516 12125
rect 6484 12075 6516 12076
rect 6484 12045 6485 12075
rect 6485 12045 6515 12075
rect 6515 12045 6516 12075
rect 6484 12044 6516 12045
rect 6484 11995 6516 11996
rect 6484 11965 6485 11995
rect 6485 11965 6515 11995
rect 6515 11965 6516 11995
rect 6484 11964 6516 11965
rect 6484 11915 6516 11916
rect 6484 11885 6485 11915
rect 6485 11885 6515 11915
rect 6515 11885 6516 11915
rect 6484 11884 6516 11885
rect 6484 11835 6516 11836
rect 6484 11805 6485 11835
rect 6485 11805 6515 11835
rect 6515 11805 6516 11835
rect 6484 11804 6516 11805
rect 6484 11755 6516 11756
rect 6484 11725 6485 11755
rect 6485 11725 6515 11755
rect 6515 11725 6516 11755
rect 6484 11724 6516 11725
rect 6484 11675 6516 11676
rect 6484 11645 6485 11675
rect 6485 11645 6515 11675
rect 6515 11645 6516 11675
rect 6484 11644 6516 11645
rect 6484 11595 6516 11596
rect 6484 11565 6485 11595
rect 6485 11565 6515 11595
rect 6515 11565 6516 11595
rect 6484 11564 6516 11565
rect 6484 11515 6516 11516
rect 6484 11485 6485 11515
rect 6485 11485 6515 11515
rect 6515 11485 6516 11515
rect 6484 11484 6516 11485
rect 6484 11435 6516 11436
rect 6484 11405 6485 11435
rect 6485 11405 6515 11435
rect 6515 11405 6516 11435
rect 6484 11404 6516 11405
rect 6484 11355 6516 11356
rect 6484 11325 6485 11355
rect 6485 11325 6515 11355
rect 6515 11325 6516 11355
rect 6484 11324 6516 11325
rect 6484 11195 6516 11196
rect 6484 11165 6485 11195
rect 6485 11165 6515 11195
rect 6515 11165 6516 11195
rect 6484 11164 6516 11165
rect 6484 11115 6516 11116
rect 6484 11085 6485 11115
rect 6485 11085 6515 11115
rect 6515 11085 6516 11115
rect 6484 11084 6516 11085
rect 6484 11035 6516 11036
rect 6484 11005 6485 11035
rect 6485 11005 6515 11035
rect 6515 11005 6516 11035
rect 6484 11004 6516 11005
rect 6484 10875 6516 10876
rect 6484 10845 6485 10875
rect 6485 10845 6515 10875
rect 6515 10845 6516 10875
rect 6484 10844 6516 10845
rect 6484 10715 6516 10716
rect 6484 10685 6485 10715
rect 6485 10685 6515 10715
rect 6515 10685 6516 10715
rect 6484 10684 6516 10685
rect 6484 10635 6516 10636
rect 6484 10605 6485 10635
rect 6485 10605 6515 10635
rect 6515 10605 6516 10635
rect 6484 10604 6516 10605
rect 6484 10475 6516 10476
rect 6484 10445 6485 10475
rect 6485 10445 6515 10475
rect 6515 10445 6516 10475
rect 6484 10444 6516 10445
rect 6484 10315 6516 10316
rect 6484 10285 6485 10315
rect 6485 10285 6515 10315
rect 6515 10285 6516 10315
rect 6484 10284 6516 10285
rect 6484 10235 6516 10236
rect 6484 10205 6485 10235
rect 6485 10205 6515 10235
rect 6515 10205 6516 10235
rect 6484 10204 6516 10205
rect 6484 10155 6516 10156
rect 6484 10125 6485 10155
rect 6485 10125 6515 10155
rect 6515 10125 6516 10155
rect 6484 10124 6516 10125
rect 6484 10075 6516 10076
rect 6484 10045 6485 10075
rect 6485 10045 6515 10075
rect 6515 10045 6516 10075
rect 6484 10044 6516 10045
rect 6484 9995 6516 9996
rect 6484 9965 6485 9995
rect 6485 9965 6515 9995
rect 6515 9965 6516 9995
rect 6484 9964 6516 9965
rect 6484 9915 6516 9916
rect 6484 9885 6485 9915
rect 6485 9885 6515 9915
rect 6515 9885 6516 9915
rect 6484 9884 6516 9885
rect 6484 9835 6516 9836
rect 6484 9805 6485 9835
rect 6485 9805 6515 9835
rect 6515 9805 6516 9835
rect 6484 9804 6516 9805
rect 6484 9755 6516 9756
rect 6484 9725 6485 9755
rect 6485 9725 6515 9755
rect 6515 9725 6516 9755
rect 6484 9724 6516 9725
rect 6484 9675 6516 9676
rect 6484 9645 6485 9675
rect 6485 9645 6515 9675
rect 6515 9645 6516 9675
rect 6484 9644 6516 9645
rect 6484 9595 6516 9596
rect 6484 9565 6485 9595
rect 6485 9565 6515 9595
rect 6515 9565 6516 9595
rect 6484 9564 6516 9565
rect 6484 9515 6516 9516
rect 6484 9485 6485 9515
rect 6485 9485 6515 9515
rect 6515 9485 6516 9515
rect 6484 9484 6516 9485
rect 6484 9435 6516 9436
rect 6484 9405 6485 9435
rect 6485 9405 6515 9435
rect 6515 9405 6516 9435
rect 6484 9404 6516 9405
rect 6484 9355 6516 9356
rect 6484 9325 6485 9355
rect 6485 9325 6515 9355
rect 6515 9325 6516 9355
rect 6484 9324 6516 9325
rect 6484 9275 6516 9276
rect 6484 9245 6485 9275
rect 6485 9245 6515 9275
rect 6515 9245 6516 9275
rect 6484 9244 6516 9245
rect 6484 9115 6516 9116
rect 6484 9085 6485 9115
rect 6485 9085 6515 9115
rect 6515 9085 6516 9115
rect 6484 9084 6516 9085
rect 6484 9035 6516 9036
rect 6484 9005 6485 9035
rect 6485 9005 6515 9035
rect 6515 9005 6516 9035
rect 6484 9004 6516 9005
rect 6484 8955 6516 8956
rect 6484 8925 6485 8955
rect 6485 8925 6515 8955
rect 6515 8925 6516 8955
rect 6484 8924 6516 8925
rect 6484 8635 6516 8636
rect 6484 8605 6485 8635
rect 6485 8605 6515 8635
rect 6515 8605 6516 8635
rect 6484 8604 6516 8605
rect 6484 8555 6516 8556
rect 6484 8525 6485 8555
rect 6485 8525 6515 8555
rect 6515 8525 6516 8555
rect 6484 8524 6516 8525
rect 6484 8395 6516 8396
rect 6484 8365 6485 8395
rect 6485 8365 6515 8395
rect 6515 8365 6516 8395
rect 6484 8364 6516 8365
rect 6484 8235 6516 8236
rect 6484 8205 6485 8235
rect 6485 8205 6515 8235
rect 6515 8205 6516 8235
rect 6484 8204 6516 8205
rect 6484 8155 6516 8156
rect 6484 8125 6485 8155
rect 6485 8125 6515 8155
rect 6515 8125 6516 8155
rect 6484 8124 6516 8125
rect 6484 8075 6516 8076
rect 6484 8045 6485 8075
rect 6485 8045 6515 8075
rect 6515 8045 6516 8075
rect 6484 8044 6516 8045
rect 6484 7995 6516 7996
rect 6484 7965 6485 7995
rect 6485 7965 6515 7995
rect 6515 7965 6516 7995
rect 6484 7964 6516 7965
rect 6484 7915 6516 7916
rect 6484 7885 6485 7915
rect 6485 7885 6515 7915
rect 6515 7885 6516 7915
rect 6484 7884 6516 7885
rect 6484 7835 6516 7836
rect 6484 7805 6485 7835
rect 6485 7805 6515 7835
rect 6515 7805 6516 7835
rect 6484 7804 6516 7805
rect 6484 7755 6516 7756
rect 6484 7725 6485 7755
rect 6485 7725 6515 7755
rect 6515 7725 6516 7755
rect 6484 7724 6516 7725
rect 6484 7675 6516 7676
rect 6484 7645 6485 7675
rect 6485 7645 6515 7675
rect 6515 7645 6516 7675
rect 6484 7644 6516 7645
rect 6484 7595 6516 7596
rect 6484 7565 6485 7595
rect 6485 7565 6515 7595
rect 6515 7565 6516 7595
rect 6484 7564 6516 7565
rect 6484 7515 6516 7516
rect 6484 7485 6485 7515
rect 6485 7485 6515 7515
rect 6515 7485 6516 7515
rect 6484 7484 6516 7485
rect 6484 7435 6516 7436
rect 6484 7405 6485 7435
rect 6485 7405 6515 7435
rect 6515 7405 6516 7435
rect 6484 7404 6516 7405
rect 6484 7355 6516 7356
rect 6484 7325 6485 7355
rect 6485 7325 6515 7355
rect 6515 7325 6516 7355
rect 6484 7324 6516 7325
rect 6484 7275 6516 7276
rect 6484 7245 6485 7275
rect 6485 7245 6515 7275
rect 6515 7245 6516 7275
rect 6484 7244 6516 7245
rect 6484 7195 6516 7196
rect 6484 7165 6485 7195
rect 6485 7165 6515 7195
rect 6515 7165 6516 7195
rect 6484 7164 6516 7165
rect 6484 7115 6516 7116
rect 6484 7085 6485 7115
rect 6485 7085 6515 7115
rect 6515 7085 6516 7115
rect 6484 7084 6516 7085
rect 6484 7035 6516 7036
rect 6484 7005 6485 7035
rect 6485 7005 6515 7035
rect 6515 7005 6516 7035
rect 6484 7004 6516 7005
rect 6484 6955 6516 6956
rect 6484 6925 6485 6955
rect 6485 6925 6515 6955
rect 6515 6925 6516 6955
rect 6484 6924 6516 6925
rect 6484 6875 6516 6876
rect 6484 6845 6485 6875
rect 6485 6845 6515 6875
rect 6515 6845 6516 6875
rect 6484 6844 6516 6845
rect 6484 6795 6516 6796
rect 6484 6765 6485 6795
rect 6485 6765 6515 6795
rect 6515 6765 6516 6795
rect 6484 6764 6516 6765
rect 6484 6715 6516 6716
rect 6484 6685 6485 6715
rect 6485 6685 6515 6715
rect 6515 6685 6516 6715
rect 6484 6684 6516 6685
rect 6484 6635 6516 6636
rect 6484 6605 6485 6635
rect 6485 6605 6515 6635
rect 6515 6605 6516 6635
rect 6484 6604 6516 6605
rect 6484 6555 6516 6556
rect 6484 6525 6485 6555
rect 6485 6525 6515 6555
rect 6515 6525 6516 6555
rect 6484 6524 6516 6525
rect 6484 6475 6516 6476
rect 6484 6445 6485 6475
rect 6485 6445 6515 6475
rect 6515 6445 6516 6475
rect 6484 6444 6516 6445
rect 6484 6315 6516 6316
rect 6484 6285 6485 6315
rect 6485 6285 6515 6315
rect 6515 6285 6516 6315
rect 6484 6284 6516 6285
rect 6484 6235 6516 6236
rect 6484 6205 6485 6235
rect 6485 6205 6515 6235
rect 6515 6205 6516 6235
rect 6484 6204 6516 6205
rect 6484 6155 6516 6156
rect 6484 6125 6485 6155
rect 6485 6125 6515 6155
rect 6515 6125 6516 6155
rect 6484 6124 6516 6125
rect 6484 5995 6516 5996
rect 6484 5965 6485 5995
rect 6485 5965 6515 5995
rect 6515 5965 6516 5995
rect 6484 5964 6516 5965
rect 6484 5835 6516 5836
rect 6484 5805 6485 5835
rect 6485 5805 6515 5835
rect 6515 5805 6516 5835
rect 6484 5804 6516 5805
rect 6484 5755 6516 5756
rect 6484 5725 6485 5755
rect 6485 5725 6515 5755
rect 6515 5725 6516 5755
rect 6484 5724 6516 5725
rect 6484 5675 6516 5676
rect 6484 5645 6485 5675
rect 6485 5645 6515 5675
rect 6515 5645 6516 5675
rect 6484 5644 6516 5645
rect 6484 5595 6516 5596
rect 6484 5565 6485 5595
rect 6485 5565 6515 5595
rect 6515 5565 6516 5595
rect 6484 5564 6516 5565
rect 6484 5515 6516 5516
rect 6484 5485 6485 5515
rect 6485 5485 6515 5515
rect 6515 5485 6516 5515
rect 6484 5484 6516 5485
rect 6484 5435 6516 5436
rect 6484 5405 6485 5435
rect 6485 5405 6515 5435
rect 6515 5405 6516 5435
rect 6484 5404 6516 5405
rect 6484 5355 6516 5356
rect 6484 5325 6485 5355
rect 6485 5325 6515 5355
rect 6515 5325 6516 5355
rect 6484 5324 6516 5325
rect 6484 5275 6516 5276
rect 6484 5245 6485 5275
rect 6485 5245 6515 5275
rect 6515 5245 6516 5275
rect 6484 5244 6516 5245
rect 6484 5195 6516 5196
rect 6484 5165 6485 5195
rect 6485 5165 6515 5195
rect 6515 5165 6516 5195
rect 6484 5164 6516 5165
rect 6484 5115 6516 5116
rect 6484 5085 6485 5115
rect 6485 5085 6515 5115
rect 6515 5085 6516 5115
rect 6484 5084 6516 5085
rect 6484 5035 6516 5036
rect 6484 5005 6485 5035
rect 6485 5005 6515 5035
rect 6515 5005 6516 5035
rect 6484 5004 6516 5005
rect 6484 4955 6516 4956
rect 6484 4925 6485 4955
rect 6485 4925 6515 4955
rect 6515 4925 6516 4955
rect 6484 4924 6516 4925
rect 6484 4875 6516 4876
rect 6484 4845 6485 4875
rect 6485 4845 6515 4875
rect 6515 4845 6516 4875
rect 6484 4844 6516 4845
rect 6484 4795 6516 4796
rect 6484 4765 6485 4795
rect 6485 4765 6515 4795
rect 6515 4765 6516 4795
rect 6484 4764 6516 4765
rect 6484 4715 6516 4716
rect 6484 4685 6485 4715
rect 6485 4685 6515 4715
rect 6515 4685 6516 4715
rect 6484 4684 6516 4685
rect 6484 4635 6516 4636
rect 6484 4605 6485 4635
rect 6485 4605 6515 4635
rect 6515 4605 6516 4635
rect 6484 4604 6516 4605
rect 6484 4555 6516 4556
rect 6484 4525 6485 4555
rect 6485 4525 6515 4555
rect 6515 4525 6516 4555
rect 6484 4524 6516 4525
rect 6484 4475 6516 4476
rect 6484 4445 6485 4475
rect 6485 4445 6515 4475
rect 6515 4445 6516 4475
rect 6484 4444 6516 4445
rect 6484 4395 6516 4396
rect 6484 4365 6485 4395
rect 6485 4365 6515 4395
rect 6515 4365 6516 4395
rect 6484 4364 6516 4365
rect 6484 4315 6516 4316
rect 6484 4285 6485 4315
rect 6485 4285 6515 4315
rect 6515 4285 6516 4315
rect 6484 4284 6516 4285
rect 6484 4235 6516 4236
rect 6484 4205 6485 4235
rect 6485 4205 6515 4235
rect 6515 4205 6516 4235
rect 6484 4204 6516 4205
rect 6484 4155 6516 4156
rect 6484 4125 6485 4155
rect 6485 4125 6515 4155
rect 6515 4125 6516 4155
rect 6484 4124 6516 4125
rect 6484 4075 6516 4076
rect 6484 4045 6485 4075
rect 6485 4045 6515 4075
rect 6515 4045 6516 4075
rect 6484 4044 6516 4045
rect 6484 3995 6516 3996
rect 6484 3965 6485 3995
rect 6485 3965 6515 3995
rect 6515 3965 6516 3995
rect 6484 3964 6516 3965
rect 6484 3915 6516 3916
rect 6484 3885 6485 3915
rect 6485 3885 6515 3915
rect 6515 3885 6516 3915
rect 6484 3884 6516 3885
rect 6484 3835 6516 3836
rect 6484 3805 6485 3835
rect 6485 3805 6515 3835
rect 6515 3805 6516 3835
rect 6484 3804 6516 3805
rect 6484 3755 6516 3756
rect 6484 3725 6485 3755
rect 6485 3725 6515 3755
rect 6515 3725 6516 3755
rect 6484 3724 6516 3725
rect 6484 3595 6516 3596
rect 6484 3565 6485 3595
rect 6485 3565 6515 3595
rect 6515 3565 6516 3595
rect 6484 3564 6516 3565
rect 6484 3435 6516 3436
rect 6484 3405 6485 3435
rect 6485 3405 6515 3435
rect 6515 3405 6516 3435
rect 6484 3404 6516 3405
rect 6484 3355 6516 3356
rect 6484 3325 6485 3355
rect 6485 3325 6515 3355
rect 6515 3325 6516 3355
rect 6484 3324 6516 3325
rect 6484 3275 6516 3276
rect 6484 3245 6485 3275
rect 6485 3245 6515 3275
rect 6515 3245 6516 3275
rect 6484 3244 6516 3245
rect 6484 3195 6516 3196
rect 6484 3165 6485 3195
rect 6485 3165 6515 3195
rect 6515 3165 6516 3195
rect 6484 3164 6516 3165
rect 6484 3115 6516 3116
rect 6484 3085 6485 3115
rect 6485 3085 6515 3115
rect 6515 3085 6516 3115
rect 6484 3084 6516 3085
rect 6484 3035 6516 3036
rect 6484 3005 6485 3035
rect 6485 3005 6515 3035
rect 6515 3005 6516 3035
rect 6484 3004 6516 3005
rect 6484 2955 6516 2956
rect 6484 2925 6485 2955
rect 6485 2925 6515 2955
rect 6515 2925 6516 2955
rect 6484 2924 6516 2925
rect 6484 2875 6516 2876
rect 6484 2845 6485 2875
rect 6485 2845 6515 2875
rect 6515 2845 6516 2875
rect 6484 2844 6516 2845
rect 6484 2795 6516 2796
rect 6484 2765 6485 2795
rect 6485 2765 6515 2795
rect 6515 2765 6516 2795
rect 6484 2764 6516 2765
rect 6484 2715 6516 2716
rect 6484 2685 6485 2715
rect 6485 2685 6515 2715
rect 6515 2685 6516 2715
rect 6484 2684 6516 2685
rect 6484 2635 6516 2636
rect 6484 2605 6485 2635
rect 6485 2605 6515 2635
rect 6515 2605 6516 2635
rect 6484 2604 6516 2605
rect 6484 2555 6516 2556
rect 6484 2525 6485 2555
rect 6485 2525 6515 2555
rect 6515 2525 6516 2555
rect 6484 2524 6516 2525
rect 6484 2475 6516 2476
rect 6484 2445 6485 2475
rect 6485 2445 6515 2475
rect 6515 2445 6516 2475
rect 6484 2444 6516 2445
rect 6484 2395 6516 2396
rect 6484 2365 6485 2395
rect 6485 2365 6515 2395
rect 6515 2365 6516 2395
rect 6484 2364 6516 2365
rect 6484 2315 6516 2316
rect 6484 2285 6485 2315
rect 6485 2285 6515 2315
rect 6515 2285 6516 2315
rect 6484 2284 6516 2285
rect 6484 2235 6516 2236
rect 6484 2205 6485 2235
rect 6485 2205 6515 2235
rect 6515 2205 6516 2235
rect 6484 2204 6516 2205
rect 6484 2155 6516 2156
rect 6484 2125 6485 2155
rect 6485 2125 6515 2155
rect 6515 2125 6516 2155
rect 6484 2124 6516 2125
rect 6484 2075 6516 2076
rect 6484 2045 6485 2075
rect 6485 2045 6515 2075
rect 6515 2045 6516 2075
rect 6484 2044 6516 2045
rect 6484 1995 6516 1996
rect 6484 1965 6485 1995
rect 6485 1965 6515 1995
rect 6515 1965 6516 1995
rect 6484 1964 6516 1965
rect 6484 1915 6516 1916
rect 6484 1885 6485 1915
rect 6485 1885 6515 1915
rect 6515 1885 6516 1915
rect 6484 1884 6516 1885
rect 6484 1835 6516 1836
rect 6484 1805 6485 1835
rect 6485 1805 6515 1835
rect 6515 1805 6516 1835
rect 6484 1804 6516 1805
rect 6484 1755 6516 1756
rect 6484 1725 6485 1755
rect 6485 1725 6515 1755
rect 6515 1725 6516 1755
rect 6484 1724 6516 1725
rect 6484 1675 6516 1676
rect 6484 1645 6485 1675
rect 6485 1645 6515 1675
rect 6515 1645 6516 1675
rect 6484 1644 6516 1645
rect 6484 1595 6516 1596
rect 6484 1565 6485 1595
rect 6485 1565 6515 1595
rect 6515 1565 6516 1595
rect 6484 1564 6516 1565
rect 6484 1515 6516 1516
rect 6484 1485 6485 1515
rect 6485 1485 6515 1515
rect 6515 1485 6516 1515
rect 6484 1484 6516 1485
rect 6484 1435 6516 1436
rect 6484 1405 6485 1435
rect 6485 1405 6515 1435
rect 6515 1405 6516 1435
rect 6484 1404 6516 1405
rect 6484 1355 6516 1356
rect 6484 1325 6485 1355
rect 6485 1325 6515 1355
rect 6515 1325 6516 1355
rect 6484 1324 6516 1325
rect 6484 1275 6516 1276
rect 6484 1245 6485 1275
rect 6485 1245 6515 1275
rect 6515 1245 6516 1275
rect 6484 1244 6516 1245
rect 6484 1195 6516 1196
rect 6484 1165 6485 1195
rect 6485 1165 6515 1195
rect 6515 1165 6516 1195
rect 6484 1164 6516 1165
rect 6484 1115 6516 1116
rect 6484 1085 6485 1115
rect 6485 1085 6515 1115
rect 6515 1085 6516 1115
rect 6484 1084 6516 1085
rect 6484 1035 6516 1036
rect 6484 1005 6485 1035
rect 6485 1005 6515 1035
rect 6515 1005 6516 1035
rect 6484 1004 6516 1005
rect 6484 955 6516 956
rect 6484 925 6485 955
rect 6485 925 6515 955
rect 6515 925 6516 955
rect 6484 924 6516 925
rect 6484 875 6516 876
rect 6484 845 6485 875
rect 6485 845 6515 875
rect 6515 845 6516 875
rect 6484 844 6516 845
rect 6484 795 6516 796
rect 6484 765 6485 795
rect 6485 765 6515 795
rect 6515 765 6516 795
rect 6484 764 6516 765
rect 6484 715 6516 716
rect 6484 685 6485 715
rect 6485 685 6515 715
rect 6515 685 6516 715
rect 6484 684 6516 685
rect 6484 595 6516 596
rect 6484 565 6485 595
rect 6485 565 6515 595
rect 6515 565 6516 595
rect 6484 564 6516 565
rect 6484 515 6516 516
rect 6484 485 6485 515
rect 6485 485 6515 515
rect 6515 485 6516 515
rect 6484 484 6516 485
rect 6484 435 6516 436
rect 6484 405 6485 435
rect 6485 405 6515 435
rect 6515 405 6516 435
rect 6484 404 6516 405
rect 6484 355 6516 356
rect 6484 325 6485 355
rect 6485 325 6515 355
rect 6515 325 6516 355
rect 6484 324 6516 325
rect 6484 275 6516 276
rect 6484 245 6485 275
rect 6485 245 6515 275
rect 6515 245 6516 275
rect 6484 244 6516 245
rect 6484 195 6516 196
rect 6484 165 6485 195
rect 6485 165 6515 195
rect 6515 165 6516 195
rect 6484 164 6516 165
rect 6484 115 6516 116
rect 6484 85 6485 115
rect 6485 85 6515 115
rect 6515 85 6516 115
rect 6484 84 6516 85
rect 6484 35 6516 36
rect 6484 5 6485 35
rect 6485 5 6515 35
rect 6515 5 6516 35
rect 6484 4 6516 5
rect 6804 16644 6836 16836
rect 6644 16595 6676 16596
rect 6644 16565 6645 16595
rect 6645 16565 6675 16595
rect 6675 16565 6676 16595
rect 6644 16564 6676 16565
rect 6644 16515 6676 16516
rect 6644 16485 6645 16515
rect 6645 16485 6675 16515
rect 6675 16485 6676 16515
rect 6644 16484 6676 16485
rect 6644 16435 6676 16436
rect 6644 16405 6645 16435
rect 6645 16405 6675 16435
rect 6675 16405 6676 16435
rect 6644 16404 6676 16405
rect 6644 16355 6676 16356
rect 6644 16325 6645 16355
rect 6645 16325 6675 16355
rect 6675 16325 6676 16355
rect 6644 16324 6676 16325
rect 6644 16275 6676 16276
rect 6644 16245 6645 16275
rect 6645 16245 6675 16275
rect 6675 16245 6676 16275
rect 6644 16244 6676 16245
rect 6644 16195 6676 16196
rect 6644 16165 6645 16195
rect 6645 16165 6675 16195
rect 6675 16165 6676 16195
rect 6644 16164 6676 16165
rect 6644 16115 6676 16116
rect 6644 16085 6645 16115
rect 6645 16085 6675 16115
rect 6675 16085 6676 16115
rect 6644 16084 6676 16085
rect 6644 16035 6676 16036
rect 6644 16005 6645 16035
rect 6645 16005 6675 16035
rect 6675 16005 6676 16035
rect 6644 16004 6676 16005
rect 6644 15955 6676 15956
rect 6644 15925 6645 15955
rect 6645 15925 6675 15955
rect 6675 15925 6676 15955
rect 6644 15924 6676 15925
rect 6644 15435 6676 15436
rect 6644 15405 6645 15435
rect 6645 15405 6675 15435
rect 6675 15405 6676 15435
rect 6644 15404 6676 15405
rect 6644 15355 6676 15356
rect 6644 15325 6645 15355
rect 6645 15325 6675 15355
rect 6675 15325 6676 15355
rect 6644 15324 6676 15325
rect 6644 15275 6676 15276
rect 6644 15245 6645 15275
rect 6645 15245 6675 15275
rect 6675 15245 6676 15275
rect 6644 15244 6676 15245
rect 6644 15195 6676 15196
rect 6644 15165 6645 15195
rect 6645 15165 6675 15195
rect 6675 15165 6676 15195
rect 6644 15164 6676 15165
rect 6644 15115 6676 15116
rect 6644 15085 6645 15115
rect 6645 15085 6675 15115
rect 6675 15085 6676 15115
rect 6644 15084 6676 15085
rect 6644 15035 6676 15036
rect 6644 15005 6645 15035
rect 6645 15005 6675 15035
rect 6675 15005 6676 15035
rect 6644 15004 6676 15005
rect 6644 14955 6676 14956
rect 6644 14925 6645 14955
rect 6645 14925 6675 14955
rect 6675 14925 6676 14955
rect 6644 14924 6676 14925
rect 6644 14875 6676 14876
rect 6644 14845 6645 14875
rect 6645 14845 6675 14875
rect 6675 14845 6676 14875
rect 6644 14844 6676 14845
rect 6644 14795 6676 14796
rect 6644 14765 6645 14795
rect 6645 14765 6675 14795
rect 6675 14765 6676 14795
rect 6644 14764 6676 14765
rect 6644 14715 6676 14716
rect 6644 14685 6645 14715
rect 6645 14685 6675 14715
rect 6675 14685 6676 14715
rect 6644 14684 6676 14685
rect 6644 14635 6676 14636
rect 6644 14605 6645 14635
rect 6645 14605 6675 14635
rect 6675 14605 6676 14635
rect 6644 14604 6676 14605
rect 6644 14555 6676 14556
rect 6644 14525 6645 14555
rect 6645 14525 6675 14555
rect 6675 14525 6676 14555
rect 6644 14524 6676 14525
rect 6644 14475 6676 14476
rect 6644 14445 6645 14475
rect 6645 14445 6675 14475
rect 6675 14445 6676 14475
rect 6644 14444 6676 14445
rect 6644 13995 6676 13996
rect 6644 13965 6645 13995
rect 6645 13965 6675 13995
rect 6675 13965 6676 13995
rect 6644 13964 6676 13965
rect 6644 13875 6676 13876
rect 6644 13845 6645 13875
rect 6645 13845 6675 13875
rect 6675 13845 6676 13875
rect 6644 13844 6676 13845
rect 6644 13795 6676 13796
rect 6644 13765 6645 13795
rect 6645 13765 6675 13795
rect 6675 13765 6676 13795
rect 6644 13764 6676 13765
rect 6644 13715 6676 13716
rect 6644 13685 6645 13715
rect 6645 13685 6675 13715
rect 6675 13685 6676 13715
rect 6644 13684 6676 13685
rect 6644 13635 6676 13636
rect 6644 13605 6645 13635
rect 6645 13605 6675 13635
rect 6675 13605 6676 13635
rect 6644 13604 6676 13605
rect 6644 13555 6676 13556
rect 6644 13525 6645 13555
rect 6645 13525 6675 13555
rect 6675 13525 6676 13555
rect 6644 13524 6676 13525
rect 6644 13475 6676 13476
rect 6644 13445 6645 13475
rect 6645 13445 6675 13475
rect 6675 13445 6676 13475
rect 6644 13444 6676 13445
rect 6644 13395 6676 13396
rect 6644 13365 6645 13395
rect 6645 13365 6675 13395
rect 6675 13365 6676 13395
rect 6644 13364 6676 13365
rect 6644 13315 6676 13316
rect 6644 13285 6645 13315
rect 6645 13285 6675 13315
rect 6675 13285 6676 13315
rect 6644 13284 6676 13285
rect 6644 13235 6676 13236
rect 6644 13205 6645 13235
rect 6645 13205 6675 13235
rect 6675 13205 6676 13235
rect 6644 13204 6676 13205
rect 6644 13155 6676 13156
rect 6644 13125 6645 13155
rect 6645 13125 6675 13155
rect 6675 13125 6676 13155
rect 6644 13124 6676 13125
rect 6644 13075 6676 13076
rect 6644 13045 6645 13075
rect 6645 13045 6675 13075
rect 6675 13045 6676 13075
rect 6644 13044 6676 13045
rect 6644 12995 6676 12996
rect 6644 12965 6645 12995
rect 6645 12965 6675 12995
rect 6675 12965 6676 12995
rect 6644 12964 6676 12965
rect 6644 12515 6676 12516
rect 6644 12485 6645 12515
rect 6645 12485 6675 12515
rect 6675 12485 6676 12515
rect 6644 12484 6676 12485
rect 6644 12435 6676 12436
rect 6644 12405 6645 12435
rect 6645 12405 6675 12435
rect 6675 12405 6676 12435
rect 6644 12404 6676 12405
rect 6644 12315 6676 12316
rect 6644 12285 6645 12315
rect 6645 12285 6675 12315
rect 6675 12285 6676 12315
rect 6644 12284 6676 12285
rect 6644 12235 6676 12236
rect 6644 12205 6645 12235
rect 6645 12205 6675 12235
rect 6675 12205 6676 12235
rect 6644 12204 6676 12205
rect 6644 12155 6676 12156
rect 6644 12125 6645 12155
rect 6645 12125 6675 12155
rect 6675 12125 6676 12155
rect 6644 12124 6676 12125
rect 6644 12075 6676 12076
rect 6644 12045 6645 12075
rect 6645 12045 6675 12075
rect 6675 12045 6676 12075
rect 6644 12044 6676 12045
rect 6644 11995 6676 11996
rect 6644 11965 6645 11995
rect 6645 11965 6675 11995
rect 6675 11965 6676 11995
rect 6644 11964 6676 11965
rect 6644 11915 6676 11916
rect 6644 11885 6645 11915
rect 6645 11885 6675 11915
rect 6675 11885 6676 11915
rect 6644 11884 6676 11885
rect 6644 11835 6676 11836
rect 6644 11805 6645 11835
rect 6645 11805 6675 11835
rect 6675 11805 6676 11835
rect 6644 11804 6676 11805
rect 6644 11755 6676 11756
rect 6644 11725 6645 11755
rect 6645 11725 6675 11755
rect 6675 11725 6676 11755
rect 6644 11724 6676 11725
rect 6644 11675 6676 11676
rect 6644 11645 6645 11675
rect 6645 11645 6675 11675
rect 6675 11645 6676 11675
rect 6644 11644 6676 11645
rect 6644 11595 6676 11596
rect 6644 11565 6645 11595
rect 6645 11565 6675 11595
rect 6675 11565 6676 11595
rect 6644 11564 6676 11565
rect 6644 11515 6676 11516
rect 6644 11485 6645 11515
rect 6645 11485 6675 11515
rect 6675 11485 6676 11515
rect 6644 11484 6676 11485
rect 6644 11435 6676 11436
rect 6644 11405 6645 11435
rect 6645 11405 6675 11435
rect 6675 11405 6676 11435
rect 6644 11404 6676 11405
rect 6644 11355 6676 11356
rect 6644 11325 6645 11355
rect 6645 11325 6675 11355
rect 6675 11325 6676 11355
rect 6644 11324 6676 11325
rect 6644 11195 6676 11196
rect 6644 11165 6645 11195
rect 6645 11165 6675 11195
rect 6675 11165 6676 11195
rect 6644 11164 6676 11165
rect 6644 11115 6676 11116
rect 6644 11085 6645 11115
rect 6645 11085 6675 11115
rect 6675 11085 6676 11115
rect 6644 11084 6676 11085
rect 6644 11035 6676 11036
rect 6644 11005 6645 11035
rect 6645 11005 6675 11035
rect 6675 11005 6676 11035
rect 6644 11004 6676 11005
rect 6644 10875 6676 10876
rect 6644 10845 6645 10875
rect 6645 10845 6675 10875
rect 6675 10845 6676 10875
rect 6644 10844 6676 10845
rect 6644 10715 6676 10716
rect 6644 10685 6645 10715
rect 6645 10685 6675 10715
rect 6675 10685 6676 10715
rect 6644 10684 6676 10685
rect 6644 10635 6676 10636
rect 6644 10605 6645 10635
rect 6645 10605 6675 10635
rect 6675 10605 6676 10635
rect 6644 10604 6676 10605
rect 6644 10475 6676 10476
rect 6644 10445 6645 10475
rect 6645 10445 6675 10475
rect 6675 10445 6676 10475
rect 6644 10444 6676 10445
rect 6644 10315 6676 10316
rect 6644 10285 6645 10315
rect 6645 10285 6675 10315
rect 6675 10285 6676 10315
rect 6644 10284 6676 10285
rect 6644 10235 6676 10236
rect 6644 10205 6645 10235
rect 6645 10205 6675 10235
rect 6675 10205 6676 10235
rect 6644 10204 6676 10205
rect 6644 10155 6676 10156
rect 6644 10125 6645 10155
rect 6645 10125 6675 10155
rect 6675 10125 6676 10155
rect 6644 10124 6676 10125
rect 6644 10075 6676 10076
rect 6644 10045 6645 10075
rect 6645 10045 6675 10075
rect 6675 10045 6676 10075
rect 6644 10044 6676 10045
rect 6644 9995 6676 9996
rect 6644 9965 6645 9995
rect 6645 9965 6675 9995
rect 6675 9965 6676 9995
rect 6644 9964 6676 9965
rect 6644 9915 6676 9916
rect 6644 9885 6645 9915
rect 6645 9885 6675 9915
rect 6675 9885 6676 9915
rect 6644 9884 6676 9885
rect 6644 9835 6676 9836
rect 6644 9805 6645 9835
rect 6645 9805 6675 9835
rect 6675 9805 6676 9835
rect 6644 9804 6676 9805
rect 6644 9755 6676 9756
rect 6644 9725 6645 9755
rect 6645 9725 6675 9755
rect 6675 9725 6676 9755
rect 6644 9724 6676 9725
rect 6644 9675 6676 9676
rect 6644 9645 6645 9675
rect 6645 9645 6675 9675
rect 6675 9645 6676 9675
rect 6644 9644 6676 9645
rect 6644 9595 6676 9596
rect 6644 9565 6645 9595
rect 6645 9565 6675 9595
rect 6675 9565 6676 9595
rect 6644 9564 6676 9565
rect 6644 9515 6676 9516
rect 6644 9485 6645 9515
rect 6645 9485 6675 9515
rect 6675 9485 6676 9515
rect 6644 9484 6676 9485
rect 6644 9435 6676 9436
rect 6644 9405 6645 9435
rect 6645 9405 6675 9435
rect 6675 9405 6676 9435
rect 6644 9404 6676 9405
rect 6644 9355 6676 9356
rect 6644 9325 6645 9355
rect 6645 9325 6675 9355
rect 6675 9325 6676 9355
rect 6644 9324 6676 9325
rect 6644 9275 6676 9276
rect 6644 9245 6645 9275
rect 6645 9245 6675 9275
rect 6675 9245 6676 9275
rect 6644 9244 6676 9245
rect 6644 9115 6676 9116
rect 6644 9085 6645 9115
rect 6645 9085 6675 9115
rect 6675 9085 6676 9115
rect 6644 9084 6676 9085
rect 6644 9035 6676 9036
rect 6644 9005 6645 9035
rect 6645 9005 6675 9035
rect 6675 9005 6676 9035
rect 6644 9004 6676 9005
rect 6644 8955 6676 8956
rect 6644 8925 6645 8955
rect 6645 8925 6675 8955
rect 6675 8925 6676 8955
rect 6644 8924 6676 8925
rect 6644 8635 6676 8636
rect 6644 8605 6645 8635
rect 6645 8605 6675 8635
rect 6675 8605 6676 8635
rect 6644 8604 6676 8605
rect 6644 8555 6676 8556
rect 6644 8525 6645 8555
rect 6645 8525 6675 8555
rect 6675 8525 6676 8555
rect 6644 8524 6676 8525
rect 6644 8395 6676 8396
rect 6644 8365 6645 8395
rect 6645 8365 6675 8395
rect 6675 8365 6676 8395
rect 6644 8364 6676 8365
rect 6644 8235 6676 8236
rect 6644 8205 6645 8235
rect 6645 8205 6675 8235
rect 6675 8205 6676 8235
rect 6644 8204 6676 8205
rect 6644 8155 6676 8156
rect 6644 8125 6645 8155
rect 6645 8125 6675 8155
rect 6675 8125 6676 8155
rect 6644 8124 6676 8125
rect 6644 8075 6676 8076
rect 6644 8045 6645 8075
rect 6645 8045 6675 8075
rect 6675 8045 6676 8075
rect 6644 8044 6676 8045
rect 6644 7995 6676 7996
rect 6644 7965 6645 7995
rect 6645 7965 6675 7995
rect 6675 7965 6676 7995
rect 6644 7964 6676 7965
rect 6644 7915 6676 7916
rect 6644 7885 6645 7915
rect 6645 7885 6675 7915
rect 6675 7885 6676 7915
rect 6644 7884 6676 7885
rect 6644 7835 6676 7836
rect 6644 7805 6645 7835
rect 6645 7805 6675 7835
rect 6675 7805 6676 7835
rect 6644 7804 6676 7805
rect 6644 7755 6676 7756
rect 6644 7725 6645 7755
rect 6645 7725 6675 7755
rect 6675 7725 6676 7755
rect 6644 7724 6676 7725
rect 6644 7675 6676 7676
rect 6644 7645 6645 7675
rect 6645 7645 6675 7675
rect 6675 7645 6676 7675
rect 6644 7644 6676 7645
rect 6644 7595 6676 7596
rect 6644 7565 6645 7595
rect 6645 7565 6675 7595
rect 6675 7565 6676 7595
rect 6644 7564 6676 7565
rect 6644 7515 6676 7516
rect 6644 7485 6645 7515
rect 6645 7485 6675 7515
rect 6675 7485 6676 7515
rect 6644 7484 6676 7485
rect 6644 7435 6676 7436
rect 6644 7405 6645 7435
rect 6645 7405 6675 7435
rect 6675 7405 6676 7435
rect 6644 7404 6676 7405
rect 6644 7355 6676 7356
rect 6644 7325 6645 7355
rect 6645 7325 6675 7355
rect 6675 7325 6676 7355
rect 6644 7324 6676 7325
rect 6644 7275 6676 7276
rect 6644 7245 6645 7275
rect 6645 7245 6675 7275
rect 6675 7245 6676 7275
rect 6644 7244 6676 7245
rect 6644 7195 6676 7196
rect 6644 7165 6645 7195
rect 6645 7165 6675 7195
rect 6675 7165 6676 7195
rect 6644 7164 6676 7165
rect 6644 7115 6676 7116
rect 6644 7085 6645 7115
rect 6645 7085 6675 7115
rect 6675 7085 6676 7115
rect 6644 7084 6676 7085
rect 6644 7035 6676 7036
rect 6644 7005 6645 7035
rect 6645 7005 6675 7035
rect 6675 7005 6676 7035
rect 6644 7004 6676 7005
rect 6644 6955 6676 6956
rect 6644 6925 6645 6955
rect 6645 6925 6675 6955
rect 6675 6925 6676 6955
rect 6644 6924 6676 6925
rect 6644 6875 6676 6876
rect 6644 6845 6645 6875
rect 6645 6845 6675 6875
rect 6675 6845 6676 6875
rect 6644 6844 6676 6845
rect 6644 6795 6676 6796
rect 6644 6765 6645 6795
rect 6645 6765 6675 6795
rect 6675 6765 6676 6795
rect 6644 6764 6676 6765
rect 6644 6715 6676 6716
rect 6644 6685 6645 6715
rect 6645 6685 6675 6715
rect 6675 6685 6676 6715
rect 6644 6684 6676 6685
rect 6644 6635 6676 6636
rect 6644 6605 6645 6635
rect 6645 6605 6675 6635
rect 6675 6605 6676 6635
rect 6644 6604 6676 6605
rect 6644 6555 6676 6556
rect 6644 6525 6645 6555
rect 6645 6525 6675 6555
rect 6675 6525 6676 6555
rect 6644 6524 6676 6525
rect 6644 6475 6676 6476
rect 6644 6445 6645 6475
rect 6645 6445 6675 6475
rect 6675 6445 6676 6475
rect 6644 6444 6676 6445
rect 6644 6395 6676 6396
rect 6644 6365 6645 6395
rect 6645 6365 6675 6395
rect 6675 6365 6676 6395
rect 6644 6364 6676 6365
rect 6644 6315 6676 6316
rect 6644 6285 6645 6315
rect 6645 6285 6675 6315
rect 6675 6285 6676 6315
rect 6644 6284 6676 6285
rect 6644 6235 6676 6236
rect 6644 6205 6645 6235
rect 6645 6205 6675 6235
rect 6675 6205 6676 6235
rect 6644 6204 6676 6205
rect 6644 6155 6676 6156
rect 6644 6125 6645 6155
rect 6645 6125 6675 6155
rect 6675 6125 6676 6155
rect 6644 6124 6676 6125
rect 6644 5995 6676 5996
rect 6644 5965 6645 5995
rect 6645 5965 6675 5995
rect 6675 5965 6676 5995
rect 6644 5964 6676 5965
rect 6644 5835 6676 5836
rect 6644 5805 6645 5835
rect 6645 5805 6675 5835
rect 6675 5805 6676 5835
rect 6644 5804 6676 5805
rect 6644 5755 6676 5756
rect 6644 5725 6645 5755
rect 6645 5725 6675 5755
rect 6675 5725 6676 5755
rect 6644 5724 6676 5725
rect 6644 5675 6676 5676
rect 6644 5645 6645 5675
rect 6645 5645 6675 5675
rect 6675 5645 6676 5675
rect 6644 5644 6676 5645
rect 6644 5595 6676 5596
rect 6644 5565 6645 5595
rect 6645 5565 6675 5595
rect 6675 5565 6676 5595
rect 6644 5564 6676 5565
rect 6644 5515 6676 5516
rect 6644 5485 6645 5515
rect 6645 5485 6675 5515
rect 6675 5485 6676 5515
rect 6644 5484 6676 5485
rect 6644 5435 6676 5436
rect 6644 5405 6645 5435
rect 6645 5405 6675 5435
rect 6675 5405 6676 5435
rect 6644 5404 6676 5405
rect 6644 5355 6676 5356
rect 6644 5325 6645 5355
rect 6645 5325 6675 5355
rect 6675 5325 6676 5355
rect 6644 5324 6676 5325
rect 6644 5275 6676 5276
rect 6644 5245 6645 5275
rect 6645 5245 6675 5275
rect 6675 5245 6676 5275
rect 6644 5244 6676 5245
rect 6644 5195 6676 5196
rect 6644 5165 6645 5195
rect 6645 5165 6675 5195
rect 6675 5165 6676 5195
rect 6644 5164 6676 5165
rect 6644 5115 6676 5116
rect 6644 5085 6645 5115
rect 6645 5085 6675 5115
rect 6675 5085 6676 5115
rect 6644 5084 6676 5085
rect 6644 5035 6676 5036
rect 6644 5005 6645 5035
rect 6645 5005 6675 5035
rect 6675 5005 6676 5035
rect 6644 5004 6676 5005
rect 6644 4955 6676 4956
rect 6644 4925 6645 4955
rect 6645 4925 6675 4955
rect 6675 4925 6676 4955
rect 6644 4924 6676 4925
rect 6644 4875 6676 4876
rect 6644 4845 6645 4875
rect 6645 4845 6675 4875
rect 6675 4845 6676 4875
rect 6644 4844 6676 4845
rect 6644 4795 6676 4796
rect 6644 4765 6645 4795
rect 6645 4765 6675 4795
rect 6675 4765 6676 4795
rect 6644 4764 6676 4765
rect 6644 4715 6676 4716
rect 6644 4685 6645 4715
rect 6645 4685 6675 4715
rect 6675 4685 6676 4715
rect 6644 4684 6676 4685
rect 6644 4635 6676 4636
rect 6644 4605 6645 4635
rect 6645 4605 6675 4635
rect 6675 4605 6676 4635
rect 6644 4604 6676 4605
rect 6644 4555 6676 4556
rect 6644 4525 6645 4555
rect 6645 4525 6675 4555
rect 6675 4525 6676 4555
rect 6644 4524 6676 4525
rect 6644 4475 6676 4476
rect 6644 4445 6645 4475
rect 6645 4445 6675 4475
rect 6675 4445 6676 4475
rect 6644 4444 6676 4445
rect 6644 4395 6676 4396
rect 6644 4365 6645 4395
rect 6645 4365 6675 4395
rect 6675 4365 6676 4395
rect 6644 4364 6676 4365
rect 6644 4315 6676 4316
rect 6644 4285 6645 4315
rect 6645 4285 6675 4315
rect 6675 4285 6676 4315
rect 6644 4284 6676 4285
rect 6644 4235 6676 4236
rect 6644 4205 6645 4235
rect 6645 4205 6675 4235
rect 6675 4205 6676 4235
rect 6644 4204 6676 4205
rect 6644 4155 6676 4156
rect 6644 4125 6645 4155
rect 6645 4125 6675 4155
rect 6675 4125 6676 4155
rect 6644 4124 6676 4125
rect 6644 4075 6676 4076
rect 6644 4045 6645 4075
rect 6645 4045 6675 4075
rect 6675 4045 6676 4075
rect 6644 4044 6676 4045
rect 6644 3995 6676 3996
rect 6644 3965 6645 3995
rect 6645 3965 6675 3995
rect 6675 3965 6676 3995
rect 6644 3964 6676 3965
rect 6644 3915 6676 3916
rect 6644 3885 6645 3915
rect 6645 3885 6675 3915
rect 6675 3885 6676 3915
rect 6644 3884 6676 3885
rect 6644 3835 6676 3836
rect 6644 3805 6645 3835
rect 6645 3805 6675 3835
rect 6675 3805 6676 3835
rect 6644 3804 6676 3805
rect 6644 3755 6676 3756
rect 6644 3725 6645 3755
rect 6645 3725 6675 3755
rect 6675 3725 6676 3755
rect 6644 3724 6676 3725
rect 6644 3595 6676 3596
rect 6644 3565 6645 3595
rect 6645 3565 6675 3595
rect 6675 3565 6676 3595
rect 6644 3564 6676 3565
rect 6644 3435 6676 3436
rect 6644 3405 6645 3435
rect 6645 3405 6675 3435
rect 6675 3405 6676 3435
rect 6644 3404 6676 3405
rect 6644 3355 6676 3356
rect 6644 3325 6645 3355
rect 6645 3325 6675 3355
rect 6675 3325 6676 3355
rect 6644 3324 6676 3325
rect 6644 3275 6676 3276
rect 6644 3245 6645 3275
rect 6645 3245 6675 3275
rect 6675 3245 6676 3275
rect 6644 3244 6676 3245
rect 6644 3195 6676 3196
rect 6644 3165 6645 3195
rect 6645 3165 6675 3195
rect 6675 3165 6676 3195
rect 6644 3164 6676 3165
rect 6644 3115 6676 3116
rect 6644 3085 6645 3115
rect 6645 3085 6675 3115
rect 6675 3085 6676 3115
rect 6644 3084 6676 3085
rect 6644 3035 6676 3036
rect 6644 3005 6645 3035
rect 6645 3005 6675 3035
rect 6675 3005 6676 3035
rect 6644 3004 6676 3005
rect 6644 2955 6676 2956
rect 6644 2925 6645 2955
rect 6645 2925 6675 2955
rect 6675 2925 6676 2955
rect 6644 2924 6676 2925
rect 6644 2875 6676 2876
rect 6644 2845 6645 2875
rect 6645 2845 6675 2875
rect 6675 2845 6676 2875
rect 6644 2844 6676 2845
rect 6644 2795 6676 2796
rect 6644 2765 6645 2795
rect 6645 2765 6675 2795
rect 6675 2765 6676 2795
rect 6644 2764 6676 2765
rect 6644 2715 6676 2716
rect 6644 2685 6645 2715
rect 6645 2685 6675 2715
rect 6675 2685 6676 2715
rect 6644 2684 6676 2685
rect 6644 2635 6676 2636
rect 6644 2605 6645 2635
rect 6645 2605 6675 2635
rect 6675 2605 6676 2635
rect 6644 2604 6676 2605
rect 6644 2555 6676 2556
rect 6644 2525 6645 2555
rect 6645 2525 6675 2555
rect 6675 2525 6676 2555
rect 6644 2524 6676 2525
rect 6644 2475 6676 2476
rect 6644 2445 6645 2475
rect 6645 2445 6675 2475
rect 6675 2445 6676 2475
rect 6644 2444 6676 2445
rect 6644 2395 6676 2396
rect 6644 2365 6645 2395
rect 6645 2365 6675 2395
rect 6675 2365 6676 2395
rect 6644 2364 6676 2365
rect 6644 2315 6676 2316
rect 6644 2285 6645 2315
rect 6645 2285 6675 2315
rect 6675 2285 6676 2315
rect 6644 2284 6676 2285
rect 6644 2235 6676 2236
rect 6644 2205 6645 2235
rect 6645 2205 6675 2235
rect 6675 2205 6676 2235
rect 6644 2204 6676 2205
rect 6644 2155 6676 2156
rect 6644 2125 6645 2155
rect 6645 2125 6675 2155
rect 6675 2125 6676 2155
rect 6644 2124 6676 2125
rect 6644 2075 6676 2076
rect 6644 2045 6645 2075
rect 6645 2045 6675 2075
rect 6675 2045 6676 2075
rect 6644 2044 6676 2045
rect 6644 1995 6676 1996
rect 6644 1965 6645 1995
rect 6645 1965 6675 1995
rect 6675 1965 6676 1995
rect 6644 1964 6676 1965
rect 6644 1915 6676 1916
rect 6644 1885 6645 1915
rect 6645 1885 6675 1915
rect 6675 1885 6676 1915
rect 6644 1884 6676 1885
rect 6644 1835 6676 1836
rect 6644 1805 6645 1835
rect 6645 1805 6675 1835
rect 6675 1805 6676 1835
rect 6644 1804 6676 1805
rect 6644 1755 6676 1756
rect 6644 1725 6645 1755
rect 6645 1725 6675 1755
rect 6675 1725 6676 1755
rect 6644 1724 6676 1725
rect 6644 1675 6676 1676
rect 6644 1645 6645 1675
rect 6645 1645 6675 1675
rect 6675 1645 6676 1675
rect 6644 1644 6676 1645
rect 6644 1595 6676 1596
rect 6644 1565 6645 1595
rect 6645 1565 6675 1595
rect 6675 1565 6676 1595
rect 6644 1564 6676 1565
rect 6644 1515 6676 1516
rect 6644 1485 6645 1515
rect 6645 1485 6675 1515
rect 6675 1485 6676 1515
rect 6644 1484 6676 1485
rect 6644 1435 6676 1436
rect 6644 1405 6645 1435
rect 6645 1405 6675 1435
rect 6675 1405 6676 1435
rect 6644 1404 6676 1405
rect 6644 1355 6676 1356
rect 6644 1325 6645 1355
rect 6645 1325 6675 1355
rect 6675 1325 6676 1355
rect 6644 1324 6676 1325
rect 6644 1275 6676 1276
rect 6644 1245 6645 1275
rect 6645 1245 6675 1275
rect 6675 1245 6676 1275
rect 6644 1244 6676 1245
rect 6644 1195 6676 1196
rect 6644 1165 6645 1195
rect 6645 1165 6675 1195
rect 6675 1165 6676 1195
rect 6644 1164 6676 1165
rect 6644 1115 6676 1116
rect 6644 1085 6645 1115
rect 6645 1085 6675 1115
rect 6675 1085 6676 1115
rect 6644 1084 6676 1085
rect 6644 1035 6676 1036
rect 6644 1005 6645 1035
rect 6645 1005 6675 1035
rect 6675 1005 6676 1035
rect 6644 1004 6676 1005
rect 6644 955 6676 956
rect 6644 925 6645 955
rect 6645 925 6675 955
rect 6675 925 6676 955
rect 6644 924 6676 925
rect 6644 875 6676 876
rect 6644 845 6645 875
rect 6645 845 6675 875
rect 6675 845 6676 875
rect 6644 844 6676 845
rect 6644 795 6676 796
rect 6644 765 6645 795
rect 6645 765 6675 795
rect 6675 765 6676 795
rect 6644 764 6676 765
rect 6644 715 6676 716
rect 6644 685 6645 715
rect 6645 685 6675 715
rect 6675 685 6676 715
rect 6644 684 6676 685
rect 6644 595 6676 596
rect 6644 565 6645 595
rect 6645 565 6675 595
rect 6675 565 6676 595
rect 6644 564 6676 565
rect 6644 515 6676 516
rect 6644 485 6645 515
rect 6645 485 6675 515
rect 6675 485 6676 515
rect 6644 484 6676 485
rect 6644 435 6676 436
rect 6644 405 6645 435
rect 6645 405 6675 435
rect 6675 405 6676 435
rect 6644 404 6676 405
rect 6644 355 6676 356
rect 6644 325 6645 355
rect 6645 325 6675 355
rect 6675 325 6676 355
rect 6644 324 6676 325
rect 6644 275 6676 276
rect 6644 245 6645 275
rect 6645 245 6675 275
rect 6675 245 6676 275
rect 6644 244 6676 245
rect 6644 195 6676 196
rect 6644 165 6645 195
rect 6645 165 6675 195
rect 6675 165 6676 195
rect 6644 164 6676 165
rect 6644 115 6676 116
rect 6644 85 6645 115
rect 6645 85 6675 115
rect 6675 85 6676 115
rect 6644 84 6676 85
rect 6644 35 6676 36
rect 6644 5 6645 35
rect 6645 5 6675 35
rect 6675 5 6676 35
rect 6644 4 6676 5
rect 6964 16644 6996 16836
rect 6804 16595 6836 16596
rect 6804 16565 6805 16595
rect 6805 16565 6835 16595
rect 6835 16565 6836 16595
rect 6804 16564 6836 16565
rect 6804 16515 6836 16516
rect 6804 16485 6805 16515
rect 6805 16485 6835 16515
rect 6835 16485 6836 16515
rect 6804 16484 6836 16485
rect 6804 16435 6836 16436
rect 6804 16405 6805 16435
rect 6805 16405 6835 16435
rect 6835 16405 6836 16435
rect 6804 16404 6836 16405
rect 6804 16355 6836 16356
rect 6804 16325 6805 16355
rect 6805 16325 6835 16355
rect 6835 16325 6836 16355
rect 6804 16324 6836 16325
rect 6804 16275 6836 16276
rect 6804 16245 6805 16275
rect 6805 16245 6835 16275
rect 6835 16245 6836 16275
rect 6804 16244 6836 16245
rect 6804 16195 6836 16196
rect 6804 16165 6805 16195
rect 6805 16165 6835 16195
rect 6835 16165 6836 16195
rect 6804 16164 6836 16165
rect 6804 16115 6836 16116
rect 6804 16085 6805 16115
rect 6805 16085 6835 16115
rect 6835 16085 6836 16115
rect 6804 16084 6836 16085
rect 6804 16035 6836 16036
rect 6804 16005 6805 16035
rect 6805 16005 6835 16035
rect 6835 16005 6836 16035
rect 6804 16004 6836 16005
rect 6804 15955 6836 15956
rect 6804 15925 6805 15955
rect 6805 15925 6835 15955
rect 6835 15925 6836 15955
rect 6804 15924 6836 15925
rect 6804 15435 6836 15436
rect 6804 15405 6805 15435
rect 6805 15405 6835 15435
rect 6835 15405 6836 15435
rect 6804 15404 6836 15405
rect 6804 15355 6836 15356
rect 6804 15325 6805 15355
rect 6805 15325 6835 15355
rect 6835 15325 6836 15355
rect 6804 15324 6836 15325
rect 6804 15275 6836 15276
rect 6804 15245 6805 15275
rect 6805 15245 6835 15275
rect 6835 15245 6836 15275
rect 6804 15244 6836 15245
rect 6804 15195 6836 15196
rect 6804 15165 6805 15195
rect 6805 15165 6835 15195
rect 6835 15165 6836 15195
rect 6804 15164 6836 15165
rect 6804 15115 6836 15116
rect 6804 15085 6805 15115
rect 6805 15085 6835 15115
rect 6835 15085 6836 15115
rect 6804 15084 6836 15085
rect 6804 15035 6836 15036
rect 6804 15005 6805 15035
rect 6805 15005 6835 15035
rect 6835 15005 6836 15035
rect 6804 15004 6836 15005
rect 6804 14955 6836 14956
rect 6804 14925 6805 14955
rect 6805 14925 6835 14955
rect 6835 14925 6836 14955
rect 6804 14924 6836 14925
rect 6804 14875 6836 14876
rect 6804 14845 6805 14875
rect 6805 14845 6835 14875
rect 6835 14845 6836 14875
rect 6804 14844 6836 14845
rect 6804 14795 6836 14796
rect 6804 14765 6805 14795
rect 6805 14765 6835 14795
rect 6835 14765 6836 14795
rect 6804 14764 6836 14765
rect 6804 14715 6836 14716
rect 6804 14685 6805 14715
rect 6805 14685 6835 14715
rect 6835 14685 6836 14715
rect 6804 14684 6836 14685
rect 6804 14635 6836 14636
rect 6804 14605 6805 14635
rect 6805 14605 6835 14635
rect 6835 14605 6836 14635
rect 6804 14604 6836 14605
rect 6804 14555 6836 14556
rect 6804 14525 6805 14555
rect 6805 14525 6835 14555
rect 6835 14525 6836 14555
rect 6804 14524 6836 14525
rect 6804 14475 6836 14476
rect 6804 14445 6805 14475
rect 6805 14445 6835 14475
rect 6835 14445 6836 14475
rect 6804 14444 6836 14445
rect 6804 13995 6836 13996
rect 6804 13965 6805 13995
rect 6805 13965 6835 13995
rect 6835 13965 6836 13995
rect 6804 13964 6836 13965
rect 6804 13875 6836 13876
rect 6804 13845 6805 13875
rect 6805 13845 6835 13875
rect 6835 13845 6836 13875
rect 6804 13844 6836 13845
rect 6804 13795 6836 13796
rect 6804 13765 6805 13795
rect 6805 13765 6835 13795
rect 6835 13765 6836 13795
rect 6804 13764 6836 13765
rect 6804 13715 6836 13716
rect 6804 13685 6805 13715
rect 6805 13685 6835 13715
rect 6835 13685 6836 13715
rect 6804 13684 6836 13685
rect 6804 13635 6836 13636
rect 6804 13605 6805 13635
rect 6805 13605 6835 13635
rect 6835 13605 6836 13635
rect 6804 13604 6836 13605
rect 6804 13555 6836 13556
rect 6804 13525 6805 13555
rect 6805 13525 6835 13555
rect 6835 13525 6836 13555
rect 6804 13524 6836 13525
rect 6804 13475 6836 13476
rect 6804 13445 6805 13475
rect 6805 13445 6835 13475
rect 6835 13445 6836 13475
rect 6804 13444 6836 13445
rect 6804 13395 6836 13396
rect 6804 13365 6805 13395
rect 6805 13365 6835 13395
rect 6835 13365 6836 13395
rect 6804 13364 6836 13365
rect 6804 13315 6836 13316
rect 6804 13285 6805 13315
rect 6805 13285 6835 13315
rect 6835 13285 6836 13315
rect 6804 13284 6836 13285
rect 6804 13235 6836 13236
rect 6804 13205 6805 13235
rect 6805 13205 6835 13235
rect 6835 13205 6836 13235
rect 6804 13204 6836 13205
rect 6804 13155 6836 13156
rect 6804 13125 6805 13155
rect 6805 13125 6835 13155
rect 6835 13125 6836 13155
rect 6804 13124 6836 13125
rect 6804 13075 6836 13076
rect 6804 13045 6805 13075
rect 6805 13045 6835 13075
rect 6835 13045 6836 13075
rect 6804 13044 6836 13045
rect 6804 12995 6836 12996
rect 6804 12965 6805 12995
rect 6805 12965 6835 12995
rect 6835 12965 6836 12995
rect 6804 12964 6836 12965
rect 6804 12515 6836 12516
rect 6804 12485 6805 12515
rect 6805 12485 6835 12515
rect 6835 12485 6836 12515
rect 6804 12484 6836 12485
rect 6804 12435 6836 12436
rect 6804 12405 6805 12435
rect 6805 12405 6835 12435
rect 6835 12405 6836 12435
rect 6804 12404 6836 12405
rect 6804 12315 6836 12316
rect 6804 12285 6805 12315
rect 6805 12285 6835 12315
rect 6835 12285 6836 12315
rect 6804 12284 6836 12285
rect 6804 12235 6836 12236
rect 6804 12205 6805 12235
rect 6805 12205 6835 12235
rect 6835 12205 6836 12235
rect 6804 12204 6836 12205
rect 6804 12155 6836 12156
rect 6804 12125 6805 12155
rect 6805 12125 6835 12155
rect 6835 12125 6836 12155
rect 6804 12124 6836 12125
rect 6804 12075 6836 12076
rect 6804 12045 6805 12075
rect 6805 12045 6835 12075
rect 6835 12045 6836 12075
rect 6804 12044 6836 12045
rect 6804 11995 6836 11996
rect 6804 11965 6805 11995
rect 6805 11965 6835 11995
rect 6835 11965 6836 11995
rect 6804 11964 6836 11965
rect 6804 11915 6836 11916
rect 6804 11885 6805 11915
rect 6805 11885 6835 11915
rect 6835 11885 6836 11915
rect 6804 11884 6836 11885
rect 6804 11835 6836 11836
rect 6804 11805 6805 11835
rect 6805 11805 6835 11835
rect 6835 11805 6836 11835
rect 6804 11804 6836 11805
rect 6804 11755 6836 11756
rect 6804 11725 6805 11755
rect 6805 11725 6835 11755
rect 6835 11725 6836 11755
rect 6804 11724 6836 11725
rect 6804 11675 6836 11676
rect 6804 11645 6805 11675
rect 6805 11645 6835 11675
rect 6835 11645 6836 11675
rect 6804 11644 6836 11645
rect 6804 11595 6836 11596
rect 6804 11565 6805 11595
rect 6805 11565 6835 11595
rect 6835 11565 6836 11595
rect 6804 11564 6836 11565
rect 6804 11515 6836 11516
rect 6804 11485 6805 11515
rect 6805 11485 6835 11515
rect 6835 11485 6836 11515
rect 6804 11484 6836 11485
rect 6804 11435 6836 11436
rect 6804 11405 6805 11435
rect 6805 11405 6835 11435
rect 6835 11405 6836 11435
rect 6804 11404 6836 11405
rect 6804 11355 6836 11356
rect 6804 11325 6805 11355
rect 6805 11325 6835 11355
rect 6835 11325 6836 11355
rect 6804 11324 6836 11325
rect 6804 11195 6836 11196
rect 6804 11165 6805 11195
rect 6805 11165 6835 11195
rect 6835 11165 6836 11195
rect 6804 11164 6836 11165
rect 6804 11115 6836 11116
rect 6804 11085 6805 11115
rect 6805 11085 6835 11115
rect 6835 11085 6836 11115
rect 6804 11084 6836 11085
rect 6804 11035 6836 11036
rect 6804 11005 6805 11035
rect 6805 11005 6835 11035
rect 6835 11005 6836 11035
rect 6804 11004 6836 11005
rect 6804 10875 6836 10876
rect 6804 10845 6805 10875
rect 6805 10845 6835 10875
rect 6835 10845 6836 10875
rect 6804 10844 6836 10845
rect 6804 10715 6836 10716
rect 6804 10685 6805 10715
rect 6805 10685 6835 10715
rect 6835 10685 6836 10715
rect 6804 10684 6836 10685
rect 6804 10635 6836 10636
rect 6804 10605 6805 10635
rect 6805 10605 6835 10635
rect 6835 10605 6836 10635
rect 6804 10604 6836 10605
rect 6804 10475 6836 10476
rect 6804 10445 6805 10475
rect 6805 10445 6835 10475
rect 6835 10445 6836 10475
rect 6804 10444 6836 10445
rect 6804 10315 6836 10316
rect 6804 10285 6805 10315
rect 6805 10285 6835 10315
rect 6835 10285 6836 10315
rect 6804 10284 6836 10285
rect 6804 10235 6836 10236
rect 6804 10205 6805 10235
rect 6805 10205 6835 10235
rect 6835 10205 6836 10235
rect 6804 10204 6836 10205
rect 6804 10155 6836 10156
rect 6804 10125 6805 10155
rect 6805 10125 6835 10155
rect 6835 10125 6836 10155
rect 6804 10124 6836 10125
rect 6804 10075 6836 10076
rect 6804 10045 6805 10075
rect 6805 10045 6835 10075
rect 6835 10045 6836 10075
rect 6804 10044 6836 10045
rect 6804 9995 6836 9996
rect 6804 9965 6805 9995
rect 6805 9965 6835 9995
rect 6835 9965 6836 9995
rect 6804 9964 6836 9965
rect 6804 9915 6836 9916
rect 6804 9885 6805 9915
rect 6805 9885 6835 9915
rect 6835 9885 6836 9915
rect 6804 9884 6836 9885
rect 6804 9835 6836 9836
rect 6804 9805 6805 9835
rect 6805 9805 6835 9835
rect 6835 9805 6836 9835
rect 6804 9804 6836 9805
rect 6804 9755 6836 9756
rect 6804 9725 6805 9755
rect 6805 9725 6835 9755
rect 6835 9725 6836 9755
rect 6804 9724 6836 9725
rect 6804 9675 6836 9676
rect 6804 9645 6805 9675
rect 6805 9645 6835 9675
rect 6835 9645 6836 9675
rect 6804 9644 6836 9645
rect 6804 9595 6836 9596
rect 6804 9565 6805 9595
rect 6805 9565 6835 9595
rect 6835 9565 6836 9595
rect 6804 9564 6836 9565
rect 6804 9515 6836 9516
rect 6804 9485 6805 9515
rect 6805 9485 6835 9515
rect 6835 9485 6836 9515
rect 6804 9484 6836 9485
rect 6804 9435 6836 9436
rect 6804 9405 6805 9435
rect 6805 9405 6835 9435
rect 6835 9405 6836 9435
rect 6804 9404 6836 9405
rect 6804 9355 6836 9356
rect 6804 9325 6805 9355
rect 6805 9325 6835 9355
rect 6835 9325 6836 9355
rect 6804 9324 6836 9325
rect 6804 9275 6836 9276
rect 6804 9245 6805 9275
rect 6805 9245 6835 9275
rect 6835 9245 6836 9275
rect 6804 9244 6836 9245
rect 6804 9115 6836 9116
rect 6804 9085 6805 9115
rect 6805 9085 6835 9115
rect 6835 9085 6836 9115
rect 6804 9084 6836 9085
rect 6804 9035 6836 9036
rect 6804 9005 6805 9035
rect 6805 9005 6835 9035
rect 6835 9005 6836 9035
rect 6804 9004 6836 9005
rect 6804 8955 6836 8956
rect 6804 8925 6805 8955
rect 6805 8925 6835 8955
rect 6835 8925 6836 8955
rect 6804 8924 6836 8925
rect 6804 8635 6836 8636
rect 6804 8605 6805 8635
rect 6805 8605 6835 8635
rect 6835 8605 6836 8635
rect 6804 8604 6836 8605
rect 6804 8555 6836 8556
rect 6804 8525 6805 8555
rect 6805 8525 6835 8555
rect 6835 8525 6836 8555
rect 6804 8524 6836 8525
rect 6804 8395 6836 8396
rect 6804 8365 6805 8395
rect 6805 8365 6835 8395
rect 6835 8365 6836 8395
rect 6804 8364 6836 8365
rect 6804 8315 6836 8316
rect 6804 8285 6805 8315
rect 6805 8285 6835 8315
rect 6835 8285 6836 8315
rect 6804 8284 6836 8285
rect 6804 8235 6836 8236
rect 6804 8205 6805 8235
rect 6805 8205 6835 8235
rect 6835 8205 6836 8235
rect 6804 8204 6836 8205
rect 6804 8155 6836 8156
rect 6804 8125 6805 8155
rect 6805 8125 6835 8155
rect 6835 8125 6836 8155
rect 6804 8124 6836 8125
rect 6804 8075 6836 8076
rect 6804 8045 6805 8075
rect 6805 8045 6835 8075
rect 6835 8045 6836 8075
rect 6804 8044 6836 8045
rect 6804 7995 6836 7996
rect 6804 7965 6805 7995
rect 6805 7965 6835 7995
rect 6835 7965 6836 7995
rect 6804 7964 6836 7965
rect 6804 7915 6836 7916
rect 6804 7885 6805 7915
rect 6805 7885 6835 7915
rect 6835 7885 6836 7915
rect 6804 7884 6836 7885
rect 6804 7835 6836 7836
rect 6804 7805 6805 7835
rect 6805 7805 6835 7835
rect 6835 7805 6836 7835
rect 6804 7804 6836 7805
rect 6804 7755 6836 7756
rect 6804 7725 6805 7755
rect 6805 7725 6835 7755
rect 6835 7725 6836 7755
rect 6804 7724 6836 7725
rect 6804 7675 6836 7676
rect 6804 7645 6805 7675
rect 6805 7645 6835 7675
rect 6835 7645 6836 7675
rect 6804 7644 6836 7645
rect 6804 7595 6836 7596
rect 6804 7565 6805 7595
rect 6805 7565 6835 7595
rect 6835 7565 6836 7595
rect 6804 7564 6836 7565
rect 6804 7515 6836 7516
rect 6804 7485 6805 7515
rect 6805 7485 6835 7515
rect 6835 7485 6836 7515
rect 6804 7484 6836 7485
rect 6804 7435 6836 7436
rect 6804 7405 6805 7435
rect 6805 7405 6835 7435
rect 6835 7405 6836 7435
rect 6804 7404 6836 7405
rect 6804 7355 6836 7356
rect 6804 7325 6805 7355
rect 6805 7325 6835 7355
rect 6835 7325 6836 7355
rect 6804 7324 6836 7325
rect 6804 7275 6836 7276
rect 6804 7245 6805 7275
rect 6805 7245 6835 7275
rect 6835 7245 6836 7275
rect 6804 7244 6836 7245
rect 6804 7195 6836 7196
rect 6804 7165 6805 7195
rect 6805 7165 6835 7195
rect 6835 7165 6836 7195
rect 6804 7164 6836 7165
rect 6804 7115 6836 7116
rect 6804 7085 6805 7115
rect 6805 7085 6835 7115
rect 6835 7085 6836 7115
rect 6804 7084 6836 7085
rect 6804 7035 6836 7036
rect 6804 7005 6805 7035
rect 6805 7005 6835 7035
rect 6835 7005 6836 7035
rect 6804 7004 6836 7005
rect 6804 6955 6836 6956
rect 6804 6925 6805 6955
rect 6805 6925 6835 6955
rect 6835 6925 6836 6955
rect 6804 6924 6836 6925
rect 6804 6875 6836 6876
rect 6804 6845 6805 6875
rect 6805 6845 6835 6875
rect 6835 6845 6836 6875
rect 6804 6844 6836 6845
rect 6804 6795 6836 6796
rect 6804 6765 6805 6795
rect 6805 6765 6835 6795
rect 6835 6765 6836 6795
rect 6804 6764 6836 6765
rect 6804 6715 6836 6716
rect 6804 6685 6805 6715
rect 6805 6685 6835 6715
rect 6835 6685 6836 6715
rect 6804 6684 6836 6685
rect 6804 6635 6836 6636
rect 6804 6605 6805 6635
rect 6805 6605 6835 6635
rect 6835 6605 6836 6635
rect 6804 6604 6836 6605
rect 6804 6555 6836 6556
rect 6804 6525 6805 6555
rect 6805 6525 6835 6555
rect 6835 6525 6836 6555
rect 6804 6524 6836 6525
rect 6804 6475 6836 6476
rect 6804 6445 6805 6475
rect 6805 6445 6835 6475
rect 6835 6445 6836 6475
rect 6804 6444 6836 6445
rect 6804 6395 6836 6396
rect 6804 6365 6805 6395
rect 6805 6365 6835 6395
rect 6835 6365 6836 6395
rect 6804 6364 6836 6365
rect 6804 6315 6836 6316
rect 6804 6285 6805 6315
rect 6805 6285 6835 6315
rect 6835 6285 6836 6315
rect 6804 6284 6836 6285
rect 6804 6235 6836 6236
rect 6804 6205 6805 6235
rect 6805 6205 6835 6235
rect 6835 6205 6836 6235
rect 6804 6204 6836 6205
rect 6804 6155 6836 6156
rect 6804 6125 6805 6155
rect 6805 6125 6835 6155
rect 6835 6125 6836 6155
rect 6804 6124 6836 6125
rect 6804 5995 6836 5996
rect 6804 5965 6805 5995
rect 6805 5965 6835 5995
rect 6835 5965 6836 5995
rect 6804 5964 6836 5965
rect 6804 5835 6836 5836
rect 6804 5805 6805 5835
rect 6805 5805 6835 5835
rect 6835 5805 6836 5835
rect 6804 5804 6836 5805
rect 6804 5755 6836 5756
rect 6804 5725 6805 5755
rect 6805 5725 6835 5755
rect 6835 5725 6836 5755
rect 6804 5724 6836 5725
rect 6804 5675 6836 5676
rect 6804 5645 6805 5675
rect 6805 5645 6835 5675
rect 6835 5645 6836 5675
rect 6804 5644 6836 5645
rect 6804 5595 6836 5596
rect 6804 5565 6805 5595
rect 6805 5565 6835 5595
rect 6835 5565 6836 5595
rect 6804 5564 6836 5565
rect 6804 5515 6836 5516
rect 6804 5485 6805 5515
rect 6805 5485 6835 5515
rect 6835 5485 6836 5515
rect 6804 5484 6836 5485
rect 6804 5435 6836 5436
rect 6804 5405 6805 5435
rect 6805 5405 6835 5435
rect 6835 5405 6836 5435
rect 6804 5404 6836 5405
rect 6804 5355 6836 5356
rect 6804 5325 6805 5355
rect 6805 5325 6835 5355
rect 6835 5325 6836 5355
rect 6804 5324 6836 5325
rect 6804 5275 6836 5276
rect 6804 5245 6805 5275
rect 6805 5245 6835 5275
rect 6835 5245 6836 5275
rect 6804 5244 6836 5245
rect 6804 5195 6836 5196
rect 6804 5165 6805 5195
rect 6805 5165 6835 5195
rect 6835 5165 6836 5195
rect 6804 5164 6836 5165
rect 6804 5115 6836 5116
rect 6804 5085 6805 5115
rect 6805 5085 6835 5115
rect 6835 5085 6836 5115
rect 6804 5084 6836 5085
rect 6804 5035 6836 5036
rect 6804 5005 6805 5035
rect 6805 5005 6835 5035
rect 6835 5005 6836 5035
rect 6804 5004 6836 5005
rect 6804 4955 6836 4956
rect 6804 4925 6805 4955
rect 6805 4925 6835 4955
rect 6835 4925 6836 4955
rect 6804 4924 6836 4925
rect 6804 4875 6836 4876
rect 6804 4845 6805 4875
rect 6805 4845 6835 4875
rect 6835 4845 6836 4875
rect 6804 4844 6836 4845
rect 6804 4795 6836 4796
rect 6804 4765 6805 4795
rect 6805 4765 6835 4795
rect 6835 4765 6836 4795
rect 6804 4764 6836 4765
rect 6804 4715 6836 4716
rect 6804 4685 6805 4715
rect 6805 4685 6835 4715
rect 6835 4685 6836 4715
rect 6804 4684 6836 4685
rect 6804 4635 6836 4636
rect 6804 4605 6805 4635
rect 6805 4605 6835 4635
rect 6835 4605 6836 4635
rect 6804 4604 6836 4605
rect 6804 4555 6836 4556
rect 6804 4525 6805 4555
rect 6805 4525 6835 4555
rect 6835 4525 6836 4555
rect 6804 4524 6836 4525
rect 6804 4475 6836 4476
rect 6804 4445 6805 4475
rect 6805 4445 6835 4475
rect 6835 4445 6836 4475
rect 6804 4444 6836 4445
rect 6804 4395 6836 4396
rect 6804 4365 6805 4395
rect 6805 4365 6835 4395
rect 6835 4365 6836 4395
rect 6804 4364 6836 4365
rect 6804 4315 6836 4316
rect 6804 4285 6805 4315
rect 6805 4285 6835 4315
rect 6835 4285 6836 4315
rect 6804 4284 6836 4285
rect 6804 4235 6836 4236
rect 6804 4205 6805 4235
rect 6805 4205 6835 4235
rect 6835 4205 6836 4235
rect 6804 4204 6836 4205
rect 6804 4155 6836 4156
rect 6804 4125 6805 4155
rect 6805 4125 6835 4155
rect 6835 4125 6836 4155
rect 6804 4124 6836 4125
rect 6804 4075 6836 4076
rect 6804 4045 6805 4075
rect 6805 4045 6835 4075
rect 6835 4045 6836 4075
rect 6804 4044 6836 4045
rect 6804 3995 6836 3996
rect 6804 3965 6805 3995
rect 6805 3965 6835 3995
rect 6835 3965 6836 3995
rect 6804 3964 6836 3965
rect 6804 3915 6836 3916
rect 6804 3885 6805 3915
rect 6805 3885 6835 3915
rect 6835 3885 6836 3915
rect 6804 3884 6836 3885
rect 6804 3835 6836 3836
rect 6804 3805 6805 3835
rect 6805 3805 6835 3835
rect 6835 3805 6836 3835
rect 6804 3804 6836 3805
rect 6804 3755 6836 3756
rect 6804 3725 6805 3755
rect 6805 3725 6835 3755
rect 6835 3725 6836 3755
rect 6804 3724 6836 3725
rect 6804 3595 6836 3596
rect 6804 3565 6805 3595
rect 6805 3565 6835 3595
rect 6835 3565 6836 3595
rect 6804 3564 6836 3565
rect 6804 3515 6836 3516
rect 6804 3485 6805 3515
rect 6805 3485 6835 3515
rect 6835 3485 6836 3515
rect 6804 3484 6836 3485
rect 6804 3435 6836 3436
rect 6804 3405 6805 3435
rect 6805 3405 6835 3435
rect 6835 3405 6836 3435
rect 6804 3404 6836 3405
rect 6804 3355 6836 3356
rect 6804 3325 6805 3355
rect 6805 3325 6835 3355
rect 6835 3325 6836 3355
rect 6804 3324 6836 3325
rect 6804 3275 6836 3276
rect 6804 3245 6805 3275
rect 6805 3245 6835 3275
rect 6835 3245 6836 3275
rect 6804 3244 6836 3245
rect 6804 3195 6836 3196
rect 6804 3165 6805 3195
rect 6805 3165 6835 3195
rect 6835 3165 6836 3195
rect 6804 3164 6836 3165
rect 6804 3115 6836 3116
rect 6804 3085 6805 3115
rect 6805 3085 6835 3115
rect 6835 3085 6836 3115
rect 6804 3084 6836 3085
rect 6804 3035 6836 3036
rect 6804 3005 6805 3035
rect 6805 3005 6835 3035
rect 6835 3005 6836 3035
rect 6804 3004 6836 3005
rect 6804 2955 6836 2956
rect 6804 2925 6805 2955
rect 6805 2925 6835 2955
rect 6835 2925 6836 2955
rect 6804 2924 6836 2925
rect 6804 2875 6836 2876
rect 6804 2845 6805 2875
rect 6805 2845 6835 2875
rect 6835 2845 6836 2875
rect 6804 2844 6836 2845
rect 6804 2795 6836 2796
rect 6804 2765 6805 2795
rect 6805 2765 6835 2795
rect 6835 2765 6836 2795
rect 6804 2764 6836 2765
rect 6804 2715 6836 2716
rect 6804 2685 6805 2715
rect 6805 2685 6835 2715
rect 6835 2685 6836 2715
rect 6804 2684 6836 2685
rect 6804 2635 6836 2636
rect 6804 2605 6805 2635
rect 6805 2605 6835 2635
rect 6835 2605 6836 2635
rect 6804 2604 6836 2605
rect 6804 2555 6836 2556
rect 6804 2525 6805 2555
rect 6805 2525 6835 2555
rect 6835 2525 6836 2555
rect 6804 2524 6836 2525
rect 6804 2475 6836 2476
rect 6804 2445 6805 2475
rect 6805 2445 6835 2475
rect 6835 2445 6836 2475
rect 6804 2444 6836 2445
rect 6804 2395 6836 2396
rect 6804 2365 6805 2395
rect 6805 2365 6835 2395
rect 6835 2365 6836 2395
rect 6804 2364 6836 2365
rect 6804 2315 6836 2316
rect 6804 2285 6805 2315
rect 6805 2285 6835 2315
rect 6835 2285 6836 2315
rect 6804 2284 6836 2285
rect 6804 2235 6836 2236
rect 6804 2205 6805 2235
rect 6805 2205 6835 2235
rect 6835 2205 6836 2235
rect 6804 2204 6836 2205
rect 6804 2155 6836 2156
rect 6804 2125 6805 2155
rect 6805 2125 6835 2155
rect 6835 2125 6836 2155
rect 6804 2124 6836 2125
rect 6804 2075 6836 2076
rect 6804 2045 6805 2075
rect 6805 2045 6835 2075
rect 6835 2045 6836 2075
rect 6804 2044 6836 2045
rect 6804 1995 6836 1996
rect 6804 1965 6805 1995
rect 6805 1965 6835 1995
rect 6835 1965 6836 1995
rect 6804 1964 6836 1965
rect 6804 1915 6836 1916
rect 6804 1885 6805 1915
rect 6805 1885 6835 1915
rect 6835 1885 6836 1915
rect 6804 1884 6836 1885
rect 6804 1835 6836 1836
rect 6804 1805 6805 1835
rect 6805 1805 6835 1835
rect 6835 1805 6836 1835
rect 6804 1804 6836 1805
rect 6804 1755 6836 1756
rect 6804 1725 6805 1755
rect 6805 1725 6835 1755
rect 6835 1725 6836 1755
rect 6804 1724 6836 1725
rect 6804 1675 6836 1676
rect 6804 1645 6805 1675
rect 6805 1645 6835 1675
rect 6835 1645 6836 1675
rect 6804 1644 6836 1645
rect 6804 1595 6836 1596
rect 6804 1565 6805 1595
rect 6805 1565 6835 1595
rect 6835 1565 6836 1595
rect 6804 1564 6836 1565
rect 6804 1515 6836 1516
rect 6804 1485 6805 1515
rect 6805 1485 6835 1515
rect 6835 1485 6836 1515
rect 6804 1484 6836 1485
rect 6804 1435 6836 1436
rect 6804 1405 6805 1435
rect 6805 1405 6835 1435
rect 6835 1405 6836 1435
rect 6804 1404 6836 1405
rect 6804 1355 6836 1356
rect 6804 1325 6805 1355
rect 6805 1325 6835 1355
rect 6835 1325 6836 1355
rect 6804 1324 6836 1325
rect 6804 1275 6836 1276
rect 6804 1245 6805 1275
rect 6805 1245 6835 1275
rect 6835 1245 6836 1275
rect 6804 1244 6836 1245
rect 6804 1195 6836 1196
rect 6804 1165 6805 1195
rect 6805 1165 6835 1195
rect 6835 1165 6836 1195
rect 6804 1164 6836 1165
rect 6804 1115 6836 1116
rect 6804 1085 6805 1115
rect 6805 1085 6835 1115
rect 6835 1085 6836 1115
rect 6804 1084 6836 1085
rect 6804 1035 6836 1036
rect 6804 1005 6805 1035
rect 6805 1005 6835 1035
rect 6835 1005 6836 1035
rect 6804 1004 6836 1005
rect 6804 955 6836 956
rect 6804 925 6805 955
rect 6805 925 6835 955
rect 6835 925 6836 955
rect 6804 924 6836 925
rect 6804 875 6836 876
rect 6804 845 6805 875
rect 6805 845 6835 875
rect 6835 845 6836 875
rect 6804 844 6836 845
rect 6804 795 6836 796
rect 6804 765 6805 795
rect 6805 765 6835 795
rect 6835 765 6836 795
rect 6804 764 6836 765
rect 6804 715 6836 716
rect 6804 685 6805 715
rect 6805 685 6835 715
rect 6835 685 6836 715
rect 6804 684 6836 685
rect 6804 595 6836 596
rect 6804 565 6805 595
rect 6805 565 6835 595
rect 6835 565 6836 595
rect 6804 564 6836 565
rect 6804 515 6836 516
rect 6804 485 6805 515
rect 6805 485 6835 515
rect 6835 485 6836 515
rect 6804 484 6836 485
rect 6804 435 6836 436
rect 6804 405 6805 435
rect 6805 405 6835 435
rect 6835 405 6836 435
rect 6804 404 6836 405
rect 6804 355 6836 356
rect 6804 325 6805 355
rect 6805 325 6835 355
rect 6835 325 6836 355
rect 6804 324 6836 325
rect 6804 275 6836 276
rect 6804 245 6805 275
rect 6805 245 6835 275
rect 6835 245 6836 275
rect 6804 244 6836 245
rect 6804 195 6836 196
rect 6804 165 6805 195
rect 6805 165 6835 195
rect 6835 165 6836 195
rect 6804 164 6836 165
rect 6804 115 6836 116
rect 6804 85 6805 115
rect 6805 85 6835 115
rect 6835 85 6836 115
rect 6804 84 6836 85
rect 6804 35 6836 36
rect 6804 5 6805 35
rect 6805 5 6835 35
rect 6835 5 6836 35
rect 6804 4 6836 5
rect 7124 16644 7156 16836
rect 6964 16595 6996 16596
rect 6964 16565 6965 16595
rect 6965 16565 6995 16595
rect 6995 16565 6996 16595
rect 6964 16564 6996 16565
rect 6964 16515 6996 16516
rect 6964 16485 6965 16515
rect 6965 16485 6995 16515
rect 6995 16485 6996 16515
rect 6964 16484 6996 16485
rect 6964 16435 6996 16436
rect 6964 16405 6965 16435
rect 6965 16405 6995 16435
rect 6995 16405 6996 16435
rect 6964 16404 6996 16405
rect 6964 16355 6996 16356
rect 6964 16325 6965 16355
rect 6965 16325 6995 16355
rect 6995 16325 6996 16355
rect 6964 16324 6996 16325
rect 6964 16275 6996 16276
rect 6964 16245 6965 16275
rect 6965 16245 6995 16275
rect 6995 16245 6996 16275
rect 6964 16244 6996 16245
rect 6964 16195 6996 16196
rect 6964 16165 6965 16195
rect 6965 16165 6995 16195
rect 6995 16165 6996 16195
rect 6964 16164 6996 16165
rect 6964 16115 6996 16116
rect 6964 16085 6965 16115
rect 6965 16085 6995 16115
rect 6995 16085 6996 16115
rect 6964 16084 6996 16085
rect 6964 16035 6996 16036
rect 6964 16005 6965 16035
rect 6965 16005 6995 16035
rect 6995 16005 6996 16035
rect 6964 16004 6996 16005
rect 6964 15955 6996 15956
rect 6964 15925 6965 15955
rect 6965 15925 6995 15955
rect 6995 15925 6996 15955
rect 6964 15924 6996 15925
rect 6964 15435 6996 15436
rect 6964 15405 6965 15435
rect 6965 15405 6995 15435
rect 6995 15405 6996 15435
rect 6964 15404 6996 15405
rect 6964 15355 6996 15356
rect 6964 15325 6965 15355
rect 6965 15325 6995 15355
rect 6995 15325 6996 15355
rect 6964 15324 6996 15325
rect 6964 15275 6996 15276
rect 6964 15245 6965 15275
rect 6965 15245 6995 15275
rect 6995 15245 6996 15275
rect 6964 15244 6996 15245
rect 6964 15195 6996 15196
rect 6964 15165 6965 15195
rect 6965 15165 6995 15195
rect 6995 15165 6996 15195
rect 6964 15164 6996 15165
rect 6964 15115 6996 15116
rect 6964 15085 6965 15115
rect 6965 15085 6995 15115
rect 6995 15085 6996 15115
rect 6964 15084 6996 15085
rect 6964 15035 6996 15036
rect 6964 15005 6965 15035
rect 6965 15005 6995 15035
rect 6995 15005 6996 15035
rect 6964 15004 6996 15005
rect 6964 14955 6996 14956
rect 6964 14925 6965 14955
rect 6965 14925 6995 14955
rect 6995 14925 6996 14955
rect 6964 14924 6996 14925
rect 6964 14875 6996 14876
rect 6964 14845 6965 14875
rect 6965 14845 6995 14875
rect 6995 14845 6996 14875
rect 6964 14844 6996 14845
rect 6964 14795 6996 14796
rect 6964 14765 6965 14795
rect 6965 14765 6995 14795
rect 6995 14765 6996 14795
rect 6964 14764 6996 14765
rect 6964 14715 6996 14716
rect 6964 14685 6965 14715
rect 6965 14685 6995 14715
rect 6995 14685 6996 14715
rect 6964 14684 6996 14685
rect 6964 14635 6996 14636
rect 6964 14605 6965 14635
rect 6965 14605 6995 14635
rect 6995 14605 6996 14635
rect 6964 14604 6996 14605
rect 6964 14555 6996 14556
rect 6964 14525 6965 14555
rect 6965 14525 6995 14555
rect 6995 14525 6996 14555
rect 6964 14524 6996 14525
rect 6964 14475 6996 14476
rect 6964 14445 6965 14475
rect 6965 14445 6995 14475
rect 6995 14445 6996 14475
rect 6964 14444 6996 14445
rect 6964 13995 6996 13996
rect 6964 13965 6965 13995
rect 6965 13965 6995 13995
rect 6995 13965 6996 13995
rect 6964 13964 6996 13965
rect 6964 13875 6996 13876
rect 6964 13845 6965 13875
rect 6965 13845 6995 13875
rect 6995 13845 6996 13875
rect 6964 13844 6996 13845
rect 6964 13795 6996 13796
rect 6964 13765 6965 13795
rect 6965 13765 6995 13795
rect 6995 13765 6996 13795
rect 6964 13764 6996 13765
rect 6964 13715 6996 13716
rect 6964 13685 6965 13715
rect 6965 13685 6995 13715
rect 6995 13685 6996 13715
rect 6964 13684 6996 13685
rect 6964 13635 6996 13636
rect 6964 13605 6965 13635
rect 6965 13605 6995 13635
rect 6995 13605 6996 13635
rect 6964 13604 6996 13605
rect 6964 13555 6996 13556
rect 6964 13525 6965 13555
rect 6965 13525 6995 13555
rect 6995 13525 6996 13555
rect 6964 13524 6996 13525
rect 6964 13475 6996 13476
rect 6964 13445 6965 13475
rect 6965 13445 6995 13475
rect 6995 13445 6996 13475
rect 6964 13444 6996 13445
rect 6964 13395 6996 13396
rect 6964 13365 6965 13395
rect 6965 13365 6995 13395
rect 6995 13365 6996 13395
rect 6964 13364 6996 13365
rect 6964 13315 6996 13316
rect 6964 13285 6965 13315
rect 6965 13285 6995 13315
rect 6995 13285 6996 13315
rect 6964 13284 6996 13285
rect 6964 13235 6996 13236
rect 6964 13205 6965 13235
rect 6965 13205 6995 13235
rect 6995 13205 6996 13235
rect 6964 13204 6996 13205
rect 6964 13155 6996 13156
rect 6964 13125 6965 13155
rect 6965 13125 6995 13155
rect 6995 13125 6996 13155
rect 6964 13124 6996 13125
rect 6964 13075 6996 13076
rect 6964 13045 6965 13075
rect 6965 13045 6995 13075
rect 6995 13045 6996 13075
rect 6964 13044 6996 13045
rect 6964 12995 6996 12996
rect 6964 12965 6965 12995
rect 6965 12965 6995 12995
rect 6995 12965 6996 12995
rect 6964 12964 6996 12965
rect 6964 12515 6996 12516
rect 6964 12485 6965 12515
rect 6965 12485 6995 12515
rect 6995 12485 6996 12515
rect 6964 12484 6996 12485
rect 6964 12435 6996 12436
rect 6964 12405 6965 12435
rect 6965 12405 6995 12435
rect 6995 12405 6996 12435
rect 6964 12404 6996 12405
rect 6964 12315 6996 12316
rect 6964 12285 6965 12315
rect 6965 12285 6995 12315
rect 6995 12285 6996 12315
rect 6964 12284 6996 12285
rect 6964 12235 6996 12236
rect 6964 12205 6965 12235
rect 6965 12205 6995 12235
rect 6995 12205 6996 12235
rect 6964 12204 6996 12205
rect 6964 12155 6996 12156
rect 6964 12125 6965 12155
rect 6965 12125 6995 12155
rect 6995 12125 6996 12155
rect 6964 12124 6996 12125
rect 6964 12075 6996 12076
rect 6964 12045 6965 12075
rect 6965 12045 6995 12075
rect 6995 12045 6996 12075
rect 6964 12044 6996 12045
rect 6964 11995 6996 11996
rect 6964 11965 6965 11995
rect 6965 11965 6995 11995
rect 6995 11965 6996 11995
rect 6964 11964 6996 11965
rect 6964 11915 6996 11916
rect 6964 11885 6965 11915
rect 6965 11885 6995 11915
rect 6995 11885 6996 11915
rect 6964 11884 6996 11885
rect 6964 11835 6996 11836
rect 6964 11805 6965 11835
rect 6965 11805 6995 11835
rect 6995 11805 6996 11835
rect 6964 11804 6996 11805
rect 6964 11755 6996 11756
rect 6964 11725 6965 11755
rect 6965 11725 6995 11755
rect 6995 11725 6996 11755
rect 6964 11724 6996 11725
rect 6964 11675 6996 11676
rect 6964 11645 6965 11675
rect 6965 11645 6995 11675
rect 6995 11645 6996 11675
rect 6964 11644 6996 11645
rect 6964 11595 6996 11596
rect 6964 11565 6965 11595
rect 6965 11565 6995 11595
rect 6995 11565 6996 11595
rect 6964 11564 6996 11565
rect 6964 11515 6996 11516
rect 6964 11485 6965 11515
rect 6965 11485 6995 11515
rect 6995 11485 6996 11515
rect 6964 11484 6996 11485
rect 6964 11435 6996 11436
rect 6964 11405 6965 11435
rect 6965 11405 6995 11435
rect 6995 11405 6996 11435
rect 6964 11404 6996 11405
rect 6964 11355 6996 11356
rect 6964 11325 6965 11355
rect 6965 11325 6995 11355
rect 6995 11325 6996 11355
rect 6964 11324 6996 11325
rect 6964 11195 6996 11196
rect 6964 11165 6965 11195
rect 6965 11165 6995 11195
rect 6995 11165 6996 11195
rect 6964 11164 6996 11165
rect 6964 11115 6996 11116
rect 6964 11085 6965 11115
rect 6965 11085 6995 11115
rect 6995 11085 6996 11115
rect 6964 11084 6996 11085
rect 6964 11035 6996 11036
rect 6964 11005 6965 11035
rect 6965 11005 6995 11035
rect 6995 11005 6996 11035
rect 6964 11004 6996 11005
rect 6964 10875 6996 10876
rect 6964 10845 6965 10875
rect 6965 10845 6995 10875
rect 6995 10845 6996 10875
rect 6964 10844 6996 10845
rect 6964 10715 6996 10716
rect 6964 10685 6965 10715
rect 6965 10685 6995 10715
rect 6995 10685 6996 10715
rect 6964 10684 6996 10685
rect 6964 10635 6996 10636
rect 6964 10605 6965 10635
rect 6965 10605 6995 10635
rect 6995 10605 6996 10635
rect 6964 10604 6996 10605
rect 6964 10475 6996 10476
rect 6964 10445 6965 10475
rect 6965 10445 6995 10475
rect 6995 10445 6996 10475
rect 6964 10444 6996 10445
rect 6964 10395 6996 10396
rect 6964 10365 6965 10395
rect 6965 10365 6995 10395
rect 6995 10365 6996 10395
rect 6964 10364 6996 10365
rect 6964 10315 6996 10316
rect 6964 10285 6965 10315
rect 6965 10285 6995 10315
rect 6995 10285 6996 10315
rect 6964 10284 6996 10285
rect 6964 10235 6996 10236
rect 6964 10205 6965 10235
rect 6965 10205 6995 10235
rect 6995 10205 6996 10235
rect 6964 10204 6996 10205
rect 6964 10155 6996 10156
rect 6964 10125 6965 10155
rect 6965 10125 6995 10155
rect 6995 10125 6996 10155
rect 6964 10124 6996 10125
rect 6964 10075 6996 10076
rect 6964 10045 6965 10075
rect 6965 10045 6995 10075
rect 6995 10045 6996 10075
rect 6964 10044 6996 10045
rect 6964 9995 6996 9996
rect 6964 9965 6965 9995
rect 6965 9965 6995 9995
rect 6995 9965 6996 9995
rect 6964 9964 6996 9965
rect 6964 9915 6996 9916
rect 6964 9885 6965 9915
rect 6965 9885 6995 9915
rect 6995 9885 6996 9915
rect 6964 9884 6996 9885
rect 6964 9835 6996 9836
rect 6964 9805 6965 9835
rect 6965 9805 6995 9835
rect 6995 9805 6996 9835
rect 6964 9804 6996 9805
rect 6964 9755 6996 9756
rect 6964 9725 6965 9755
rect 6965 9725 6995 9755
rect 6995 9725 6996 9755
rect 6964 9724 6996 9725
rect 6964 9675 6996 9676
rect 6964 9645 6965 9675
rect 6965 9645 6995 9675
rect 6995 9645 6996 9675
rect 6964 9644 6996 9645
rect 6964 9595 6996 9596
rect 6964 9565 6965 9595
rect 6965 9565 6995 9595
rect 6995 9565 6996 9595
rect 6964 9564 6996 9565
rect 6964 9515 6996 9516
rect 6964 9485 6965 9515
rect 6965 9485 6995 9515
rect 6995 9485 6996 9515
rect 6964 9484 6996 9485
rect 6964 9435 6996 9436
rect 6964 9405 6965 9435
rect 6965 9405 6995 9435
rect 6995 9405 6996 9435
rect 6964 9404 6996 9405
rect 6964 9355 6996 9356
rect 6964 9325 6965 9355
rect 6965 9325 6995 9355
rect 6995 9325 6996 9355
rect 6964 9324 6996 9325
rect 6964 9275 6996 9276
rect 6964 9245 6965 9275
rect 6965 9245 6995 9275
rect 6995 9245 6996 9275
rect 6964 9244 6996 9245
rect 6964 9115 6996 9116
rect 6964 9085 6965 9115
rect 6965 9085 6995 9115
rect 6995 9085 6996 9115
rect 6964 9084 6996 9085
rect 6964 9035 6996 9036
rect 6964 9005 6965 9035
rect 6965 9005 6995 9035
rect 6995 9005 6996 9035
rect 6964 9004 6996 9005
rect 6964 8955 6996 8956
rect 6964 8925 6965 8955
rect 6965 8925 6995 8955
rect 6995 8925 6996 8955
rect 6964 8924 6996 8925
rect 6964 8635 6996 8636
rect 6964 8605 6965 8635
rect 6965 8605 6995 8635
rect 6995 8605 6996 8635
rect 6964 8604 6996 8605
rect 6964 8555 6996 8556
rect 6964 8525 6965 8555
rect 6965 8525 6995 8555
rect 6995 8525 6996 8555
rect 6964 8524 6996 8525
rect 6964 8395 6996 8396
rect 6964 8365 6965 8395
rect 6965 8365 6995 8395
rect 6995 8365 6996 8395
rect 6964 8364 6996 8365
rect 6964 8315 6996 8316
rect 6964 8285 6965 8315
rect 6965 8285 6995 8315
rect 6995 8285 6996 8315
rect 6964 8284 6996 8285
rect 6964 8235 6996 8236
rect 6964 8205 6965 8235
rect 6965 8205 6995 8235
rect 6995 8205 6996 8235
rect 6964 8204 6996 8205
rect 6964 8155 6996 8156
rect 6964 8125 6965 8155
rect 6965 8125 6995 8155
rect 6995 8125 6996 8155
rect 6964 8124 6996 8125
rect 6964 8075 6996 8076
rect 6964 8045 6965 8075
rect 6965 8045 6995 8075
rect 6995 8045 6996 8075
rect 6964 8044 6996 8045
rect 6964 7995 6996 7996
rect 6964 7965 6965 7995
rect 6965 7965 6995 7995
rect 6995 7965 6996 7995
rect 6964 7964 6996 7965
rect 6964 7915 6996 7916
rect 6964 7885 6965 7915
rect 6965 7885 6995 7915
rect 6995 7885 6996 7915
rect 6964 7884 6996 7885
rect 6964 7835 6996 7836
rect 6964 7805 6965 7835
rect 6965 7805 6995 7835
rect 6995 7805 6996 7835
rect 6964 7804 6996 7805
rect 6964 7755 6996 7756
rect 6964 7725 6965 7755
rect 6965 7725 6995 7755
rect 6995 7725 6996 7755
rect 6964 7724 6996 7725
rect 6964 7675 6996 7676
rect 6964 7645 6965 7675
rect 6965 7645 6995 7675
rect 6995 7645 6996 7675
rect 6964 7644 6996 7645
rect 6964 7595 6996 7596
rect 6964 7565 6965 7595
rect 6965 7565 6995 7595
rect 6995 7565 6996 7595
rect 6964 7564 6996 7565
rect 6964 7515 6996 7516
rect 6964 7485 6965 7515
rect 6965 7485 6995 7515
rect 6995 7485 6996 7515
rect 6964 7484 6996 7485
rect 6964 7435 6996 7436
rect 6964 7405 6965 7435
rect 6965 7405 6995 7435
rect 6995 7405 6996 7435
rect 6964 7404 6996 7405
rect 6964 7355 6996 7356
rect 6964 7325 6965 7355
rect 6965 7325 6995 7355
rect 6995 7325 6996 7355
rect 6964 7324 6996 7325
rect 6964 7275 6996 7276
rect 6964 7245 6965 7275
rect 6965 7245 6995 7275
rect 6995 7245 6996 7275
rect 6964 7244 6996 7245
rect 6964 7195 6996 7196
rect 6964 7165 6965 7195
rect 6965 7165 6995 7195
rect 6995 7165 6996 7195
rect 6964 7164 6996 7165
rect 6964 7115 6996 7116
rect 6964 7085 6965 7115
rect 6965 7085 6995 7115
rect 6995 7085 6996 7115
rect 6964 7084 6996 7085
rect 6964 7035 6996 7036
rect 6964 7005 6965 7035
rect 6965 7005 6995 7035
rect 6995 7005 6996 7035
rect 6964 7004 6996 7005
rect 6964 6955 6996 6956
rect 6964 6925 6965 6955
rect 6965 6925 6995 6955
rect 6995 6925 6996 6955
rect 6964 6924 6996 6925
rect 6964 6875 6996 6876
rect 6964 6845 6965 6875
rect 6965 6845 6995 6875
rect 6995 6845 6996 6875
rect 6964 6844 6996 6845
rect 6964 6795 6996 6796
rect 6964 6765 6965 6795
rect 6965 6765 6995 6795
rect 6995 6765 6996 6795
rect 6964 6764 6996 6765
rect 6964 6715 6996 6716
rect 6964 6685 6965 6715
rect 6965 6685 6995 6715
rect 6995 6685 6996 6715
rect 6964 6684 6996 6685
rect 6964 6635 6996 6636
rect 6964 6605 6965 6635
rect 6965 6605 6995 6635
rect 6995 6605 6996 6635
rect 6964 6604 6996 6605
rect 6964 6555 6996 6556
rect 6964 6525 6965 6555
rect 6965 6525 6995 6555
rect 6995 6525 6996 6555
rect 6964 6524 6996 6525
rect 6964 6475 6996 6476
rect 6964 6445 6965 6475
rect 6965 6445 6995 6475
rect 6995 6445 6996 6475
rect 6964 6444 6996 6445
rect 6964 6395 6996 6396
rect 6964 6365 6965 6395
rect 6965 6365 6995 6395
rect 6995 6365 6996 6395
rect 6964 6364 6996 6365
rect 6964 6315 6996 6316
rect 6964 6285 6965 6315
rect 6965 6285 6995 6315
rect 6995 6285 6996 6315
rect 6964 6284 6996 6285
rect 6964 6235 6996 6236
rect 6964 6205 6965 6235
rect 6965 6205 6995 6235
rect 6995 6205 6996 6235
rect 6964 6204 6996 6205
rect 6964 6155 6996 6156
rect 6964 6125 6965 6155
rect 6965 6125 6995 6155
rect 6995 6125 6996 6155
rect 6964 6124 6996 6125
rect 6964 5995 6996 5996
rect 6964 5965 6965 5995
rect 6965 5965 6995 5995
rect 6995 5965 6996 5995
rect 6964 5964 6996 5965
rect 6964 5915 6996 5916
rect 6964 5885 6965 5915
rect 6965 5885 6995 5915
rect 6995 5885 6996 5915
rect 6964 5884 6996 5885
rect 6964 5835 6996 5836
rect 6964 5805 6965 5835
rect 6965 5805 6995 5835
rect 6995 5805 6996 5835
rect 6964 5804 6996 5805
rect 6964 5755 6996 5756
rect 6964 5725 6965 5755
rect 6965 5725 6995 5755
rect 6995 5725 6996 5755
rect 6964 5724 6996 5725
rect 6964 5675 6996 5676
rect 6964 5645 6965 5675
rect 6965 5645 6995 5675
rect 6995 5645 6996 5675
rect 6964 5644 6996 5645
rect 6964 5595 6996 5596
rect 6964 5565 6965 5595
rect 6965 5565 6995 5595
rect 6995 5565 6996 5595
rect 6964 5564 6996 5565
rect 6964 5515 6996 5516
rect 6964 5485 6965 5515
rect 6965 5485 6995 5515
rect 6995 5485 6996 5515
rect 6964 5484 6996 5485
rect 6964 5435 6996 5436
rect 6964 5405 6965 5435
rect 6965 5405 6995 5435
rect 6995 5405 6996 5435
rect 6964 5404 6996 5405
rect 6964 5355 6996 5356
rect 6964 5325 6965 5355
rect 6965 5325 6995 5355
rect 6995 5325 6996 5355
rect 6964 5324 6996 5325
rect 6964 5275 6996 5276
rect 6964 5245 6965 5275
rect 6965 5245 6995 5275
rect 6995 5245 6996 5275
rect 6964 5244 6996 5245
rect 6964 5195 6996 5196
rect 6964 5165 6965 5195
rect 6965 5165 6995 5195
rect 6995 5165 6996 5195
rect 6964 5164 6996 5165
rect 6964 5115 6996 5116
rect 6964 5085 6965 5115
rect 6965 5085 6995 5115
rect 6995 5085 6996 5115
rect 6964 5084 6996 5085
rect 6964 5035 6996 5036
rect 6964 5005 6965 5035
rect 6965 5005 6995 5035
rect 6995 5005 6996 5035
rect 6964 5004 6996 5005
rect 6964 4955 6996 4956
rect 6964 4925 6965 4955
rect 6965 4925 6995 4955
rect 6995 4925 6996 4955
rect 6964 4924 6996 4925
rect 6964 4875 6996 4876
rect 6964 4845 6965 4875
rect 6965 4845 6995 4875
rect 6995 4845 6996 4875
rect 6964 4844 6996 4845
rect 6964 4795 6996 4796
rect 6964 4765 6965 4795
rect 6965 4765 6995 4795
rect 6995 4765 6996 4795
rect 6964 4764 6996 4765
rect 6964 4715 6996 4716
rect 6964 4685 6965 4715
rect 6965 4685 6995 4715
rect 6995 4685 6996 4715
rect 6964 4684 6996 4685
rect 6964 4635 6996 4636
rect 6964 4605 6965 4635
rect 6965 4605 6995 4635
rect 6995 4605 6996 4635
rect 6964 4604 6996 4605
rect 6964 4555 6996 4556
rect 6964 4525 6965 4555
rect 6965 4525 6995 4555
rect 6995 4525 6996 4555
rect 6964 4524 6996 4525
rect 6964 4475 6996 4476
rect 6964 4445 6965 4475
rect 6965 4445 6995 4475
rect 6995 4445 6996 4475
rect 6964 4444 6996 4445
rect 6964 4395 6996 4396
rect 6964 4365 6965 4395
rect 6965 4365 6995 4395
rect 6995 4365 6996 4395
rect 6964 4364 6996 4365
rect 6964 4315 6996 4316
rect 6964 4285 6965 4315
rect 6965 4285 6995 4315
rect 6995 4285 6996 4315
rect 6964 4284 6996 4285
rect 6964 4235 6996 4236
rect 6964 4205 6965 4235
rect 6965 4205 6995 4235
rect 6995 4205 6996 4235
rect 6964 4204 6996 4205
rect 6964 4155 6996 4156
rect 6964 4125 6965 4155
rect 6965 4125 6995 4155
rect 6995 4125 6996 4155
rect 6964 4124 6996 4125
rect 6964 4075 6996 4076
rect 6964 4045 6965 4075
rect 6965 4045 6995 4075
rect 6995 4045 6996 4075
rect 6964 4044 6996 4045
rect 6964 3995 6996 3996
rect 6964 3965 6965 3995
rect 6965 3965 6995 3995
rect 6995 3965 6996 3995
rect 6964 3964 6996 3965
rect 6964 3915 6996 3916
rect 6964 3885 6965 3915
rect 6965 3885 6995 3915
rect 6995 3885 6996 3915
rect 6964 3884 6996 3885
rect 6964 3835 6996 3836
rect 6964 3805 6965 3835
rect 6965 3805 6995 3835
rect 6995 3805 6996 3835
rect 6964 3804 6996 3805
rect 6964 3755 6996 3756
rect 6964 3725 6965 3755
rect 6965 3725 6995 3755
rect 6995 3725 6996 3755
rect 6964 3724 6996 3725
rect 6964 3595 6996 3596
rect 6964 3565 6965 3595
rect 6965 3565 6995 3595
rect 6995 3565 6996 3595
rect 6964 3564 6996 3565
rect 6964 3515 6996 3516
rect 6964 3485 6965 3515
rect 6965 3485 6995 3515
rect 6995 3485 6996 3515
rect 6964 3484 6996 3485
rect 6964 3435 6996 3436
rect 6964 3405 6965 3435
rect 6965 3405 6995 3435
rect 6995 3405 6996 3435
rect 6964 3404 6996 3405
rect 6964 3355 6996 3356
rect 6964 3325 6965 3355
rect 6965 3325 6995 3355
rect 6995 3325 6996 3355
rect 6964 3324 6996 3325
rect 6964 3275 6996 3276
rect 6964 3245 6965 3275
rect 6965 3245 6995 3275
rect 6995 3245 6996 3275
rect 6964 3244 6996 3245
rect 6964 3195 6996 3196
rect 6964 3165 6965 3195
rect 6965 3165 6995 3195
rect 6995 3165 6996 3195
rect 6964 3164 6996 3165
rect 6964 3115 6996 3116
rect 6964 3085 6965 3115
rect 6965 3085 6995 3115
rect 6995 3085 6996 3115
rect 6964 3084 6996 3085
rect 6964 3035 6996 3036
rect 6964 3005 6965 3035
rect 6965 3005 6995 3035
rect 6995 3005 6996 3035
rect 6964 3004 6996 3005
rect 6964 2955 6996 2956
rect 6964 2925 6965 2955
rect 6965 2925 6995 2955
rect 6995 2925 6996 2955
rect 6964 2924 6996 2925
rect 6964 2875 6996 2876
rect 6964 2845 6965 2875
rect 6965 2845 6995 2875
rect 6995 2845 6996 2875
rect 6964 2844 6996 2845
rect 6964 2795 6996 2796
rect 6964 2765 6965 2795
rect 6965 2765 6995 2795
rect 6995 2765 6996 2795
rect 6964 2764 6996 2765
rect 6964 2715 6996 2716
rect 6964 2685 6965 2715
rect 6965 2685 6995 2715
rect 6995 2685 6996 2715
rect 6964 2684 6996 2685
rect 6964 2635 6996 2636
rect 6964 2605 6965 2635
rect 6965 2605 6995 2635
rect 6995 2605 6996 2635
rect 6964 2604 6996 2605
rect 6964 2555 6996 2556
rect 6964 2525 6965 2555
rect 6965 2525 6995 2555
rect 6995 2525 6996 2555
rect 6964 2524 6996 2525
rect 6964 2475 6996 2476
rect 6964 2445 6965 2475
rect 6965 2445 6995 2475
rect 6995 2445 6996 2475
rect 6964 2444 6996 2445
rect 6964 2395 6996 2396
rect 6964 2365 6965 2395
rect 6965 2365 6995 2395
rect 6995 2365 6996 2395
rect 6964 2364 6996 2365
rect 6964 2315 6996 2316
rect 6964 2285 6965 2315
rect 6965 2285 6995 2315
rect 6995 2285 6996 2315
rect 6964 2284 6996 2285
rect 6964 2235 6996 2236
rect 6964 2205 6965 2235
rect 6965 2205 6995 2235
rect 6995 2205 6996 2235
rect 6964 2204 6996 2205
rect 6964 2155 6996 2156
rect 6964 2125 6965 2155
rect 6965 2125 6995 2155
rect 6995 2125 6996 2155
rect 6964 2124 6996 2125
rect 6964 2075 6996 2076
rect 6964 2045 6965 2075
rect 6965 2045 6995 2075
rect 6995 2045 6996 2075
rect 6964 2044 6996 2045
rect 6964 1995 6996 1996
rect 6964 1965 6965 1995
rect 6965 1965 6995 1995
rect 6995 1965 6996 1995
rect 6964 1964 6996 1965
rect 6964 1915 6996 1916
rect 6964 1885 6965 1915
rect 6965 1885 6995 1915
rect 6995 1885 6996 1915
rect 6964 1884 6996 1885
rect 6964 1835 6996 1836
rect 6964 1805 6965 1835
rect 6965 1805 6995 1835
rect 6995 1805 6996 1835
rect 6964 1804 6996 1805
rect 6964 1755 6996 1756
rect 6964 1725 6965 1755
rect 6965 1725 6995 1755
rect 6995 1725 6996 1755
rect 6964 1724 6996 1725
rect 6964 1675 6996 1676
rect 6964 1645 6965 1675
rect 6965 1645 6995 1675
rect 6995 1645 6996 1675
rect 6964 1644 6996 1645
rect 6964 1595 6996 1596
rect 6964 1565 6965 1595
rect 6965 1565 6995 1595
rect 6995 1565 6996 1595
rect 6964 1564 6996 1565
rect 6964 1515 6996 1516
rect 6964 1485 6965 1515
rect 6965 1485 6995 1515
rect 6995 1485 6996 1515
rect 6964 1484 6996 1485
rect 6964 1435 6996 1436
rect 6964 1405 6965 1435
rect 6965 1405 6995 1435
rect 6995 1405 6996 1435
rect 6964 1404 6996 1405
rect 6964 1355 6996 1356
rect 6964 1325 6965 1355
rect 6965 1325 6995 1355
rect 6995 1325 6996 1355
rect 6964 1324 6996 1325
rect 6964 1275 6996 1276
rect 6964 1245 6965 1275
rect 6965 1245 6995 1275
rect 6995 1245 6996 1275
rect 6964 1244 6996 1245
rect 6964 1195 6996 1196
rect 6964 1165 6965 1195
rect 6965 1165 6995 1195
rect 6995 1165 6996 1195
rect 6964 1164 6996 1165
rect 6964 1115 6996 1116
rect 6964 1085 6965 1115
rect 6965 1085 6995 1115
rect 6995 1085 6996 1115
rect 6964 1084 6996 1085
rect 6964 1035 6996 1036
rect 6964 1005 6965 1035
rect 6965 1005 6995 1035
rect 6995 1005 6996 1035
rect 6964 1004 6996 1005
rect 6964 955 6996 956
rect 6964 925 6965 955
rect 6965 925 6995 955
rect 6995 925 6996 955
rect 6964 924 6996 925
rect 6964 875 6996 876
rect 6964 845 6965 875
rect 6965 845 6995 875
rect 6995 845 6996 875
rect 6964 844 6996 845
rect 6964 795 6996 796
rect 6964 765 6965 795
rect 6965 765 6995 795
rect 6995 765 6996 795
rect 6964 764 6996 765
rect 6964 715 6996 716
rect 6964 685 6965 715
rect 6965 685 6995 715
rect 6995 685 6996 715
rect 6964 684 6996 685
rect 6964 595 6996 596
rect 6964 565 6965 595
rect 6965 565 6995 595
rect 6995 565 6996 595
rect 6964 564 6996 565
rect 6964 515 6996 516
rect 6964 485 6965 515
rect 6965 485 6995 515
rect 6995 485 6996 515
rect 6964 484 6996 485
rect 6964 435 6996 436
rect 6964 405 6965 435
rect 6965 405 6995 435
rect 6995 405 6996 435
rect 6964 404 6996 405
rect 6964 355 6996 356
rect 6964 325 6965 355
rect 6965 325 6995 355
rect 6995 325 6996 355
rect 6964 324 6996 325
rect 6964 275 6996 276
rect 6964 245 6965 275
rect 6965 245 6995 275
rect 6995 245 6996 275
rect 6964 244 6996 245
rect 6964 195 6996 196
rect 6964 165 6965 195
rect 6965 165 6995 195
rect 6995 165 6996 195
rect 6964 164 6996 165
rect 6964 115 6996 116
rect 6964 85 6965 115
rect 6965 85 6995 115
rect 6995 85 6996 115
rect 6964 84 6996 85
rect 6964 35 6996 36
rect 6964 5 6965 35
rect 6965 5 6995 35
rect 6995 5 6996 35
rect 6964 4 6996 5
rect 7284 16644 7316 16836
rect 7124 16595 7156 16596
rect 7124 16565 7125 16595
rect 7125 16565 7155 16595
rect 7155 16565 7156 16595
rect 7124 16564 7156 16565
rect 7124 16515 7156 16516
rect 7124 16485 7125 16515
rect 7125 16485 7155 16515
rect 7155 16485 7156 16515
rect 7124 16484 7156 16485
rect 7124 16435 7156 16436
rect 7124 16405 7125 16435
rect 7125 16405 7155 16435
rect 7155 16405 7156 16435
rect 7124 16404 7156 16405
rect 7124 16355 7156 16356
rect 7124 16325 7125 16355
rect 7125 16325 7155 16355
rect 7155 16325 7156 16355
rect 7124 16324 7156 16325
rect 7124 16275 7156 16276
rect 7124 16245 7125 16275
rect 7125 16245 7155 16275
rect 7155 16245 7156 16275
rect 7124 16244 7156 16245
rect 7124 16195 7156 16196
rect 7124 16165 7125 16195
rect 7125 16165 7155 16195
rect 7155 16165 7156 16195
rect 7124 16164 7156 16165
rect 7124 16115 7156 16116
rect 7124 16085 7125 16115
rect 7125 16085 7155 16115
rect 7155 16085 7156 16115
rect 7124 16084 7156 16085
rect 7124 16035 7156 16036
rect 7124 16005 7125 16035
rect 7125 16005 7155 16035
rect 7155 16005 7156 16035
rect 7124 16004 7156 16005
rect 7124 15955 7156 15956
rect 7124 15925 7125 15955
rect 7125 15925 7155 15955
rect 7155 15925 7156 15955
rect 7124 15924 7156 15925
rect 7124 15435 7156 15436
rect 7124 15405 7125 15435
rect 7125 15405 7155 15435
rect 7155 15405 7156 15435
rect 7124 15404 7156 15405
rect 7124 15355 7156 15356
rect 7124 15325 7125 15355
rect 7125 15325 7155 15355
rect 7155 15325 7156 15355
rect 7124 15324 7156 15325
rect 7124 15275 7156 15276
rect 7124 15245 7125 15275
rect 7125 15245 7155 15275
rect 7155 15245 7156 15275
rect 7124 15244 7156 15245
rect 7124 15195 7156 15196
rect 7124 15165 7125 15195
rect 7125 15165 7155 15195
rect 7155 15165 7156 15195
rect 7124 15164 7156 15165
rect 7124 15115 7156 15116
rect 7124 15085 7125 15115
rect 7125 15085 7155 15115
rect 7155 15085 7156 15115
rect 7124 15084 7156 15085
rect 7124 15035 7156 15036
rect 7124 15005 7125 15035
rect 7125 15005 7155 15035
rect 7155 15005 7156 15035
rect 7124 15004 7156 15005
rect 7124 14955 7156 14956
rect 7124 14925 7125 14955
rect 7125 14925 7155 14955
rect 7155 14925 7156 14955
rect 7124 14924 7156 14925
rect 7124 14875 7156 14876
rect 7124 14845 7125 14875
rect 7125 14845 7155 14875
rect 7155 14845 7156 14875
rect 7124 14844 7156 14845
rect 7124 14795 7156 14796
rect 7124 14765 7125 14795
rect 7125 14765 7155 14795
rect 7155 14765 7156 14795
rect 7124 14764 7156 14765
rect 7124 14715 7156 14716
rect 7124 14685 7125 14715
rect 7125 14685 7155 14715
rect 7155 14685 7156 14715
rect 7124 14684 7156 14685
rect 7124 14635 7156 14636
rect 7124 14605 7125 14635
rect 7125 14605 7155 14635
rect 7155 14605 7156 14635
rect 7124 14604 7156 14605
rect 7124 14555 7156 14556
rect 7124 14525 7125 14555
rect 7125 14525 7155 14555
rect 7155 14525 7156 14555
rect 7124 14524 7156 14525
rect 7124 14475 7156 14476
rect 7124 14445 7125 14475
rect 7125 14445 7155 14475
rect 7155 14445 7156 14475
rect 7124 14444 7156 14445
rect 7124 13995 7156 13996
rect 7124 13965 7125 13995
rect 7125 13965 7155 13995
rect 7155 13965 7156 13995
rect 7124 13964 7156 13965
rect 7124 13875 7156 13876
rect 7124 13845 7125 13875
rect 7125 13845 7155 13875
rect 7155 13845 7156 13875
rect 7124 13844 7156 13845
rect 7124 13795 7156 13796
rect 7124 13765 7125 13795
rect 7125 13765 7155 13795
rect 7155 13765 7156 13795
rect 7124 13764 7156 13765
rect 7124 13715 7156 13716
rect 7124 13685 7125 13715
rect 7125 13685 7155 13715
rect 7155 13685 7156 13715
rect 7124 13684 7156 13685
rect 7124 13635 7156 13636
rect 7124 13605 7125 13635
rect 7125 13605 7155 13635
rect 7155 13605 7156 13635
rect 7124 13604 7156 13605
rect 7124 13555 7156 13556
rect 7124 13525 7125 13555
rect 7125 13525 7155 13555
rect 7155 13525 7156 13555
rect 7124 13524 7156 13525
rect 7124 13475 7156 13476
rect 7124 13445 7125 13475
rect 7125 13445 7155 13475
rect 7155 13445 7156 13475
rect 7124 13444 7156 13445
rect 7124 13395 7156 13396
rect 7124 13365 7125 13395
rect 7125 13365 7155 13395
rect 7155 13365 7156 13395
rect 7124 13364 7156 13365
rect 7124 13315 7156 13316
rect 7124 13285 7125 13315
rect 7125 13285 7155 13315
rect 7155 13285 7156 13315
rect 7124 13284 7156 13285
rect 7124 13235 7156 13236
rect 7124 13205 7125 13235
rect 7125 13205 7155 13235
rect 7155 13205 7156 13235
rect 7124 13204 7156 13205
rect 7124 13155 7156 13156
rect 7124 13125 7125 13155
rect 7125 13125 7155 13155
rect 7155 13125 7156 13155
rect 7124 13124 7156 13125
rect 7124 13075 7156 13076
rect 7124 13045 7125 13075
rect 7125 13045 7155 13075
rect 7155 13045 7156 13075
rect 7124 13044 7156 13045
rect 7124 12995 7156 12996
rect 7124 12965 7125 12995
rect 7125 12965 7155 12995
rect 7155 12965 7156 12995
rect 7124 12964 7156 12965
rect 7124 12515 7156 12516
rect 7124 12485 7125 12515
rect 7125 12485 7155 12515
rect 7155 12485 7156 12515
rect 7124 12484 7156 12485
rect 7124 12435 7156 12436
rect 7124 12405 7125 12435
rect 7125 12405 7155 12435
rect 7155 12405 7156 12435
rect 7124 12404 7156 12405
rect 7124 12315 7156 12316
rect 7124 12285 7125 12315
rect 7125 12285 7155 12315
rect 7155 12285 7156 12315
rect 7124 12284 7156 12285
rect 7124 12235 7156 12236
rect 7124 12205 7125 12235
rect 7125 12205 7155 12235
rect 7155 12205 7156 12235
rect 7124 12204 7156 12205
rect 7124 12155 7156 12156
rect 7124 12125 7125 12155
rect 7125 12125 7155 12155
rect 7155 12125 7156 12155
rect 7124 12124 7156 12125
rect 7124 12075 7156 12076
rect 7124 12045 7125 12075
rect 7125 12045 7155 12075
rect 7155 12045 7156 12075
rect 7124 12044 7156 12045
rect 7124 11995 7156 11996
rect 7124 11965 7125 11995
rect 7125 11965 7155 11995
rect 7155 11965 7156 11995
rect 7124 11964 7156 11965
rect 7124 11915 7156 11916
rect 7124 11885 7125 11915
rect 7125 11885 7155 11915
rect 7155 11885 7156 11915
rect 7124 11884 7156 11885
rect 7124 11835 7156 11836
rect 7124 11805 7125 11835
rect 7125 11805 7155 11835
rect 7155 11805 7156 11835
rect 7124 11804 7156 11805
rect 7124 11755 7156 11756
rect 7124 11725 7125 11755
rect 7125 11725 7155 11755
rect 7155 11725 7156 11755
rect 7124 11724 7156 11725
rect 7124 11675 7156 11676
rect 7124 11645 7125 11675
rect 7125 11645 7155 11675
rect 7155 11645 7156 11675
rect 7124 11644 7156 11645
rect 7124 11595 7156 11596
rect 7124 11565 7125 11595
rect 7125 11565 7155 11595
rect 7155 11565 7156 11595
rect 7124 11564 7156 11565
rect 7124 11515 7156 11516
rect 7124 11485 7125 11515
rect 7125 11485 7155 11515
rect 7155 11485 7156 11515
rect 7124 11484 7156 11485
rect 7124 11435 7156 11436
rect 7124 11405 7125 11435
rect 7125 11405 7155 11435
rect 7155 11405 7156 11435
rect 7124 11404 7156 11405
rect 7124 11355 7156 11356
rect 7124 11325 7125 11355
rect 7125 11325 7155 11355
rect 7155 11325 7156 11355
rect 7124 11324 7156 11325
rect 7124 11195 7156 11196
rect 7124 11165 7125 11195
rect 7125 11165 7155 11195
rect 7155 11165 7156 11195
rect 7124 11164 7156 11165
rect 7124 11115 7156 11116
rect 7124 11085 7125 11115
rect 7125 11085 7155 11115
rect 7155 11085 7156 11115
rect 7124 11084 7156 11085
rect 7124 11035 7156 11036
rect 7124 11005 7125 11035
rect 7125 11005 7155 11035
rect 7155 11005 7156 11035
rect 7124 11004 7156 11005
rect 7124 10875 7156 10876
rect 7124 10845 7125 10875
rect 7125 10845 7155 10875
rect 7155 10845 7156 10875
rect 7124 10844 7156 10845
rect 7124 10795 7156 10796
rect 7124 10765 7125 10795
rect 7125 10765 7155 10795
rect 7155 10765 7156 10795
rect 7124 10764 7156 10765
rect 7124 10715 7156 10716
rect 7124 10685 7125 10715
rect 7125 10685 7155 10715
rect 7155 10685 7156 10715
rect 7124 10684 7156 10685
rect 7124 10635 7156 10636
rect 7124 10605 7125 10635
rect 7125 10605 7155 10635
rect 7155 10605 7156 10635
rect 7124 10604 7156 10605
rect 7124 10555 7156 10556
rect 7124 10525 7125 10555
rect 7125 10525 7155 10555
rect 7155 10525 7156 10555
rect 7124 10524 7156 10525
rect 7124 10475 7156 10476
rect 7124 10445 7125 10475
rect 7125 10445 7155 10475
rect 7155 10445 7156 10475
rect 7124 10444 7156 10445
rect 7124 10395 7156 10396
rect 7124 10365 7125 10395
rect 7125 10365 7155 10395
rect 7155 10365 7156 10395
rect 7124 10364 7156 10365
rect 7124 10315 7156 10316
rect 7124 10285 7125 10315
rect 7125 10285 7155 10315
rect 7155 10285 7156 10315
rect 7124 10284 7156 10285
rect 7124 10235 7156 10236
rect 7124 10205 7125 10235
rect 7125 10205 7155 10235
rect 7155 10205 7156 10235
rect 7124 10204 7156 10205
rect 7124 10155 7156 10156
rect 7124 10125 7125 10155
rect 7125 10125 7155 10155
rect 7155 10125 7156 10155
rect 7124 10124 7156 10125
rect 7124 10075 7156 10076
rect 7124 10045 7125 10075
rect 7125 10045 7155 10075
rect 7155 10045 7156 10075
rect 7124 10044 7156 10045
rect 7124 9995 7156 9996
rect 7124 9965 7125 9995
rect 7125 9965 7155 9995
rect 7155 9965 7156 9995
rect 7124 9964 7156 9965
rect 7124 9915 7156 9916
rect 7124 9885 7125 9915
rect 7125 9885 7155 9915
rect 7155 9885 7156 9915
rect 7124 9884 7156 9885
rect 7124 9835 7156 9836
rect 7124 9805 7125 9835
rect 7125 9805 7155 9835
rect 7155 9805 7156 9835
rect 7124 9804 7156 9805
rect 7124 9755 7156 9756
rect 7124 9725 7125 9755
rect 7125 9725 7155 9755
rect 7155 9725 7156 9755
rect 7124 9724 7156 9725
rect 7124 9675 7156 9676
rect 7124 9645 7125 9675
rect 7125 9645 7155 9675
rect 7155 9645 7156 9675
rect 7124 9644 7156 9645
rect 7124 9595 7156 9596
rect 7124 9565 7125 9595
rect 7125 9565 7155 9595
rect 7155 9565 7156 9595
rect 7124 9564 7156 9565
rect 7124 9515 7156 9516
rect 7124 9485 7125 9515
rect 7125 9485 7155 9515
rect 7155 9485 7156 9515
rect 7124 9484 7156 9485
rect 7124 9435 7156 9436
rect 7124 9405 7125 9435
rect 7125 9405 7155 9435
rect 7155 9405 7156 9435
rect 7124 9404 7156 9405
rect 7124 9355 7156 9356
rect 7124 9325 7125 9355
rect 7125 9325 7155 9355
rect 7155 9325 7156 9355
rect 7124 9324 7156 9325
rect 7124 9275 7156 9276
rect 7124 9245 7125 9275
rect 7125 9245 7155 9275
rect 7155 9245 7156 9275
rect 7124 9244 7156 9245
rect 7124 9115 7156 9116
rect 7124 9085 7125 9115
rect 7125 9085 7155 9115
rect 7155 9085 7156 9115
rect 7124 9084 7156 9085
rect 7124 9035 7156 9036
rect 7124 9005 7125 9035
rect 7125 9005 7155 9035
rect 7155 9005 7156 9035
rect 7124 9004 7156 9005
rect 7124 8955 7156 8956
rect 7124 8925 7125 8955
rect 7125 8925 7155 8955
rect 7155 8925 7156 8955
rect 7124 8924 7156 8925
rect 7124 8635 7156 8636
rect 7124 8605 7125 8635
rect 7125 8605 7155 8635
rect 7155 8605 7156 8635
rect 7124 8604 7156 8605
rect 7124 8555 7156 8556
rect 7124 8525 7125 8555
rect 7125 8525 7155 8555
rect 7155 8525 7156 8555
rect 7124 8524 7156 8525
rect 7124 8475 7156 8476
rect 7124 8445 7125 8475
rect 7125 8445 7155 8475
rect 7155 8445 7156 8475
rect 7124 8444 7156 8445
rect 7124 8395 7156 8396
rect 7124 8365 7125 8395
rect 7125 8365 7155 8395
rect 7155 8365 7156 8395
rect 7124 8364 7156 8365
rect 7124 8315 7156 8316
rect 7124 8285 7125 8315
rect 7125 8285 7155 8315
rect 7155 8285 7156 8315
rect 7124 8284 7156 8285
rect 7124 8235 7156 8236
rect 7124 8205 7125 8235
rect 7125 8205 7155 8235
rect 7155 8205 7156 8235
rect 7124 8204 7156 8205
rect 7124 8155 7156 8156
rect 7124 8125 7125 8155
rect 7125 8125 7155 8155
rect 7155 8125 7156 8155
rect 7124 8124 7156 8125
rect 7124 8075 7156 8076
rect 7124 8045 7125 8075
rect 7125 8045 7155 8075
rect 7155 8045 7156 8075
rect 7124 8044 7156 8045
rect 7124 7995 7156 7996
rect 7124 7965 7125 7995
rect 7125 7965 7155 7995
rect 7155 7965 7156 7995
rect 7124 7964 7156 7965
rect 7124 7915 7156 7916
rect 7124 7885 7125 7915
rect 7125 7885 7155 7915
rect 7155 7885 7156 7915
rect 7124 7884 7156 7885
rect 7124 7835 7156 7836
rect 7124 7805 7125 7835
rect 7125 7805 7155 7835
rect 7155 7805 7156 7835
rect 7124 7804 7156 7805
rect 7124 7755 7156 7756
rect 7124 7725 7125 7755
rect 7125 7725 7155 7755
rect 7155 7725 7156 7755
rect 7124 7724 7156 7725
rect 7124 7675 7156 7676
rect 7124 7645 7125 7675
rect 7125 7645 7155 7675
rect 7155 7645 7156 7675
rect 7124 7644 7156 7645
rect 7124 7595 7156 7596
rect 7124 7565 7125 7595
rect 7125 7565 7155 7595
rect 7155 7565 7156 7595
rect 7124 7564 7156 7565
rect 7124 7515 7156 7516
rect 7124 7485 7125 7515
rect 7125 7485 7155 7515
rect 7155 7485 7156 7515
rect 7124 7484 7156 7485
rect 7124 7435 7156 7436
rect 7124 7405 7125 7435
rect 7125 7405 7155 7435
rect 7155 7405 7156 7435
rect 7124 7404 7156 7405
rect 7124 7355 7156 7356
rect 7124 7325 7125 7355
rect 7125 7325 7155 7355
rect 7155 7325 7156 7355
rect 7124 7324 7156 7325
rect 7124 7275 7156 7276
rect 7124 7245 7125 7275
rect 7125 7245 7155 7275
rect 7155 7245 7156 7275
rect 7124 7244 7156 7245
rect 7124 7195 7156 7196
rect 7124 7165 7125 7195
rect 7125 7165 7155 7195
rect 7155 7165 7156 7195
rect 7124 7164 7156 7165
rect 7124 7115 7156 7116
rect 7124 7085 7125 7115
rect 7125 7085 7155 7115
rect 7155 7085 7156 7115
rect 7124 7084 7156 7085
rect 7124 7035 7156 7036
rect 7124 7005 7125 7035
rect 7125 7005 7155 7035
rect 7155 7005 7156 7035
rect 7124 7004 7156 7005
rect 7124 6955 7156 6956
rect 7124 6925 7125 6955
rect 7125 6925 7155 6955
rect 7155 6925 7156 6955
rect 7124 6924 7156 6925
rect 7124 6875 7156 6876
rect 7124 6845 7125 6875
rect 7125 6845 7155 6875
rect 7155 6845 7156 6875
rect 7124 6844 7156 6845
rect 7124 6795 7156 6796
rect 7124 6765 7125 6795
rect 7125 6765 7155 6795
rect 7155 6765 7156 6795
rect 7124 6764 7156 6765
rect 7124 6715 7156 6716
rect 7124 6685 7125 6715
rect 7125 6685 7155 6715
rect 7155 6685 7156 6715
rect 7124 6684 7156 6685
rect 7124 6635 7156 6636
rect 7124 6605 7125 6635
rect 7125 6605 7155 6635
rect 7155 6605 7156 6635
rect 7124 6604 7156 6605
rect 7124 6555 7156 6556
rect 7124 6525 7125 6555
rect 7125 6525 7155 6555
rect 7155 6525 7156 6555
rect 7124 6524 7156 6525
rect 7124 6475 7156 6476
rect 7124 6445 7125 6475
rect 7125 6445 7155 6475
rect 7155 6445 7156 6475
rect 7124 6444 7156 6445
rect 7124 6395 7156 6396
rect 7124 6365 7125 6395
rect 7125 6365 7155 6395
rect 7155 6365 7156 6395
rect 7124 6364 7156 6365
rect 7124 6315 7156 6316
rect 7124 6285 7125 6315
rect 7125 6285 7155 6315
rect 7155 6285 7156 6315
rect 7124 6284 7156 6285
rect 7124 6235 7156 6236
rect 7124 6205 7125 6235
rect 7125 6205 7155 6235
rect 7155 6205 7156 6235
rect 7124 6204 7156 6205
rect 7124 6155 7156 6156
rect 7124 6125 7125 6155
rect 7125 6125 7155 6155
rect 7155 6125 7156 6155
rect 7124 6124 7156 6125
rect 7124 6075 7156 6076
rect 7124 6045 7125 6075
rect 7125 6045 7155 6075
rect 7155 6045 7156 6075
rect 7124 6044 7156 6045
rect 7124 5995 7156 5996
rect 7124 5965 7125 5995
rect 7125 5965 7155 5995
rect 7155 5965 7156 5995
rect 7124 5964 7156 5965
rect 7124 5915 7156 5916
rect 7124 5885 7125 5915
rect 7125 5885 7155 5915
rect 7155 5885 7156 5915
rect 7124 5884 7156 5885
rect 7124 5835 7156 5836
rect 7124 5805 7125 5835
rect 7125 5805 7155 5835
rect 7155 5805 7156 5835
rect 7124 5804 7156 5805
rect 7124 5755 7156 5756
rect 7124 5725 7125 5755
rect 7125 5725 7155 5755
rect 7155 5725 7156 5755
rect 7124 5724 7156 5725
rect 7124 5675 7156 5676
rect 7124 5645 7125 5675
rect 7125 5645 7155 5675
rect 7155 5645 7156 5675
rect 7124 5644 7156 5645
rect 7124 5595 7156 5596
rect 7124 5565 7125 5595
rect 7125 5565 7155 5595
rect 7155 5565 7156 5595
rect 7124 5564 7156 5565
rect 7124 5515 7156 5516
rect 7124 5485 7125 5515
rect 7125 5485 7155 5515
rect 7155 5485 7156 5515
rect 7124 5484 7156 5485
rect 7124 5435 7156 5436
rect 7124 5405 7125 5435
rect 7125 5405 7155 5435
rect 7155 5405 7156 5435
rect 7124 5404 7156 5405
rect 7124 5355 7156 5356
rect 7124 5325 7125 5355
rect 7125 5325 7155 5355
rect 7155 5325 7156 5355
rect 7124 5324 7156 5325
rect 7124 5275 7156 5276
rect 7124 5245 7125 5275
rect 7125 5245 7155 5275
rect 7155 5245 7156 5275
rect 7124 5244 7156 5245
rect 7124 5195 7156 5196
rect 7124 5165 7125 5195
rect 7125 5165 7155 5195
rect 7155 5165 7156 5195
rect 7124 5164 7156 5165
rect 7124 5115 7156 5116
rect 7124 5085 7125 5115
rect 7125 5085 7155 5115
rect 7155 5085 7156 5115
rect 7124 5084 7156 5085
rect 7124 5035 7156 5036
rect 7124 5005 7125 5035
rect 7125 5005 7155 5035
rect 7155 5005 7156 5035
rect 7124 5004 7156 5005
rect 7124 4955 7156 4956
rect 7124 4925 7125 4955
rect 7125 4925 7155 4955
rect 7155 4925 7156 4955
rect 7124 4924 7156 4925
rect 7124 4875 7156 4876
rect 7124 4845 7125 4875
rect 7125 4845 7155 4875
rect 7155 4845 7156 4875
rect 7124 4844 7156 4845
rect 7124 4795 7156 4796
rect 7124 4765 7125 4795
rect 7125 4765 7155 4795
rect 7155 4765 7156 4795
rect 7124 4764 7156 4765
rect 7124 4715 7156 4716
rect 7124 4685 7125 4715
rect 7125 4685 7155 4715
rect 7155 4685 7156 4715
rect 7124 4684 7156 4685
rect 7124 4635 7156 4636
rect 7124 4605 7125 4635
rect 7125 4605 7155 4635
rect 7155 4605 7156 4635
rect 7124 4604 7156 4605
rect 7124 4555 7156 4556
rect 7124 4525 7125 4555
rect 7125 4525 7155 4555
rect 7155 4525 7156 4555
rect 7124 4524 7156 4525
rect 7124 4475 7156 4476
rect 7124 4445 7125 4475
rect 7125 4445 7155 4475
rect 7155 4445 7156 4475
rect 7124 4444 7156 4445
rect 7124 4395 7156 4396
rect 7124 4365 7125 4395
rect 7125 4365 7155 4395
rect 7155 4365 7156 4395
rect 7124 4364 7156 4365
rect 7124 4315 7156 4316
rect 7124 4285 7125 4315
rect 7125 4285 7155 4315
rect 7155 4285 7156 4315
rect 7124 4284 7156 4285
rect 7124 4235 7156 4236
rect 7124 4205 7125 4235
rect 7125 4205 7155 4235
rect 7155 4205 7156 4235
rect 7124 4204 7156 4205
rect 7124 4155 7156 4156
rect 7124 4125 7125 4155
rect 7125 4125 7155 4155
rect 7155 4125 7156 4155
rect 7124 4124 7156 4125
rect 7124 4075 7156 4076
rect 7124 4045 7125 4075
rect 7125 4045 7155 4075
rect 7155 4045 7156 4075
rect 7124 4044 7156 4045
rect 7124 3995 7156 3996
rect 7124 3965 7125 3995
rect 7125 3965 7155 3995
rect 7155 3965 7156 3995
rect 7124 3964 7156 3965
rect 7124 3915 7156 3916
rect 7124 3885 7125 3915
rect 7125 3885 7155 3915
rect 7155 3885 7156 3915
rect 7124 3884 7156 3885
rect 7124 3835 7156 3836
rect 7124 3805 7125 3835
rect 7125 3805 7155 3835
rect 7155 3805 7156 3835
rect 7124 3804 7156 3805
rect 7124 3755 7156 3756
rect 7124 3725 7125 3755
rect 7125 3725 7155 3755
rect 7155 3725 7156 3755
rect 7124 3724 7156 3725
rect 7124 3675 7156 3676
rect 7124 3645 7125 3675
rect 7125 3645 7155 3675
rect 7155 3645 7156 3675
rect 7124 3644 7156 3645
rect 7124 3595 7156 3596
rect 7124 3565 7125 3595
rect 7125 3565 7155 3595
rect 7155 3565 7156 3595
rect 7124 3564 7156 3565
rect 7124 3515 7156 3516
rect 7124 3485 7125 3515
rect 7125 3485 7155 3515
rect 7155 3485 7156 3515
rect 7124 3484 7156 3485
rect 7124 3435 7156 3436
rect 7124 3405 7125 3435
rect 7125 3405 7155 3435
rect 7155 3405 7156 3435
rect 7124 3404 7156 3405
rect 7124 3355 7156 3356
rect 7124 3325 7125 3355
rect 7125 3325 7155 3355
rect 7155 3325 7156 3355
rect 7124 3324 7156 3325
rect 7124 3275 7156 3276
rect 7124 3245 7125 3275
rect 7125 3245 7155 3275
rect 7155 3245 7156 3275
rect 7124 3244 7156 3245
rect 7124 3195 7156 3196
rect 7124 3165 7125 3195
rect 7125 3165 7155 3195
rect 7155 3165 7156 3195
rect 7124 3164 7156 3165
rect 7124 3115 7156 3116
rect 7124 3085 7125 3115
rect 7125 3085 7155 3115
rect 7155 3085 7156 3115
rect 7124 3084 7156 3085
rect 7124 3035 7156 3036
rect 7124 3005 7125 3035
rect 7125 3005 7155 3035
rect 7155 3005 7156 3035
rect 7124 3004 7156 3005
rect 7124 2955 7156 2956
rect 7124 2925 7125 2955
rect 7125 2925 7155 2955
rect 7155 2925 7156 2955
rect 7124 2924 7156 2925
rect 7124 2875 7156 2876
rect 7124 2845 7125 2875
rect 7125 2845 7155 2875
rect 7155 2845 7156 2875
rect 7124 2844 7156 2845
rect 7124 2795 7156 2796
rect 7124 2765 7125 2795
rect 7125 2765 7155 2795
rect 7155 2765 7156 2795
rect 7124 2764 7156 2765
rect 7124 2715 7156 2716
rect 7124 2685 7125 2715
rect 7125 2685 7155 2715
rect 7155 2685 7156 2715
rect 7124 2684 7156 2685
rect 7124 2635 7156 2636
rect 7124 2605 7125 2635
rect 7125 2605 7155 2635
rect 7155 2605 7156 2635
rect 7124 2604 7156 2605
rect 7124 2555 7156 2556
rect 7124 2525 7125 2555
rect 7125 2525 7155 2555
rect 7155 2525 7156 2555
rect 7124 2524 7156 2525
rect 7124 2475 7156 2476
rect 7124 2445 7125 2475
rect 7125 2445 7155 2475
rect 7155 2445 7156 2475
rect 7124 2444 7156 2445
rect 7124 2395 7156 2396
rect 7124 2365 7125 2395
rect 7125 2365 7155 2395
rect 7155 2365 7156 2395
rect 7124 2364 7156 2365
rect 7124 2315 7156 2316
rect 7124 2285 7125 2315
rect 7125 2285 7155 2315
rect 7155 2285 7156 2315
rect 7124 2284 7156 2285
rect 7124 2235 7156 2236
rect 7124 2205 7125 2235
rect 7125 2205 7155 2235
rect 7155 2205 7156 2235
rect 7124 2204 7156 2205
rect 7124 2155 7156 2156
rect 7124 2125 7125 2155
rect 7125 2125 7155 2155
rect 7155 2125 7156 2155
rect 7124 2124 7156 2125
rect 7124 2075 7156 2076
rect 7124 2045 7125 2075
rect 7125 2045 7155 2075
rect 7155 2045 7156 2075
rect 7124 2044 7156 2045
rect 7124 1995 7156 1996
rect 7124 1965 7125 1995
rect 7125 1965 7155 1995
rect 7155 1965 7156 1995
rect 7124 1964 7156 1965
rect 7124 1915 7156 1916
rect 7124 1885 7125 1915
rect 7125 1885 7155 1915
rect 7155 1885 7156 1915
rect 7124 1884 7156 1885
rect 7124 1835 7156 1836
rect 7124 1805 7125 1835
rect 7125 1805 7155 1835
rect 7155 1805 7156 1835
rect 7124 1804 7156 1805
rect 7124 1755 7156 1756
rect 7124 1725 7125 1755
rect 7125 1725 7155 1755
rect 7155 1725 7156 1755
rect 7124 1724 7156 1725
rect 7124 1675 7156 1676
rect 7124 1645 7125 1675
rect 7125 1645 7155 1675
rect 7155 1645 7156 1675
rect 7124 1644 7156 1645
rect 7124 1595 7156 1596
rect 7124 1565 7125 1595
rect 7125 1565 7155 1595
rect 7155 1565 7156 1595
rect 7124 1564 7156 1565
rect 7124 1515 7156 1516
rect 7124 1485 7125 1515
rect 7125 1485 7155 1515
rect 7155 1485 7156 1515
rect 7124 1484 7156 1485
rect 7124 1435 7156 1436
rect 7124 1405 7125 1435
rect 7125 1405 7155 1435
rect 7155 1405 7156 1435
rect 7124 1404 7156 1405
rect 7124 1355 7156 1356
rect 7124 1325 7125 1355
rect 7125 1325 7155 1355
rect 7155 1325 7156 1355
rect 7124 1324 7156 1325
rect 7124 1275 7156 1276
rect 7124 1245 7125 1275
rect 7125 1245 7155 1275
rect 7155 1245 7156 1275
rect 7124 1244 7156 1245
rect 7124 1195 7156 1196
rect 7124 1165 7125 1195
rect 7125 1165 7155 1195
rect 7155 1165 7156 1195
rect 7124 1164 7156 1165
rect 7124 1115 7156 1116
rect 7124 1085 7125 1115
rect 7125 1085 7155 1115
rect 7155 1085 7156 1115
rect 7124 1084 7156 1085
rect 7124 1035 7156 1036
rect 7124 1005 7125 1035
rect 7125 1005 7155 1035
rect 7155 1005 7156 1035
rect 7124 1004 7156 1005
rect 7124 955 7156 956
rect 7124 925 7125 955
rect 7125 925 7155 955
rect 7155 925 7156 955
rect 7124 924 7156 925
rect 7124 875 7156 876
rect 7124 845 7125 875
rect 7125 845 7155 875
rect 7155 845 7156 875
rect 7124 844 7156 845
rect 7124 795 7156 796
rect 7124 765 7125 795
rect 7125 765 7155 795
rect 7155 765 7156 795
rect 7124 764 7156 765
rect 7124 715 7156 716
rect 7124 685 7125 715
rect 7125 685 7155 715
rect 7155 685 7156 715
rect 7124 684 7156 685
rect 7124 595 7156 596
rect 7124 565 7125 595
rect 7125 565 7155 595
rect 7155 565 7156 595
rect 7124 564 7156 565
rect 7124 515 7156 516
rect 7124 485 7125 515
rect 7125 485 7155 515
rect 7155 485 7156 515
rect 7124 484 7156 485
rect 7124 435 7156 436
rect 7124 405 7125 435
rect 7125 405 7155 435
rect 7155 405 7156 435
rect 7124 404 7156 405
rect 7124 355 7156 356
rect 7124 325 7125 355
rect 7125 325 7155 355
rect 7155 325 7156 355
rect 7124 324 7156 325
rect 7124 275 7156 276
rect 7124 245 7125 275
rect 7125 245 7155 275
rect 7155 245 7156 275
rect 7124 244 7156 245
rect 7124 195 7156 196
rect 7124 165 7125 195
rect 7125 165 7155 195
rect 7155 165 7156 195
rect 7124 164 7156 165
rect 7124 115 7156 116
rect 7124 85 7125 115
rect 7125 85 7155 115
rect 7155 85 7156 115
rect 7124 84 7156 85
rect 7124 35 7156 36
rect 7124 5 7125 35
rect 7125 5 7155 35
rect 7155 5 7156 35
rect 7124 4 7156 5
rect 7284 16595 7316 16596
rect 7284 16565 7285 16595
rect 7285 16565 7315 16595
rect 7315 16565 7316 16595
rect 7284 16564 7316 16565
rect 7284 16515 7316 16516
rect 7284 16485 7285 16515
rect 7285 16485 7315 16515
rect 7315 16485 7316 16515
rect 7284 16484 7316 16485
rect 7284 16435 7316 16436
rect 7284 16405 7285 16435
rect 7285 16405 7315 16435
rect 7315 16405 7316 16435
rect 7284 16404 7316 16405
rect 7284 16355 7316 16356
rect 7284 16325 7285 16355
rect 7285 16325 7315 16355
rect 7315 16325 7316 16355
rect 7284 16324 7316 16325
rect 7284 16275 7316 16276
rect 7284 16245 7285 16275
rect 7285 16245 7315 16275
rect 7315 16245 7316 16275
rect 7284 16244 7316 16245
rect 7284 16195 7316 16196
rect 7284 16165 7285 16195
rect 7285 16165 7315 16195
rect 7315 16165 7316 16195
rect 7284 16164 7316 16165
rect 7284 16115 7316 16116
rect 7284 16085 7285 16115
rect 7285 16085 7315 16115
rect 7315 16085 7316 16115
rect 7284 16084 7316 16085
rect 7284 16035 7316 16036
rect 7284 16005 7285 16035
rect 7285 16005 7315 16035
rect 7315 16005 7316 16035
rect 7284 16004 7316 16005
rect 7284 15955 7316 15956
rect 7284 15925 7285 15955
rect 7285 15925 7315 15955
rect 7315 15925 7316 15955
rect 7284 15924 7316 15925
rect 7284 15435 7316 15436
rect 7284 15405 7285 15435
rect 7285 15405 7315 15435
rect 7315 15405 7316 15435
rect 7284 15404 7316 15405
rect 7284 15355 7316 15356
rect 7284 15325 7285 15355
rect 7285 15325 7315 15355
rect 7315 15325 7316 15355
rect 7284 15324 7316 15325
rect 7284 15275 7316 15276
rect 7284 15245 7285 15275
rect 7285 15245 7315 15275
rect 7315 15245 7316 15275
rect 7284 15244 7316 15245
rect 7284 15195 7316 15196
rect 7284 15165 7285 15195
rect 7285 15165 7315 15195
rect 7315 15165 7316 15195
rect 7284 15164 7316 15165
rect 7284 15115 7316 15116
rect 7284 15085 7285 15115
rect 7285 15085 7315 15115
rect 7315 15085 7316 15115
rect 7284 15084 7316 15085
rect 7284 15035 7316 15036
rect 7284 15005 7285 15035
rect 7285 15005 7315 15035
rect 7315 15005 7316 15035
rect 7284 15004 7316 15005
rect 7284 14955 7316 14956
rect 7284 14925 7285 14955
rect 7285 14925 7315 14955
rect 7315 14925 7316 14955
rect 7284 14924 7316 14925
rect 7284 14875 7316 14876
rect 7284 14845 7285 14875
rect 7285 14845 7315 14875
rect 7315 14845 7316 14875
rect 7284 14844 7316 14845
rect 7284 14795 7316 14796
rect 7284 14765 7285 14795
rect 7285 14765 7315 14795
rect 7315 14765 7316 14795
rect 7284 14764 7316 14765
rect 7284 14715 7316 14716
rect 7284 14685 7285 14715
rect 7285 14685 7315 14715
rect 7315 14685 7316 14715
rect 7284 14684 7316 14685
rect 7284 14635 7316 14636
rect 7284 14605 7285 14635
rect 7285 14605 7315 14635
rect 7315 14605 7316 14635
rect 7284 14604 7316 14605
rect 7284 14555 7316 14556
rect 7284 14525 7285 14555
rect 7285 14525 7315 14555
rect 7315 14525 7316 14555
rect 7284 14524 7316 14525
rect 7284 14475 7316 14476
rect 7284 14445 7285 14475
rect 7285 14445 7315 14475
rect 7315 14445 7316 14475
rect 7284 14444 7316 14445
rect 7284 13995 7316 13996
rect 7284 13965 7285 13995
rect 7285 13965 7315 13995
rect 7315 13965 7316 13995
rect 7284 13964 7316 13965
rect 7284 13875 7316 13876
rect 7284 13845 7285 13875
rect 7285 13845 7315 13875
rect 7315 13845 7316 13875
rect 7284 13844 7316 13845
rect 7284 13795 7316 13796
rect 7284 13765 7285 13795
rect 7285 13765 7315 13795
rect 7315 13765 7316 13795
rect 7284 13764 7316 13765
rect 7284 13715 7316 13716
rect 7284 13685 7285 13715
rect 7285 13685 7315 13715
rect 7315 13685 7316 13715
rect 7284 13684 7316 13685
rect 7284 13635 7316 13636
rect 7284 13605 7285 13635
rect 7285 13605 7315 13635
rect 7315 13605 7316 13635
rect 7284 13604 7316 13605
rect 7284 13555 7316 13556
rect 7284 13525 7285 13555
rect 7285 13525 7315 13555
rect 7315 13525 7316 13555
rect 7284 13524 7316 13525
rect 7284 13475 7316 13476
rect 7284 13445 7285 13475
rect 7285 13445 7315 13475
rect 7315 13445 7316 13475
rect 7284 13444 7316 13445
rect 7284 13395 7316 13396
rect 7284 13365 7285 13395
rect 7285 13365 7315 13395
rect 7315 13365 7316 13395
rect 7284 13364 7316 13365
rect 7284 13315 7316 13316
rect 7284 13285 7285 13315
rect 7285 13285 7315 13315
rect 7315 13285 7316 13315
rect 7284 13284 7316 13285
rect 7284 13235 7316 13236
rect 7284 13205 7285 13235
rect 7285 13205 7315 13235
rect 7315 13205 7316 13235
rect 7284 13204 7316 13205
rect 7284 13155 7316 13156
rect 7284 13125 7285 13155
rect 7285 13125 7315 13155
rect 7315 13125 7316 13155
rect 7284 13124 7316 13125
rect 7284 13075 7316 13076
rect 7284 13045 7285 13075
rect 7285 13045 7315 13075
rect 7315 13045 7316 13075
rect 7284 13044 7316 13045
rect 7284 12995 7316 12996
rect 7284 12965 7285 12995
rect 7285 12965 7315 12995
rect 7315 12965 7316 12995
rect 7284 12964 7316 12965
rect 7284 12515 7316 12516
rect 7284 12485 7285 12515
rect 7285 12485 7315 12515
rect 7315 12485 7316 12515
rect 7284 12484 7316 12485
rect 7284 12435 7316 12436
rect 7284 12405 7285 12435
rect 7285 12405 7315 12435
rect 7315 12405 7316 12435
rect 7284 12404 7316 12405
rect 7284 12315 7316 12316
rect 7284 12285 7285 12315
rect 7285 12285 7315 12315
rect 7315 12285 7316 12315
rect 7284 12284 7316 12285
rect 7284 12235 7316 12236
rect 7284 12205 7285 12235
rect 7285 12205 7315 12235
rect 7315 12205 7316 12235
rect 7284 12204 7316 12205
rect 7284 12155 7316 12156
rect 7284 12125 7285 12155
rect 7285 12125 7315 12155
rect 7315 12125 7316 12155
rect 7284 12124 7316 12125
rect 7284 12075 7316 12076
rect 7284 12045 7285 12075
rect 7285 12045 7315 12075
rect 7315 12045 7316 12075
rect 7284 12044 7316 12045
rect 7284 11995 7316 11996
rect 7284 11965 7285 11995
rect 7285 11965 7315 11995
rect 7315 11965 7316 11995
rect 7284 11964 7316 11965
rect 7284 11915 7316 11916
rect 7284 11885 7285 11915
rect 7285 11885 7315 11915
rect 7315 11885 7316 11915
rect 7284 11884 7316 11885
rect 7284 11835 7316 11836
rect 7284 11805 7285 11835
rect 7285 11805 7315 11835
rect 7315 11805 7316 11835
rect 7284 11804 7316 11805
rect 7284 11755 7316 11756
rect 7284 11725 7285 11755
rect 7285 11725 7315 11755
rect 7315 11725 7316 11755
rect 7284 11724 7316 11725
rect 7284 11675 7316 11676
rect 7284 11645 7285 11675
rect 7285 11645 7315 11675
rect 7315 11645 7316 11675
rect 7284 11644 7316 11645
rect 7284 11595 7316 11596
rect 7284 11565 7285 11595
rect 7285 11565 7315 11595
rect 7315 11565 7316 11595
rect 7284 11564 7316 11565
rect 7284 11515 7316 11516
rect 7284 11485 7285 11515
rect 7285 11485 7315 11515
rect 7315 11485 7316 11515
rect 7284 11484 7316 11485
rect 7284 11435 7316 11436
rect 7284 11405 7285 11435
rect 7285 11405 7315 11435
rect 7315 11405 7316 11435
rect 7284 11404 7316 11405
rect 7284 11355 7316 11356
rect 7284 11325 7285 11355
rect 7285 11325 7315 11355
rect 7315 11325 7316 11355
rect 7284 11324 7316 11325
rect 7284 11195 7316 11196
rect 7284 11165 7285 11195
rect 7285 11165 7315 11195
rect 7315 11165 7316 11195
rect 7284 11164 7316 11165
rect 7284 11115 7316 11116
rect 7284 11085 7285 11115
rect 7285 11085 7315 11115
rect 7315 11085 7316 11115
rect 7284 11084 7316 11085
rect 7284 11035 7316 11036
rect 7284 11005 7285 11035
rect 7285 11005 7315 11035
rect 7315 11005 7316 11035
rect 7284 11004 7316 11005
rect 7284 10875 7316 10876
rect 7284 10845 7285 10875
rect 7285 10845 7315 10875
rect 7315 10845 7316 10875
rect 7284 10844 7316 10845
rect 7284 10795 7316 10796
rect 7284 10765 7285 10795
rect 7285 10765 7315 10795
rect 7315 10765 7316 10795
rect 7284 10764 7316 10765
rect 7284 10715 7316 10716
rect 7284 10685 7285 10715
rect 7285 10685 7315 10715
rect 7315 10685 7316 10715
rect 7284 10684 7316 10685
rect 7284 10635 7316 10636
rect 7284 10605 7285 10635
rect 7285 10605 7315 10635
rect 7315 10605 7316 10635
rect 7284 10604 7316 10605
rect 7284 10555 7316 10556
rect 7284 10525 7285 10555
rect 7285 10525 7315 10555
rect 7315 10525 7316 10555
rect 7284 10524 7316 10525
rect 7284 10475 7316 10476
rect 7284 10445 7285 10475
rect 7285 10445 7315 10475
rect 7315 10445 7316 10475
rect 7284 10444 7316 10445
rect 7284 10395 7316 10396
rect 7284 10365 7285 10395
rect 7285 10365 7315 10395
rect 7315 10365 7316 10395
rect 7284 10364 7316 10365
rect 7284 10315 7316 10316
rect 7284 10285 7285 10315
rect 7285 10285 7315 10315
rect 7315 10285 7316 10315
rect 7284 10284 7316 10285
rect 7284 10235 7316 10236
rect 7284 10205 7285 10235
rect 7285 10205 7315 10235
rect 7315 10205 7316 10235
rect 7284 10204 7316 10205
rect 7284 10155 7316 10156
rect 7284 10125 7285 10155
rect 7285 10125 7315 10155
rect 7315 10125 7316 10155
rect 7284 10124 7316 10125
rect 7284 10075 7316 10076
rect 7284 10045 7285 10075
rect 7285 10045 7315 10075
rect 7315 10045 7316 10075
rect 7284 10044 7316 10045
rect 7284 9995 7316 9996
rect 7284 9965 7285 9995
rect 7285 9965 7315 9995
rect 7315 9965 7316 9995
rect 7284 9964 7316 9965
rect 7284 9915 7316 9916
rect 7284 9885 7285 9915
rect 7285 9885 7315 9915
rect 7315 9885 7316 9915
rect 7284 9884 7316 9885
rect 7284 9835 7316 9836
rect 7284 9805 7285 9835
rect 7285 9805 7315 9835
rect 7315 9805 7316 9835
rect 7284 9804 7316 9805
rect 7284 9755 7316 9756
rect 7284 9725 7285 9755
rect 7285 9725 7315 9755
rect 7315 9725 7316 9755
rect 7284 9724 7316 9725
rect 7284 9675 7316 9676
rect 7284 9645 7285 9675
rect 7285 9645 7315 9675
rect 7315 9645 7316 9675
rect 7284 9644 7316 9645
rect 7284 9595 7316 9596
rect 7284 9565 7285 9595
rect 7285 9565 7315 9595
rect 7315 9565 7316 9595
rect 7284 9564 7316 9565
rect 7284 9515 7316 9516
rect 7284 9485 7285 9515
rect 7285 9485 7315 9515
rect 7315 9485 7316 9515
rect 7284 9484 7316 9485
rect 7284 9435 7316 9436
rect 7284 9405 7285 9435
rect 7285 9405 7315 9435
rect 7315 9405 7316 9435
rect 7284 9404 7316 9405
rect 7284 9355 7316 9356
rect 7284 9325 7285 9355
rect 7285 9325 7315 9355
rect 7315 9325 7316 9355
rect 7284 9324 7316 9325
rect 7284 9275 7316 9276
rect 7284 9245 7285 9275
rect 7285 9245 7315 9275
rect 7315 9245 7316 9275
rect 7284 9244 7316 9245
rect 7284 9115 7316 9116
rect 7284 9085 7285 9115
rect 7285 9085 7315 9115
rect 7315 9085 7316 9115
rect 7284 9084 7316 9085
rect 7284 9035 7316 9036
rect 7284 9005 7285 9035
rect 7285 9005 7315 9035
rect 7315 9005 7316 9035
rect 7284 9004 7316 9005
rect 7284 8955 7316 8956
rect 7284 8925 7285 8955
rect 7285 8925 7315 8955
rect 7315 8925 7316 8955
rect 7284 8924 7316 8925
rect 7284 8635 7316 8636
rect 7284 8605 7285 8635
rect 7285 8605 7315 8635
rect 7315 8605 7316 8635
rect 7284 8604 7316 8605
rect 7284 8555 7316 8556
rect 7284 8525 7285 8555
rect 7285 8525 7315 8555
rect 7315 8525 7316 8555
rect 7284 8524 7316 8525
rect 7284 8475 7316 8476
rect 7284 8445 7285 8475
rect 7285 8445 7315 8475
rect 7315 8445 7316 8475
rect 7284 8444 7316 8445
rect 7284 8395 7316 8396
rect 7284 8365 7285 8395
rect 7285 8365 7315 8395
rect 7315 8365 7316 8395
rect 7284 8364 7316 8365
rect 7284 8315 7316 8316
rect 7284 8285 7285 8315
rect 7285 8285 7315 8315
rect 7315 8285 7316 8315
rect 7284 8284 7316 8285
rect 7284 8235 7316 8236
rect 7284 8205 7285 8235
rect 7285 8205 7315 8235
rect 7315 8205 7316 8235
rect 7284 8204 7316 8205
rect 7284 8155 7316 8156
rect 7284 8125 7285 8155
rect 7285 8125 7315 8155
rect 7315 8125 7316 8155
rect 7284 8124 7316 8125
rect 7284 8075 7316 8076
rect 7284 8045 7285 8075
rect 7285 8045 7315 8075
rect 7315 8045 7316 8075
rect 7284 8044 7316 8045
rect 7284 7995 7316 7996
rect 7284 7965 7285 7995
rect 7285 7965 7315 7995
rect 7315 7965 7316 7995
rect 7284 7964 7316 7965
rect 7284 7915 7316 7916
rect 7284 7885 7285 7915
rect 7285 7885 7315 7915
rect 7315 7885 7316 7915
rect 7284 7884 7316 7885
rect 7284 7835 7316 7836
rect 7284 7805 7285 7835
rect 7285 7805 7315 7835
rect 7315 7805 7316 7835
rect 7284 7804 7316 7805
rect 7284 7755 7316 7756
rect 7284 7725 7285 7755
rect 7285 7725 7315 7755
rect 7315 7725 7316 7755
rect 7284 7724 7316 7725
rect 7284 7675 7316 7676
rect 7284 7645 7285 7675
rect 7285 7645 7315 7675
rect 7315 7645 7316 7675
rect 7284 7644 7316 7645
rect 7284 7595 7316 7596
rect 7284 7565 7285 7595
rect 7285 7565 7315 7595
rect 7315 7565 7316 7595
rect 7284 7564 7316 7565
rect 7284 7515 7316 7516
rect 7284 7485 7285 7515
rect 7285 7485 7315 7515
rect 7315 7485 7316 7515
rect 7284 7484 7316 7485
rect 7284 7435 7316 7436
rect 7284 7405 7285 7435
rect 7285 7405 7315 7435
rect 7315 7405 7316 7435
rect 7284 7404 7316 7405
rect 7284 7355 7316 7356
rect 7284 7325 7285 7355
rect 7285 7325 7315 7355
rect 7315 7325 7316 7355
rect 7284 7324 7316 7325
rect 7284 7275 7316 7276
rect 7284 7245 7285 7275
rect 7285 7245 7315 7275
rect 7315 7245 7316 7275
rect 7284 7244 7316 7245
rect 7284 7195 7316 7196
rect 7284 7165 7285 7195
rect 7285 7165 7315 7195
rect 7315 7165 7316 7195
rect 7284 7164 7316 7165
rect 7284 7115 7316 7116
rect 7284 7085 7285 7115
rect 7285 7085 7315 7115
rect 7315 7085 7316 7115
rect 7284 7084 7316 7085
rect 7284 7035 7316 7036
rect 7284 7005 7285 7035
rect 7285 7005 7315 7035
rect 7315 7005 7316 7035
rect 7284 7004 7316 7005
rect 7284 6955 7316 6956
rect 7284 6925 7285 6955
rect 7285 6925 7315 6955
rect 7315 6925 7316 6955
rect 7284 6924 7316 6925
rect 7284 6875 7316 6876
rect 7284 6845 7285 6875
rect 7285 6845 7315 6875
rect 7315 6845 7316 6875
rect 7284 6844 7316 6845
rect 7284 6795 7316 6796
rect 7284 6765 7285 6795
rect 7285 6765 7315 6795
rect 7315 6765 7316 6795
rect 7284 6764 7316 6765
rect 7284 6715 7316 6716
rect 7284 6685 7285 6715
rect 7285 6685 7315 6715
rect 7315 6685 7316 6715
rect 7284 6684 7316 6685
rect 7284 6635 7316 6636
rect 7284 6605 7285 6635
rect 7285 6605 7315 6635
rect 7315 6605 7316 6635
rect 7284 6604 7316 6605
rect 7284 6555 7316 6556
rect 7284 6525 7285 6555
rect 7285 6525 7315 6555
rect 7315 6525 7316 6555
rect 7284 6524 7316 6525
rect 7284 6475 7316 6476
rect 7284 6445 7285 6475
rect 7285 6445 7315 6475
rect 7315 6445 7316 6475
rect 7284 6444 7316 6445
rect 7284 6395 7316 6396
rect 7284 6365 7285 6395
rect 7285 6365 7315 6395
rect 7315 6365 7316 6395
rect 7284 6364 7316 6365
rect 7284 6315 7316 6316
rect 7284 6285 7285 6315
rect 7285 6285 7315 6315
rect 7315 6285 7316 6315
rect 7284 6284 7316 6285
rect 7284 6235 7316 6236
rect 7284 6205 7285 6235
rect 7285 6205 7315 6235
rect 7315 6205 7316 6235
rect 7284 6204 7316 6205
rect 7284 6155 7316 6156
rect 7284 6125 7285 6155
rect 7285 6125 7315 6155
rect 7315 6125 7316 6155
rect 7284 6124 7316 6125
rect 7284 6075 7316 6076
rect 7284 6045 7285 6075
rect 7285 6045 7315 6075
rect 7315 6045 7316 6075
rect 7284 6044 7316 6045
rect 7284 5995 7316 5996
rect 7284 5965 7285 5995
rect 7285 5965 7315 5995
rect 7315 5965 7316 5995
rect 7284 5964 7316 5965
rect 7284 5915 7316 5916
rect 7284 5885 7285 5915
rect 7285 5885 7315 5915
rect 7315 5885 7316 5915
rect 7284 5884 7316 5885
rect 7284 5835 7316 5836
rect 7284 5805 7285 5835
rect 7285 5805 7315 5835
rect 7315 5805 7316 5835
rect 7284 5804 7316 5805
rect 7284 5755 7316 5756
rect 7284 5725 7285 5755
rect 7285 5725 7315 5755
rect 7315 5725 7316 5755
rect 7284 5724 7316 5725
rect 7284 5675 7316 5676
rect 7284 5645 7285 5675
rect 7285 5645 7315 5675
rect 7315 5645 7316 5675
rect 7284 5644 7316 5645
rect 7284 5595 7316 5596
rect 7284 5565 7285 5595
rect 7285 5565 7315 5595
rect 7315 5565 7316 5595
rect 7284 5564 7316 5565
rect 7284 5515 7316 5516
rect 7284 5485 7285 5515
rect 7285 5485 7315 5515
rect 7315 5485 7316 5515
rect 7284 5484 7316 5485
rect 7284 5435 7316 5436
rect 7284 5405 7285 5435
rect 7285 5405 7315 5435
rect 7315 5405 7316 5435
rect 7284 5404 7316 5405
rect 7284 5355 7316 5356
rect 7284 5325 7285 5355
rect 7285 5325 7315 5355
rect 7315 5325 7316 5355
rect 7284 5324 7316 5325
rect 7284 5275 7316 5276
rect 7284 5245 7285 5275
rect 7285 5245 7315 5275
rect 7315 5245 7316 5275
rect 7284 5244 7316 5245
rect 7284 5195 7316 5196
rect 7284 5165 7285 5195
rect 7285 5165 7315 5195
rect 7315 5165 7316 5195
rect 7284 5164 7316 5165
rect 7284 5115 7316 5116
rect 7284 5085 7285 5115
rect 7285 5085 7315 5115
rect 7315 5085 7316 5115
rect 7284 5084 7316 5085
rect 7284 5035 7316 5036
rect 7284 5005 7285 5035
rect 7285 5005 7315 5035
rect 7315 5005 7316 5035
rect 7284 5004 7316 5005
rect 7284 4955 7316 4956
rect 7284 4925 7285 4955
rect 7285 4925 7315 4955
rect 7315 4925 7316 4955
rect 7284 4924 7316 4925
rect 7284 4875 7316 4876
rect 7284 4845 7285 4875
rect 7285 4845 7315 4875
rect 7315 4845 7316 4875
rect 7284 4844 7316 4845
rect 7284 4795 7316 4796
rect 7284 4765 7285 4795
rect 7285 4765 7315 4795
rect 7315 4765 7316 4795
rect 7284 4764 7316 4765
rect 7284 4715 7316 4716
rect 7284 4685 7285 4715
rect 7285 4685 7315 4715
rect 7315 4685 7316 4715
rect 7284 4684 7316 4685
rect 7284 4635 7316 4636
rect 7284 4605 7285 4635
rect 7285 4605 7315 4635
rect 7315 4605 7316 4635
rect 7284 4604 7316 4605
rect 7284 4555 7316 4556
rect 7284 4525 7285 4555
rect 7285 4525 7315 4555
rect 7315 4525 7316 4555
rect 7284 4524 7316 4525
rect 7284 4475 7316 4476
rect 7284 4445 7285 4475
rect 7285 4445 7315 4475
rect 7315 4445 7316 4475
rect 7284 4444 7316 4445
rect 7284 4395 7316 4396
rect 7284 4365 7285 4395
rect 7285 4365 7315 4395
rect 7315 4365 7316 4395
rect 7284 4364 7316 4365
rect 7284 4315 7316 4316
rect 7284 4285 7285 4315
rect 7285 4285 7315 4315
rect 7315 4285 7316 4315
rect 7284 4284 7316 4285
rect 7284 4235 7316 4236
rect 7284 4205 7285 4235
rect 7285 4205 7315 4235
rect 7315 4205 7316 4235
rect 7284 4204 7316 4205
rect 7284 4155 7316 4156
rect 7284 4125 7285 4155
rect 7285 4125 7315 4155
rect 7315 4125 7316 4155
rect 7284 4124 7316 4125
rect 7284 4075 7316 4076
rect 7284 4045 7285 4075
rect 7285 4045 7315 4075
rect 7315 4045 7316 4075
rect 7284 4044 7316 4045
rect 7284 3995 7316 3996
rect 7284 3965 7285 3995
rect 7285 3965 7315 3995
rect 7315 3965 7316 3995
rect 7284 3964 7316 3965
rect 7284 3915 7316 3916
rect 7284 3885 7285 3915
rect 7285 3885 7315 3915
rect 7315 3885 7316 3915
rect 7284 3884 7316 3885
rect 7284 3835 7316 3836
rect 7284 3805 7285 3835
rect 7285 3805 7315 3835
rect 7315 3805 7316 3835
rect 7284 3804 7316 3805
rect 7284 3755 7316 3756
rect 7284 3725 7285 3755
rect 7285 3725 7315 3755
rect 7315 3725 7316 3755
rect 7284 3724 7316 3725
rect 7284 3675 7316 3676
rect 7284 3645 7285 3675
rect 7285 3645 7315 3675
rect 7315 3645 7316 3675
rect 7284 3644 7316 3645
rect 7284 3595 7316 3596
rect 7284 3565 7285 3595
rect 7285 3565 7315 3595
rect 7315 3565 7316 3595
rect 7284 3564 7316 3565
rect 7284 3515 7316 3516
rect 7284 3485 7285 3515
rect 7285 3485 7315 3515
rect 7315 3485 7316 3515
rect 7284 3484 7316 3485
rect 7284 3435 7316 3436
rect 7284 3405 7285 3435
rect 7285 3405 7315 3435
rect 7315 3405 7316 3435
rect 7284 3404 7316 3405
rect 7284 3355 7316 3356
rect 7284 3325 7285 3355
rect 7285 3325 7315 3355
rect 7315 3325 7316 3355
rect 7284 3324 7316 3325
rect 7284 3275 7316 3276
rect 7284 3245 7285 3275
rect 7285 3245 7315 3275
rect 7315 3245 7316 3275
rect 7284 3244 7316 3245
rect 7284 3195 7316 3196
rect 7284 3165 7285 3195
rect 7285 3165 7315 3195
rect 7315 3165 7316 3195
rect 7284 3164 7316 3165
rect 7284 3115 7316 3116
rect 7284 3085 7285 3115
rect 7285 3085 7315 3115
rect 7315 3085 7316 3115
rect 7284 3084 7316 3085
rect 7284 3035 7316 3036
rect 7284 3005 7285 3035
rect 7285 3005 7315 3035
rect 7315 3005 7316 3035
rect 7284 3004 7316 3005
rect 7284 2955 7316 2956
rect 7284 2925 7285 2955
rect 7285 2925 7315 2955
rect 7315 2925 7316 2955
rect 7284 2924 7316 2925
rect 7284 2875 7316 2876
rect 7284 2845 7285 2875
rect 7285 2845 7315 2875
rect 7315 2845 7316 2875
rect 7284 2844 7316 2845
rect 7284 2795 7316 2796
rect 7284 2765 7285 2795
rect 7285 2765 7315 2795
rect 7315 2765 7316 2795
rect 7284 2764 7316 2765
rect 7284 2715 7316 2716
rect 7284 2685 7285 2715
rect 7285 2685 7315 2715
rect 7315 2685 7316 2715
rect 7284 2684 7316 2685
rect 7284 2635 7316 2636
rect 7284 2605 7285 2635
rect 7285 2605 7315 2635
rect 7315 2605 7316 2635
rect 7284 2604 7316 2605
rect 7284 2555 7316 2556
rect 7284 2525 7285 2555
rect 7285 2525 7315 2555
rect 7315 2525 7316 2555
rect 7284 2524 7316 2525
rect 7284 2475 7316 2476
rect 7284 2445 7285 2475
rect 7285 2445 7315 2475
rect 7315 2445 7316 2475
rect 7284 2444 7316 2445
rect 7284 2395 7316 2396
rect 7284 2365 7285 2395
rect 7285 2365 7315 2395
rect 7315 2365 7316 2395
rect 7284 2364 7316 2365
rect 7284 2315 7316 2316
rect 7284 2285 7285 2315
rect 7285 2285 7315 2315
rect 7315 2285 7316 2315
rect 7284 2284 7316 2285
rect 7284 2235 7316 2236
rect 7284 2205 7285 2235
rect 7285 2205 7315 2235
rect 7315 2205 7316 2235
rect 7284 2204 7316 2205
rect 7284 2155 7316 2156
rect 7284 2125 7285 2155
rect 7285 2125 7315 2155
rect 7315 2125 7316 2155
rect 7284 2124 7316 2125
rect 7284 2075 7316 2076
rect 7284 2045 7285 2075
rect 7285 2045 7315 2075
rect 7315 2045 7316 2075
rect 7284 2044 7316 2045
rect 7284 1995 7316 1996
rect 7284 1965 7285 1995
rect 7285 1965 7315 1995
rect 7315 1965 7316 1995
rect 7284 1964 7316 1965
rect 7284 1915 7316 1916
rect 7284 1885 7285 1915
rect 7285 1885 7315 1915
rect 7315 1885 7316 1915
rect 7284 1884 7316 1885
rect 7284 1835 7316 1836
rect 7284 1805 7285 1835
rect 7285 1805 7315 1835
rect 7315 1805 7316 1835
rect 7284 1804 7316 1805
rect 7284 1755 7316 1756
rect 7284 1725 7285 1755
rect 7285 1725 7315 1755
rect 7315 1725 7316 1755
rect 7284 1724 7316 1725
rect 7284 1675 7316 1676
rect 7284 1645 7285 1675
rect 7285 1645 7315 1675
rect 7315 1645 7316 1675
rect 7284 1644 7316 1645
rect 7284 1595 7316 1596
rect 7284 1565 7285 1595
rect 7285 1565 7315 1595
rect 7315 1565 7316 1595
rect 7284 1564 7316 1565
rect 7284 1515 7316 1516
rect 7284 1485 7285 1515
rect 7285 1485 7315 1515
rect 7315 1485 7316 1515
rect 7284 1484 7316 1485
rect 7284 1435 7316 1436
rect 7284 1405 7285 1435
rect 7285 1405 7315 1435
rect 7315 1405 7316 1435
rect 7284 1404 7316 1405
rect 7284 1355 7316 1356
rect 7284 1325 7285 1355
rect 7285 1325 7315 1355
rect 7315 1325 7316 1355
rect 7284 1324 7316 1325
rect 7284 1275 7316 1276
rect 7284 1245 7285 1275
rect 7285 1245 7315 1275
rect 7315 1245 7316 1275
rect 7284 1244 7316 1245
rect 7284 1195 7316 1196
rect 7284 1165 7285 1195
rect 7285 1165 7315 1195
rect 7315 1165 7316 1195
rect 7284 1164 7316 1165
rect 7284 1115 7316 1116
rect 7284 1085 7285 1115
rect 7285 1085 7315 1115
rect 7315 1085 7316 1115
rect 7284 1084 7316 1085
rect 7284 1035 7316 1036
rect 7284 1005 7285 1035
rect 7285 1005 7315 1035
rect 7315 1005 7316 1035
rect 7284 1004 7316 1005
rect 7284 955 7316 956
rect 7284 925 7285 955
rect 7285 925 7315 955
rect 7315 925 7316 955
rect 7284 924 7316 925
rect 7284 875 7316 876
rect 7284 845 7285 875
rect 7285 845 7315 875
rect 7315 845 7316 875
rect 7284 844 7316 845
rect 7284 795 7316 796
rect 7284 765 7285 795
rect 7285 765 7315 795
rect 7315 765 7316 795
rect 7284 764 7316 765
rect 7284 715 7316 716
rect 7284 685 7285 715
rect 7285 685 7315 715
rect 7315 685 7316 715
rect 7284 684 7316 685
rect 7284 595 7316 596
rect 7284 565 7285 595
rect 7285 565 7315 595
rect 7315 565 7316 595
rect 7284 564 7316 565
rect 7284 515 7316 516
rect 7284 485 7285 515
rect 7285 485 7315 515
rect 7315 485 7316 515
rect 7284 484 7316 485
rect 7284 435 7316 436
rect 7284 405 7285 435
rect 7285 405 7315 435
rect 7315 405 7316 435
rect 7284 404 7316 405
rect 7284 355 7316 356
rect 7284 325 7285 355
rect 7285 325 7315 355
rect 7315 325 7316 355
rect 7284 324 7316 325
rect 7284 275 7316 276
rect 7284 245 7285 275
rect 7285 245 7315 275
rect 7315 245 7316 275
rect 7284 244 7316 245
rect 7284 195 7316 196
rect 7284 165 7285 195
rect 7285 165 7315 195
rect 7315 165 7316 195
rect 7284 164 7316 165
rect 7284 115 7316 116
rect 7284 85 7285 115
rect 7285 85 7315 115
rect 7315 85 7316 115
rect 7284 84 7316 85
rect 7284 35 7316 36
rect 7284 5 7285 35
rect 7285 5 7315 35
rect 7315 5 7316 35
rect 7284 4 7316 5
rect 7524 19684 7556 19716
rect 7364 18484 7396 18516
rect 7364 18404 7396 18436
rect 7364 16595 7396 16596
rect 7364 16565 7365 16595
rect 7365 16565 7395 16595
rect 7395 16565 7396 16595
rect 7364 16564 7396 16565
rect 7364 16515 7396 16516
rect 7364 16485 7365 16515
rect 7365 16485 7395 16515
rect 7395 16485 7396 16515
rect 7364 16484 7396 16485
rect 7364 16435 7396 16436
rect 7364 16405 7365 16435
rect 7365 16405 7395 16435
rect 7395 16405 7396 16435
rect 7364 16404 7396 16405
rect 7364 16355 7396 16356
rect 7364 16325 7365 16355
rect 7365 16325 7395 16355
rect 7395 16325 7396 16355
rect 7364 16324 7396 16325
rect 7364 16275 7396 16276
rect 7364 16245 7365 16275
rect 7365 16245 7395 16275
rect 7395 16245 7396 16275
rect 7364 16244 7396 16245
rect 7364 16195 7396 16196
rect 7364 16165 7365 16195
rect 7365 16165 7395 16195
rect 7395 16165 7396 16195
rect 7364 16164 7396 16165
rect 7364 16115 7396 16116
rect 7364 16085 7365 16115
rect 7365 16085 7395 16115
rect 7395 16085 7396 16115
rect 7364 16084 7396 16085
rect 7364 16035 7396 16036
rect 7364 16005 7365 16035
rect 7365 16005 7395 16035
rect 7395 16005 7396 16035
rect 7364 16004 7396 16005
rect 7364 15955 7396 15956
rect 7364 15925 7365 15955
rect 7365 15925 7395 15955
rect 7395 15925 7396 15955
rect 7364 15924 7396 15925
rect 7364 15435 7396 15436
rect 7364 15405 7365 15435
rect 7365 15405 7395 15435
rect 7395 15405 7396 15435
rect 7364 15404 7396 15405
rect 7364 15355 7396 15356
rect 7364 15325 7365 15355
rect 7365 15325 7395 15355
rect 7395 15325 7396 15355
rect 7364 15324 7396 15325
rect 7364 15275 7396 15276
rect 7364 15245 7365 15275
rect 7365 15245 7395 15275
rect 7395 15245 7396 15275
rect 7364 15244 7396 15245
rect 7364 15195 7396 15196
rect 7364 15165 7365 15195
rect 7365 15165 7395 15195
rect 7395 15165 7396 15195
rect 7364 15164 7396 15165
rect 7364 15115 7396 15116
rect 7364 15085 7365 15115
rect 7365 15085 7395 15115
rect 7395 15085 7396 15115
rect 7364 15084 7396 15085
rect 7364 15035 7396 15036
rect 7364 15005 7365 15035
rect 7365 15005 7395 15035
rect 7395 15005 7396 15035
rect 7364 15004 7396 15005
rect 7364 14955 7396 14956
rect 7364 14925 7365 14955
rect 7365 14925 7395 14955
rect 7395 14925 7396 14955
rect 7364 14924 7396 14925
rect 7364 14875 7396 14876
rect 7364 14845 7365 14875
rect 7365 14845 7395 14875
rect 7395 14845 7396 14875
rect 7364 14844 7396 14845
rect 7364 14795 7396 14796
rect 7364 14765 7365 14795
rect 7365 14765 7395 14795
rect 7395 14765 7396 14795
rect 7364 14764 7396 14765
rect 7364 14715 7396 14716
rect 7364 14685 7365 14715
rect 7365 14685 7395 14715
rect 7395 14685 7396 14715
rect 7364 14684 7396 14685
rect 7364 14635 7396 14636
rect 7364 14605 7365 14635
rect 7365 14605 7395 14635
rect 7395 14605 7396 14635
rect 7364 14604 7396 14605
rect 7364 14555 7396 14556
rect 7364 14525 7365 14555
rect 7365 14525 7395 14555
rect 7395 14525 7396 14555
rect 7364 14524 7396 14525
rect 7364 14475 7396 14476
rect 7364 14445 7365 14475
rect 7365 14445 7395 14475
rect 7395 14445 7396 14475
rect 7364 14444 7396 14445
rect 7364 14395 7396 14396
rect 7364 14365 7365 14395
rect 7365 14365 7395 14395
rect 7395 14365 7396 14395
rect 7364 14364 7396 14365
rect 7364 14315 7396 14316
rect 7364 14285 7365 14315
rect 7365 14285 7395 14315
rect 7395 14285 7396 14315
rect 7364 14284 7396 14285
rect 7364 14235 7396 14236
rect 7364 14205 7365 14235
rect 7365 14205 7395 14235
rect 7395 14205 7396 14235
rect 7364 14204 7396 14205
rect 7364 14155 7396 14156
rect 7364 14125 7365 14155
rect 7365 14125 7395 14155
rect 7395 14125 7396 14155
rect 7364 14124 7396 14125
rect 7364 14075 7396 14076
rect 7364 14045 7365 14075
rect 7365 14045 7395 14075
rect 7395 14045 7396 14075
rect 7364 14044 7396 14045
rect 7364 13995 7396 13996
rect 7364 13965 7365 13995
rect 7365 13965 7395 13995
rect 7395 13965 7396 13995
rect 7364 13964 7396 13965
rect 7364 13875 7396 13876
rect 7364 13845 7365 13875
rect 7365 13845 7395 13875
rect 7395 13845 7396 13875
rect 7364 13844 7396 13845
rect 7364 13795 7396 13796
rect 7364 13765 7365 13795
rect 7365 13765 7395 13795
rect 7395 13765 7396 13795
rect 7364 13764 7396 13765
rect 7364 13715 7396 13716
rect 7364 13685 7365 13715
rect 7365 13685 7395 13715
rect 7395 13685 7396 13715
rect 7364 13684 7396 13685
rect 7364 13635 7396 13636
rect 7364 13605 7365 13635
rect 7365 13605 7395 13635
rect 7395 13605 7396 13635
rect 7364 13604 7396 13605
rect 7364 13555 7396 13556
rect 7364 13525 7365 13555
rect 7365 13525 7395 13555
rect 7395 13525 7396 13555
rect 7364 13524 7396 13525
rect 7364 13475 7396 13476
rect 7364 13445 7365 13475
rect 7365 13445 7395 13475
rect 7395 13445 7396 13475
rect 7364 13444 7396 13445
rect 7364 13395 7396 13396
rect 7364 13365 7365 13395
rect 7365 13365 7395 13395
rect 7395 13365 7396 13395
rect 7364 13364 7396 13365
rect 7364 13315 7396 13316
rect 7364 13285 7365 13315
rect 7365 13285 7395 13315
rect 7395 13285 7396 13315
rect 7364 13284 7396 13285
rect 7364 13235 7396 13236
rect 7364 13205 7365 13235
rect 7365 13205 7395 13235
rect 7395 13205 7396 13235
rect 7364 13204 7396 13205
rect 7364 13155 7396 13156
rect 7364 13125 7365 13155
rect 7365 13125 7395 13155
rect 7395 13125 7396 13155
rect 7364 13124 7396 13125
rect 7364 13075 7396 13076
rect 7364 13045 7365 13075
rect 7365 13045 7395 13075
rect 7395 13045 7396 13075
rect 7364 13044 7396 13045
rect 7364 12995 7396 12996
rect 7364 12965 7365 12995
rect 7365 12965 7395 12995
rect 7395 12965 7396 12995
rect 7364 12964 7396 12965
rect 7364 12475 7396 12476
rect 7364 12445 7365 12475
rect 7365 12445 7395 12475
rect 7395 12445 7396 12475
rect 7364 12444 7396 12445
rect 7364 12395 7396 12396
rect 7364 12365 7365 12395
rect 7365 12365 7395 12395
rect 7395 12365 7396 12395
rect 7364 12364 7396 12365
rect 7364 12315 7396 12316
rect 7364 12285 7365 12315
rect 7365 12285 7395 12315
rect 7395 12285 7396 12315
rect 7364 12284 7396 12285
rect 7364 12235 7396 12236
rect 7364 12205 7365 12235
rect 7365 12205 7395 12235
rect 7395 12205 7396 12235
rect 7364 12204 7396 12205
rect 7364 12155 7396 12156
rect 7364 12125 7365 12155
rect 7365 12125 7395 12155
rect 7395 12125 7396 12155
rect 7364 12124 7396 12125
rect 7364 12075 7396 12076
rect 7364 12045 7365 12075
rect 7365 12045 7395 12075
rect 7395 12045 7396 12075
rect 7364 12044 7396 12045
rect 7364 11995 7396 11996
rect 7364 11965 7365 11995
rect 7365 11965 7395 11995
rect 7395 11965 7396 11995
rect 7364 11964 7396 11965
rect 7364 11915 7396 11916
rect 7364 11885 7365 11915
rect 7365 11885 7395 11915
rect 7395 11885 7396 11915
rect 7364 11884 7396 11885
rect 7364 11835 7396 11836
rect 7364 11805 7365 11835
rect 7365 11805 7395 11835
rect 7395 11805 7396 11835
rect 7364 11804 7396 11805
rect 7364 11755 7396 11756
rect 7364 11725 7365 11755
rect 7365 11725 7395 11755
rect 7395 11725 7396 11755
rect 7364 11724 7396 11725
rect 7364 11675 7396 11676
rect 7364 11645 7365 11675
rect 7365 11645 7395 11675
rect 7395 11645 7396 11675
rect 7364 11644 7396 11645
rect 7364 11595 7396 11596
rect 7364 11565 7365 11595
rect 7365 11565 7395 11595
rect 7395 11565 7396 11595
rect 7364 11564 7396 11565
rect 7364 11515 7396 11516
rect 7364 11485 7365 11515
rect 7365 11485 7395 11515
rect 7395 11485 7396 11515
rect 7364 11484 7396 11485
rect 7364 11435 7396 11436
rect 7364 11405 7365 11435
rect 7365 11405 7395 11435
rect 7395 11405 7396 11435
rect 7364 11404 7396 11405
rect 7364 11355 7396 11356
rect 7364 11325 7365 11355
rect 7365 11325 7395 11355
rect 7395 11325 7396 11355
rect 7364 11324 7396 11325
rect 7364 11275 7396 11276
rect 7364 11245 7365 11275
rect 7365 11245 7395 11275
rect 7395 11245 7396 11275
rect 7364 11244 7396 11245
rect 7364 11195 7396 11196
rect 7364 11165 7365 11195
rect 7365 11165 7395 11195
rect 7395 11165 7396 11195
rect 7364 11164 7396 11165
rect 7364 11115 7396 11116
rect 7364 11085 7365 11115
rect 7365 11085 7395 11115
rect 7395 11085 7396 11115
rect 7364 11084 7396 11085
rect 7364 11035 7396 11036
rect 7364 11005 7365 11035
rect 7365 11005 7395 11035
rect 7395 11005 7396 11035
rect 7364 11004 7396 11005
rect 7364 10955 7396 10956
rect 7364 10925 7365 10955
rect 7365 10925 7395 10955
rect 7395 10925 7396 10955
rect 7364 10924 7396 10925
rect 7364 10875 7396 10876
rect 7364 10845 7365 10875
rect 7365 10845 7395 10875
rect 7395 10845 7396 10875
rect 7364 10844 7396 10845
rect 7364 10795 7396 10796
rect 7364 10765 7365 10795
rect 7365 10765 7395 10795
rect 7395 10765 7396 10795
rect 7364 10764 7396 10765
rect 7364 10715 7396 10716
rect 7364 10685 7365 10715
rect 7365 10685 7395 10715
rect 7395 10685 7396 10715
rect 7364 10684 7396 10685
rect 7364 10635 7396 10636
rect 7364 10605 7365 10635
rect 7365 10605 7395 10635
rect 7395 10605 7396 10635
rect 7364 10604 7396 10605
rect 7364 10555 7396 10556
rect 7364 10525 7365 10555
rect 7365 10525 7395 10555
rect 7395 10525 7396 10555
rect 7364 10524 7396 10525
rect 7364 10475 7396 10476
rect 7364 10445 7365 10475
rect 7365 10445 7395 10475
rect 7395 10445 7396 10475
rect 7364 10444 7396 10445
rect 7364 10395 7396 10396
rect 7364 10365 7365 10395
rect 7365 10365 7395 10395
rect 7395 10365 7396 10395
rect 7364 10364 7396 10365
rect 7364 10315 7396 10316
rect 7364 10285 7365 10315
rect 7365 10285 7395 10315
rect 7395 10285 7396 10315
rect 7364 10284 7396 10285
rect 7364 10235 7396 10236
rect 7364 10205 7365 10235
rect 7365 10205 7395 10235
rect 7395 10205 7396 10235
rect 7364 10204 7396 10205
rect 7364 10155 7396 10156
rect 7364 10125 7365 10155
rect 7365 10125 7395 10155
rect 7395 10125 7396 10155
rect 7364 10124 7396 10125
rect 7364 10075 7396 10076
rect 7364 10045 7365 10075
rect 7365 10045 7395 10075
rect 7395 10045 7396 10075
rect 7364 10044 7396 10045
rect 7364 9995 7396 9996
rect 7364 9965 7365 9995
rect 7365 9965 7395 9995
rect 7395 9965 7396 9995
rect 7364 9964 7396 9965
rect 7364 9915 7396 9916
rect 7364 9885 7365 9915
rect 7365 9885 7395 9915
rect 7395 9885 7396 9915
rect 7364 9884 7396 9885
rect 7364 9835 7396 9836
rect 7364 9805 7365 9835
rect 7365 9805 7395 9835
rect 7395 9805 7396 9835
rect 7364 9804 7396 9805
rect 7364 9755 7396 9756
rect 7364 9725 7365 9755
rect 7365 9725 7395 9755
rect 7395 9725 7396 9755
rect 7364 9724 7396 9725
rect 7364 9675 7396 9676
rect 7364 9645 7365 9675
rect 7365 9645 7395 9675
rect 7395 9645 7396 9675
rect 7364 9644 7396 9645
rect 7364 9595 7396 9596
rect 7364 9565 7365 9595
rect 7365 9565 7395 9595
rect 7395 9565 7396 9595
rect 7364 9564 7396 9565
rect 7364 9515 7396 9516
rect 7364 9485 7365 9515
rect 7365 9485 7395 9515
rect 7395 9485 7396 9515
rect 7364 9484 7396 9485
rect 7364 9435 7396 9436
rect 7364 9405 7365 9435
rect 7365 9405 7395 9435
rect 7395 9405 7396 9435
rect 7364 9404 7396 9405
rect 7364 9355 7396 9356
rect 7364 9325 7365 9355
rect 7365 9325 7395 9355
rect 7395 9325 7396 9355
rect 7364 9324 7396 9325
rect 7364 9275 7396 9276
rect 7364 9245 7365 9275
rect 7365 9245 7395 9275
rect 7395 9245 7396 9275
rect 7364 9244 7396 9245
rect 7364 9195 7396 9196
rect 7364 9165 7365 9195
rect 7365 9165 7395 9195
rect 7395 9165 7396 9195
rect 7364 9164 7396 9165
rect 7364 9115 7396 9116
rect 7364 9085 7365 9115
rect 7365 9085 7395 9115
rect 7395 9085 7396 9115
rect 7364 9084 7396 9085
rect 7364 9035 7396 9036
rect 7364 9005 7365 9035
rect 7365 9005 7395 9035
rect 7395 9005 7396 9035
rect 7364 9004 7396 9005
rect 7364 8955 7396 8956
rect 7364 8925 7365 8955
rect 7365 8925 7395 8955
rect 7395 8925 7396 8955
rect 7364 8924 7396 8925
rect 7364 8635 7396 8636
rect 7364 8605 7365 8635
rect 7365 8605 7395 8635
rect 7395 8605 7396 8635
rect 7364 8604 7396 8605
rect 7364 8555 7396 8556
rect 7364 8525 7365 8555
rect 7365 8525 7395 8555
rect 7395 8525 7396 8555
rect 7364 8524 7396 8525
rect 7364 8475 7396 8476
rect 7364 8445 7365 8475
rect 7365 8445 7395 8475
rect 7395 8445 7396 8475
rect 7364 8444 7396 8445
rect 7364 8395 7396 8396
rect 7364 8365 7365 8395
rect 7365 8365 7395 8395
rect 7395 8365 7396 8395
rect 7364 8364 7396 8365
rect 7364 8315 7396 8316
rect 7364 8285 7365 8315
rect 7365 8285 7395 8315
rect 7395 8285 7396 8315
rect 7364 8284 7396 8285
rect 7364 8235 7396 8236
rect 7364 8205 7365 8235
rect 7365 8205 7395 8235
rect 7395 8205 7396 8235
rect 7364 8204 7396 8205
rect 7364 8155 7396 8156
rect 7364 8125 7365 8155
rect 7365 8125 7395 8155
rect 7395 8125 7396 8155
rect 7364 8124 7396 8125
rect 7364 8075 7396 8076
rect 7364 8045 7365 8075
rect 7365 8045 7395 8075
rect 7395 8045 7396 8075
rect 7364 8044 7396 8045
rect 7364 7995 7396 7996
rect 7364 7965 7365 7995
rect 7365 7965 7395 7995
rect 7395 7965 7396 7995
rect 7364 7964 7396 7965
rect 7364 7915 7396 7916
rect 7364 7885 7365 7915
rect 7365 7885 7395 7915
rect 7395 7885 7396 7915
rect 7364 7884 7396 7885
rect 7364 7835 7396 7836
rect 7364 7805 7365 7835
rect 7365 7805 7395 7835
rect 7395 7805 7396 7835
rect 7364 7804 7396 7805
rect 7364 7755 7396 7756
rect 7364 7725 7365 7755
rect 7365 7725 7395 7755
rect 7395 7725 7396 7755
rect 7364 7724 7396 7725
rect 7364 7675 7396 7676
rect 7364 7645 7365 7675
rect 7365 7645 7395 7675
rect 7395 7645 7396 7675
rect 7364 7644 7396 7645
rect 7364 7595 7396 7596
rect 7364 7565 7365 7595
rect 7365 7565 7395 7595
rect 7395 7565 7396 7595
rect 7364 7564 7396 7565
rect 7364 7515 7396 7516
rect 7364 7485 7365 7515
rect 7365 7485 7395 7515
rect 7395 7485 7396 7515
rect 7364 7484 7396 7485
rect 7364 7435 7396 7436
rect 7364 7405 7365 7435
rect 7365 7405 7395 7435
rect 7395 7405 7396 7435
rect 7364 7404 7396 7405
rect 7364 7355 7396 7356
rect 7364 7325 7365 7355
rect 7365 7325 7395 7355
rect 7395 7325 7396 7355
rect 7364 7324 7396 7325
rect 7364 7275 7396 7276
rect 7364 7245 7365 7275
rect 7365 7245 7395 7275
rect 7395 7245 7396 7275
rect 7364 7244 7396 7245
rect 7364 7195 7396 7196
rect 7364 7165 7365 7195
rect 7365 7165 7395 7195
rect 7395 7165 7396 7195
rect 7364 7164 7396 7165
rect 7364 7115 7396 7116
rect 7364 7085 7365 7115
rect 7365 7085 7395 7115
rect 7395 7085 7396 7115
rect 7364 7084 7396 7085
rect 7364 7035 7396 7036
rect 7364 7005 7365 7035
rect 7365 7005 7395 7035
rect 7395 7005 7396 7035
rect 7364 7004 7396 7005
rect 7364 6955 7396 6956
rect 7364 6925 7365 6955
rect 7365 6925 7395 6955
rect 7395 6925 7396 6955
rect 7364 6924 7396 6925
rect 7364 6875 7396 6876
rect 7364 6845 7365 6875
rect 7365 6845 7395 6875
rect 7395 6845 7396 6875
rect 7364 6844 7396 6845
rect 7364 6795 7396 6796
rect 7364 6765 7365 6795
rect 7365 6765 7395 6795
rect 7395 6765 7396 6795
rect 7364 6764 7396 6765
rect 7364 6715 7396 6716
rect 7364 6685 7365 6715
rect 7365 6685 7395 6715
rect 7395 6685 7396 6715
rect 7364 6684 7396 6685
rect 7364 6635 7396 6636
rect 7364 6605 7365 6635
rect 7365 6605 7395 6635
rect 7395 6605 7396 6635
rect 7364 6604 7396 6605
rect 7364 6555 7396 6556
rect 7364 6525 7365 6555
rect 7365 6525 7395 6555
rect 7395 6525 7396 6555
rect 7364 6524 7396 6525
rect 7364 6475 7396 6476
rect 7364 6445 7365 6475
rect 7365 6445 7395 6475
rect 7395 6445 7396 6475
rect 7364 6444 7396 6445
rect 7364 6395 7396 6396
rect 7364 6365 7365 6395
rect 7365 6365 7395 6395
rect 7395 6365 7396 6395
rect 7364 6364 7396 6365
rect 7364 6315 7396 6316
rect 7364 6285 7365 6315
rect 7365 6285 7395 6315
rect 7395 6285 7396 6315
rect 7364 6284 7396 6285
rect 7364 6235 7396 6236
rect 7364 6205 7365 6235
rect 7365 6205 7395 6235
rect 7395 6205 7396 6235
rect 7364 6204 7396 6205
rect 7364 6155 7396 6156
rect 7364 6125 7365 6155
rect 7365 6125 7395 6155
rect 7395 6125 7396 6155
rect 7364 6124 7396 6125
rect 7364 6075 7396 6076
rect 7364 6045 7365 6075
rect 7365 6045 7395 6075
rect 7395 6045 7396 6075
rect 7364 6044 7396 6045
rect 7364 5995 7396 5996
rect 7364 5965 7365 5995
rect 7365 5965 7395 5995
rect 7395 5965 7396 5995
rect 7364 5964 7396 5965
rect 7364 5915 7396 5916
rect 7364 5885 7365 5915
rect 7365 5885 7395 5915
rect 7395 5885 7396 5915
rect 7364 5884 7396 5885
rect 7364 5835 7396 5836
rect 7364 5805 7365 5835
rect 7365 5805 7395 5835
rect 7395 5805 7396 5835
rect 7364 5804 7396 5805
rect 7364 5755 7396 5756
rect 7364 5725 7365 5755
rect 7365 5725 7395 5755
rect 7395 5725 7396 5755
rect 7364 5724 7396 5725
rect 7364 5675 7396 5676
rect 7364 5645 7365 5675
rect 7365 5645 7395 5675
rect 7395 5645 7396 5675
rect 7364 5644 7396 5645
rect 7364 5595 7396 5596
rect 7364 5565 7365 5595
rect 7365 5565 7395 5595
rect 7395 5565 7396 5595
rect 7364 5564 7396 5565
rect 7364 5515 7396 5516
rect 7364 5485 7365 5515
rect 7365 5485 7395 5515
rect 7395 5485 7396 5515
rect 7364 5484 7396 5485
rect 7364 5435 7396 5436
rect 7364 5405 7365 5435
rect 7365 5405 7395 5435
rect 7395 5405 7396 5435
rect 7364 5404 7396 5405
rect 7364 5355 7396 5356
rect 7364 5325 7365 5355
rect 7365 5325 7395 5355
rect 7395 5325 7396 5355
rect 7364 5324 7396 5325
rect 7364 5275 7396 5276
rect 7364 5245 7365 5275
rect 7365 5245 7395 5275
rect 7395 5245 7396 5275
rect 7364 5244 7396 5245
rect 7364 5195 7396 5196
rect 7364 5165 7365 5195
rect 7365 5165 7395 5195
rect 7395 5165 7396 5195
rect 7364 5164 7396 5165
rect 7364 5115 7396 5116
rect 7364 5085 7365 5115
rect 7365 5085 7395 5115
rect 7395 5085 7396 5115
rect 7364 5084 7396 5085
rect 7364 5035 7396 5036
rect 7364 5005 7365 5035
rect 7365 5005 7395 5035
rect 7395 5005 7396 5035
rect 7364 5004 7396 5005
rect 7364 4955 7396 4956
rect 7364 4925 7365 4955
rect 7365 4925 7395 4955
rect 7395 4925 7396 4955
rect 7364 4924 7396 4925
rect 7364 4875 7396 4876
rect 7364 4845 7365 4875
rect 7365 4845 7395 4875
rect 7395 4845 7396 4875
rect 7364 4844 7396 4845
rect 7364 4795 7396 4796
rect 7364 4765 7365 4795
rect 7365 4765 7395 4795
rect 7395 4765 7396 4795
rect 7364 4764 7396 4765
rect 7364 4715 7396 4716
rect 7364 4685 7365 4715
rect 7365 4685 7395 4715
rect 7395 4685 7396 4715
rect 7364 4684 7396 4685
rect 7364 4635 7396 4636
rect 7364 4605 7365 4635
rect 7365 4605 7395 4635
rect 7395 4605 7396 4635
rect 7364 4604 7396 4605
rect 7364 4555 7396 4556
rect 7364 4525 7365 4555
rect 7365 4525 7395 4555
rect 7395 4525 7396 4555
rect 7364 4524 7396 4525
rect 7364 4475 7396 4476
rect 7364 4445 7365 4475
rect 7365 4445 7395 4475
rect 7395 4445 7396 4475
rect 7364 4444 7396 4445
rect 7364 4395 7396 4396
rect 7364 4365 7365 4395
rect 7365 4365 7395 4395
rect 7395 4365 7396 4395
rect 7364 4364 7396 4365
rect 7364 4315 7396 4316
rect 7364 4285 7365 4315
rect 7365 4285 7395 4315
rect 7395 4285 7396 4315
rect 7364 4284 7396 4285
rect 7364 4235 7396 4236
rect 7364 4205 7365 4235
rect 7365 4205 7395 4235
rect 7395 4205 7396 4235
rect 7364 4204 7396 4205
rect 7364 4155 7396 4156
rect 7364 4125 7365 4155
rect 7365 4125 7395 4155
rect 7395 4125 7396 4155
rect 7364 4124 7396 4125
rect 7364 4075 7396 4076
rect 7364 4045 7365 4075
rect 7365 4045 7395 4075
rect 7395 4045 7396 4075
rect 7364 4044 7396 4045
rect 7364 3995 7396 3996
rect 7364 3965 7365 3995
rect 7365 3965 7395 3995
rect 7395 3965 7396 3995
rect 7364 3964 7396 3965
rect 7364 3915 7396 3916
rect 7364 3885 7365 3915
rect 7365 3885 7395 3915
rect 7395 3885 7396 3915
rect 7364 3884 7396 3885
rect 7364 3835 7396 3836
rect 7364 3805 7365 3835
rect 7365 3805 7395 3835
rect 7395 3805 7396 3835
rect 7364 3804 7396 3805
rect 7364 3755 7396 3756
rect 7364 3725 7365 3755
rect 7365 3725 7395 3755
rect 7395 3725 7396 3755
rect 7364 3724 7396 3725
rect 7364 3675 7396 3676
rect 7364 3645 7365 3675
rect 7365 3645 7395 3675
rect 7395 3645 7396 3675
rect 7364 3644 7396 3645
rect 7364 3595 7396 3596
rect 7364 3565 7365 3595
rect 7365 3565 7395 3595
rect 7395 3565 7396 3595
rect 7364 3564 7396 3565
rect 7364 3515 7396 3516
rect 7364 3485 7365 3515
rect 7365 3485 7395 3515
rect 7395 3485 7396 3515
rect 7364 3484 7396 3485
rect 7364 3435 7396 3436
rect 7364 3405 7365 3435
rect 7365 3405 7395 3435
rect 7395 3405 7396 3435
rect 7364 3404 7396 3405
rect 7364 3355 7396 3356
rect 7364 3325 7365 3355
rect 7365 3325 7395 3355
rect 7395 3325 7396 3355
rect 7364 3324 7396 3325
rect 7364 3275 7396 3276
rect 7364 3245 7365 3275
rect 7365 3245 7395 3275
rect 7395 3245 7396 3275
rect 7364 3244 7396 3245
rect 7364 3195 7396 3196
rect 7364 3165 7365 3195
rect 7365 3165 7395 3195
rect 7395 3165 7396 3195
rect 7364 3164 7396 3165
rect 7364 3115 7396 3116
rect 7364 3085 7365 3115
rect 7365 3085 7395 3115
rect 7395 3085 7396 3115
rect 7364 3084 7396 3085
rect 7364 3035 7396 3036
rect 7364 3005 7365 3035
rect 7365 3005 7395 3035
rect 7395 3005 7396 3035
rect 7364 3004 7396 3005
rect 7364 2955 7396 2956
rect 7364 2925 7365 2955
rect 7365 2925 7395 2955
rect 7395 2925 7396 2955
rect 7364 2924 7396 2925
rect 7364 2875 7396 2876
rect 7364 2845 7365 2875
rect 7365 2845 7395 2875
rect 7395 2845 7396 2875
rect 7364 2844 7396 2845
rect 7364 2795 7396 2796
rect 7364 2765 7365 2795
rect 7365 2765 7395 2795
rect 7395 2765 7396 2795
rect 7364 2764 7396 2765
rect 7364 2715 7396 2716
rect 7364 2685 7365 2715
rect 7365 2685 7395 2715
rect 7395 2685 7396 2715
rect 7364 2684 7396 2685
rect 7364 2635 7396 2636
rect 7364 2605 7365 2635
rect 7365 2605 7395 2635
rect 7395 2605 7396 2635
rect 7364 2604 7396 2605
rect 7364 2555 7396 2556
rect 7364 2525 7365 2555
rect 7365 2525 7395 2555
rect 7395 2525 7396 2555
rect 7364 2524 7396 2525
rect 7364 2475 7396 2476
rect 7364 2445 7365 2475
rect 7365 2445 7395 2475
rect 7395 2445 7396 2475
rect 7364 2444 7396 2445
rect 7364 2395 7396 2396
rect 7364 2365 7365 2395
rect 7365 2365 7395 2395
rect 7395 2365 7396 2395
rect 7364 2364 7396 2365
rect 7364 2315 7396 2316
rect 7364 2285 7365 2315
rect 7365 2285 7395 2315
rect 7395 2285 7396 2315
rect 7364 2284 7396 2285
rect 7364 2235 7396 2236
rect 7364 2205 7365 2235
rect 7365 2205 7395 2235
rect 7395 2205 7396 2235
rect 7364 2204 7396 2205
rect 7364 2155 7396 2156
rect 7364 2125 7365 2155
rect 7365 2125 7395 2155
rect 7395 2125 7396 2155
rect 7364 2124 7396 2125
rect 7364 2075 7396 2076
rect 7364 2045 7365 2075
rect 7365 2045 7395 2075
rect 7395 2045 7396 2075
rect 7364 2044 7396 2045
rect 7364 1995 7396 1996
rect 7364 1965 7365 1995
rect 7365 1965 7395 1995
rect 7395 1965 7396 1995
rect 7364 1964 7396 1965
rect 7364 1915 7396 1916
rect 7364 1885 7365 1915
rect 7365 1885 7395 1915
rect 7395 1885 7396 1915
rect 7364 1884 7396 1885
rect 7364 1835 7396 1836
rect 7364 1805 7365 1835
rect 7365 1805 7395 1835
rect 7395 1805 7396 1835
rect 7364 1804 7396 1805
rect 7364 1755 7396 1756
rect 7364 1725 7365 1755
rect 7365 1725 7395 1755
rect 7395 1725 7396 1755
rect 7364 1724 7396 1725
rect 7364 1675 7396 1676
rect 7364 1645 7365 1675
rect 7365 1645 7395 1675
rect 7395 1645 7396 1675
rect 7364 1644 7396 1645
rect 7364 1595 7396 1596
rect 7364 1565 7365 1595
rect 7365 1565 7395 1595
rect 7395 1565 7396 1595
rect 7364 1564 7396 1565
rect 7364 1515 7396 1516
rect 7364 1485 7365 1515
rect 7365 1485 7395 1515
rect 7395 1485 7396 1515
rect 7364 1484 7396 1485
rect 7364 1435 7396 1436
rect 7364 1405 7365 1435
rect 7365 1405 7395 1435
rect 7395 1405 7396 1435
rect 7364 1404 7396 1405
rect 7364 1355 7396 1356
rect 7364 1325 7365 1355
rect 7365 1325 7395 1355
rect 7395 1325 7396 1355
rect 7364 1324 7396 1325
rect 7364 1275 7396 1276
rect 7364 1245 7365 1275
rect 7365 1245 7395 1275
rect 7395 1245 7396 1275
rect 7364 1244 7396 1245
rect 7364 1195 7396 1196
rect 7364 1165 7365 1195
rect 7365 1165 7395 1195
rect 7395 1165 7396 1195
rect 7364 1164 7396 1165
rect 7364 1115 7396 1116
rect 7364 1085 7365 1115
rect 7365 1085 7395 1115
rect 7395 1085 7396 1115
rect 7364 1084 7396 1085
rect 7364 1035 7396 1036
rect 7364 1005 7365 1035
rect 7365 1005 7395 1035
rect 7395 1005 7396 1035
rect 7364 1004 7396 1005
rect 7364 955 7396 956
rect 7364 925 7365 955
rect 7365 925 7395 955
rect 7395 925 7396 955
rect 7364 924 7396 925
rect 7364 875 7396 876
rect 7364 845 7365 875
rect 7365 845 7395 875
rect 7395 845 7396 875
rect 7364 844 7396 845
rect 7364 795 7396 796
rect 7364 765 7365 795
rect 7365 765 7395 795
rect 7395 765 7396 795
rect 7364 764 7396 765
rect 7364 715 7396 716
rect 7364 685 7365 715
rect 7365 685 7395 715
rect 7395 685 7396 715
rect 7364 684 7396 685
rect 7364 595 7396 596
rect 7364 565 7365 595
rect 7365 565 7395 595
rect 7395 565 7396 595
rect 7364 564 7396 565
rect 7364 515 7396 516
rect 7364 485 7365 515
rect 7365 485 7395 515
rect 7395 485 7396 515
rect 7364 484 7396 485
rect 7364 435 7396 436
rect 7364 405 7365 435
rect 7365 405 7395 435
rect 7395 405 7396 435
rect 7364 404 7396 405
rect 7364 355 7396 356
rect 7364 325 7365 355
rect 7365 325 7395 355
rect 7395 325 7396 355
rect 7364 324 7396 325
rect 7364 275 7396 276
rect 7364 245 7365 275
rect 7365 245 7395 275
rect 7395 245 7396 275
rect 7364 244 7396 245
rect 7364 195 7396 196
rect 7364 165 7365 195
rect 7365 165 7395 195
rect 7395 165 7396 195
rect 7364 164 7396 165
rect 7364 115 7396 116
rect 7364 85 7365 115
rect 7365 85 7395 115
rect 7395 85 7396 115
rect 7364 84 7396 85
rect 7364 35 7396 36
rect 7364 5 7365 35
rect 7365 5 7395 35
rect 7395 5 7396 35
rect 7364 4 7396 5
rect 7444 19604 7476 19636
rect 7524 18484 7556 18516
rect 7524 18404 7556 18436
rect 7684 19684 7716 19716
rect 7684 18484 7716 18516
rect 7684 18404 7716 18436
rect 7604 17284 7636 17316
rect 7524 16595 7556 16596
rect 7524 16565 7525 16595
rect 7525 16565 7555 16595
rect 7555 16565 7556 16595
rect 7524 16564 7556 16565
rect 7524 16515 7556 16516
rect 7524 16485 7525 16515
rect 7525 16485 7555 16515
rect 7555 16485 7556 16515
rect 7524 16484 7556 16485
rect 7524 16435 7556 16436
rect 7524 16405 7525 16435
rect 7525 16405 7555 16435
rect 7555 16405 7556 16435
rect 7524 16404 7556 16405
rect 7524 16355 7556 16356
rect 7524 16325 7525 16355
rect 7525 16325 7555 16355
rect 7555 16325 7556 16355
rect 7524 16324 7556 16325
rect 7524 16275 7556 16276
rect 7524 16245 7525 16275
rect 7525 16245 7555 16275
rect 7555 16245 7556 16275
rect 7524 16244 7556 16245
rect 7524 16195 7556 16196
rect 7524 16165 7525 16195
rect 7525 16165 7555 16195
rect 7555 16165 7556 16195
rect 7524 16164 7556 16165
rect 7524 16115 7556 16116
rect 7524 16085 7525 16115
rect 7525 16085 7555 16115
rect 7555 16085 7556 16115
rect 7524 16084 7556 16085
rect 7524 16035 7556 16036
rect 7524 16005 7525 16035
rect 7525 16005 7555 16035
rect 7555 16005 7556 16035
rect 7524 16004 7556 16005
rect 7524 15955 7556 15956
rect 7524 15925 7525 15955
rect 7525 15925 7555 15955
rect 7555 15925 7556 15955
rect 7524 15924 7556 15925
rect 7524 15435 7556 15436
rect 7524 15405 7525 15435
rect 7525 15405 7555 15435
rect 7555 15405 7556 15435
rect 7524 15404 7556 15405
rect 7524 15355 7556 15356
rect 7524 15325 7525 15355
rect 7525 15325 7555 15355
rect 7555 15325 7556 15355
rect 7524 15324 7556 15325
rect 7524 15275 7556 15276
rect 7524 15245 7525 15275
rect 7525 15245 7555 15275
rect 7555 15245 7556 15275
rect 7524 15244 7556 15245
rect 7524 15195 7556 15196
rect 7524 15165 7525 15195
rect 7525 15165 7555 15195
rect 7555 15165 7556 15195
rect 7524 15164 7556 15165
rect 7524 15115 7556 15116
rect 7524 15085 7525 15115
rect 7525 15085 7555 15115
rect 7555 15085 7556 15115
rect 7524 15084 7556 15085
rect 7524 15035 7556 15036
rect 7524 15005 7525 15035
rect 7525 15005 7555 15035
rect 7555 15005 7556 15035
rect 7524 15004 7556 15005
rect 7524 14955 7556 14956
rect 7524 14925 7525 14955
rect 7525 14925 7555 14955
rect 7555 14925 7556 14955
rect 7524 14924 7556 14925
rect 7524 14875 7556 14876
rect 7524 14845 7525 14875
rect 7525 14845 7555 14875
rect 7555 14845 7556 14875
rect 7524 14844 7556 14845
rect 7524 14795 7556 14796
rect 7524 14765 7525 14795
rect 7525 14765 7555 14795
rect 7555 14765 7556 14795
rect 7524 14764 7556 14765
rect 7524 14715 7556 14716
rect 7524 14685 7525 14715
rect 7525 14685 7555 14715
rect 7555 14685 7556 14715
rect 7524 14684 7556 14685
rect 7524 14635 7556 14636
rect 7524 14605 7525 14635
rect 7525 14605 7555 14635
rect 7555 14605 7556 14635
rect 7524 14604 7556 14605
rect 7524 14555 7556 14556
rect 7524 14525 7525 14555
rect 7525 14525 7555 14555
rect 7555 14525 7556 14555
rect 7524 14524 7556 14525
rect 7524 14475 7556 14476
rect 7524 14445 7525 14475
rect 7525 14445 7555 14475
rect 7555 14445 7556 14475
rect 7524 14444 7556 14445
rect 7524 14395 7556 14396
rect 7524 14365 7525 14395
rect 7525 14365 7555 14395
rect 7555 14365 7556 14395
rect 7524 14364 7556 14365
rect 7524 14315 7556 14316
rect 7524 14285 7525 14315
rect 7525 14285 7555 14315
rect 7555 14285 7556 14315
rect 7524 14284 7556 14285
rect 7524 14235 7556 14236
rect 7524 14205 7525 14235
rect 7525 14205 7555 14235
rect 7555 14205 7556 14235
rect 7524 14204 7556 14205
rect 7524 14155 7556 14156
rect 7524 14125 7525 14155
rect 7525 14125 7555 14155
rect 7555 14125 7556 14155
rect 7524 14124 7556 14125
rect 7524 14075 7556 14076
rect 7524 14045 7525 14075
rect 7525 14045 7555 14075
rect 7555 14045 7556 14075
rect 7524 14044 7556 14045
rect 7524 13995 7556 13996
rect 7524 13965 7525 13995
rect 7525 13965 7555 13995
rect 7555 13965 7556 13995
rect 7524 13964 7556 13965
rect 7524 13875 7556 13876
rect 7524 13845 7525 13875
rect 7525 13845 7555 13875
rect 7555 13845 7556 13875
rect 7524 13844 7556 13845
rect 7524 13795 7556 13796
rect 7524 13765 7525 13795
rect 7525 13765 7555 13795
rect 7555 13765 7556 13795
rect 7524 13764 7556 13765
rect 7524 13715 7556 13716
rect 7524 13685 7525 13715
rect 7525 13685 7555 13715
rect 7555 13685 7556 13715
rect 7524 13684 7556 13685
rect 7524 13635 7556 13636
rect 7524 13605 7525 13635
rect 7525 13605 7555 13635
rect 7555 13605 7556 13635
rect 7524 13604 7556 13605
rect 7524 13555 7556 13556
rect 7524 13525 7525 13555
rect 7525 13525 7555 13555
rect 7555 13525 7556 13555
rect 7524 13524 7556 13525
rect 7524 13475 7556 13476
rect 7524 13445 7525 13475
rect 7525 13445 7555 13475
rect 7555 13445 7556 13475
rect 7524 13444 7556 13445
rect 7524 13395 7556 13396
rect 7524 13365 7525 13395
rect 7525 13365 7555 13395
rect 7555 13365 7556 13395
rect 7524 13364 7556 13365
rect 7524 13315 7556 13316
rect 7524 13285 7525 13315
rect 7525 13285 7555 13315
rect 7555 13285 7556 13315
rect 7524 13284 7556 13285
rect 7524 13235 7556 13236
rect 7524 13205 7525 13235
rect 7525 13205 7555 13235
rect 7555 13205 7556 13235
rect 7524 13204 7556 13205
rect 7524 13155 7556 13156
rect 7524 13125 7525 13155
rect 7525 13125 7555 13155
rect 7555 13125 7556 13155
rect 7524 13124 7556 13125
rect 7524 13075 7556 13076
rect 7524 13045 7525 13075
rect 7525 13045 7555 13075
rect 7555 13045 7556 13075
rect 7524 13044 7556 13045
rect 7524 12995 7556 12996
rect 7524 12965 7525 12995
rect 7525 12965 7555 12995
rect 7555 12965 7556 12995
rect 7524 12964 7556 12965
rect 7524 12475 7556 12476
rect 7524 12445 7525 12475
rect 7525 12445 7555 12475
rect 7555 12445 7556 12475
rect 7524 12444 7556 12445
rect 7524 12395 7556 12396
rect 7524 12365 7525 12395
rect 7525 12365 7555 12395
rect 7555 12365 7556 12395
rect 7524 12364 7556 12365
rect 7524 12315 7556 12316
rect 7524 12285 7525 12315
rect 7525 12285 7555 12315
rect 7555 12285 7556 12315
rect 7524 12284 7556 12285
rect 7524 12235 7556 12236
rect 7524 12205 7525 12235
rect 7525 12205 7555 12235
rect 7555 12205 7556 12235
rect 7524 12204 7556 12205
rect 7524 12155 7556 12156
rect 7524 12125 7525 12155
rect 7525 12125 7555 12155
rect 7555 12125 7556 12155
rect 7524 12124 7556 12125
rect 7524 12075 7556 12076
rect 7524 12045 7525 12075
rect 7525 12045 7555 12075
rect 7555 12045 7556 12075
rect 7524 12044 7556 12045
rect 7524 11995 7556 11996
rect 7524 11965 7525 11995
rect 7525 11965 7555 11995
rect 7555 11965 7556 11995
rect 7524 11964 7556 11965
rect 7524 11915 7556 11916
rect 7524 11885 7525 11915
rect 7525 11885 7555 11915
rect 7555 11885 7556 11915
rect 7524 11884 7556 11885
rect 7524 11835 7556 11836
rect 7524 11805 7525 11835
rect 7525 11805 7555 11835
rect 7555 11805 7556 11835
rect 7524 11804 7556 11805
rect 7524 11755 7556 11756
rect 7524 11725 7525 11755
rect 7525 11725 7555 11755
rect 7555 11725 7556 11755
rect 7524 11724 7556 11725
rect 7524 11675 7556 11676
rect 7524 11645 7525 11675
rect 7525 11645 7555 11675
rect 7555 11645 7556 11675
rect 7524 11644 7556 11645
rect 7524 11595 7556 11596
rect 7524 11565 7525 11595
rect 7525 11565 7555 11595
rect 7555 11565 7556 11595
rect 7524 11564 7556 11565
rect 7524 11515 7556 11516
rect 7524 11485 7525 11515
rect 7525 11485 7555 11515
rect 7555 11485 7556 11515
rect 7524 11484 7556 11485
rect 7524 11435 7556 11436
rect 7524 11405 7525 11435
rect 7525 11405 7555 11435
rect 7555 11405 7556 11435
rect 7524 11404 7556 11405
rect 7524 11355 7556 11356
rect 7524 11325 7525 11355
rect 7525 11325 7555 11355
rect 7555 11325 7556 11355
rect 7524 11324 7556 11325
rect 7524 11275 7556 11276
rect 7524 11245 7525 11275
rect 7525 11245 7555 11275
rect 7555 11245 7556 11275
rect 7524 11244 7556 11245
rect 7524 11195 7556 11196
rect 7524 11165 7525 11195
rect 7525 11165 7555 11195
rect 7555 11165 7556 11195
rect 7524 11164 7556 11165
rect 7524 11115 7556 11116
rect 7524 11085 7525 11115
rect 7525 11085 7555 11115
rect 7555 11085 7556 11115
rect 7524 11084 7556 11085
rect 7524 11035 7556 11036
rect 7524 11005 7525 11035
rect 7525 11005 7555 11035
rect 7555 11005 7556 11035
rect 7524 11004 7556 11005
rect 7524 10955 7556 10956
rect 7524 10925 7525 10955
rect 7525 10925 7555 10955
rect 7555 10925 7556 10955
rect 7524 10924 7556 10925
rect 7524 10875 7556 10876
rect 7524 10845 7525 10875
rect 7525 10845 7555 10875
rect 7555 10845 7556 10875
rect 7524 10844 7556 10845
rect 7524 10795 7556 10796
rect 7524 10765 7525 10795
rect 7525 10765 7555 10795
rect 7555 10765 7556 10795
rect 7524 10764 7556 10765
rect 7524 10715 7556 10716
rect 7524 10685 7525 10715
rect 7525 10685 7555 10715
rect 7555 10685 7556 10715
rect 7524 10684 7556 10685
rect 7524 10635 7556 10636
rect 7524 10605 7525 10635
rect 7525 10605 7555 10635
rect 7555 10605 7556 10635
rect 7524 10604 7556 10605
rect 7524 10555 7556 10556
rect 7524 10525 7525 10555
rect 7525 10525 7555 10555
rect 7555 10525 7556 10555
rect 7524 10524 7556 10525
rect 7524 10475 7556 10476
rect 7524 10445 7525 10475
rect 7525 10445 7555 10475
rect 7555 10445 7556 10475
rect 7524 10444 7556 10445
rect 7524 10395 7556 10396
rect 7524 10365 7525 10395
rect 7525 10365 7555 10395
rect 7555 10365 7556 10395
rect 7524 10364 7556 10365
rect 7524 10315 7556 10316
rect 7524 10285 7525 10315
rect 7525 10285 7555 10315
rect 7555 10285 7556 10315
rect 7524 10284 7556 10285
rect 7524 10235 7556 10236
rect 7524 10205 7525 10235
rect 7525 10205 7555 10235
rect 7555 10205 7556 10235
rect 7524 10204 7556 10205
rect 7524 10155 7556 10156
rect 7524 10125 7525 10155
rect 7525 10125 7555 10155
rect 7555 10125 7556 10155
rect 7524 10124 7556 10125
rect 7524 10075 7556 10076
rect 7524 10045 7525 10075
rect 7525 10045 7555 10075
rect 7555 10045 7556 10075
rect 7524 10044 7556 10045
rect 7524 9995 7556 9996
rect 7524 9965 7525 9995
rect 7525 9965 7555 9995
rect 7555 9965 7556 9995
rect 7524 9964 7556 9965
rect 7524 9915 7556 9916
rect 7524 9885 7525 9915
rect 7525 9885 7555 9915
rect 7555 9885 7556 9915
rect 7524 9884 7556 9885
rect 7524 9835 7556 9836
rect 7524 9805 7525 9835
rect 7525 9805 7555 9835
rect 7555 9805 7556 9835
rect 7524 9804 7556 9805
rect 7524 9755 7556 9756
rect 7524 9725 7525 9755
rect 7525 9725 7555 9755
rect 7555 9725 7556 9755
rect 7524 9724 7556 9725
rect 7524 9675 7556 9676
rect 7524 9645 7525 9675
rect 7525 9645 7555 9675
rect 7555 9645 7556 9675
rect 7524 9644 7556 9645
rect 7524 9595 7556 9596
rect 7524 9565 7525 9595
rect 7525 9565 7555 9595
rect 7555 9565 7556 9595
rect 7524 9564 7556 9565
rect 7524 9515 7556 9516
rect 7524 9485 7525 9515
rect 7525 9485 7555 9515
rect 7555 9485 7556 9515
rect 7524 9484 7556 9485
rect 7524 9435 7556 9436
rect 7524 9405 7525 9435
rect 7525 9405 7555 9435
rect 7555 9405 7556 9435
rect 7524 9404 7556 9405
rect 7524 9355 7556 9356
rect 7524 9325 7525 9355
rect 7525 9325 7555 9355
rect 7555 9325 7556 9355
rect 7524 9324 7556 9325
rect 7524 9275 7556 9276
rect 7524 9245 7525 9275
rect 7525 9245 7555 9275
rect 7555 9245 7556 9275
rect 7524 9244 7556 9245
rect 7524 9195 7556 9196
rect 7524 9165 7525 9195
rect 7525 9165 7555 9195
rect 7555 9165 7556 9195
rect 7524 9164 7556 9165
rect 7524 9115 7556 9116
rect 7524 9085 7525 9115
rect 7525 9085 7555 9115
rect 7555 9085 7556 9115
rect 7524 9084 7556 9085
rect 7524 9035 7556 9036
rect 7524 9005 7525 9035
rect 7525 9005 7555 9035
rect 7555 9005 7556 9035
rect 7524 9004 7556 9005
rect 7524 8955 7556 8956
rect 7524 8925 7525 8955
rect 7525 8925 7555 8955
rect 7555 8925 7556 8955
rect 7524 8924 7556 8925
rect 7524 8635 7556 8636
rect 7524 8605 7525 8635
rect 7525 8605 7555 8635
rect 7555 8605 7556 8635
rect 7524 8604 7556 8605
rect 7524 8555 7556 8556
rect 7524 8525 7525 8555
rect 7525 8525 7555 8555
rect 7555 8525 7556 8555
rect 7524 8524 7556 8525
rect 7524 8475 7556 8476
rect 7524 8445 7525 8475
rect 7525 8445 7555 8475
rect 7555 8445 7556 8475
rect 7524 8444 7556 8445
rect 7524 8395 7556 8396
rect 7524 8365 7525 8395
rect 7525 8365 7555 8395
rect 7555 8365 7556 8395
rect 7524 8364 7556 8365
rect 7524 8315 7556 8316
rect 7524 8285 7525 8315
rect 7525 8285 7555 8315
rect 7555 8285 7556 8315
rect 7524 8284 7556 8285
rect 7524 8235 7556 8236
rect 7524 8205 7525 8235
rect 7525 8205 7555 8235
rect 7555 8205 7556 8235
rect 7524 8204 7556 8205
rect 7524 8155 7556 8156
rect 7524 8125 7525 8155
rect 7525 8125 7555 8155
rect 7555 8125 7556 8155
rect 7524 8124 7556 8125
rect 7524 8075 7556 8076
rect 7524 8045 7525 8075
rect 7525 8045 7555 8075
rect 7555 8045 7556 8075
rect 7524 8044 7556 8045
rect 7524 7995 7556 7996
rect 7524 7965 7525 7995
rect 7525 7965 7555 7995
rect 7555 7965 7556 7995
rect 7524 7964 7556 7965
rect 7524 7915 7556 7916
rect 7524 7885 7525 7915
rect 7525 7885 7555 7915
rect 7555 7885 7556 7915
rect 7524 7884 7556 7885
rect 7524 7835 7556 7836
rect 7524 7805 7525 7835
rect 7525 7805 7555 7835
rect 7555 7805 7556 7835
rect 7524 7804 7556 7805
rect 7524 7755 7556 7756
rect 7524 7725 7525 7755
rect 7525 7725 7555 7755
rect 7555 7725 7556 7755
rect 7524 7724 7556 7725
rect 7524 7675 7556 7676
rect 7524 7645 7525 7675
rect 7525 7645 7555 7675
rect 7555 7645 7556 7675
rect 7524 7644 7556 7645
rect 7524 7595 7556 7596
rect 7524 7565 7525 7595
rect 7525 7565 7555 7595
rect 7555 7565 7556 7595
rect 7524 7564 7556 7565
rect 7524 7515 7556 7516
rect 7524 7485 7525 7515
rect 7525 7485 7555 7515
rect 7555 7485 7556 7515
rect 7524 7484 7556 7485
rect 7524 7435 7556 7436
rect 7524 7405 7525 7435
rect 7525 7405 7555 7435
rect 7555 7405 7556 7435
rect 7524 7404 7556 7405
rect 7524 7355 7556 7356
rect 7524 7325 7525 7355
rect 7525 7325 7555 7355
rect 7555 7325 7556 7355
rect 7524 7324 7556 7325
rect 7524 7275 7556 7276
rect 7524 7245 7525 7275
rect 7525 7245 7555 7275
rect 7555 7245 7556 7275
rect 7524 7244 7556 7245
rect 7524 7195 7556 7196
rect 7524 7165 7525 7195
rect 7525 7165 7555 7195
rect 7555 7165 7556 7195
rect 7524 7164 7556 7165
rect 7524 7115 7556 7116
rect 7524 7085 7525 7115
rect 7525 7085 7555 7115
rect 7555 7085 7556 7115
rect 7524 7084 7556 7085
rect 7524 7035 7556 7036
rect 7524 7005 7525 7035
rect 7525 7005 7555 7035
rect 7555 7005 7556 7035
rect 7524 7004 7556 7005
rect 7524 6955 7556 6956
rect 7524 6925 7525 6955
rect 7525 6925 7555 6955
rect 7555 6925 7556 6955
rect 7524 6924 7556 6925
rect 7524 6875 7556 6876
rect 7524 6845 7525 6875
rect 7525 6845 7555 6875
rect 7555 6845 7556 6875
rect 7524 6844 7556 6845
rect 7524 6795 7556 6796
rect 7524 6765 7525 6795
rect 7525 6765 7555 6795
rect 7555 6765 7556 6795
rect 7524 6764 7556 6765
rect 7524 6715 7556 6716
rect 7524 6685 7525 6715
rect 7525 6685 7555 6715
rect 7555 6685 7556 6715
rect 7524 6684 7556 6685
rect 7524 6635 7556 6636
rect 7524 6605 7525 6635
rect 7525 6605 7555 6635
rect 7555 6605 7556 6635
rect 7524 6604 7556 6605
rect 7524 6555 7556 6556
rect 7524 6525 7525 6555
rect 7525 6525 7555 6555
rect 7555 6525 7556 6555
rect 7524 6524 7556 6525
rect 7524 6475 7556 6476
rect 7524 6445 7525 6475
rect 7525 6445 7555 6475
rect 7555 6445 7556 6475
rect 7524 6444 7556 6445
rect 7524 6395 7556 6396
rect 7524 6365 7525 6395
rect 7525 6365 7555 6395
rect 7555 6365 7556 6395
rect 7524 6364 7556 6365
rect 7524 6315 7556 6316
rect 7524 6285 7525 6315
rect 7525 6285 7555 6315
rect 7555 6285 7556 6315
rect 7524 6284 7556 6285
rect 7524 6235 7556 6236
rect 7524 6205 7525 6235
rect 7525 6205 7555 6235
rect 7555 6205 7556 6235
rect 7524 6204 7556 6205
rect 7524 6155 7556 6156
rect 7524 6125 7525 6155
rect 7525 6125 7555 6155
rect 7555 6125 7556 6155
rect 7524 6124 7556 6125
rect 7524 6075 7556 6076
rect 7524 6045 7525 6075
rect 7525 6045 7555 6075
rect 7555 6045 7556 6075
rect 7524 6044 7556 6045
rect 7524 5995 7556 5996
rect 7524 5965 7525 5995
rect 7525 5965 7555 5995
rect 7555 5965 7556 5995
rect 7524 5964 7556 5965
rect 7524 5915 7556 5916
rect 7524 5885 7525 5915
rect 7525 5885 7555 5915
rect 7555 5885 7556 5915
rect 7524 5884 7556 5885
rect 7524 5835 7556 5836
rect 7524 5805 7525 5835
rect 7525 5805 7555 5835
rect 7555 5805 7556 5835
rect 7524 5804 7556 5805
rect 7524 5755 7556 5756
rect 7524 5725 7525 5755
rect 7525 5725 7555 5755
rect 7555 5725 7556 5755
rect 7524 5724 7556 5725
rect 7524 5675 7556 5676
rect 7524 5645 7525 5675
rect 7525 5645 7555 5675
rect 7555 5645 7556 5675
rect 7524 5644 7556 5645
rect 7524 5595 7556 5596
rect 7524 5565 7525 5595
rect 7525 5565 7555 5595
rect 7555 5565 7556 5595
rect 7524 5564 7556 5565
rect 7524 5515 7556 5516
rect 7524 5485 7525 5515
rect 7525 5485 7555 5515
rect 7555 5485 7556 5515
rect 7524 5484 7556 5485
rect 7524 5435 7556 5436
rect 7524 5405 7525 5435
rect 7525 5405 7555 5435
rect 7555 5405 7556 5435
rect 7524 5404 7556 5405
rect 7524 5355 7556 5356
rect 7524 5325 7525 5355
rect 7525 5325 7555 5355
rect 7555 5325 7556 5355
rect 7524 5324 7556 5325
rect 7524 5275 7556 5276
rect 7524 5245 7525 5275
rect 7525 5245 7555 5275
rect 7555 5245 7556 5275
rect 7524 5244 7556 5245
rect 7524 5195 7556 5196
rect 7524 5165 7525 5195
rect 7525 5165 7555 5195
rect 7555 5165 7556 5195
rect 7524 5164 7556 5165
rect 7524 5115 7556 5116
rect 7524 5085 7525 5115
rect 7525 5085 7555 5115
rect 7555 5085 7556 5115
rect 7524 5084 7556 5085
rect 7524 5035 7556 5036
rect 7524 5005 7525 5035
rect 7525 5005 7555 5035
rect 7555 5005 7556 5035
rect 7524 5004 7556 5005
rect 7524 4955 7556 4956
rect 7524 4925 7525 4955
rect 7525 4925 7555 4955
rect 7555 4925 7556 4955
rect 7524 4924 7556 4925
rect 7524 4875 7556 4876
rect 7524 4845 7525 4875
rect 7525 4845 7555 4875
rect 7555 4845 7556 4875
rect 7524 4844 7556 4845
rect 7524 4795 7556 4796
rect 7524 4765 7525 4795
rect 7525 4765 7555 4795
rect 7555 4765 7556 4795
rect 7524 4764 7556 4765
rect 7524 4715 7556 4716
rect 7524 4685 7525 4715
rect 7525 4685 7555 4715
rect 7555 4685 7556 4715
rect 7524 4684 7556 4685
rect 7524 4635 7556 4636
rect 7524 4605 7525 4635
rect 7525 4605 7555 4635
rect 7555 4605 7556 4635
rect 7524 4604 7556 4605
rect 7524 4555 7556 4556
rect 7524 4525 7525 4555
rect 7525 4525 7555 4555
rect 7555 4525 7556 4555
rect 7524 4524 7556 4525
rect 7524 4475 7556 4476
rect 7524 4445 7525 4475
rect 7525 4445 7555 4475
rect 7555 4445 7556 4475
rect 7524 4444 7556 4445
rect 7524 4395 7556 4396
rect 7524 4365 7525 4395
rect 7525 4365 7555 4395
rect 7555 4365 7556 4395
rect 7524 4364 7556 4365
rect 7524 4315 7556 4316
rect 7524 4285 7525 4315
rect 7525 4285 7555 4315
rect 7555 4285 7556 4315
rect 7524 4284 7556 4285
rect 7524 4235 7556 4236
rect 7524 4205 7525 4235
rect 7525 4205 7555 4235
rect 7555 4205 7556 4235
rect 7524 4204 7556 4205
rect 7524 4155 7556 4156
rect 7524 4125 7525 4155
rect 7525 4125 7555 4155
rect 7555 4125 7556 4155
rect 7524 4124 7556 4125
rect 7524 4075 7556 4076
rect 7524 4045 7525 4075
rect 7525 4045 7555 4075
rect 7555 4045 7556 4075
rect 7524 4044 7556 4045
rect 7524 3995 7556 3996
rect 7524 3965 7525 3995
rect 7525 3965 7555 3995
rect 7555 3965 7556 3995
rect 7524 3964 7556 3965
rect 7524 3915 7556 3916
rect 7524 3885 7525 3915
rect 7525 3885 7555 3915
rect 7555 3885 7556 3915
rect 7524 3884 7556 3885
rect 7524 3835 7556 3836
rect 7524 3805 7525 3835
rect 7525 3805 7555 3835
rect 7555 3805 7556 3835
rect 7524 3804 7556 3805
rect 7524 3755 7556 3756
rect 7524 3725 7525 3755
rect 7525 3725 7555 3755
rect 7555 3725 7556 3755
rect 7524 3724 7556 3725
rect 7524 3675 7556 3676
rect 7524 3645 7525 3675
rect 7525 3645 7555 3675
rect 7555 3645 7556 3675
rect 7524 3644 7556 3645
rect 7524 3595 7556 3596
rect 7524 3565 7525 3595
rect 7525 3565 7555 3595
rect 7555 3565 7556 3595
rect 7524 3564 7556 3565
rect 7524 3515 7556 3516
rect 7524 3485 7525 3515
rect 7525 3485 7555 3515
rect 7555 3485 7556 3515
rect 7524 3484 7556 3485
rect 7524 3435 7556 3436
rect 7524 3405 7525 3435
rect 7525 3405 7555 3435
rect 7555 3405 7556 3435
rect 7524 3404 7556 3405
rect 7524 3355 7556 3356
rect 7524 3325 7525 3355
rect 7525 3325 7555 3355
rect 7555 3325 7556 3355
rect 7524 3324 7556 3325
rect 7524 3275 7556 3276
rect 7524 3245 7525 3275
rect 7525 3245 7555 3275
rect 7555 3245 7556 3275
rect 7524 3244 7556 3245
rect 7524 3195 7556 3196
rect 7524 3165 7525 3195
rect 7525 3165 7555 3195
rect 7555 3165 7556 3195
rect 7524 3164 7556 3165
rect 7524 3115 7556 3116
rect 7524 3085 7525 3115
rect 7525 3085 7555 3115
rect 7555 3085 7556 3115
rect 7524 3084 7556 3085
rect 7524 3035 7556 3036
rect 7524 3005 7525 3035
rect 7525 3005 7555 3035
rect 7555 3005 7556 3035
rect 7524 3004 7556 3005
rect 7524 2955 7556 2956
rect 7524 2925 7525 2955
rect 7525 2925 7555 2955
rect 7555 2925 7556 2955
rect 7524 2924 7556 2925
rect 7524 2875 7556 2876
rect 7524 2845 7525 2875
rect 7525 2845 7555 2875
rect 7555 2845 7556 2875
rect 7524 2844 7556 2845
rect 7524 2795 7556 2796
rect 7524 2765 7525 2795
rect 7525 2765 7555 2795
rect 7555 2765 7556 2795
rect 7524 2764 7556 2765
rect 7524 2715 7556 2716
rect 7524 2685 7525 2715
rect 7525 2685 7555 2715
rect 7555 2685 7556 2715
rect 7524 2684 7556 2685
rect 7524 2635 7556 2636
rect 7524 2605 7525 2635
rect 7525 2605 7555 2635
rect 7555 2605 7556 2635
rect 7524 2604 7556 2605
rect 7524 2555 7556 2556
rect 7524 2525 7525 2555
rect 7525 2525 7555 2555
rect 7555 2525 7556 2555
rect 7524 2524 7556 2525
rect 7524 2475 7556 2476
rect 7524 2445 7525 2475
rect 7525 2445 7555 2475
rect 7555 2445 7556 2475
rect 7524 2444 7556 2445
rect 7524 2395 7556 2396
rect 7524 2365 7525 2395
rect 7525 2365 7555 2395
rect 7555 2365 7556 2395
rect 7524 2364 7556 2365
rect 7524 2315 7556 2316
rect 7524 2285 7525 2315
rect 7525 2285 7555 2315
rect 7555 2285 7556 2315
rect 7524 2284 7556 2285
rect 7524 2235 7556 2236
rect 7524 2205 7525 2235
rect 7525 2205 7555 2235
rect 7555 2205 7556 2235
rect 7524 2204 7556 2205
rect 7524 2155 7556 2156
rect 7524 2125 7525 2155
rect 7525 2125 7555 2155
rect 7555 2125 7556 2155
rect 7524 2124 7556 2125
rect 7524 2075 7556 2076
rect 7524 2045 7525 2075
rect 7525 2045 7555 2075
rect 7555 2045 7556 2075
rect 7524 2044 7556 2045
rect 7524 1995 7556 1996
rect 7524 1965 7525 1995
rect 7525 1965 7555 1995
rect 7555 1965 7556 1995
rect 7524 1964 7556 1965
rect 7524 1915 7556 1916
rect 7524 1885 7525 1915
rect 7525 1885 7555 1915
rect 7555 1885 7556 1915
rect 7524 1884 7556 1885
rect 7524 1835 7556 1836
rect 7524 1805 7525 1835
rect 7525 1805 7555 1835
rect 7555 1805 7556 1835
rect 7524 1804 7556 1805
rect 7524 1755 7556 1756
rect 7524 1725 7525 1755
rect 7525 1725 7555 1755
rect 7555 1725 7556 1755
rect 7524 1724 7556 1725
rect 7524 1675 7556 1676
rect 7524 1645 7525 1675
rect 7525 1645 7555 1675
rect 7555 1645 7556 1675
rect 7524 1644 7556 1645
rect 7524 1595 7556 1596
rect 7524 1565 7525 1595
rect 7525 1565 7555 1595
rect 7555 1565 7556 1595
rect 7524 1564 7556 1565
rect 7524 1515 7556 1516
rect 7524 1485 7525 1515
rect 7525 1485 7555 1515
rect 7555 1485 7556 1515
rect 7524 1484 7556 1485
rect 7524 1435 7556 1436
rect 7524 1405 7525 1435
rect 7525 1405 7555 1435
rect 7555 1405 7556 1435
rect 7524 1404 7556 1405
rect 7524 1355 7556 1356
rect 7524 1325 7525 1355
rect 7525 1325 7555 1355
rect 7555 1325 7556 1355
rect 7524 1324 7556 1325
rect 7524 1275 7556 1276
rect 7524 1245 7525 1275
rect 7525 1245 7555 1275
rect 7555 1245 7556 1275
rect 7524 1244 7556 1245
rect 7524 1195 7556 1196
rect 7524 1165 7525 1195
rect 7525 1165 7555 1195
rect 7555 1165 7556 1195
rect 7524 1164 7556 1165
rect 7524 1115 7556 1116
rect 7524 1085 7525 1115
rect 7525 1085 7555 1115
rect 7555 1085 7556 1115
rect 7524 1084 7556 1085
rect 7524 1035 7556 1036
rect 7524 1005 7525 1035
rect 7525 1005 7555 1035
rect 7555 1005 7556 1035
rect 7524 1004 7556 1005
rect 7524 955 7556 956
rect 7524 925 7525 955
rect 7525 925 7555 955
rect 7555 925 7556 955
rect 7524 924 7556 925
rect 7524 875 7556 876
rect 7524 845 7525 875
rect 7525 845 7555 875
rect 7555 845 7556 875
rect 7524 844 7556 845
rect 7524 795 7556 796
rect 7524 765 7525 795
rect 7525 765 7555 795
rect 7555 765 7556 795
rect 7524 764 7556 765
rect 7524 715 7556 716
rect 7524 685 7525 715
rect 7525 685 7555 715
rect 7555 685 7556 715
rect 7524 684 7556 685
rect 7524 595 7556 596
rect 7524 565 7525 595
rect 7525 565 7555 595
rect 7555 565 7556 595
rect 7524 564 7556 565
rect 7524 515 7556 516
rect 7524 485 7525 515
rect 7525 485 7555 515
rect 7555 485 7556 515
rect 7524 484 7556 485
rect 7524 435 7556 436
rect 7524 405 7525 435
rect 7525 405 7555 435
rect 7555 405 7556 435
rect 7524 404 7556 405
rect 7524 355 7556 356
rect 7524 325 7525 355
rect 7525 325 7555 355
rect 7555 325 7556 355
rect 7524 324 7556 325
rect 7524 275 7556 276
rect 7524 245 7525 275
rect 7525 245 7555 275
rect 7555 245 7556 275
rect 7524 244 7556 245
rect 7524 195 7556 196
rect 7524 165 7525 195
rect 7525 165 7555 195
rect 7555 165 7556 195
rect 7524 164 7556 165
rect 7524 115 7556 116
rect 7524 85 7525 115
rect 7525 85 7555 115
rect 7555 85 7556 115
rect 7524 84 7556 85
rect 7524 35 7556 36
rect 7524 5 7525 35
rect 7525 5 7555 35
rect 7555 5 7556 35
rect 7524 4 7556 5
rect 7764 16644 7796 16836
rect 7684 16595 7716 16596
rect 7684 16565 7685 16595
rect 7685 16565 7715 16595
rect 7715 16565 7716 16595
rect 7684 16564 7716 16565
rect 7684 16515 7716 16516
rect 7684 16485 7685 16515
rect 7685 16485 7715 16515
rect 7715 16485 7716 16515
rect 7684 16484 7716 16485
rect 7684 16435 7716 16436
rect 7684 16405 7685 16435
rect 7685 16405 7715 16435
rect 7715 16405 7716 16435
rect 7684 16404 7716 16405
rect 7684 16355 7716 16356
rect 7684 16325 7685 16355
rect 7685 16325 7715 16355
rect 7715 16325 7716 16355
rect 7684 16324 7716 16325
rect 7684 16275 7716 16276
rect 7684 16245 7685 16275
rect 7685 16245 7715 16275
rect 7715 16245 7716 16275
rect 7684 16244 7716 16245
rect 7684 16195 7716 16196
rect 7684 16165 7685 16195
rect 7685 16165 7715 16195
rect 7715 16165 7716 16195
rect 7684 16164 7716 16165
rect 7684 16115 7716 16116
rect 7684 16085 7685 16115
rect 7685 16085 7715 16115
rect 7715 16085 7716 16115
rect 7684 16084 7716 16085
rect 7684 16035 7716 16036
rect 7684 16005 7685 16035
rect 7685 16005 7715 16035
rect 7715 16005 7716 16035
rect 7684 16004 7716 16005
rect 7684 15955 7716 15956
rect 7684 15925 7685 15955
rect 7685 15925 7715 15955
rect 7715 15925 7716 15955
rect 7684 15924 7716 15925
rect 7684 15435 7716 15436
rect 7684 15405 7685 15435
rect 7685 15405 7715 15435
rect 7715 15405 7716 15435
rect 7684 15404 7716 15405
rect 7684 15355 7716 15356
rect 7684 15325 7685 15355
rect 7685 15325 7715 15355
rect 7715 15325 7716 15355
rect 7684 15324 7716 15325
rect 7684 15275 7716 15276
rect 7684 15245 7685 15275
rect 7685 15245 7715 15275
rect 7715 15245 7716 15275
rect 7684 15244 7716 15245
rect 7684 15195 7716 15196
rect 7684 15165 7685 15195
rect 7685 15165 7715 15195
rect 7715 15165 7716 15195
rect 7684 15164 7716 15165
rect 7684 15115 7716 15116
rect 7684 15085 7685 15115
rect 7685 15085 7715 15115
rect 7715 15085 7716 15115
rect 7684 15084 7716 15085
rect 7684 15035 7716 15036
rect 7684 15005 7685 15035
rect 7685 15005 7715 15035
rect 7715 15005 7716 15035
rect 7684 15004 7716 15005
rect 7684 14955 7716 14956
rect 7684 14925 7685 14955
rect 7685 14925 7715 14955
rect 7715 14925 7716 14955
rect 7684 14924 7716 14925
rect 7684 14875 7716 14876
rect 7684 14845 7685 14875
rect 7685 14845 7715 14875
rect 7715 14845 7716 14875
rect 7684 14844 7716 14845
rect 7684 14795 7716 14796
rect 7684 14765 7685 14795
rect 7685 14765 7715 14795
rect 7715 14765 7716 14795
rect 7684 14764 7716 14765
rect 7684 14715 7716 14716
rect 7684 14685 7685 14715
rect 7685 14685 7715 14715
rect 7715 14685 7716 14715
rect 7684 14684 7716 14685
rect 7684 14635 7716 14636
rect 7684 14605 7685 14635
rect 7685 14605 7715 14635
rect 7715 14605 7716 14635
rect 7684 14604 7716 14605
rect 7684 14555 7716 14556
rect 7684 14525 7685 14555
rect 7685 14525 7715 14555
rect 7715 14525 7716 14555
rect 7684 14524 7716 14525
rect 7684 14475 7716 14476
rect 7684 14445 7685 14475
rect 7685 14445 7715 14475
rect 7715 14445 7716 14475
rect 7684 14444 7716 14445
rect 7684 14395 7716 14396
rect 7684 14365 7685 14395
rect 7685 14365 7715 14395
rect 7715 14365 7716 14395
rect 7684 14364 7716 14365
rect 7684 14315 7716 14316
rect 7684 14285 7685 14315
rect 7685 14285 7715 14315
rect 7715 14285 7716 14315
rect 7684 14284 7716 14285
rect 7684 14235 7716 14236
rect 7684 14205 7685 14235
rect 7685 14205 7715 14235
rect 7715 14205 7716 14235
rect 7684 14204 7716 14205
rect 7684 14155 7716 14156
rect 7684 14125 7685 14155
rect 7685 14125 7715 14155
rect 7715 14125 7716 14155
rect 7684 14124 7716 14125
rect 7684 14075 7716 14076
rect 7684 14045 7685 14075
rect 7685 14045 7715 14075
rect 7715 14045 7716 14075
rect 7684 14044 7716 14045
rect 7684 13995 7716 13996
rect 7684 13965 7685 13995
rect 7685 13965 7715 13995
rect 7715 13965 7716 13995
rect 7684 13964 7716 13965
rect 7684 13875 7716 13876
rect 7684 13845 7685 13875
rect 7685 13845 7715 13875
rect 7715 13845 7716 13875
rect 7684 13844 7716 13845
rect 7684 13795 7716 13796
rect 7684 13765 7685 13795
rect 7685 13765 7715 13795
rect 7715 13765 7716 13795
rect 7684 13764 7716 13765
rect 7684 13715 7716 13716
rect 7684 13685 7685 13715
rect 7685 13685 7715 13715
rect 7715 13685 7716 13715
rect 7684 13684 7716 13685
rect 7684 13635 7716 13636
rect 7684 13605 7685 13635
rect 7685 13605 7715 13635
rect 7715 13605 7716 13635
rect 7684 13604 7716 13605
rect 7684 13555 7716 13556
rect 7684 13525 7685 13555
rect 7685 13525 7715 13555
rect 7715 13525 7716 13555
rect 7684 13524 7716 13525
rect 7684 13475 7716 13476
rect 7684 13445 7685 13475
rect 7685 13445 7715 13475
rect 7715 13445 7716 13475
rect 7684 13444 7716 13445
rect 7684 13395 7716 13396
rect 7684 13365 7685 13395
rect 7685 13365 7715 13395
rect 7715 13365 7716 13395
rect 7684 13364 7716 13365
rect 7684 13315 7716 13316
rect 7684 13285 7685 13315
rect 7685 13285 7715 13315
rect 7715 13285 7716 13315
rect 7684 13284 7716 13285
rect 7684 13235 7716 13236
rect 7684 13205 7685 13235
rect 7685 13205 7715 13235
rect 7715 13205 7716 13235
rect 7684 13204 7716 13205
rect 7684 13155 7716 13156
rect 7684 13125 7685 13155
rect 7685 13125 7715 13155
rect 7715 13125 7716 13155
rect 7684 13124 7716 13125
rect 7684 13075 7716 13076
rect 7684 13045 7685 13075
rect 7685 13045 7715 13075
rect 7715 13045 7716 13075
rect 7684 13044 7716 13045
rect 7684 12995 7716 12996
rect 7684 12965 7685 12995
rect 7685 12965 7715 12995
rect 7715 12965 7716 12995
rect 7684 12964 7716 12965
rect 7684 12475 7716 12476
rect 7684 12445 7685 12475
rect 7685 12445 7715 12475
rect 7715 12445 7716 12475
rect 7684 12444 7716 12445
rect 7684 12395 7716 12396
rect 7684 12365 7685 12395
rect 7685 12365 7715 12395
rect 7715 12365 7716 12395
rect 7684 12364 7716 12365
rect 7684 12315 7716 12316
rect 7684 12285 7685 12315
rect 7685 12285 7715 12315
rect 7715 12285 7716 12315
rect 7684 12284 7716 12285
rect 7684 12235 7716 12236
rect 7684 12205 7685 12235
rect 7685 12205 7715 12235
rect 7715 12205 7716 12235
rect 7684 12204 7716 12205
rect 7684 12155 7716 12156
rect 7684 12125 7685 12155
rect 7685 12125 7715 12155
rect 7715 12125 7716 12155
rect 7684 12124 7716 12125
rect 7684 12075 7716 12076
rect 7684 12045 7685 12075
rect 7685 12045 7715 12075
rect 7715 12045 7716 12075
rect 7684 12044 7716 12045
rect 7684 11995 7716 11996
rect 7684 11965 7685 11995
rect 7685 11965 7715 11995
rect 7715 11965 7716 11995
rect 7684 11964 7716 11965
rect 7684 11915 7716 11916
rect 7684 11885 7685 11915
rect 7685 11885 7715 11915
rect 7715 11885 7716 11915
rect 7684 11884 7716 11885
rect 7684 11835 7716 11836
rect 7684 11805 7685 11835
rect 7685 11805 7715 11835
rect 7715 11805 7716 11835
rect 7684 11804 7716 11805
rect 7684 11755 7716 11756
rect 7684 11725 7685 11755
rect 7685 11725 7715 11755
rect 7715 11725 7716 11755
rect 7684 11724 7716 11725
rect 7684 11675 7716 11676
rect 7684 11645 7685 11675
rect 7685 11645 7715 11675
rect 7715 11645 7716 11675
rect 7684 11644 7716 11645
rect 7684 11595 7716 11596
rect 7684 11565 7685 11595
rect 7685 11565 7715 11595
rect 7715 11565 7716 11595
rect 7684 11564 7716 11565
rect 7684 11515 7716 11516
rect 7684 11485 7685 11515
rect 7685 11485 7715 11515
rect 7715 11485 7716 11515
rect 7684 11484 7716 11485
rect 7684 11435 7716 11436
rect 7684 11405 7685 11435
rect 7685 11405 7715 11435
rect 7715 11405 7716 11435
rect 7684 11404 7716 11405
rect 7684 11355 7716 11356
rect 7684 11325 7685 11355
rect 7685 11325 7715 11355
rect 7715 11325 7716 11355
rect 7684 11324 7716 11325
rect 7684 11275 7716 11276
rect 7684 11245 7685 11275
rect 7685 11245 7715 11275
rect 7715 11245 7716 11275
rect 7684 11244 7716 11245
rect 7684 11195 7716 11196
rect 7684 11165 7685 11195
rect 7685 11165 7715 11195
rect 7715 11165 7716 11195
rect 7684 11164 7716 11165
rect 7684 11115 7716 11116
rect 7684 11085 7685 11115
rect 7685 11085 7715 11115
rect 7715 11085 7716 11115
rect 7684 11084 7716 11085
rect 7684 11035 7716 11036
rect 7684 11005 7685 11035
rect 7685 11005 7715 11035
rect 7715 11005 7716 11035
rect 7684 11004 7716 11005
rect 7684 10955 7716 10956
rect 7684 10925 7685 10955
rect 7685 10925 7715 10955
rect 7715 10925 7716 10955
rect 7684 10924 7716 10925
rect 7684 10875 7716 10876
rect 7684 10845 7685 10875
rect 7685 10845 7715 10875
rect 7715 10845 7716 10875
rect 7684 10844 7716 10845
rect 7684 10795 7716 10796
rect 7684 10765 7685 10795
rect 7685 10765 7715 10795
rect 7715 10765 7716 10795
rect 7684 10764 7716 10765
rect 7684 10715 7716 10716
rect 7684 10685 7685 10715
rect 7685 10685 7715 10715
rect 7715 10685 7716 10715
rect 7684 10684 7716 10685
rect 7684 10635 7716 10636
rect 7684 10605 7685 10635
rect 7685 10605 7715 10635
rect 7715 10605 7716 10635
rect 7684 10604 7716 10605
rect 7684 10555 7716 10556
rect 7684 10525 7685 10555
rect 7685 10525 7715 10555
rect 7715 10525 7716 10555
rect 7684 10524 7716 10525
rect 7684 10475 7716 10476
rect 7684 10445 7685 10475
rect 7685 10445 7715 10475
rect 7715 10445 7716 10475
rect 7684 10444 7716 10445
rect 7684 10395 7716 10396
rect 7684 10365 7685 10395
rect 7685 10365 7715 10395
rect 7715 10365 7716 10395
rect 7684 10364 7716 10365
rect 7684 10315 7716 10316
rect 7684 10285 7685 10315
rect 7685 10285 7715 10315
rect 7715 10285 7716 10315
rect 7684 10284 7716 10285
rect 7684 10235 7716 10236
rect 7684 10205 7685 10235
rect 7685 10205 7715 10235
rect 7715 10205 7716 10235
rect 7684 10204 7716 10205
rect 7684 10155 7716 10156
rect 7684 10125 7685 10155
rect 7685 10125 7715 10155
rect 7715 10125 7716 10155
rect 7684 10124 7716 10125
rect 7684 10075 7716 10076
rect 7684 10045 7685 10075
rect 7685 10045 7715 10075
rect 7715 10045 7716 10075
rect 7684 10044 7716 10045
rect 7684 9995 7716 9996
rect 7684 9965 7685 9995
rect 7685 9965 7715 9995
rect 7715 9965 7716 9995
rect 7684 9964 7716 9965
rect 7684 9915 7716 9916
rect 7684 9885 7685 9915
rect 7685 9885 7715 9915
rect 7715 9885 7716 9915
rect 7684 9884 7716 9885
rect 7684 9835 7716 9836
rect 7684 9805 7685 9835
rect 7685 9805 7715 9835
rect 7715 9805 7716 9835
rect 7684 9804 7716 9805
rect 7684 9755 7716 9756
rect 7684 9725 7685 9755
rect 7685 9725 7715 9755
rect 7715 9725 7716 9755
rect 7684 9724 7716 9725
rect 7684 9675 7716 9676
rect 7684 9645 7685 9675
rect 7685 9645 7715 9675
rect 7715 9645 7716 9675
rect 7684 9644 7716 9645
rect 7684 9595 7716 9596
rect 7684 9565 7685 9595
rect 7685 9565 7715 9595
rect 7715 9565 7716 9595
rect 7684 9564 7716 9565
rect 7684 9515 7716 9516
rect 7684 9485 7685 9515
rect 7685 9485 7715 9515
rect 7715 9485 7716 9515
rect 7684 9484 7716 9485
rect 7684 9435 7716 9436
rect 7684 9405 7685 9435
rect 7685 9405 7715 9435
rect 7715 9405 7716 9435
rect 7684 9404 7716 9405
rect 7684 9355 7716 9356
rect 7684 9325 7685 9355
rect 7685 9325 7715 9355
rect 7715 9325 7716 9355
rect 7684 9324 7716 9325
rect 7684 9275 7716 9276
rect 7684 9245 7685 9275
rect 7685 9245 7715 9275
rect 7715 9245 7716 9275
rect 7684 9244 7716 9245
rect 7684 9195 7716 9196
rect 7684 9165 7685 9195
rect 7685 9165 7715 9195
rect 7715 9165 7716 9195
rect 7684 9164 7716 9165
rect 7684 9115 7716 9116
rect 7684 9085 7685 9115
rect 7685 9085 7715 9115
rect 7715 9085 7716 9115
rect 7684 9084 7716 9085
rect 7684 9035 7716 9036
rect 7684 9005 7685 9035
rect 7685 9005 7715 9035
rect 7715 9005 7716 9035
rect 7684 9004 7716 9005
rect 7684 8955 7716 8956
rect 7684 8925 7685 8955
rect 7685 8925 7715 8955
rect 7715 8925 7716 8955
rect 7684 8924 7716 8925
rect 7684 8635 7716 8636
rect 7684 8605 7685 8635
rect 7685 8605 7715 8635
rect 7715 8605 7716 8635
rect 7684 8604 7716 8605
rect 7684 8555 7716 8556
rect 7684 8525 7685 8555
rect 7685 8525 7715 8555
rect 7715 8525 7716 8555
rect 7684 8524 7716 8525
rect 7684 8475 7716 8476
rect 7684 8445 7685 8475
rect 7685 8445 7715 8475
rect 7715 8445 7716 8475
rect 7684 8444 7716 8445
rect 7684 8395 7716 8396
rect 7684 8365 7685 8395
rect 7685 8365 7715 8395
rect 7715 8365 7716 8395
rect 7684 8364 7716 8365
rect 7684 8315 7716 8316
rect 7684 8285 7685 8315
rect 7685 8285 7715 8315
rect 7715 8285 7716 8315
rect 7684 8284 7716 8285
rect 7684 8235 7716 8236
rect 7684 8205 7685 8235
rect 7685 8205 7715 8235
rect 7715 8205 7716 8235
rect 7684 8204 7716 8205
rect 7684 8155 7716 8156
rect 7684 8125 7685 8155
rect 7685 8125 7715 8155
rect 7715 8125 7716 8155
rect 7684 8124 7716 8125
rect 7684 8075 7716 8076
rect 7684 8045 7685 8075
rect 7685 8045 7715 8075
rect 7715 8045 7716 8075
rect 7684 8044 7716 8045
rect 7684 7995 7716 7996
rect 7684 7965 7685 7995
rect 7685 7965 7715 7995
rect 7715 7965 7716 7995
rect 7684 7964 7716 7965
rect 7684 7915 7716 7916
rect 7684 7885 7685 7915
rect 7685 7885 7715 7915
rect 7715 7885 7716 7915
rect 7684 7884 7716 7885
rect 7684 7835 7716 7836
rect 7684 7805 7685 7835
rect 7685 7805 7715 7835
rect 7715 7805 7716 7835
rect 7684 7804 7716 7805
rect 7684 7755 7716 7756
rect 7684 7725 7685 7755
rect 7685 7725 7715 7755
rect 7715 7725 7716 7755
rect 7684 7724 7716 7725
rect 7684 7675 7716 7676
rect 7684 7645 7685 7675
rect 7685 7645 7715 7675
rect 7715 7645 7716 7675
rect 7684 7644 7716 7645
rect 7684 7595 7716 7596
rect 7684 7565 7685 7595
rect 7685 7565 7715 7595
rect 7715 7565 7716 7595
rect 7684 7564 7716 7565
rect 7684 7515 7716 7516
rect 7684 7485 7685 7515
rect 7685 7485 7715 7515
rect 7715 7485 7716 7515
rect 7684 7484 7716 7485
rect 7684 7435 7716 7436
rect 7684 7405 7685 7435
rect 7685 7405 7715 7435
rect 7715 7405 7716 7435
rect 7684 7404 7716 7405
rect 7684 7355 7716 7356
rect 7684 7325 7685 7355
rect 7685 7325 7715 7355
rect 7715 7325 7716 7355
rect 7684 7324 7716 7325
rect 7684 7275 7716 7276
rect 7684 7245 7685 7275
rect 7685 7245 7715 7275
rect 7715 7245 7716 7275
rect 7684 7244 7716 7245
rect 7684 7195 7716 7196
rect 7684 7165 7685 7195
rect 7685 7165 7715 7195
rect 7715 7165 7716 7195
rect 7684 7164 7716 7165
rect 7684 7115 7716 7116
rect 7684 7085 7685 7115
rect 7685 7085 7715 7115
rect 7715 7085 7716 7115
rect 7684 7084 7716 7085
rect 7684 7035 7716 7036
rect 7684 7005 7685 7035
rect 7685 7005 7715 7035
rect 7715 7005 7716 7035
rect 7684 7004 7716 7005
rect 7684 6955 7716 6956
rect 7684 6925 7685 6955
rect 7685 6925 7715 6955
rect 7715 6925 7716 6955
rect 7684 6924 7716 6925
rect 7684 6875 7716 6876
rect 7684 6845 7685 6875
rect 7685 6845 7715 6875
rect 7715 6845 7716 6875
rect 7684 6844 7716 6845
rect 7684 6795 7716 6796
rect 7684 6765 7685 6795
rect 7685 6765 7715 6795
rect 7715 6765 7716 6795
rect 7684 6764 7716 6765
rect 7684 6715 7716 6716
rect 7684 6685 7685 6715
rect 7685 6685 7715 6715
rect 7715 6685 7716 6715
rect 7684 6684 7716 6685
rect 7684 6635 7716 6636
rect 7684 6605 7685 6635
rect 7685 6605 7715 6635
rect 7715 6605 7716 6635
rect 7684 6604 7716 6605
rect 7684 6555 7716 6556
rect 7684 6525 7685 6555
rect 7685 6525 7715 6555
rect 7715 6525 7716 6555
rect 7684 6524 7716 6525
rect 7684 6475 7716 6476
rect 7684 6445 7685 6475
rect 7685 6445 7715 6475
rect 7715 6445 7716 6475
rect 7684 6444 7716 6445
rect 7684 6395 7716 6396
rect 7684 6365 7685 6395
rect 7685 6365 7715 6395
rect 7715 6365 7716 6395
rect 7684 6364 7716 6365
rect 7684 6315 7716 6316
rect 7684 6285 7685 6315
rect 7685 6285 7715 6315
rect 7715 6285 7716 6315
rect 7684 6284 7716 6285
rect 7684 6235 7716 6236
rect 7684 6205 7685 6235
rect 7685 6205 7715 6235
rect 7715 6205 7716 6235
rect 7684 6204 7716 6205
rect 7684 6155 7716 6156
rect 7684 6125 7685 6155
rect 7685 6125 7715 6155
rect 7715 6125 7716 6155
rect 7684 6124 7716 6125
rect 7684 6075 7716 6076
rect 7684 6045 7685 6075
rect 7685 6045 7715 6075
rect 7715 6045 7716 6075
rect 7684 6044 7716 6045
rect 7684 5995 7716 5996
rect 7684 5965 7685 5995
rect 7685 5965 7715 5995
rect 7715 5965 7716 5995
rect 7684 5964 7716 5965
rect 7684 5915 7716 5916
rect 7684 5885 7685 5915
rect 7685 5885 7715 5915
rect 7715 5885 7716 5915
rect 7684 5884 7716 5885
rect 7684 5835 7716 5836
rect 7684 5805 7685 5835
rect 7685 5805 7715 5835
rect 7715 5805 7716 5835
rect 7684 5804 7716 5805
rect 7684 5755 7716 5756
rect 7684 5725 7685 5755
rect 7685 5725 7715 5755
rect 7715 5725 7716 5755
rect 7684 5724 7716 5725
rect 7684 5675 7716 5676
rect 7684 5645 7685 5675
rect 7685 5645 7715 5675
rect 7715 5645 7716 5675
rect 7684 5644 7716 5645
rect 7684 5595 7716 5596
rect 7684 5565 7685 5595
rect 7685 5565 7715 5595
rect 7715 5565 7716 5595
rect 7684 5564 7716 5565
rect 7684 5515 7716 5516
rect 7684 5485 7685 5515
rect 7685 5485 7715 5515
rect 7715 5485 7716 5515
rect 7684 5484 7716 5485
rect 7684 5435 7716 5436
rect 7684 5405 7685 5435
rect 7685 5405 7715 5435
rect 7715 5405 7716 5435
rect 7684 5404 7716 5405
rect 7684 5355 7716 5356
rect 7684 5325 7685 5355
rect 7685 5325 7715 5355
rect 7715 5325 7716 5355
rect 7684 5324 7716 5325
rect 7684 5275 7716 5276
rect 7684 5245 7685 5275
rect 7685 5245 7715 5275
rect 7715 5245 7716 5275
rect 7684 5244 7716 5245
rect 7684 5195 7716 5196
rect 7684 5165 7685 5195
rect 7685 5165 7715 5195
rect 7715 5165 7716 5195
rect 7684 5164 7716 5165
rect 7684 5115 7716 5116
rect 7684 5085 7685 5115
rect 7685 5085 7715 5115
rect 7715 5085 7716 5115
rect 7684 5084 7716 5085
rect 7684 5035 7716 5036
rect 7684 5005 7685 5035
rect 7685 5005 7715 5035
rect 7715 5005 7716 5035
rect 7684 5004 7716 5005
rect 7684 4955 7716 4956
rect 7684 4925 7685 4955
rect 7685 4925 7715 4955
rect 7715 4925 7716 4955
rect 7684 4924 7716 4925
rect 7684 4875 7716 4876
rect 7684 4845 7685 4875
rect 7685 4845 7715 4875
rect 7715 4845 7716 4875
rect 7684 4844 7716 4845
rect 7684 4795 7716 4796
rect 7684 4765 7685 4795
rect 7685 4765 7715 4795
rect 7715 4765 7716 4795
rect 7684 4764 7716 4765
rect 7684 4715 7716 4716
rect 7684 4685 7685 4715
rect 7685 4685 7715 4715
rect 7715 4685 7716 4715
rect 7684 4684 7716 4685
rect 7684 4635 7716 4636
rect 7684 4605 7685 4635
rect 7685 4605 7715 4635
rect 7715 4605 7716 4635
rect 7684 4604 7716 4605
rect 7684 4555 7716 4556
rect 7684 4525 7685 4555
rect 7685 4525 7715 4555
rect 7715 4525 7716 4555
rect 7684 4524 7716 4525
rect 7684 4475 7716 4476
rect 7684 4445 7685 4475
rect 7685 4445 7715 4475
rect 7715 4445 7716 4475
rect 7684 4444 7716 4445
rect 7684 4395 7716 4396
rect 7684 4365 7685 4395
rect 7685 4365 7715 4395
rect 7715 4365 7716 4395
rect 7684 4364 7716 4365
rect 7684 4315 7716 4316
rect 7684 4285 7685 4315
rect 7685 4285 7715 4315
rect 7715 4285 7716 4315
rect 7684 4284 7716 4285
rect 7684 4235 7716 4236
rect 7684 4205 7685 4235
rect 7685 4205 7715 4235
rect 7715 4205 7716 4235
rect 7684 4204 7716 4205
rect 7684 4155 7716 4156
rect 7684 4125 7685 4155
rect 7685 4125 7715 4155
rect 7715 4125 7716 4155
rect 7684 4124 7716 4125
rect 7684 4075 7716 4076
rect 7684 4045 7685 4075
rect 7685 4045 7715 4075
rect 7715 4045 7716 4075
rect 7684 4044 7716 4045
rect 7684 3995 7716 3996
rect 7684 3965 7685 3995
rect 7685 3965 7715 3995
rect 7715 3965 7716 3995
rect 7684 3964 7716 3965
rect 7684 3915 7716 3916
rect 7684 3885 7685 3915
rect 7685 3885 7715 3915
rect 7715 3885 7716 3915
rect 7684 3884 7716 3885
rect 7684 3835 7716 3836
rect 7684 3805 7685 3835
rect 7685 3805 7715 3835
rect 7715 3805 7716 3835
rect 7684 3804 7716 3805
rect 7684 3755 7716 3756
rect 7684 3725 7685 3755
rect 7685 3725 7715 3755
rect 7715 3725 7716 3755
rect 7684 3724 7716 3725
rect 7684 3675 7716 3676
rect 7684 3645 7685 3675
rect 7685 3645 7715 3675
rect 7715 3645 7716 3675
rect 7684 3644 7716 3645
rect 7684 3595 7716 3596
rect 7684 3565 7685 3595
rect 7685 3565 7715 3595
rect 7715 3565 7716 3595
rect 7684 3564 7716 3565
rect 7684 3515 7716 3516
rect 7684 3485 7685 3515
rect 7685 3485 7715 3515
rect 7715 3485 7716 3515
rect 7684 3484 7716 3485
rect 7684 3435 7716 3436
rect 7684 3405 7685 3435
rect 7685 3405 7715 3435
rect 7715 3405 7716 3435
rect 7684 3404 7716 3405
rect 7684 3355 7716 3356
rect 7684 3325 7685 3355
rect 7685 3325 7715 3355
rect 7715 3325 7716 3355
rect 7684 3324 7716 3325
rect 7684 3275 7716 3276
rect 7684 3245 7685 3275
rect 7685 3245 7715 3275
rect 7715 3245 7716 3275
rect 7684 3244 7716 3245
rect 7684 3195 7716 3196
rect 7684 3165 7685 3195
rect 7685 3165 7715 3195
rect 7715 3165 7716 3195
rect 7684 3164 7716 3165
rect 7684 3115 7716 3116
rect 7684 3085 7685 3115
rect 7685 3085 7715 3115
rect 7715 3085 7716 3115
rect 7684 3084 7716 3085
rect 7684 3035 7716 3036
rect 7684 3005 7685 3035
rect 7685 3005 7715 3035
rect 7715 3005 7716 3035
rect 7684 3004 7716 3005
rect 7684 2955 7716 2956
rect 7684 2925 7685 2955
rect 7685 2925 7715 2955
rect 7715 2925 7716 2955
rect 7684 2924 7716 2925
rect 7684 2875 7716 2876
rect 7684 2845 7685 2875
rect 7685 2845 7715 2875
rect 7715 2845 7716 2875
rect 7684 2844 7716 2845
rect 7684 2795 7716 2796
rect 7684 2765 7685 2795
rect 7685 2765 7715 2795
rect 7715 2765 7716 2795
rect 7684 2764 7716 2765
rect 7684 2715 7716 2716
rect 7684 2685 7685 2715
rect 7685 2685 7715 2715
rect 7715 2685 7716 2715
rect 7684 2684 7716 2685
rect 7684 2635 7716 2636
rect 7684 2605 7685 2635
rect 7685 2605 7715 2635
rect 7715 2605 7716 2635
rect 7684 2604 7716 2605
rect 7684 2555 7716 2556
rect 7684 2525 7685 2555
rect 7685 2525 7715 2555
rect 7715 2525 7716 2555
rect 7684 2524 7716 2525
rect 7684 2475 7716 2476
rect 7684 2445 7685 2475
rect 7685 2445 7715 2475
rect 7715 2445 7716 2475
rect 7684 2444 7716 2445
rect 7684 2395 7716 2396
rect 7684 2365 7685 2395
rect 7685 2365 7715 2395
rect 7715 2365 7716 2395
rect 7684 2364 7716 2365
rect 7684 2315 7716 2316
rect 7684 2285 7685 2315
rect 7685 2285 7715 2315
rect 7715 2285 7716 2315
rect 7684 2284 7716 2285
rect 7684 2235 7716 2236
rect 7684 2205 7685 2235
rect 7685 2205 7715 2235
rect 7715 2205 7716 2235
rect 7684 2204 7716 2205
rect 7684 2155 7716 2156
rect 7684 2125 7685 2155
rect 7685 2125 7715 2155
rect 7715 2125 7716 2155
rect 7684 2124 7716 2125
rect 7684 2075 7716 2076
rect 7684 2045 7685 2075
rect 7685 2045 7715 2075
rect 7715 2045 7716 2075
rect 7684 2044 7716 2045
rect 7684 1995 7716 1996
rect 7684 1965 7685 1995
rect 7685 1965 7715 1995
rect 7715 1965 7716 1995
rect 7684 1964 7716 1965
rect 7684 1915 7716 1916
rect 7684 1885 7685 1915
rect 7685 1885 7715 1915
rect 7715 1885 7716 1915
rect 7684 1884 7716 1885
rect 7684 1835 7716 1836
rect 7684 1805 7685 1835
rect 7685 1805 7715 1835
rect 7715 1805 7716 1835
rect 7684 1804 7716 1805
rect 7684 1755 7716 1756
rect 7684 1725 7685 1755
rect 7685 1725 7715 1755
rect 7715 1725 7716 1755
rect 7684 1724 7716 1725
rect 7684 1675 7716 1676
rect 7684 1645 7685 1675
rect 7685 1645 7715 1675
rect 7715 1645 7716 1675
rect 7684 1644 7716 1645
rect 7684 1595 7716 1596
rect 7684 1565 7685 1595
rect 7685 1565 7715 1595
rect 7715 1565 7716 1595
rect 7684 1564 7716 1565
rect 7684 1515 7716 1516
rect 7684 1485 7685 1515
rect 7685 1485 7715 1515
rect 7715 1485 7716 1515
rect 7684 1484 7716 1485
rect 7684 1435 7716 1436
rect 7684 1405 7685 1435
rect 7685 1405 7715 1435
rect 7715 1405 7716 1435
rect 7684 1404 7716 1405
rect 7684 1355 7716 1356
rect 7684 1325 7685 1355
rect 7685 1325 7715 1355
rect 7715 1325 7716 1355
rect 7684 1324 7716 1325
rect 7684 1275 7716 1276
rect 7684 1245 7685 1275
rect 7685 1245 7715 1275
rect 7715 1245 7716 1275
rect 7684 1244 7716 1245
rect 7684 1195 7716 1196
rect 7684 1165 7685 1195
rect 7685 1165 7715 1195
rect 7715 1165 7716 1195
rect 7684 1164 7716 1165
rect 7684 1115 7716 1116
rect 7684 1085 7685 1115
rect 7685 1085 7715 1115
rect 7715 1085 7716 1115
rect 7684 1084 7716 1085
rect 7684 1035 7716 1036
rect 7684 1005 7685 1035
rect 7685 1005 7715 1035
rect 7715 1005 7716 1035
rect 7684 1004 7716 1005
rect 7684 955 7716 956
rect 7684 925 7685 955
rect 7685 925 7715 955
rect 7715 925 7716 955
rect 7684 924 7716 925
rect 7684 875 7716 876
rect 7684 845 7685 875
rect 7685 845 7715 875
rect 7715 845 7716 875
rect 7684 844 7716 845
rect 7684 795 7716 796
rect 7684 765 7685 795
rect 7685 765 7715 795
rect 7715 765 7716 795
rect 7684 764 7716 765
rect 7684 715 7716 716
rect 7684 685 7685 715
rect 7685 685 7715 715
rect 7715 685 7716 715
rect 7684 684 7716 685
rect 7684 595 7716 596
rect 7684 565 7685 595
rect 7685 565 7715 595
rect 7715 565 7716 595
rect 7684 564 7716 565
rect 7684 515 7716 516
rect 7684 485 7685 515
rect 7685 485 7715 515
rect 7715 485 7716 515
rect 7684 484 7716 485
rect 7684 435 7716 436
rect 7684 405 7685 435
rect 7685 405 7715 435
rect 7715 405 7716 435
rect 7684 404 7716 405
rect 7684 355 7716 356
rect 7684 325 7685 355
rect 7685 325 7715 355
rect 7715 325 7716 355
rect 7684 324 7716 325
rect 7684 275 7716 276
rect 7684 245 7685 275
rect 7685 245 7715 275
rect 7715 245 7716 275
rect 7684 244 7716 245
rect 7684 195 7716 196
rect 7684 165 7685 195
rect 7685 165 7715 195
rect 7715 165 7716 195
rect 7684 164 7716 165
rect 7684 115 7716 116
rect 7684 85 7685 115
rect 7685 85 7715 115
rect 7715 85 7716 115
rect 7684 84 7716 85
rect 7684 35 7716 36
rect 7684 5 7685 35
rect 7685 5 7715 35
rect 7715 5 7716 35
rect 7684 4 7716 5
<< mimcap >>
rect 600 19480 1600 19520
rect 600 18560 640 19480
rect 1560 18560 1600 19480
rect 600 18520 1600 18560
rect 1720 19480 2720 19520
rect 1720 18560 1760 19480
rect 2680 18560 2720 19480
rect 1720 18520 2720 18560
rect 2840 19480 3840 19520
rect 2840 18560 2880 19480
rect 3800 18560 3840 19480
rect 2840 18520 3840 18560
rect 3960 19480 4960 19520
rect 3960 18560 4000 19480
rect 4920 18560 4960 19480
rect 3960 18520 4960 18560
rect 5080 19480 6080 19520
rect 5080 18560 5120 19480
rect 6040 18560 6080 19480
rect 5080 18520 6080 18560
rect 6200 19480 7200 19520
rect 6200 18560 6240 19480
rect 7160 18560 7200 19480
rect 6200 18520 7200 18560
rect 600 18360 1600 18400
rect 600 17440 640 18360
rect 1560 17440 1600 18360
rect 600 17400 1600 17440
rect 1720 18360 2720 18400
rect 1720 17440 1760 18360
rect 2680 17440 2720 18360
rect 1720 17400 2720 17440
rect 2840 18360 3840 18400
rect 2840 17440 2880 18360
rect 3800 17440 3840 18360
rect 2840 17400 3840 17440
rect 3960 18360 4960 18400
rect 3960 17440 4000 18360
rect 4920 17440 4960 18360
rect 3960 17400 4960 17440
rect 5080 18360 6080 18400
rect 5080 17440 5120 18360
rect 6040 17440 6080 18360
rect 5080 17400 6080 17440
rect 6200 18360 7200 18400
rect 6200 17440 6240 18360
rect 7160 17440 7200 18360
rect 6200 17400 7200 17440
<< mimcapcontact >>
rect 640 18560 1560 19480
rect 1760 18560 2680 19480
rect 2880 18560 3800 19480
rect 4000 18560 4920 19480
rect 5120 18560 6040 19480
rect 6240 18560 7160 19480
rect 640 17440 1560 18360
rect 1760 17440 2680 18360
rect 2880 17440 3800 18360
rect 4000 17440 4920 18360
rect 5120 17440 6040 18360
rect 6240 17440 7160 18360
<< metal4 >>
rect 400 19760 7800 19800
rect 400 17160 440 19760
rect 480 19716 7800 19720
rect 480 19684 7364 19716
rect 7396 19684 7524 19716
rect 7556 19684 7684 19716
rect 7716 19684 7800 19716
rect 480 19680 7800 19684
rect 480 17240 520 19680
rect 560 19636 7480 19640
rect 560 19604 564 19636
rect 1636 19604 1684 19636
rect 2756 19604 2804 19636
rect 3876 19604 3924 19636
rect 4996 19604 5044 19636
rect 6116 19604 6164 19636
rect 7236 19604 7444 19636
rect 7476 19604 7480 19636
rect 560 19600 7480 19604
rect 560 19480 1640 19560
rect 560 18560 640 19480
rect 1560 18560 1640 19480
rect 560 18520 1640 18560
rect 1680 19480 2760 19560
rect 1680 18560 1760 19480
rect 2680 18560 2760 19480
rect 1680 18520 2760 18560
rect 2800 19480 3880 19560
rect 2800 18560 2880 19480
rect 3800 18560 3880 19480
rect 2800 18520 3880 18560
rect 3920 19480 5000 19560
rect 3920 18560 4000 19480
rect 4920 18560 5000 19480
rect 3920 18520 5000 18560
rect 5040 19480 6120 19560
rect 5040 18560 5120 19480
rect 6040 18560 6120 19480
rect 5040 18520 6120 18560
rect 6160 19480 7240 19560
rect 6160 18560 6240 19480
rect 7160 18560 7240 19480
rect 6160 18520 7240 18560
rect 560 18516 7720 18520
rect 560 18484 7364 18516
rect 7396 18484 7524 18516
rect 7556 18484 7684 18516
rect 7716 18484 7720 18516
rect 560 18480 7720 18484
rect 560 18440 600 18480
rect 1600 18440 1640 18480
rect 1680 18440 1720 18480
rect 2720 18440 2760 18480
rect 2800 18440 2840 18480
rect 3840 18440 3880 18480
rect 3920 18440 3960 18480
rect 4960 18440 5000 18480
rect 5040 18440 5080 18480
rect 6080 18440 6120 18480
rect 6160 18440 6200 18480
rect 7200 18440 7240 18480
rect 560 18436 7720 18440
rect 560 18404 7364 18436
rect 7396 18404 7524 18436
rect 7556 18404 7684 18436
rect 7716 18404 7720 18436
rect 560 18400 7720 18404
rect 560 18360 1640 18400
rect 560 17440 640 18360
rect 1560 17440 1640 18360
rect 560 17360 1640 17440
rect 1680 18360 2760 18400
rect 1680 17440 1760 18360
rect 2680 17440 2760 18360
rect 1680 17360 2760 17440
rect 2800 18360 3880 18400
rect 2800 17440 2880 18360
rect 3800 17440 3880 18360
rect 2800 17360 3880 17440
rect 3920 18360 5000 18400
rect 3920 17440 4000 18360
rect 4920 17440 5000 18360
rect 3920 17360 5000 17440
rect 5040 18360 6120 18400
rect 5040 17440 5120 18360
rect 6040 17440 6120 18360
rect 5040 17360 6120 17440
rect 6160 18360 7240 18400
rect 6160 17440 6240 18360
rect 7160 17440 7240 18360
rect 6160 17360 7240 17440
rect 560 17316 7640 17320
rect 560 17284 564 17316
rect 1636 17284 1684 17316
rect 2756 17284 2804 17316
rect 3876 17284 3924 17316
rect 4996 17284 5044 17316
rect 6116 17284 6164 17316
rect 7236 17284 7604 17316
rect 7636 17284 7640 17316
rect 560 17280 7640 17284
rect 480 17200 7800 17240
rect 400 17156 7800 17160
rect 400 17124 7284 17156
rect 7316 17124 7800 17156
rect 400 17120 7800 17124
rect 0 17040 7800 17080
rect 0 16920 120 17040
rect 240 16920 7800 17040
rect 0 16880 7800 16920
rect 0 16836 7800 16840
rect 0 16800 5524 16836
rect 0 16680 760 16800
rect 880 16680 5524 16800
rect 0 16644 5524 16680
rect 5556 16644 5684 16836
rect 5716 16644 5844 16836
rect 5876 16644 6004 16836
rect 6036 16644 6164 16836
rect 6196 16644 6324 16836
rect 6356 16644 6484 16836
rect 6516 16644 6644 16836
rect 6676 16644 6804 16836
rect 6836 16644 6964 16836
rect 6996 16644 7124 16836
rect 7156 16644 7284 16836
rect 7316 16644 7764 16836
rect 7796 16644 7800 16836
rect 0 16640 7800 16644
rect 5520 16596 7320 16600
rect 5520 16564 5524 16596
rect 5556 16564 5684 16596
rect 5716 16564 5844 16596
rect 5876 16564 6004 16596
rect 6036 16564 6164 16596
rect 6196 16564 6324 16596
rect 6356 16564 6484 16596
rect 6516 16564 6644 16596
rect 6676 16564 6804 16596
rect 6836 16564 6964 16596
rect 6996 16564 7124 16596
rect 7156 16564 7284 16596
rect 7316 16564 7320 16596
rect 5520 16560 7320 16564
rect 7360 16596 7720 16600
rect 7360 16564 7364 16596
rect 7396 16564 7524 16596
rect 7556 16564 7684 16596
rect 7716 16564 7720 16596
rect 7360 16560 7720 16564
rect 5520 16516 7320 16520
rect 5520 16484 5524 16516
rect 5556 16484 5684 16516
rect 5716 16484 5844 16516
rect 5876 16484 6004 16516
rect 6036 16484 6164 16516
rect 6196 16484 6324 16516
rect 6356 16484 6484 16516
rect 6516 16484 6644 16516
rect 6676 16484 6804 16516
rect 6836 16484 6964 16516
rect 6996 16484 7124 16516
rect 7156 16484 7284 16516
rect 7316 16484 7320 16516
rect 5520 16480 7320 16484
rect 7360 16516 7720 16520
rect 7360 16484 7364 16516
rect 7396 16484 7524 16516
rect 7556 16484 7684 16516
rect 7716 16484 7720 16516
rect 7360 16480 7720 16484
rect 5520 16436 7320 16440
rect 5520 16404 5524 16436
rect 5556 16404 5684 16436
rect 5716 16404 5844 16436
rect 5876 16404 6004 16436
rect 6036 16404 6164 16436
rect 6196 16404 6324 16436
rect 6356 16404 6484 16436
rect 6516 16404 6644 16436
rect 6676 16404 6804 16436
rect 6836 16404 6964 16436
rect 6996 16404 7124 16436
rect 7156 16404 7284 16436
rect 7316 16404 7320 16436
rect 5520 16400 7320 16404
rect 7360 16436 7720 16440
rect 7360 16404 7364 16436
rect 7396 16404 7524 16436
rect 7556 16404 7684 16436
rect 7716 16404 7720 16436
rect 7360 16400 7720 16404
rect 5520 16356 7320 16360
rect 5520 16324 5524 16356
rect 5556 16324 5684 16356
rect 5716 16324 5844 16356
rect 5876 16324 6004 16356
rect 6036 16324 6164 16356
rect 6196 16324 6324 16356
rect 6356 16324 6484 16356
rect 6516 16324 6644 16356
rect 6676 16324 6804 16356
rect 6836 16324 6964 16356
rect 6996 16324 7124 16356
rect 7156 16324 7284 16356
rect 7316 16324 7320 16356
rect 5520 16320 7320 16324
rect 7360 16356 7720 16360
rect 7360 16324 7364 16356
rect 7396 16324 7524 16356
rect 7556 16324 7684 16356
rect 7716 16324 7720 16356
rect 7360 16320 7720 16324
rect 5520 16276 7320 16280
rect 5520 16244 5524 16276
rect 5556 16244 5684 16276
rect 5716 16244 5844 16276
rect 5876 16244 6004 16276
rect 6036 16244 6164 16276
rect 6196 16244 6324 16276
rect 6356 16244 6484 16276
rect 6516 16244 6644 16276
rect 6676 16244 6804 16276
rect 6836 16244 6964 16276
rect 6996 16244 7124 16276
rect 7156 16244 7284 16276
rect 7316 16244 7320 16276
rect 5520 16240 7320 16244
rect 7360 16276 7720 16280
rect 7360 16244 7364 16276
rect 7396 16244 7524 16276
rect 7556 16244 7684 16276
rect 7716 16244 7720 16276
rect 7360 16240 7720 16244
rect 5520 16196 7320 16200
rect 5520 16164 5524 16196
rect 5556 16164 5684 16196
rect 5716 16164 5844 16196
rect 5876 16164 6004 16196
rect 6036 16164 6164 16196
rect 6196 16164 6324 16196
rect 6356 16164 6484 16196
rect 6516 16164 6644 16196
rect 6676 16164 6804 16196
rect 6836 16164 6964 16196
rect 6996 16164 7124 16196
rect 7156 16164 7284 16196
rect 7316 16164 7320 16196
rect 5520 16160 7320 16164
rect 7360 16196 7720 16200
rect 7360 16164 7364 16196
rect 7396 16164 7524 16196
rect 7556 16164 7684 16196
rect 7716 16164 7720 16196
rect 7360 16160 7720 16164
rect 5520 16116 7320 16120
rect 5520 16084 5524 16116
rect 5556 16084 5684 16116
rect 5716 16084 5844 16116
rect 5876 16084 6004 16116
rect 6036 16084 6164 16116
rect 6196 16084 6324 16116
rect 6356 16084 6484 16116
rect 6516 16084 6644 16116
rect 6676 16084 6804 16116
rect 6836 16084 6964 16116
rect 6996 16084 7124 16116
rect 7156 16084 7284 16116
rect 7316 16084 7320 16116
rect 5520 16080 7320 16084
rect 7360 16116 7720 16120
rect 7360 16084 7364 16116
rect 7396 16084 7524 16116
rect 7556 16084 7684 16116
rect 7716 16084 7720 16116
rect 7360 16080 7720 16084
rect 5520 16036 7320 16040
rect 5520 16004 5524 16036
rect 5556 16004 5684 16036
rect 5716 16004 5844 16036
rect 5876 16004 6004 16036
rect 6036 16004 6164 16036
rect 6196 16004 6324 16036
rect 6356 16004 6484 16036
rect 6516 16004 6644 16036
rect 6676 16004 6804 16036
rect 6836 16004 6964 16036
rect 6996 16004 7124 16036
rect 7156 16004 7284 16036
rect 7316 16004 7320 16036
rect 5520 16000 7320 16004
rect 7360 16036 7720 16040
rect 7360 16004 7364 16036
rect 7396 16004 7524 16036
rect 7556 16004 7684 16036
rect 7716 16004 7720 16036
rect 7360 16000 7720 16004
rect 5520 15956 7320 15960
rect 5520 15924 5524 15956
rect 5556 15924 5684 15956
rect 5716 15924 5844 15956
rect 5876 15924 6004 15956
rect 6036 15924 6164 15956
rect 6196 15924 6324 15956
rect 6356 15924 6484 15956
rect 6516 15924 6644 15956
rect 6676 15924 6804 15956
rect 6836 15924 6964 15956
rect 6996 15924 7124 15956
rect 7156 15924 7284 15956
rect 7316 15924 7320 15956
rect 5520 15920 7320 15924
rect 7360 15956 7720 15960
rect 7360 15924 7364 15956
rect 7396 15924 7524 15956
rect 7556 15924 7684 15956
rect 7716 15924 7720 15956
rect 7360 15920 7720 15924
rect 5520 15436 7320 15440
rect 5520 15404 5524 15436
rect 5556 15404 5684 15436
rect 5716 15404 5844 15436
rect 5876 15404 6004 15436
rect 6036 15404 6164 15436
rect 6196 15404 6324 15436
rect 6356 15404 6484 15436
rect 6516 15404 6644 15436
rect 6676 15404 6804 15436
rect 6836 15404 6964 15436
rect 6996 15404 7124 15436
rect 7156 15404 7284 15436
rect 7316 15404 7320 15436
rect 5520 15400 7320 15404
rect 7360 15436 7720 15440
rect 7360 15404 7364 15436
rect 7396 15404 7524 15436
rect 7556 15404 7684 15436
rect 7716 15404 7720 15436
rect 7360 15400 7720 15404
rect 5520 15356 7320 15360
rect 5520 15324 5524 15356
rect 5556 15324 5684 15356
rect 5716 15324 5844 15356
rect 5876 15324 6004 15356
rect 6036 15324 6164 15356
rect 6196 15324 6324 15356
rect 6356 15324 6484 15356
rect 6516 15324 6644 15356
rect 6676 15324 6804 15356
rect 6836 15324 6964 15356
rect 6996 15324 7124 15356
rect 7156 15324 7284 15356
rect 7316 15324 7320 15356
rect 5520 15320 7320 15324
rect 7360 15356 7720 15360
rect 7360 15324 7364 15356
rect 7396 15324 7524 15356
rect 7556 15324 7684 15356
rect 7716 15324 7720 15356
rect 7360 15320 7720 15324
rect 5520 15276 7320 15280
rect 5520 15244 5524 15276
rect 5556 15244 5684 15276
rect 5716 15244 5844 15276
rect 5876 15244 6004 15276
rect 6036 15244 6164 15276
rect 6196 15244 6324 15276
rect 6356 15244 6484 15276
rect 6516 15244 6644 15276
rect 6676 15244 6804 15276
rect 6836 15244 6964 15276
rect 6996 15244 7124 15276
rect 7156 15244 7284 15276
rect 7316 15244 7320 15276
rect 5520 15240 7320 15244
rect 7360 15276 7720 15280
rect 7360 15244 7364 15276
rect 7396 15244 7524 15276
rect 7556 15244 7684 15276
rect 7716 15244 7720 15276
rect 7360 15240 7720 15244
rect 5520 15196 7320 15200
rect 5520 15164 5524 15196
rect 5556 15164 5684 15196
rect 5716 15164 5844 15196
rect 5876 15164 6004 15196
rect 6036 15164 6164 15196
rect 6196 15164 6324 15196
rect 6356 15164 6484 15196
rect 6516 15164 6644 15196
rect 6676 15164 6804 15196
rect 6836 15164 6964 15196
rect 6996 15164 7124 15196
rect 7156 15164 7284 15196
rect 7316 15164 7320 15196
rect 5520 15160 7320 15164
rect 7360 15196 7720 15200
rect 7360 15164 7364 15196
rect 7396 15164 7524 15196
rect 7556 15164 7684 15196
rect 7716 15164 7720 15196
rect 7360 15160 7720 15164
rect 5520 15116 7320 15120
rect 5520 15084 5524 15116
rect 5556 15084 5684 15116
rect 5716 15084 5844 15116
rect 5876 15084 6004 15116
rect 6036 15084 6164 15116
rect 6196 15084 6324 15116
rect 6356 15084 6484 15116
rect 6516 15084 6644 15116
rect 6676 15084 6804 15116
rect 6836 15084 6964 15116
rect 6996 15084 7124 15116
rect 7156 15084 7284 15116
rect 7316 15084 7320 15116
rect 5520 15080 7320 15084
rect 7360 15116 7720 15120
rect 7360 15084 7364 15116
rect 7396 15084 7524 15116
rect 7556 15084 7684 15116
rect 7716 15084 7720 15116
rect 7360 15080 7720 15084
rect 6160 15036 7320 15040
rect 6160 15004 6164 15036
rect 6196 15004 6324 15036
rect 6356 15004 6484 15036
rect 6516 15004 6644 15036
rect 6676 15004 6804 15036
rect 6836 15004 6964 15036
rect 6996 15004 7124 15036
rect 7156 15004 7284 15036
rect 7316 15004 7320 15036
rect 6160 15000 7320 15004
rect 7360 15036 7720 15040
rect 7360 15004 7364 15036
rect 7396 15004 7524 15036
rect 7556 15004 7684 15036
rect 7716 15004 7720 15036
rect 7360 15000 7720 15004
rect 5520 14956 7320 14960
rect 5520 14924 5524 14956
rect 5556 14924 5684 14956
rect 5716 14924 5844 14956
rect 5876 14924 6004 14956
rect 6036 14924 6164 14956
rect 6196 14924 6324 14956
rect 6356 14924 6484 14956
rect 6516 14924 6644 14956
rect 6676 14924 6804 14956
rect 6836 14924 6964 14956
rect 6996 14924 7124 14956
rect 7156 14924 7284 14956
rect 7316 14924 7320 14956
rect 5520 14920 7320 14924
rect 7360 14956 7720 14960
rect 7360 14924 7364 14956
rect 7396 14924 7524 14956
rect 7556 14924 7684 14956
rect 7716 14924 7720 14956
rect 7360 14920 7720 14924
rect 5520 14876 7320 14880
rect 5520 14844 5524 14876
rect 5556 14844 5684 14876
rect 5716 14844 5844 14876
rect 5876 14844 6004 14876
rect 6036 14844 6164 14876
rect 6196 14844 6324 14876
rect 6356 14844 6484 14876
rect 6516 14844 6644 14876
rect 6676 14844 6804 14876
rect 6836 14844 6964 14876
rect 6996 14844 7124 14876
rect 7156 14844 7284 14876
rect 7316 14844 7320 14876
rect 5520 14840 7320 14844
rect 7360 14876 7720 14880
rect 7360 14844 7364 14876
rect 7396 14844 7524 14876
rect 7556 14844 7684 14876
rect 7716 14844 7720 14876
rect 7360 14840 7720 14844
rect 5520 14796 7320 14800
rect 5520 14764 5524 14796
rect 5556 14764 5684 14796
rect 5716 14764 5844 14796
rect 5876 14764 6004 14796
rect 6036 14764 6164 14796
rect 6196 14764 6324 14796
rect 6356 14764 6484 14796
rect 6516 14764 6644 14796
rect 6676 14764 6804 14796
rect 6836 14764 6964 14796
rect 6996 14764 7124 14796
rect 7156 14764 7284 14796
rect 7316 14764 7320 14796
rect 5520 14760 7320 14764
rect 7360 14796 7720 14800
rect 7360 14764 7364 14796
rect 7396 14764 7524 14796
rect 7556 14764 7684 14796
rect 7716 14764 7720 14796
rect 7360 14760 7720 14764
rect 5520 14716 7320 14720
rect 5520 14684 5524 14716
rect 5556 14684 5684 14716
rect 5716 14684 5844 14716
rect 5876 14684 6004 14716
rect 6036 14684 6164 14716
rect 6196 14684 6324 14716
rect 6356 14684 6484 14716
rect 6516 14684 6644 14716
rect 6676 14684 6804 14716
rect 6836 14684 6964 14716
rect 6996 14684 7124 14716
rect 7156 14684 7284 14716
rect 7316 14684 7320 14716
rect 5520 14680 7320 14684
rect 7360 14716 7720 14720
rect 7360 14684 7364 14716
rect 7396 14684 7524 14716
rect 7556 14684 7684 14716
rect 7716 14684 7720 14716
rect 7360 14680 7720 14684
rect 6000 14636 7320 14640
rect 6000 14604 6004 14636
rect 6036 14604 6164 14636
rect 6196 14604 6324 14636
rect 6356 14604 6484 14636
rect 6516 14604 6644 14636
rect 6676 14604 6804 14636
rect 6836 14604 6964 14636
rect 6996 14604 7124 14636
rect 7156 14604 7284 14636
rect 7316 14604 7320 14636
rect 6000 14600 7320 14604
rect 7360 14636 7720 14640
rect 7360 14604 7364 14636
rect 7396 14604 7524 14636
rect 7556 14604 7684 14636
rect 7716 14604 7720 14636
rect 7360 14600 7720 14604
rect 5520 14556 7320 14560
rect 5520 14524 5524 14556
rect 5556 14524 5684 14556
rect 5716 14524 5844 14556
rect 5876 14524 6004 14556
rect 6036 14524 6164 14556
rect 6196 14524 6324 14556
rect 6356 14524 6484 14556
rect 6516 14524 6644 14556
rect 6676 14524 6804 14556
rect 6836 14524 6964 14556
rect 6996 14524 7124 14556
rect 7156 14524 7284 14556
rect 7316 14524 7320 14556
rect 5520 14520 7320 14524
rect 7360 14556 7720 14560
rect 7360 14524 7364 14556
rect 7396 14524 7524 14556
rect 7556 14524 7684 14556
rect 7716 14524 7720 14556
rect 7360 14520 7720 14524
rect 5520 14476 7320 14480
rect 5520 14444 5524 14476
rect 5556 14444 5684 14476
rect 5716 14444 5844 14476
rect 5876 14444 6004 14476
rect 6036 14444 6164 14476
rect 6196 14444 6324 14476
rect 6356 14444 6484 14476
rect 6516 14444 6644 14476
rect 6676 14444 6804 14476
rect 6836 14444 6964 14476
rect 6996 14444 7124 14476
rect 7156 14444 7284 14476
rect 7316 14444 7320 14476
rect 5520 14440 7320 14444
rect 7360 14476 7720 14480
rect 7360 14444 7364 14476
rect 7396 14444 7524 14476
rect 7556 14444 7684 14476
rect 7716 14444 7720 14476
rect 7360 14440 7720 14444
rect 7360 14396 7720 14400
rect 7360 14364 7364 14396
rect 7396 14364 7524 14396
rect 7556 14364 7684 14396
rect 7716 14364 7720 14396
rect 7360 14360 7720 14364
rect 7360 14316 7720 14320
rect 7360 14284 7364 14316
rect 7396 14284 7524 14316
rect 7556 14284 7684 14316
rect 7716 14284 7720 14316
rect 7360 14280 7720 14284
rect 7360 14236 7720 14240
rect 7360 14204 7364 14236
rect 7396 14204 7524 14236
rect 7556 14204 7684 14236
rect 7716 14204 7720 14236
rect 7360 14200 7720 14204
rect 7360 14156 7720 14160
rect 7360 14124 7364 14156
rect 7396 14124 7524 14156
rect 7556 14124 7684 14156
rect 7716 14124 7720 14156
rect 7360 14120 7720 14124
rect 7360 14076 7720 14080
rect 7360 14044 7364 14076
rect 7396 14044 7524 14076
rect 7556 14044 7684 14076
rect 7716 14044 7720 14076
rect 7360 14040 7720 14044
rect 5520 13996 7320 14000
rect 5520 13964 5524 13996
rect 5556 13964 5684 13996
rect 5716 13964 5844 13996
rect 5876 13964 6004 13996
rect 6036 13964 6164 13996
rect 6196 13964 6324 13996
rect 6356 13964 6484 13996
rect 6516 13964 6644 13996
rect 6676 13964 6804 13996
rect 6836 13964 6964 13996
rect 6996 13964 7124 13996
rect 7156 13964 7284 13996
rect 7316 13964 7320 13996
rect 5520 13960 7320 13964
rect 7360 13996 7720 14000
rect 7360 13964 7364 13996
rect 7396 13964 7524 13996
rect 7556 13964 7684 13996
rect 7716 13964 7720 13996
rect 7360 13960 7720 13964
rect 5840 13876 7320 13880
rect 5840 13844 5844 13876
rect 5876 13844 6004 13876
rect 6036 13844 6164 13876
rect 6196 13844 6324 13876
rect 6356 13844 6484 13876
rect 6516 13844 6644 13876
rect 6676 13844 6804 13876
rect 6836 13844 6964 13876
rect 6996 13844 7124 13876
rect 7156 13844 7284 13876
rect 7316 13844 7320 13876
rect 5840 13840 7320 13844
rect 7360 13876 7720 13880
rect 7360 13844 7364 13876
rect 7396 13844 7524 13876
rect 7556 13844 7684 13876
rect 7716 13844 7720 13876
rect 7360 13840 7720 13844
rect 5520 13796 7320 13800
rect 5520 13764 5524 13796
rect 5556 13764 5684 13796
rect 5716 13764 5844 13796
rect 5876 13764 6004 13796
rect 6036 13764 6164 13796
rect 6196 13764 6324 13796
rect 6356 13764 6484 13796
rect 6516 13764 6644 13796
rect 6676 13764 6804 13796
rect 6836 13764 6964 13796
rect 6996 13764 7124 13796
rect 7156 13764 7284 13796
rect 7316 13764 7320 13796
rect 5520 13760 7320 13764
rect 7360 13796 7720 13800
rect 7360 13764 7364 13796
rect 7396 13764 7524 13796
rect 7556 13764 7684 13796
rect 7716 13764 7720 13796
rect 7360 13760 7720 13764
rect 5520 13716 7320 13720
rect 5520 13684 5524 13716
rect 5556 13684 5684 13716
rect 5716 13684 5844 13716
rect 5876 13684 6004 13716
rect 6036 13684 6164 13716
rect 6196 13684 6324 13716
rect 6356 13684 6484 13716
rect 6516 13684 6644 13716
rect 6676 13684 6804 13716
rect 6836 13684 6964 13716
rect 6996 13684 7124 13716
rect 7156 13684 7284 13716
rect 7316 13684 7320 13716
rect 5520 13680 7320 13684
rect 7360 13716 7720 13720
rect 7360 13684 7364 13716
rect 7396 13684 7524 13716
rect 7556 13684 7684 13716
rect 7716 13684 7720 13716
rect 7360 13680 7720 13684
rect 5520 13636 7320 13640
rect 5520 13604 5524 13636
rect 5556 13604 5684 13636
rect 5716 13604 5844 13636
rect 5876 13604 6004 13636
rect 6036 13604 6164 13636
rect 6196 13604 6324 13636
rect 6356 13604 6484 13636
rect 6516 13604 6644 13636
rect 6676 13604 6804 13636
rect 6836 13604 6964 13636
rect 6996 13604 7124 13636
rect 7156 13604 7284 13636
rect 7316 13604 7320 13636
rect 5520 13600 7320 13604
rect 7360 13636 7720 13640
rect 7360 13604 7364 13636
rect 7396 13604 7524 13636
rect 7556 13604 7684 13636
rect 7716 13604 7720 13636
rect 7360 13600 7720 13604
rect 6160 13556 7320 13560
rect 6160 13524 6164 13556
rect 6196 13524 6324 13556
rect 6356 13524 6484 13556
rect 6516 13524 6644 13556
rect 6676 13524 6804 13556
rect 6836 13524 6964 13556
rect 6996 13524 7124 13556
rect 7156 13524 7284 13556
rect 7316 13524 7320 13556
rect 6160 13520 7320 13524
rect 7360 13556 7720 13560
rect 7360 13524 7364 13556
rect 7396 13524 7524 13556
rect 7556 13524 7684 13556
rect 7716 13524 7720 13556
rect 7360 13520 7720 13524
rect 5520 13476 7320 13480
rect 5520 13444 5524 13476
rect 5556 13444 5684 13476
rect 5716 13444 5844 13476
rect 5876 13444 6004 13476
rect 6036 13444 6164 13476
rect 6196 13444 6324 13476
rect 6356 13444 6484 13476
rect 6516 13444 6644 13476
rect 6676 13444 6804 13476
rect 6836 13444 6964 13476
rect 6996 13444 7124 13476
rect 7156 13444 7284 13476
rect 7316 13444 7320 13476
rect 5520 13440 7320 13444
rect 7360 13476 7720 13480
rect 7360 13444 7364 13476
rect 7396 13444 7524 13476
rect 7556 13444 7684 13476
rect 7716 13444 7720 13476
rect 7360 13440 7720 13444
rect 5520 13396 7320 13400
rect 5520 13364 5524 13396
rect 5556 13364 5684 13396
rect 5716 13364 5844 13396
rect 5876 13364 6004 13396
rect 6036 13364 6164 13396
rect 6196 13364 6324 13396
rect 6356 13364 6484 13396
rect 6516 13364 6644 13396
rect 6676 13364 6804 13396
rect 6836 13364 6964 13396
rect 6996 13364 7124 13396
rect 7156 13364 7284 13396
rect 7316 13364 7320 13396
rect 5520 13360 7320 13364
rect 7360 13396 7720 13400
rect 7360 13364 7364 13396
rect 7396 13364 7524 13396
rect 7556 13364 7684 13396
rect 7716 13364 7720 13396
rect 7360 13360 7720 13364
rect 5520 13316 7320 13320
rect 5520 13284 5524 13316
rect 5556 13284 5684 13316
rect 5716 13284 5844 13316
rect 5876 13284 6004 13316
rect 6036 13284 6164 13316
rect 6196 13284 6324 13316
rect 6356 13284 6484 13316
rect 6516 13284 6644 13316
rect 6676 13284 6804 13316
rect 6836 13284 6964 13316
rect 6996 13284 7124 13316
rect 7156 13284 7284 13316
rect 7316 13284 7320 13316
rect 5520 13280 7320 13284
rect 7360 13316 7720 13320
rect 7360 13284 7364 13316
rect 7396 13284 7524 13316
rect 7556 13284 7684 13316
rect 7716 13284 7720 13316
rect 7360 13280 7720 13284
rect 5520 13236 7320 13240
rect 5520 13204 5524 13236
rect 5556 13204 5684 13236
rect 5716 13204 5844 13236
rect 5876 13204 6004 13236
rect 6036 13204 6164 13236
rect 6196 13204 6324 13236
rect 6356 13204 6484 13236
rect 6516 13204 6644 13236
rect 6676 13204 6804 13236
rect 6836 13204 6964 13236
rect 6996 13204 7124 13236
rect 7156 13204 7284 13236
rect 7316 13204 7320 13236
rect 5520 13200 7320 13204
rect 7360 13236 7720 13240
rect 7360 13204 7364 13236
rect 7396 13204 7524 13236
rect 7556 13204 7684 13236
rect 7716 13204 7720 13236
rect 7360 13200 7720 13204
rect 6000 13156 7320 13160
rect 6000 13124 6004 13156
rect 6036 13124 6164 13156
rect 6196 13124 6324 13156
rect 6356 13124 6484 13156
rect 6516 13124 6644 13156
rect 6676 13124 6804 13156
rect 6836 13124 6964 13156
rect 6996 13124 7124 13156
rect 7156 13124 7284 13156
rect 7316 13124 7320 13156
rect 6000 13120 7320 13124
rect 7360 13156 7720 13160
rect 7360 13124 7364 13156
rect 7396 13124 7524 13156
rect 7556 13124 7684 13156
rect 7716 13124 7720 13156
rect 7360 13120 7720 13124
rect 5520 13076 7320 13080
rect 5520 13044 5524 13076
rect 5556 13044 5684 13076
rect 5716 13044 5844 13076
rect 5876 13044 6004 13076
rect 6036 13044 6164 13076
rect 6196 13044 6324 13076
rect 6356 13044 6484 13076
rect 6516 13044 6644 13076
rect 6676 13044 6804 13076
rect 6836 13044 6964 13076
rect 6996 13044 7124 13076
rect 7156 13044 7284 13076
rect 7316 13044 7320 13076
rect 5520 13040 7320 13044
rect 7360 13076 7720 13080
rect 7360 13044 7364 13076
rect 7396 13044 7524 13076
rect 7556 13044 7684 13076
rect 7716 13044 7720 13076
rect 7360 13040 7720 13044
rect 5520 12996 7320 13000
rect 5520 12964 5524 12996
rect 5556 12964 5684 12996
rect 5716 12964 5844 12996
rect 5876 12964 6004 12996
rect 6036 12964 6164 12996
rect 6196 12964 6324 12996
rect 6356 12964 6484 12996
rect 6516 12964 6644 12996
rect 6676 12964 6804 12996
rect 6836 12964 6964 12996
rect 6996 12964 7124 12996
rect 7156 12964 7284 12996
rect 7316 12964 7320 12996
rect 5520 12960 7320 12964
rect 7360 12996 7720 13000
rect 7360 12964 7364 12996
rect 7396 12964 7524 12996
rect 7556 12964 7684 12996
rect 7716 12964 7720 12996
rect 7360 12960 7720 12964
rect 5520 12516 7320 12520
rect 5520 12484 5524 12516
rect 5556 12484 5684 12516
rect 5716 12484 5844 12516
rect 5876 12484 6004 12516
rect 6036 12484 6164 12516
rect 6196 12484 6324 12516
rect 6356 12484 6484 12516
rect 6516 12484 6644 12516
rect 6676 12484 6804 12516
rect 6836 12484 6964 12516
rect 6996 12484 7124 12516
rect 7156 12484 7284 12516
rect 7316 12484 7320 12516
rect 5520 12480 7320 12484
rect 7360 12476 7720 12480
rect 7360 12444 7364 12476
rect 7396 12444 7524 12476
rect 7556 12444 7684 12476
rect 7716 12444 7720 12476
rect 7360 12440 7720 12444
rect 5840 12436 7320 12440
rect 5840 12404 5844 12436
rect 5876 12404 6004 12436
rect 6036 12404 6164 12436
rect 6196 12404 6324 12436
rect 6356 12404 6484 12436
rect 6516 12404 6644 12436
rect 6676 12404 6804 12436
rect 6836 12404 6964 12436
rect 6996 12404 7124 12436
rect 7156 12404 7284 12436
rect 7316 12404 7320 12436
rect 5840 12400 7320 12404
rect 7360 12396 7720 12400
rect 7360 12364 7364 12396
rect 7396 12364 7524 12396
rect 7556 12364 7684 12396
rect 7716 12364 7720 12396
rect 7360 12360 7720 12364
rect 5520 12316 7320 12320
rect 5520 12284 5524 12316
rect 5556 12284 5684 12316
rect 5716 12284 5844 12316
rect 5876 12284 6004 12316
rect 6036 12284 6164 12316
rect 6196 12284 6324 12316
rect 6356 12284 6484 12316
rect 6516 12284 6644 12316
rect 6676 12284 6804 12316
rect 6836 12284 6964 12316
rect 6996 12284 7124 12316
rect 7156 12284 7284 12316
rect 7316 12284 7320 12316
rect 5520 12280 7320 12284
rect 7360 12316 7720 12320
rect 7360 12284 7364 12316
rect 7396 12284 7524 12316
rect 7556 12284 7684 12316
rect 7716 12284 7720 12316
rect 7360 12280 7720 12284
rect 5520 12236 7320 12240
rect 5520 12204 5524 12236
rect 5556 12204 5684 12236
rect 5716 12204 5844 12236
rect 5876 12204 6004 12236
rect 6036 12204 6164 12236
rect 6196 12204 6324 12236
rect 6356 12204 6484 12236
rect 6516 12204 6644 12236
rect 6676 12204 6804 12236
rect 6836 12204 6964 12236
rect 6996 12204 7124 12236
rect 7156 12204 7284 12236
rect 7316 12204 7320 12236
rect 5520 12200 7320 12204
rect 7360 12236 7720 12240
rect 7360 12204 7364 12236
rect 7396 12204 7524 12236
rect 7556 12204 7684 12236
rect 7716 12204 7720 12236
rect 7360 12200 7720 12204
rect 5520 12156 7320 12160
rect 5520 12124 5524 12156
rect 5556 12124 5684 12156
rect 5716 12124 5844 12156
rect 5876 12124 6004 12156
rect 6036 12124 6164 12156
rect 6196 12124 6324 12156
rect 6356 12124 6484 12156
rect 6516 12124 6644 12156
rect 6676 12124 6804 12156
rect 6836 12124 6964 12156
rect 6996 12124 7124 12156
rect 7156 12124 7284 12156
rect 7316 12124 7320 12156
rect 5520 12120 7320 12124
rect 7360 12156 7720 12160
rect 7360 12124 7364 12156
rect 7396 12124 7524 12156
rect 7556 12124 7684 12156
rect 7716 12124 7720 12156
rect 7360 12120 7720 12124
rect 5520 12076 7320 12080
rect 5520 12044 5524 12076
rect 5556 12044 5684 12076
rect 5716 12044 5844 12076
rect 5876 12044 6004 12076
rect 6036 12044 6164 12076
rect 6196 12044 6324 12076
rect 6356 12044 6484 12076
rect 6516 12044 6644 12076
rect 6676 12044 6804 12076
rect 6836 12044 6964 12076
rect 6996 12044 7124 12076
rect 7156 12044 7284 12076
rect 7316 12044 7320 12076
rect 5520 12040 7320 12044
rect 7360 12076 7720 12080
rect 7360 12044 7364 12076
rect 7396 12044 7524 12076
rect 7556 12044 7684 12076
rect 7716 12044 7720 12076
rect 7360 12040 7720 12044
rect 5520 11996 7320 12000
rect 5520 11964 5524 11996
rect 5556 11964 5684 11996
rect 5716 11964 5844 11996
rect 5876 11964 6004 11996
rect 6036 11964 6164 11996
rect 6196 11964 6324 11996
rect 6356 11964 6484 11996
rect 6516 11964 6644 11996
rect 6676 11964 6804 11996
rect 6836 11964 6964 11996
rect 6996 11964 7124 11996
rect 7156 11964 7284 11996
rect 7316 11964 7320 11996
rect 5520 11960 7320 11964
rect 7360 11996 7720 12000
rect 7360 11964 7364 11996
rect 7396 11964 7524 11996
rect 7556 11964 7684 11996
rect 7716 11964 7720 11996
rect 7360 11960 7720 11964
rect 5520 11916 7320 11920
rect 5520 11884 5524 11916
rect 5556 11884 5684 11916
rect 5716 11884 5844 11916
rect 5876 11884 6004 11916
rect 6036 11884 6164 11916
rect 6196 11884 6324 11916
rect 6356 11884 6484 11916
rect 6516 11884 6644 11916
rect 6676 11884 6804 11916
rect 6836 11884 6964 11916
rect 6996 11884 7124 11916
rect 7156 11884 7284 11916
rect 7316 11884 7320 11916
rect 5520 11880 7320 11884
rect 7360 11916 7720 11920
rect 7360 11884 7364 11916
rect 7396 11884 7524 11916
rect 7556 11884 7684 11916
rect 7716 11884 7720 11916
rect 7360 11880 7720 11884
rect 5520 11836 7320 11840
rect 5520 11804 5524 11836
rect 5556 11804 5684 11836
rect 5716 11804 5844 11836
rect 5876 11804 6004 11836
rect 6036 11804 6164 11836
rect 6196 11804 6324 11836
rect 6356 11804 6484 11836
rect 6516 11804 6644 11836
rect 6676 11804 6804 11836
rect 6836 11804 6964 11836
rect 6996 11804 7124 11836
rect 7156 11804 7284 11836
rect 7316 11804 7320 11836
rect 5520 11800 7320 11804
rect 7360 11836 7720 11840
rect 7360 11804 7364 11836
rect 7396 11804 7524 11836
rect 7556 11804 7684 11836
rect 7716 11804 7720 11836
rect 7360 11800 7720 11804
rect 5520 11756 7320 11760
rect 5520 11724 5524 11756
rect 5556 11724 5684 11756
rect 5716 11724 5844 11756
rect 5876 11724 6004 11756
rect 6036 11724 6164 11756
rect 6196 11724 6324 11756
rect 6356 11724 6484 11756
rect 6516 11724 6644 11756
rect 6676 11724 6804 11756
rect 6836 11724 6964 11756
rect 6996 11724 7124 11756
rect 7156 11724 7284 11756
rect 7316 11724 7320 11756
rect 5520 11720 7320 11724
rect 7360 11756 7720 11760
rect 7360 11724 7364 11756
rect 7396 11724 7524 11756
rect 7556 11724 7684 11756
rect 7716 11724 7720 11756
rect 7360 11720 7720 11724
rect 5520 11676 7320 11680
rect 5520 11644 5524 11676
rect 5556 11644 5684 11676
rect 5716 11644 5844 11676
rect 5876 11644 6004 11676
rect 6036 11644 6164 11676
rect 6196 11644 6324 11676
rect 6356 11644 6484 11676
rect 6516 11644 6644 11676
rect 6676 11644 6804 11676
rect 6836 11644 6964 11676
rect 6996 11644 7124 11676
rect 7156 11644 7284 11676
rect 7316 11644 7320 11676
rect 5520 11640 7320 11644
rect 7360 11676 7720 11680
rect 7360 11644 7364 11676
rect 7396 11644 7524 11676
rect 7556 11644 7684 11676
rect 7716 11644 7720 11676
rect 7360 11640 7720 11644
rect 5520 11596 7320 11600
rect 5520 11564 5524 11596
rect 5556 11564 5684 11596
rect 5716 11564 5844 11596
rect 5876 11564 6004 11596
rect 6036 11564 6164 11596
rect 6196 11564 6324 11596
rect 6356 11564 6484 11596
rect 6516 11564 6644 11596
rect 6676 11564 6804 11596
rect 6836 11564 6964 11596
rect 6996 11564 7124 11596
rect 7156 11564 7284 11596
rect 7316 11564 7320 11596
rect 5520 11560 7320 11564
rect 7360 11596 7720 11600
rect 7360 11564 7364 11596
rect 7396 11564 7524 11596
rect 7556 11564 7684 11596
rect 7716 11564 7720 11596
rect 7360 11560 7720 11564
rect 5520 11516 7320 11520
rect 5520 11484 5524 11516
rect 5556 11484 5684 11516
rect 5716 11484 5844 11516
rect 5876 11484 6004 11516
rect 6036 11484 6164 11516
rect 6196 11484 6324 11516
rect 6356 11484 6484 11516
rect 6516 11484 6644 11516
rect 6676 11484 6804 11516
rect 6836 11484 6964 11516
rect 6996 11484 7124 11516
rect 7156 11484 7284 11516
rect 7316 11484 7320 11516
rect 5520 11480 7320 11484
rect 7360 11516 7720 11520
rect 7360 11484 7364 11516
rect 7396 11484 7524 11516
rect 7556 11484 7684 11516
rect 7716 11484 7720 11516
rect 7360 11480 7720 11484
rect 5520 11436 7320 11440
rect 5520 11404 5524 11436
rect 5556 11404 5684 11436
rect 5716 11404 5844 11436
rect 5876 11404 6004 11436
rect 6036 11404 6164 11436
rect 6196 11404 6324 11436
rect 6356 11404 6484 11436
rect 6516 11404 6644 11436
rect 6676 11404 6804 11436
rect 6836 11404 6964 11436
rect 6996 11404 7124 11436
rect 7156 11404 7284 11436
rect 7316 11404 7320 11436
rect 5520 11400 7320 11404
rect 7360 11436 7720 11440
rect 7360 11404 7364 11436
rect 7396 11404 7524 11436
rect 7556 11404 7684 11436
rect 7716 11404 7720 11436
rect 7360 11400 7720 11404
rect 5520 11356 7320 11360
rect 5520 11324 5524 11356
rect 5556 11324 5684 11356
rect 5716 11324 5844 11356
rect 5876 11324 6004 11356
rect 6036 11324 6164 11356
rect 6196 11324 6324 11356
rect 6356 11324 6484 11356
rect 6516 11324 6644 11356
rect 6676 11324 6804 11356
rect 6836 11324 6964 11356
rect 6996 11324 7124 11356
rect 7156 11324 7284 11356
rect 7316 11324 7320 11356
rect 5520 11320 7320 11324
rect 7360 11356 7720 11360
rect 7360 11324 7364 11356
rect 7396 11324 7524 11356
rect 7556 11324 7684 11356
rect 7716 11324 7720 11356
rect 7360 11320 7720 11324
rect 7360 11276 7720 11280
rect 7360 11244 7364 11276
rect 7396 11244 7524 11276
rect 7556 11244 7684 11276
rect 7716 11244 7720 11276
rect 7360 11240 7720 11244
rect 5520 11196 7320 11200
rect 5520 11164 5524 11196
rect 5556 11164 5684 11196
rect 5716 11164 5844 11196
rect 5876 11164 6004 11196
rect 6036 11164 6164 11196
rect 6196 11164 6324 11196
rect 6356 11164 6484 11196
rect 6516 11164 6644 11196
rect 6676 11164 6804 11196
rect 6836 11164 6964 11196
rect 6996 11164 7124 11196
rect 7156 11164 7284 11196
rect 7316 11164 7320 11196
rect 5520 11160 7320 11164
rect 7360 11196 7720 11200
rect 7360 11164 7364 11196
rect 7396 11164 7524 11196
rect 7556 11164 7684 11196
rect 7716 11164 7720 11196
rect 7360 11160 7720 11164
rect 5520 11116 7320 11120
rect 5520 11084 5524 11116
rect 5556 11084 5684 11116
rect 5716 11084 5844 11116
rect 5876 11084 6004 11116
rect 6036 11084 6164 11116
rect 6196 11084 6324 11116
rect 6356 11084 6484 11116
rect 6516 11084 6644 11116
rect 6676 11084 6804 11116
rect 6836 11084 6964 11116
rect 6996 11084 7124 11116
rect 7156 11084 7284 11116
rect 7316 11084 7320 11116
rect 5520 11080 7320 11084
rect 7360 11116 7720 11120
rect 7360 11084 7364 11116
rect 7396 11084 7524 11116
rect 7556 11084 7684 11116
rect 7716 11084 7720 11116
rect 7360 11080 7720 11084
rect 5520 11036 7320 11040
rect 5520 11004 5524 11036
rect 5556 11004 5684 11036
rect 5716 11004 5844 11036
rect 5876 11004 6004 11036
rect 6036 11004 6164 11036
rect 6196 11004 6324 11036
rect 6356 11004 6484 11036
rect 6516 11004 6644 11036
rect 6676 11004 6804 11036
rect 6836 11004 6964 11036
rect 6996 11004 7124 11036
rect 7156 11004 7284 11036
rect 7316 11004 7320 11036
rect 5520 11000 7320 11004
rect 7360 11036 7720 11040
rect 7360 11004 7364 11036
rect 7396 11004 7524 11036
rect 7556 11004 7684 11036
rect 7716 11004 7720 11036
rect 7360 11000 7720 11004
rect 7360 10956 7720 10960
rect 7360 10924 7364 10956
rect 7396 10924 7524 10956
rect 7556 10924 7684 10956
rect 7716 10924 7720 10956
rect 7360 10920 7720 10924
rect 5520 10876 7320 10880
rect 5520 10844 5524 10876
rect 5556 10844 5684 10876
rect 5716 10844 5844 10876
rect 5876 10844 6004 10876
rect 6036 10844 6164 10876
rect 6196 10844 6324 10876
rect 6356 10844 6484 10876
rect 6516 10844 6644 10876
rect 6676 10844 6804 10876
rect 6836 10844 6964 10876
rect 6996 10844 7124 10876
rect 7156 10844 7284 10876
rect 7316 10844 7320 10876
rect 5520 10840 7320 10844
rect 7360 10876 7720 10880
rect 7360 10844 7364 10876
rect 7396 10844 7524 10876
rect 7556 10844 7684 10876
rect 7716 10844 7720 10876
rect 7360 10840 7720 10844
rect 7120 10796 7320 10800
rect 7120 10764 7124 10796
rect 7156 10764 7284 10796
rect 7316 10764 7320 10796
rect 7120 10760 7320 10764
rect 7360 10796 7720 10800
rect 7360 10764 7364 10796
rect 7396 10764 7524 10796
rect 7556 10764 7684 10796
rect 7716 10764 7720 10796
rect 7360 10760 7720 10764
rect 5520 10716 7320 10720
rect 5520 10684 5524 10716
rect 5556 10684 5684 10716
rect 5716 10684 5844 10716
rect 5876 10684 6004 10716
rect 6036 10684 6164 10716
rect 6196 10684 6324 10716
rect 6356 10684 6484 10716
rect 6516 10684 6644 10716
rect 6676 10684 6804 10716
rect 6836 10684 6964 10716
rect 6996 10684 7124 10716
rect 7156 10684 7284 10716
rect 7316 10684 7320 10716
rect 5520 10680 7320 10684
rect 7360 10716 7720 10720
rect 7360 10684 7364 10716
rect 7396 10684 7524 10716
rect 7556 10684 7684 10716
rect 7716 10684 7720 10716
rect 7360 10680 7720 10684
rect 5520 10636 7320 10640
rect 5520 10604 5524 10636
rect 5556 10604 5684 10636
rect 5716 10604 5844 10636
rect 5876 10604 6004 10636
rect 6036 10604 6164 10636
rect 6196 10604 6324 10636
rect 6356 10604 6484 10636
rect 6516 10604 6644 10636
rect 6676 10604 6804 10636
rect 6836 10604 6964 10636
rect 6996 10604 7124 10636
rect 7156 10604 7284 10636
rect 7316 10604 7320 10636
rect 5520 10600 7320 10604
rect 7360 10636 7720 10640
rect 7360 10604 7364 10636
rect 7396 10604 7524 10636
rect 7556 10604 7684 10636
rect 7716 10604 7720 10636
rect 7360 10600 7720 10604
rect 7120 10556 7320 10560
rect 7120 10524 7124 10556
rect 7156 10524 7284 10556
rect 7316 10524 7320 10556
rect 7120 10520 7320 10524
rect 7360 10556 7720 10560
rect 7360 10524 7364 10556
rect 7396 10524 7524 10556
rect 7556 10524 7684 10556
rect 7716 10524 7720 10556
rect 7360 10520 7720 10524
rect 5520 10476 7320 10480
rect 5520 10444 5524 10476
rect 5556 10444 5684 10476
rect 5716 10444 5844 10476
rect 5876 10444 6004 10476
rect 6036 10444 6164 10476
rect 6196 10444 6324 10476
rect 6356 10444 6484 10476
rect 6516 10444 6644 10476
rect 6676 10444 6804 10476
rect 6836 10444 6964 10476
rect 6996 10444 7124 10476
rect 7156 10444 7284 10476
rect 7316 10444 7320 10476
rect 5520 10440 7320 10444
rect 7360 10476 7720 10480
rect 7360 10444 7364 10476
rect 7396 10444 7524 10476
rect 7556 10444 7684 10476
rect 7716 10444 7720 10476
rect 7360 10440 7720 10444
rect 6960 10396 7320 10400
rect 6960 10364 6964 10396
rect 6996 10364 7124 10396
rect 7156 10364 7284 10396
rect 7316 10364 7320 10396
rect 6960 10360 7320 10364
rect 7360 10396 7720 10400
rect 7360 10364 7364 10396
rect 7396 10364 7524 10396
rect 7556 10364 7684 10396
rect 7716 10364 7720 10396
rect 7360 10360 7720 10364
rect 5520 10316 7320 10320
rect 5520 10284 5524 10316
rect 5556 10284 5684 10316
rect 5716 10284 5844 10316
rect 5876 10284 6004 10316
rect 6036 10284 6164 10316
rect 6196 10284 6324 10316
rect 6356 10284 6484 10316
rect 6516 10284 6644 10316
rect 6676 10284 6804 10316
rect 6836 10284 6964 10316
rect 6996 10284 7124 10316
rect 7156 10284 7284 10316
rect 7316 10284 7320 10316
rect 5520 10280 7320 10284
rect 7360 10316 7720 10320
rect 7360 10284 7364 10316
rect 7396 10284 7524 10316
rect 7556 10284 7684 10316
rect 7716 10284 7720 10316
rect 7360 10280 7720 10284
rect 5520 10236 7320 10240
rect 5520 10204 5524 10236
rect 5556 10204 5684 10236
rect 5716 10204 5844 10236
rect 5876 10204 6004 10236
rect 6036 10204 6164 10236
rect 6196 10204 6324 10236
rect 6356 10204 6484 10236
rect 6516 10204 6644 10236
rect 6676 10204 6804 10236
rect 6836 10204 6964 10236
rect 6996 10204 7124 10236
rect 7156 10204 7284 10236
rect 7316 10204 7320 10236
rect 5520 10200 7320 10204
rect 7360 10236 7720 10240
rect 7360 10204 7364 10236
rect 7396 10204 7524 10236
rect 7556 10204 7684 10236
rect 7716 10204 7720 10236
rect 7360 10200 7720 10204
rect 5520 10156 7320 10160
rect 5520 10124 5524 10156
rect 5556 10124 5684 10156
rect 5716 10124 5844 10156
rect 5876 10124 6004 10156
rect 6036 10124 6164 10156
rect 6196 10124 6324 10156
rect 6356 10124 6484 10156
rect 6516 10124 6644 10156
rect 6676 10124 6804 10156
rect 6836 10124 6964 10156
rect 6996 10124 7124 10156
rect 7156 10124 7284 10156
rect 7316 10124 7320 10156
rect 5520 10120 7320 10124
rect 7360 10156 7720 10160
rect 7360 10124 7364 10156
rect 7396 10124 7524 10156
rect 7556 10124 7684 10156
rect 7716 10124 7720 10156
rect 7360 10120 7720 10124
rect 5520 10076 7320 10080
rect 5520 10044 5524 10076
rect 5556 10044 5684 10076
rect 5716 10044 5844 10076
rect 5876 10044 6004 10076
rect 6036 10044 6164 10076
rect 6196 10044 6324 10076
rect 6356 10044 6484 10076
rect 6516 10044 6644 10076
rect 6676 10044 6804 10076
rect 6836 10044 6964 10076
rect 6996 10044 7124 10076
rect 7156 10044 7284 10076
rect 7316 10044 7320 10076
rect 5520 10040 7320 10044
rect 7360 10076 7720 10080
rect 7360 10044 7364 10076
rect 7396 10044 7524 10076
rect 7556 10044 7684 10076
rect 7716 10044 7720 10076
rect 7360 10040 7720 10044
rect 5520 9996 7320 10000
rect 5520 9964 5524 9996
rect 5556 9964 5684 9996
rect 5716 9964 5844 9996
rect 5876 9964 6004 9996
rect 6036 9964 6164 9996
rect 6196 9964 6324 9996
rect 6356 9964 6484 9996
rect 6516 9964 6644 9996
rect 6676 9964 6804 9996
rect 6836 9964 6964 9996
rect 6996 9964 7124 9996
rect 7156 9964 7284 9996
rect 7316 9964 7320 9996
rect 5520 9960 7320 9964
rect 7360 9996 7720 10000
rect 7360 9964 7364 9996
rect 7396 9964 7524 9996
rect 7556 9964 7684 9996
rect 7716 9964 7720 9996
rect 7360 9960 7720 9964
rect 5520 9916 7320 9920
rect 5520 9884 5524 9916
rect 5556 9884 5684 9916
rect 5716 9884 5844 9916
rect 5876 9884 6004 9916
rect 6036 9884 6164 9916
rect 6196 9884 6324 9916
rect 6356 9884 6484 9916
rect 6516 9884 6644 9916
rect 6676 9884 6804 9916
rect 6836 9884 6964 9916
rect 6996 9884 7124 9916
rect 7156 9884 7284 9916
rect 7316 9884 7320 9916
rect 5520 9880 7320 9884
rect 7360 9916 7720 9920
rect 7360 9884 7364 9916
rect 7396 9884 7524 9916
rect 7556 9884 7684 9916
rect 7716 9884 7720 9916
rect 7360 9880 7720 9884
rect 5520 9836 7320 9840
rect 5520 9804 5524 9836
rect 5556 9804 5684 9836
rect 5716 9804 5844 9836
rect 5876 9804 6004 9836
rect 6036 9804 6164 9836
rect 6196 9804 6324 9836
rect 6356 9804 6484 9836
rect 6516 9804 6644 9836
rect 6676 9804 6804 9836
rect 6836 9804 6964 9836
rect 6996 9804 7124 9836
rect 7156 9804 7284 9836
rect 7316 9804 7320 9836
rect 5520 9800 7320 9804
rect 7360 9836 7720 9840
rect 7360 9804 7364 9836
rect 7396 9804 7524 9836
rect 7556 9804 7684 9836
rect 7716 9804 7720 9836
rect 7360 9800 7720 9804
rect 5520 9756 7320 9760
rect 5520 9724 5524 9756
rect 5556 9724 5684 9756
rect 5716 9724 5844 9756
rect 5876 9724 6004 9756
rect 6036 9724 6164 9756
rect 6196 9724 6324 9756
rect 6356 9724 6484 9756
rect 6516 9724 6644 9756
rect 6676 9724 6804 9756
rect 6836 9724 6964 9756
rect 6996 9724 7124 9756
rect 7156 9724 7284 9756
rect 7316 9724 7320 9756
rect 5520 9720 7320 9724
rect 7360 9756 7720 9760
rect 7360 9724 7364 9756
rect 7396 9724 7524 9756
rect 7556 9724 7684 9756
rect 7716 9724 7720 9756
rect 7360 9720 7720 9724
rect 5520 9676 7320 9680
rect 5520 9644 5524 9676
rect 5556 9644 5684 9676
rect 5716 9644 5844 9676
rect 5876 9644 6004 9676
rect 6036 9644 6164 9676
rect 6196 9644 6324 9676
rect 6356 9644 6484 9676
rect 6516 9644 6644 9676
rect 6676 9644 6804 9676
rect 6836 9644 6964 9676
rect 6996 9644 7124 9676
rect 7156 9644 7284 9676
rect 7316 9644 7320 9676
rect 5520 9640 7320 9644
rect 7360 9676 7720 9680
rect 7360 9644 7364 9676
rect 7396 9644 7524 9676
rect 7556 9644 7684 9676
rect 7716 9644 7720 9676
rect 7360 9640 7720 9644
rect 5520 9596 7320 9600
rect 5520 9564 5524 9596
rect 5556 9564 5684 9596
rect 5716 9564 5844 9596
rect 5876 9564 6004 9596
rect 6036 9564 6164 9596
rect 6196 9564 6324 9596
rect 6356 9564 6484 9596
rect 6516 9564 6644 9596
rect 6676 9564 6804 9596
rect 6836 9564 6964 9596
rect 6996 9564 7124 9596
rect 7156 9564 7284 9596
rect 7316 9564 7320 9596
rect 5520 9560 7320 9564
rect 7360 9596 7720 9600
rect 7360 9564 7364 9596
rect 7396 9564 7524 9596
rect 7556 9564 7684 9596
rect 7716 9564 7720 9596
rect 7360 9560 7720 9564
rect 5520 9516 7320 9520
rect 5520 9484 5524 9516
rect 5556 9484 5684 9516
rect 5716 9484 5844 9516
rect 5876 9484 6004 9516
rect 6036 9484 6164 9516
rect 6196 9484 6324 9516
rect 6356 9484 6484 9516
rect 6516 9484 6644 9516
rect 6676 9484 6804 9516
rect 6836 9484 6964 9516
rect 6996 9484 7124 9516
rect 7156 9484 7284 9516
rect 7316 9484 7320 9516
rect 5520 9480 7320 9484
rect 7360 9516 7720 9520
rect 7360 9484 7364 9516
rect 7396 9484 7524 9516
rect 7556 9484 7684 9516
rect 7716 9484 7720 9516
rect 7360 9480 7720 9484
rect 5520 9436 7320 9440
rect 5520 9404 5524 9436
rect 5556 9404 5684 9436
rect 5716 9404 5844 9436
rect 5876 9404 6004 9436
rect 6036 9404 6164 9436
rect 6196 9404 6324 9436
rect 6356 9404 6484 9436
rect 6516 9404 6644 9436
rect 6676 9404 6804 9436
rect 6836 9404 6964 9436
rect 6996 9404 7124 9436
rect 7156 9404 7284 9436
rect 7316 9404 7320 9436
rect 5520 9400 7320 9404
rect 7360 9436 7720 9440
rect 7360 9404 7364 9436
rect 7396 9404 7524 9436
rect 7556 9404 7684 9436
rect 7716 9404 7720 9436
rect 7360 9400 7720 9404
rect 5520 9356 7320 9360
rect 5520 9324 5524 9356
rect 5556 9324 5684 9356
rect 5716 9324 5844 9356
rect 5876 9324 6004 9356
rect 6036 9324 6164 9356
rect 6196 9324 6324 9356
rect 6356 9324 6484 9356
rect 6516 9324 6644 9356
rect 6676 9324 6804 9356
rect 6836 9324 6964 9356
rect 6996 9324 7124 9356
rect 7156 9324 7284 9356
rect 7316 9324 7320 9356
rect 5520 9320 7320 9324
rect 7360 9356 7720 9360
rect 7360 9324 7364 9356
rect 7396 9324 7524 9356
rect 7556 9324 7684 9356
rect 7716 9324 7720 9356
rect 7360 9320 7720 9324
rect 5520 9276 7320 9280
rect 5520 9244 5524 9276
rect 5556 9244 5684 9276
rect 5716 9244 5844 9276
rect 5876 9244 6004 9276
rect 6036 9244 6164 9276
rect 6196 9244 6324 9276
rect 6356 9244 6484 9276
rect 6516 9244 6644 9276
rect 6676 9244 6804 9276
rect 6836 9244 6964 9276
rect 6996 9244 7124 9276
rect 7156 9244 7284 9276
rect 7316 9244 7320 9276
rect 5520 9240 7320 9244
rect 7360 9276 7720 9280
rect 7360 9244 7364 9276
rect 7396 9244 7524 9276
rect 7556 9244 7684 9276
rect 7716 9244 7720 9276
rect 7360 9240 7720 9244
rect 7360 9196 7720 9200
rect 7360 9164 7364 9196
rect 7396 9164 7524 9196
rect 7556 9164 7684 9196
rect 7716 9164 7720 9196
rect 7360 9160 7720 9164
rect 5520 9116 7320 9120
rect 5520 9084 5524 9116
rect 5556 9084 5684 9116
rect 5716 9084 5844 9116
rect 5876 9084 6004 9116
rect 6036 9084 6164 9116
rect 6196 9084 6324 9116
rect 6356 9084 6484 9116
rect 6516 9084 6644 9116
rect 6676 9084 6804 9116
rect 6836 9084 6964 9116
rect 6996 9084 7124 9116
rect 7156 9084 7284 9116
rect 7316 9084 7320 9116
rect 5520 9080 7320 9084
rect 7360 9116 7720 9120
rect 7360 9084 7364 9116
rect 7396 9084 7524 9116
rect 7556 9084 7684 9116
rect 7716 9084 7720 9116
rect 7360 9080 7720 9084
rect 5520 9036 7320 9040
rect 5520 9004 5524 9036
rect 5556 9004 5684 9036
rect 5716 9004 5844 9036
rect 5876 9004 6004 9036
rect 6036 9004 6164 9036
rect 6196 9004 6324 9036
rect 6356 9004 6484 9036
rect 6516 9004 6644 9036
rect 6676 9004 6804 9036
rect 6836 9004 6964 9036
rect 6996 9004 7124 9036
rect 7156 9004 7284 9036
rect 7316 9004 7320 9036
rect 5520 9000 7320 9004
rect 7360 9036 7720 9040
rect 7360 9004 7364 9036
rect 7396 9004 7524 9036
rect 7556 9004 7684 9036
rect 7716 9004 7720 9036
rect 7360 9000 7720 9004
rect 5520 8956 7320 8960
rect 5520 8924 5524 8956
rect 5556 8924 5684 8956
rect 5716 8924 5844 8956
rect 5876 8924 6004 8956
rect 6036 8924 6164 8956
rect 6196 8924 6324 8956
rect 6356 8924 6484 8956
rect 6516 8924 6644 8956
rect 6676 8924 6804 8956
rect 6836 8924 6964 8956
rect 6996 8924 7124 8956
rect 7156 8924 7284 8956
rect 7316 8924 7320 8956
rect 5520 8920 7320 8924
rect 7360 8956 7720 8960
rect 7360 8924 7364 8956
rect 7396 8924 7524 8956
rect 7556 8924 7684 8956
rect 7716 8924 7720 8956
rect 7360 8920 7720 8924
rect 5520 8636 7320 8640
rect 5520 8604 5524 8636
rect 5556 8604 5684 8636
rect 5716 8604 5844 8636
rect 5876 8604 6004 8636
rect 6036 8604 6164 8636
rect 6196 8604 6324 8636
rect 6356 8604 6484 8636
rect 6516 8604 6644 8636
rect 6676 8604 6804 8636
rect 6836 8604 6964 8636
rect 6996 8604 7124 8636
rect 7156 8604 7284 8636
rect 7316 8604 7320 8636
rect 5520 8600 7320 8604
rect 7360 8636 7720 8640
rect 7360 8604 7364 8636
rect 7396 8604 7524 8636
rect 7556 8604 7684 8636
rect 7716 8604 7720 8636
rect 7360 8600 7720 8604
rect 5520 8556 7320 8560
rect 5520 8524 5524 8556
rect 5556 8524 5684 8556
rect 5716 8524 5844 8556
rect 5876 8524 6004 8556
rect 6036 8524 6164 8556
rect 6196 8524 6324 8556
rect 6356 8524 6484 8556
rect 6516 8524 6644 8556
rect 6676 8524 6804 8556
rect 6836 8524 6964 8556
rect 6996 8524 7124 8556
rect 7156 8524 7284 8556
rect 7316 8524 7320 8556
rect 5520 8520 7320 8524
rect 7360 8556 7720 8560
rect 7360 8524 7364 8556
rect 7396 8524 7524 8556
rect 7556 8524 7684 8556
rect 7716 8524 7720 8556
rect 7360 8520 7720 8524
rect 7120 8476 7320 8480
rect 7120 8444 7124 8476
rect 7156 8444 7284 8476
rect 7316 8444 7320 8476
rect 7120 8440 7320 8444
rect 7360 8476 7720 8480
rect 7360 8444 7364 8476
rect 7396 8444 7524 8476
rect 7556 8444 7684 8476
rect 7716 8444 7720 8476
rect 7360 8440 7720 8444
rect 5520 8396 7320 8400
rect 5520 8364 5524 8396
rect 5556 8364 5684 8396
rect 5716 8364 5844 8396
rect 5876 8364 6004 8396
rect 6036 8364 6164 8396
rect 6196 8364 6324 8396
rect 6356 8364 6484 8396
rect 6516 8364 6644 8396
rect 6676 8364 6804 8396
rect 6836 8364 6964 8396
rect 6996 8364 7124 8396
rect 7156 8364 7284 8396
rect 7316 8364 7320 8396
rect 5520 8360 7320 8364
rect 7360 8396 7720 8400
rect 7360 8364 7364 8396
rect 7396 8364 7524 8396
rect 7556 8364 7684 8396
rect 7716 8364 7720 8396
rect 7360 8360 7720 8364
rect 6800 8316 7320 8320
rect 6800 8284 6804 8316
rect 6836 8284 6964 8316
rect 6996 8284 7124 8316
rect 7156 8284 7284 8316
rect 7316 8284 7320 8316
rect 6800 8280 7320 8284
rect 7360 8316 7720 8320
rect 7360 8284 7364 8316
rect 7396 8284 7524 8316
rect 7556 8284 7684 8316
rect 7716 8284 7720 8316
rect 7360 8280 7720 8284
rect 5520 8236 7320 8240
rect 5520 8204 5524 8236
rect 5556 8204 5684 8236
rect 5716 8204 5844 8236
rect 5876 8204 6004 8236
rect 6036 8204 6164 8236
rect 6196 8204 6324 8236
rect 6356 8204 6484 8236
rect 6516 8204 6644 8236
rect 6676 8204 6804 8236
rect 6836 8204 6964 8236
rect 6996 8204 7124 8236
rect 7156 8204 7284 8236
rect 7316 8204 7320 8236
rect 5520 8200 7320 8204
rect 7360 8236 7720 8240
rect 7360 8204 7364 8236
rect 7396 8204 7524 8236
rect 7556 8204 7684 8236
rect 7716 8204 7720 8236
rect 7360 8200 7720 8204
rect 5520 8156 7320 8160
rect 5520 8124 5524 8156
rect 5556 8124 5684 8156
rect 5716 8124 5844 8156
rect 5876 8124 6004 8156
rect 6036 8124 6164 8156
rect 6196 8124 6324 8156
rect 6356 8124 6484 8156
rect 6516 8124 6644 8156
rect 6676 8124 6804 8156
rect 6836 8124 6964 8156
rect 6996 8124 7124 8156
rect 7156 8124 7284 8156
rect 7316 8124 7320 8156
rect 5520 8120 7320 8124
rect 7360 8156 7720 8160
rect 7360 8124 7364 8156
rect 7396 8124 7524 8156
rect 7556 8124 7684 8156
rect 7716 8124 7720 8156
rect 7360 8120 7720 8124
rect 5520 8076 7320 8080
rect 5520 8044 5524 8076
rect 5556 8044 5684 8076
rect 5716 8044 5844 8076
rect 5876 8044 6004 8076
rect 6036 8044 6164 8076
rect 6196 8044 6324 8076
rect 6356 8044 6484 8076
rect 6516 8044 6644 8076
rect 6676 8044 6804 8076
rect 6836 8044 6964 8076
rect 6996 8044 7124 8076
rect 7156 8044 7284 8076
rect 7316 8044 7320 8076
rect 5520 8040 7320 8044
rect 7360 8076 7720 8080
rect 7360 8044 7364 8076
rect 7396 8044 7524 8076
rect 7556 8044 7684 8076
rect 7716 8044 7720 8076
rect 7360 8040 7720 8044
rect 5520 7996 7320 8000
rect 5520 7964 5524 7996
rect 5556 7964 5684 7996
rect 5716 7964 5844 7996
rect 5876 7964 6004 7996
rect 6036 7964 6164 7996
rect 6196 7964 6324 7996
rect 6356 7964 6484 7996
rect 6516 7964 6644 7996
rect 6676 7964 6804 7996
rect 6836 7964 6964 7996
rect 6996 7964 7124 7996
rect 7156 7964 7284 7996
rect 7316 7964 7320 7996
rect 5520 7960 7320 7964
rect 7360 7996 7720 8000
rect 7360 7964 7364 7996
rect 7396 7964 7524 7996
rect 7556 7964 7684 7996
rect 7716 7964 7720 7996
rect 7360 7960 7720 7964
rect 5520 7916 7320 7920
rect 5520 7884 5524 7916
rect 5556 7884 5684 7916
rect 5716 7884 5844 7916
rect 5876 7884 6004 7916
rect 6036 7884 6164 7916
rect 6196 7884 6324 7916
rect 6356 7884 6484 7916
rect 6516 7884 6644 7916
rect 6676 7884 6804 7916
rect 6836 7884 6964 7916
rect 6996 7884 7124 7916
rect 7156 7884 7284 7916
rect 7316 7884 7320 7916
rect 5520 7880 7320 7884
rect 7360 7916 7720 7920
rect 7360 7884 7364 7916
rect 7396 7884 7524 7916
rect 7556 7884 7684 7916
rect 7716 7884 7720 7916
rect 7360 7880 7720 7884
rect 5520 7836 7320 7840
rect 5520 7804 5524 7836
rect 5556 7804 5684 7836
rect 5716 7804 5844 7836
rect 5876 7804 6004 7836
rect 6036 7804 6164 7836
rect 6196 7804 6324 7836
rect 6356 7804 6484 7836
rect 6516 7804 6644 7836
rect 6676 7804 6804 7836
rect 6836 7804 6964 7836
rect 6996 7804 7124 7836
rect 7156 7804 7284 7836
rect 7316 7804 7320 7836
rect 5520 7800 7320 7804
rect 7360 7836 7720 7840
rect 7360 7804 7364 7836
rect 7396 7804 7524 7836
rect 7556 7804 7684 7836
rect 7716 7804 7720 7836
rect 7360 7800 7720 7804
rect 5520 7756 7320 7760
rect 5520 7724 5524 7756
rect 5556 7724 5684 7756
rect 5716 7724 5844 7756
rect 5876 7724 6004 7756
rect 6036 7724 6164 7756
rect 6196 7724 6324 7756
rect 6356 7724 6484 7756
rect 6516 7724 6644 7756
rect 6676 7724 6804 7756
rect 6836 7724 6964 7756
rect 6996 7724 7124 7756
rect 7156 7724 7284 7756
rect 7316 7724 7320 7756
rect 5520 7720 7320 7724
rect 7360 7756 7720 7760
rect 7360 7724 7364 7756
rect 7396 7724 7524 7756
rect 7556 7724 7684 7756
rect 7716 7724 7720 7756
rect 7360 7720 7720 7724
rect 5520 7676 7320 7680
rect 5520 7644 5524 7676
rect 5556 7644 5684 7676
rect 5716 7644 5844 7676
rect 5876 7644 6004 7676
rect 6036 7644 6164 7676
rect 6196 7644 6324 7676
rect 6356 7644 6484 7676
rect 6516 7644 6644 7676
rect 6676 7644 6804 7676
rect 6836 7644 6964 7676
rect 6996 7644 7124 7676
rect 7156 7644 7284 7676
rect 7316 7644 7320 7676
rect 5520 7640 7320 7644
rect 7360 7676 7720 7680
rect 7360 7644 7364 7676
rect 7396 7644 7524 7676
rect 7556 7644 7684 7676
rect 7716 7644 7720 7676
rect 7360 7640 7720 7644
rect 5520 7596 7320 7600
rect 5520 7564 5524 7596
rect 5556 7564 5684 7596
rect 5716 7564 5844 7596
rect 5876 7564 6004 7596
rect 6036 7564 6164 7596
rect 6196 7564 6324 7596
rect 6356 7564 6484 7596
rect 6516 7564 6644 7596
rect 6676 7564 6804 7596
rect 6836 7564 6964 7596
rect 6996 7564 7124 7596
rect 7156 7564 7284 7596
rect 7316 7564 7320 7596
rect 5520 7560 7320 7564
rect 7360 7596 7720 7600
rect 7360 7564 7364 7596
rect 7396 7564 7524 7596
rect 7556 7564 7684 7596
rect 7716 7564 7720 7596
rect 7360 7560 7720 7564
rect 5520 7516 7320 7520
rect 5520 7484 5524 7516
rect 5556 7484 5684 7516
rect 5716 7484 5844 7516
rect 5876 7484 6004 7516
rect 6036 7484 6164 7516
rect 6196 7484 6324 7516
rect 6356 7484 6484 7516
rect 6516 7484 6644 7516
rect 6676 7484 6804 7516
rect 6836 7484 6964 7516
rect 6996 7484 7124 7516
rect 7156 7484 7284 7516
rect 7316 7484 7320 7516
rect 5520 7480 7320 7484
rect 7360 7516 7720 7520
rect 7360 7484 7364 7516
rect 7396 7484 7524 7516
rect 7556 7484 7684 7516
rect 7716 7484 7720 7516
rect 7360 7480 7720 7484
rect 5520 7436 7320 7440
rect 5520 7404 5524 7436
rect 5556 7404 5684 7436
rect 5716 7404 5844 7436
rect 5876 7404 6004 7436
rect 6036 7404 6164 7436
rect 6196 7404 6324 7436
rect 6356 7404 6484 7436
rect 6516 7404 6644 7436
rect 6676 7404 6804 7436
rect 6836 7404 6964 7436
rect 6996 7404 7124 7436
rect 7156 7404 7284 7436
rect 7316 7404 7320 7436
rect 5520 7400 7320 7404
rect 7360 7436 7720 7440
rect 7360 7404 7364 7436
rect 7396 7404 7524 7436
rect 7556 7404 7684 7436
rect 7716 7404 7720 7436
rect 7360 7400 7720 7404
rect 5520 7356 7320 7360
rect 5520 7324 5524 7356
rect 5556 7324 5684 7356
rect 5716 7324 5844 7356
rect 5876 7324 6004 7356
rect 6036 7324 6164 7356
rect 6196 7324 6324 7356
rect 6356 7324 6484 7356
rect 6516 7324 6644 7356
rect 6676 7324 6804 7356
rect 6836 7324 6964 7356
rect 6996 7324 7124 7356
rect 7156 7324 7284 7356
rect 7316 7324 7320 7356
rect 5520 7320 7320 7324
rect 7360 7356 7720 7360
rect 7360 7324 7364 7356
rect 7396 7324 7524 7356
rect 7556 7324 7684 7356
rect 7716 7324 7720 7356
rect 7360 7320 7720 7324
rect 5520 7276 7320 7280
rect 5520 7244 5524 7276
rect 5556 7244 5684 7276
rect 5716 7244 5844 7276
rect 5876 7244 6004 7276
rect 6036 7244 6164 7276
rect 6196 7244 6324 7276
rect 6356 7244 6484 7276
rect 6516 7244 6644 7276
rect 6676 7244 6804 7276
rect 6836 7244 6964 7276
rect 6996 7244 7124 7276
rect 7156 7244 7284 7276
rect 7316 7244 7320 7276
rect 5520 7240 7320 7244
rect 7360 7276 7720 7280
rect 7360 7244 7364 7276
rect 7396 7244 7524 7276
rect 7556 7244 7684 7276
rect 7716 7244 7720 7276
rect 7360 7240 7720 7244
rect 5520 7196 7320 7200
rect 5520 7164 5524 7196
rect 5556 7164 5684 7196
rect 5716 7164 5844 7196
rect 5876 7164 6004 7196
rect 6036 7164 6164 7196
rect 6196 7164 6324 7196
rect 6356 7164 6484 7196
rect 6516 7164 6644 7196
rect 6676 7164 6804 7196
rect 6836 7164 6964 7196
rect 6996 7164 7124 7196
rect 7156 7164 7284 7196
rect 7316 7164 7320 7196
rect 5520 7160 7320 7164
rect 7360 7196 7720 7200
rect 7360 7164 7364 7196
rect 7396 7164 7524 7196
rect 7556 7164 7684 7196
rect 7716 7164 7720 7196
rect 7360 7160 7720 7164
rect 6160 7116 7320 7120
rect 6160 7084 6164 7116
rect 6196 7084 6324 7116
rect 6356 7084 6484 7116
rect 6516 7084 6644 7116
rect 6676 7084 6804 7116
rect 6836 7084 6964 7116
rect 6996 7084 7124 7116
rect 7156 7084 7284 7116
rect 7316 7084 7320 7116
rect 6160 7080 7320 7084
rect 7360 7116 7720 7120
rect 7360 7084 7364 7116
rect 7396 7084 7524 7116
rect 7556 7084 7684 7116
rect 7716 7084 7720 7116
rect 7360 7080 7720 7084
rect 5520 7036 7320 7040
rect 5520 7004 5524 7036
rect 5556 7004 5684 7036
rect 5716 7004 5844 7036
rect 5876 7004 6004 7036
rect 6036 7004 6164 7036
rect 6196 7004 6324 7036
rect 6356 7004 6484 7036
rect 6516 7004 6644 7036
rect 6676 7004 6804 7036
rect 6836 7004 6964 7036
rect 6996 7004 7124 7036
rect 7156 7004 7284 7036
rect 7316 7004 7320 7036
rect 5520 7000 7320 7004
rect 7360 7036 7720 7040
rect 7360 7004 7364 7036
rect 7396 7004 7524 7036
rect 7556 7004 7684 7036
rect 7716 7004 7720 7036
rect 7360 7000 7720 7004
rect 5520 6956 7320 6960
rect 5520 6924 5524 6956
rect 5556 6924 5684 6956
rect 5716 6924 5844 6956
rect 5876 6924 6004 6956
rect 6036 6924 6164 6956
rect 6196 6924 6324 6956
rect 6356 6924 6484 6956
rect 6516 6924 6644 6956
rect 6676 6924 6804 6956
rect 6836 6924 6964 6956
rect 6996 6924 7124 6956
rect 7156 6924 7284 6956
rect 7316 6924 7320 6956
rect 5520 6920 7320 6924
rect 7360 6956 7720 6960
rect 7360 6924 7364 6956
rect 7396 6924 7524 6956
rect 7556 6924 7684 6956
rect 7716 6924 7720 6956
rect 7360 6920 7720 6924
rect 6320 6876 7320 6880
rect 6320 6844 6324 6876
rect 6356 6844 6484 6876
rect 6516 6844 6644 6876
rect 6676 6844 6804 6876
rect 6836 6844 6964 6876
rect 6996 6844 7124 6876
rect 7156 6844 7284 6876
rect 7316 6844 7320 6876
rect 6320 6840 7320 6844
rect 7360 6876 7720 6880
rect 7360 6844 7364 6876
rect 7396 6844 7524 6876
rect 7556 6844 7684 6876
rect 7716 6844 7720 6876
rect 7360 6840 7720 6844
rect 5520 6796 7320 6800
rect 5520 6764 5524 6796
rect 5556 6764 5684 6796
rect 5716 6764 5844 6796
rect 5876 6764 6004 6796
rect 6036 6764 6164 6796
rect 6196 6764 6324 6796
rect 6356 6764 6484 6796
rect 6516 6764 6644 6796
rect 6676 6764 6804 6796
rect 6836 6764 6964 6796
rect 6996 6764 7124 6796
rect 7156 6764 7284 6796
rect 7316 6764 7320 6796
rect 5520 6760 7320 6764
rect 7360 6796 7720 6800
rect 7360 6764 7364 6796
rect 7396 6764 7524 6796
rect 7556 6764 7684 6796
rect 7716 6764 7720 6796
rect 7360 6760 7720 6764
rect 5520 6716 7320 6720
rect 5520 6684 5524 6716
rect 5556 6684 5684 6716
rect 5716 6684 5844 6716
rect 5876 6684 6004 6716
rect 6036 6684 6164 6716
rect 6196 6684 6324 6716
rect 6356 6684 6484 6716
rect 6516 6684 6644 6716
rect 6676 6684 6804 6716
rect 6836 6684 6964 6716
rect 6996 6684 7124 6716
rect 7156 6684 7284 6716
rect 7316 6684 7320 6716
rect 5520 6680 7320 6684
rect 7360 6716 7720 6720
rect 7360 6684 7364 6716
rect 7396 6684 7524 6716
rect 7556 6684 7684 6716
rect 7716 6684 7720 6716
rect 7360 6680 7720 6684
rect 5520 6636 7320 6640
rect 5520 6604 5524 6636
rect 5556 6604 5684 6636
rect 5716 6604 5844 6636
rect 5876 6604 6004 6636
rect 6036 6604 6164 6636
rect 6196 6604 6324 6636
rect 6356 6604 6484 6636
rect 6516 6604 6644 6636
rect 6676 6604 6804 6636
rect 6836 6604 6964 6636
rect 6996 6604 7124 6636
rect 7156 6604 7284 6636
rect 7316 6604 7320 6636
rect 5520 6600 7320 6604
rect 7360 6636 7720 6640
rect 7360 6604 7364 6636
rect 7396 6604 7524 6636
rect 7556 6604 7684 6636
rect 7716 6604 7720 6636
rect 7360 6600 7720 6604
rect 5520 6556 7320 6560
rect 5520 6524 5524 6556
rect 5556 6524 5684 6556
rect 5716 6524 5844 6556
rect 5876 6524 6004 6556
rect 6036 6524 6164 6556
rect 6196 6524 6324 6556
rect 6356 6524 6484 6556
rect 6516 6524 6644 6556
rect 6676 6524 6804 6556
rect 6836 6524 6964 6556
rect 6996 6524 7124 6556
rect 7156 6524 7284 6556
rect 7316 6524 7320 6556
rect 5520 6520 7320 6524
rect 7360 6556 7720 6560
rect 7360 6524 7364 6556
rect 7396 6524 7524 6556
rect 7556 6524 7684 6556
rect 7716 6524 7720 6556
rect 7360 6520 7720 6524
rect 5520 6476 7320 6480
rect 5520 6444 5524 6476
rect 5556 6444 5684 6476
rect 5716 6444 5844 6476
rect 5876 6444 6004 6476
rect 6036 6444 6164 6476
rect 6196 6444 6324 6476
rect 6356 6444 6484 6476
rect 6516 6444 6644 6476
rect 6676 6444 6804 6476
rect 6836 6444 6964 6476
rect 6996 6444 7124 6476
rect 7156 6444 7284 6476
rect 7316 6444 7320 6476
rect 5520 6440 7320 6444
rect 7360 6476 7720 6480
rect 7360 6444 7364 6476
rect 7396 6444 7524 6476
rect 7556 6444 7684 6476
rect 7716 6444 7720 6476
rect 7360 6440 7720 6444
rect 6640 6396 7320 6400
rect 6640 6364 6644 6396
rect 6676 6364 6804 6396
rect 6836 6364 6964 6396
rect 6996 6364 7124 6396
rect 7156 6364 7284 6396
rect 7316 6364 7320 6396
rect 6640 6360 7320 6364
rect 7360 6396 7720 6400
rect 7360 6364 7364 6396
rect 7396 6364 7524 6396
rect 7556 6364 7684 6396
rect 7716 6364 7720 6396
rect 7360 6360 7720 6364
rect 5520 6316 7320 6320
rect 5520 6284 5524 6316
rect 5556 6284 5684 6316
rect 5716 6284 5844 6316
rect 5876 6284 6004 6316
rect 6036 6284 6164 6316
rect 6196 6284 6324 6316
rect 6356 6284 6484 6316
rect 6516 6284 6644 6316
rect 6676 6284 6804 6316
rect 6836 6284 6964 6316
rect 6996 6284 7124 6316
rect 7156 6284 7284 6316
rect 7316 6284 7320 6316
rect 5520 6280 7320 6284
rect 7360 6316 7720 6320
rect 7360 6284 7364 6316
rect 7396 6284 7524 6316
rect 7556 6284 7684 6316
rect 7716 6284 7720 6316
rect 7360 6280 7720 6284
rect 5520 6236 7320 6240
rect 5520 6204 5524 6236
rect 5556 6204 5684 6236
rect 5716 6204 5844 6236
rect 5876 6204 6004 6236
rect 6036 6204 6164 6236
rect 6196 6204 6324 6236
rect 6356 6204 6484 6236
rect 6516 6204 6644 6236
rect 6676 6204 6804 6236
rect 6836 6204 6964 6236
rect 6996 6204 7124 6236
rect 7156 6204 7284 6236
rect 7316 6204 7320 6236
rect 5520 6200 7320 6204
rect 7360 6236 7720 6240
rect 7360 6204 7364 6236
rect 7396 6204 7524 6236
rect 7556 6204 7684 6236
rect 7716 6204 7720 6236
rect 7360 6200 7720 6204
rect 5520 6156 7320 6160
rect 5520 6124 5524 6156
rect 5556 6124 5684 6156
rect 5716 6124 5844 6156
rect 5876 6124 6004 6156
rect 6036 6124 6164 6156
rect 6196 6124 6324 6156
rect 6356 6124 6484 6156
rect 6516 6124 6644 6156
rect 6676 6124 6804 6156
rect 6836 6124 6964 6156
rect 6996 6124 7124 6156
rect 7156 6124 7284 6156
rect 7316 6124 7320 6156
rect 5520 6120 7320 6124
rect 7360 6156 7720 6160
rect 7360 6124 7364 6156
rect 7396 6124 7524 6156
rect 7556 6124 7684 6156
rect 7716 6124 7720 6156
rect 7360 6120 7720 6124
rect 7120 6076 7320 6080
rect 7120 6044 7124 6076
rect 7156 6044 7284 6076
rect 7316 6044 7320 6076
rect 7120 6040 7320 6044
rect 7360 6076 7720 6080
rect 7360 6044 7364 6076
rect 7396 6044 7524 6076
rect 7556 6044 7684 6076
rect 7716 6044 7720 6076
rect 7360 6040 7720 6044
rect 5520 5996 7320 6000
rect 5520 5964 5524 5996
rect 5556 5964 5684 5996
rect 5716 5964 5844 5996
rect 5876 5964 6004 5996
rect 6036 5964 6164 5996
rect 6196 5964 6324 5996
rect 6356 5964 6484 5996
rect 6516 5964 6644 5996
rect 6676 5964 6804 5996
rect 6836 5964 6964 5996
rect 6996 5964 7124 5996
rect 7156 5964 7284 5996
rect 7316 5964 7320 5996
rect 5520 5960 7320 5964
rect 7360 5996 7720 6000
rect 7360 5964 7364 5996
rect 7396 5964 7524 5996
rect 7556 5964 7684 5996
rect 7716 5964 7720 5996
rect 7360 5960 7720 5964
rect 6960 5916 7320 5920
rect 6960 5884 6964 5916
rect 6996 5884 7124 5916
rect 7156 5884 7284 5916
rect 7316 5884 7320 5916
rect 6960 5880 7320 5884
rect 7360 5916 7720 5920
rect 7360 5884 7364 5916
rect 7396 5884 7524 5916
rect 7556 5884 7684 5916
rect 7716 5884 7720 5916
rect 7360 5880 7720 5884
rect 5520 5836 7320 5840
rect 5520 5804 5524 5836
rect 5556 5804 5684 5836
rect 5716 5804 5844 5836
rect 5876 5804 6004 5836
rect 6036 5804 6164 5836
rect 6196 5804 6324 5836
rect 6356 5804 6484 5836
rect 6516 5804 6644 5836
rect 6676 5804 6804 5836
rect 6836 5804 6964 5836
rect 6996 5804 7124 5836
rect 7156 5804 7284 5836
rect 7316 5804 7320 5836
rect 5520 5800 7320 5804
rect 7360 5836 7720 5840
rect 7360 5804 7364 5836
rect 7396 5804 7524 5836
rect 7556 5804 7684 5836
rect 7716 5804 7720 5836
rect 7360 5800 7720 5804
rect 5520 5756 7320 5760
rect 5520 5724 5524 5756
rect 5556 5724 5684 5756
rect 5716 5724 5844 5756
rect 5876 5724 6004 5756
rect 6036 5724 6164 5756
rect 6196 5724 6324 5756
rect 6356 5724 6484 5756
rect 6516 5724 6644 5756
rect 6676 5724 6804 5756
rect 6836 5724 6964 5756
rect 6996 5724 7124 5756
rect 7156 5724 7284 5756
rect 7316 5724 7320 5756
rect 5520 5720 7320 5724
rect 7360 5756 7720 5760
rect 7360 5724 7364 5756
rect 7396 5724 7524 5756
rect 7556 5724 7684 5756
rect 7716 5724 7720 5756
rect 7360 5720 7720 5724
rect 5520 5676 7320 5680
rect 5520 5644 5524 5676
rect 5556 5644 5684 5676
rect 5716 5644 5844 5676
rect 5876 5644 6004 5676
rect 6036 5644 6164 5676
rect 6196 5644 6324 5676
rect 6356 5644 6484 5676
rect 6516 5644 6644 5676
rect 6676 5644 6804 5676
rect 6836 5644 6964 5676
rect 6996 5644 7124 5676
rect 7156 5644 7284 5676
rect 7316 5644 7320 5676
rect 5520 5640 7320 5644
rect 7360 5676 7720 5680
rect 7360 5644 7364 5676
rect 7396 5644 7524 5676
rect 7556 5644 7684 5676
rect 7716 5644 7720 5676
rect 7360 5640 7720 5644
rect 5520 5596 7320 5600
rect 5520 5564 5524 5596
rect 5556 5564 5684 5596
rect 5716 5564 5844 5596
rect 5876 5564 6004 5596
rect 6036 5564 6164 5596
rect 6196 5564 6324 5596
rect 6356 5564 6484 5596
rect 6516 5564 6644 5596
rect 6676 5564 6804 5596
rect 6836 5564 6964 5596
rect 6996 5564 7124 5596
rect 7156 5564 7284 5596
rect 7316 5564 7320 5596
rect 5520 5560 7320 5564
rect 7360 5596 7720 5600
rect 7360 5564 7364 5596
rect 7396 5564 7524 5596
rect 7556 5564 7684 5596
rect 7716 5564 7720 5596
rect 7360 5560 7720 5564
rect 5520 5516 7320 5520
rect 5520 5484 5524 5516
rect 5556 5484 5684 5516
rect 5716 5484 5844 5516
rect 5876 5484 6004 5516
rect 6036 5484 6164 5516
rect 6196 5484 6324 5516
rect 6356 5484 6484 5516
rect 6516 5484 6644 5516
rect 6676 5484 6804 5516
rect 6836 5484 6964 5516
rect 6996 5484 7124 5516
rect 7156 5484 7284 5516
rect 7316 5484 7320 5516
rect 5520 5480 7320 5484
rect 7360 5516 7720 5520
rect 7360 5484 7364 5516
rect 7396 5484 7524 5516
rect 7556 5484 7684 5516
rect 7716 5484 7720 5516
rect 7360 5480 7720 5484
rect 5520 5436 7320 5440
rect 5520 5404 5524 5436
rect 5556 5404 5684 5436
rect 5716 5404 5844 5436
rect 5876 5404 6004 5436
rect 6036 5404 6164 5436
rect 6196 5404 6324 5436
rect 6356 5404 6484 5436
rect 6516 5404 6644 5436
rect 6676 5404 6804 5436
rect 6836 5404 6964 5436
rect 6996 5404 7124 5436
rect 7156 5404 7284 5436
rect 7316 5404 7320 5436
rect 5520 5400 7320 5404
rect 7360 5436 7720 5440
rect 7360 5404 7364 5436
rect 7396 5404 7524 5436
rect 7556 5404 7684 5436
rect 7716 5404 7720 5436
rect 7360 5400 7720 5404
rect 5520 5356 7320 5360
rect 5520 5324 5524 5356
rect 5556 5324 5684 5356
rect 5716 5324 5844 5356
rect 5876 5324 6004 5356
rect 6036 5324 6164 5356
rect 6196 5324 6324 5356
rect 6356 5324 6484 5356
rect 6516 5324 6644 5356
rect 6676 5324 6804 5356
rect 6836 5324 6964 5356
rect 6996 5324 7124 5356
rect 7156 5324 7284 5356
rect 7316 5324 7320 5356
rect 5520 5320 7320 5324
rect 7360 5356 7720 5360
rect 7360 5324 7364 5356
rect 7396 5324 7524 5356
rect 7556 5324 7684 5356
rect 7716 5324 7720 5356
rect 7360 5320 7720 5324
rect 5520 5276 7320 5280
rect 5520 5244 5524 5276
rect 5556 5244 5684 5276
rect 5716 5244 5844 5276
rect 5876 5244 6004 5276
rect 6036 5244 6164 5276
rect 6196 5244 6324 5276
rect 6356 5244 6484 5276
rect 6516 5244 6644 5276
rect 6676 5244 6804 5276
rect 6836 5244 6964 5276
rect 6996 5244 7124 5276
rect 7156 5244 7284 5276
rect 7316 5244 7320 5276
rect 5520 5240 7320 5244
rect 7360 5276 7720 5280
rect 7360 5244 7364 5276
rect 7396 5244 7524 5276
rect 7556 5244 7684 5276
rect 7716 5244 7720 5276
rect 7360 5240 7720 5244
rect 5520 5196 7320 5200
rect 5520 5164 5524 5196
rect 5556 5164 5684 5196
rect 5716 5164 5844 5196
rect 5876 5164 6004 5196
rect 6036 5164 6164 5196
rect 6196 5164 6324 5196
rect 6356 5164 6484 5196
rect 6516 5164 6644 5196
rect 6676 5164 6804 5196
rect 6836 5164 6964 5196
rect 6996 5164 7124 5196
rect 7156 5164 7284 5196
rect 7316 5164 7320 5196
rect 5520 5160 7320 5164
rect 7360 5196 7720 5200
rect 7360 5164 7364 5196
rect 7396 5164 7524 5196
rect 7556 5164 7684 5196
rect 7716 5164 7720 5196
rect 7360 5160 7720 5164
rect 5520 5116 7320 5120
rect 5520 5084 5524 5116
rect 5556 5084 5684 5116
rect 5716 5084 5844 5116
rect 5876 5084 6004 5116
rect 6036 5084 6164 5116
rect 6196 5084 6324 5116
rect 6356 5084 6484 5116
rect 6516 5084 6644 5116
rect 6676 5084 6804 5116
rect 6836 5084 6964 5116
rect 6996 5084 7124 5116
rect 7156 5084 7284 5116
rect 7316 5084 7320 5116
rect 5520 5080 7320 5084
rect 7360 5116 7720 5120
rect 7360 5084 7364 5116
rect 7396 5084 7524 5116
rect 7556 5084 7684 5116
rect 7716 5084 7720 5116
rect 7360 5080 7720 5084
rect 5520 5036 7320 5040
rect 5520 5004 5524 5036
rect 5556 5004 5684 5036
rect 5716 5004 5844 5036
rect 5876 5004 6004 5036
rect 6036 5004 6164 5036
rect 6196 5004 6324 5036
rect 6356 5004 6484 5036
rect 6516 5004 6644 5036
rect 6676 5004 6804 5036
rect 6836 5004 6964 5036
rect 6996 5004 7124 5036
rect 7156 5004 7284 5036
rect 7316 5004 7320 5036
rect 5520 5000 7320 5004
rect 7360 5036 7720 5040
rect 7360 5004 7364 5036
rect 7396 5004 7524 5036
rect 7556 5004 7684 5036
rect 7716 5004 7720 5036
rect 7360 5000 7720 5004
rect 5520 4956 7320 4960
rect 5520 4924 5524 4956
rect 5556 4924 5684 4956
rect 5716 4924 5844 4956
rect 5876 4924 6004 4956
rect 6036 4924 6164 4956
rect 6196 4924 6324 4956
rect 6356 4924 6484 4956
rect 6516 4924 6644 4956
rect 6676 4924 6804 4956
rect 6836 4924 6964 4956
rect 6996 4924 7124 4956
rect 7156 4924 7284 4956
rect 7316 4924 7320 4956
rect 5520 4920 7320 4924
rect 7360 4956 7720 4960
rect 7360 4924 7364 4956
rect 7396 4924 7524 4956
rect 7556 4924 7684 4956
rect 7716 4924 7720 4956
rect 7360 4920 7720 4924
rect 5520 4876 7320 4880
rect 5520 4844 5524 4876
rect 5556 4844 5684 4876
rect 5716 4844 5844 4876
rect 5876 4844 6004 4876
rect 6036 4844 6164 4876
rect 6196 4844 6324 4876
rect 6356 4844 6484 4876
rect 6516 4844 6644 4876
rect 6676 4844 6804 4876
rect 6836 4844 6964 4876
rect 6996 4844 7124 4876
rect 7156 4844 7284 4876
rect 7316 4844 7320 4876
rect 5520 4840 7320 4844
rect 7360 4876 7720 4880
rect 7360 4844 7364 4876
rect 7396 4844 7524 4876
rect 7556 4844 7684 4876
rect 7716 4844 7720 4876
rect 7360 4840 7720 4844
rect 5520 4796 7320 4800
rect 5520 4764 5524 4796
rect 5556 4764 5684 4796
rect 5716 4764 5844 4796
rect 5876 4764 6004 4796
rect 6036 4764 6164 4796
rect 6196 4764 6324 4796
rect 6356 4764 6484 4796
rect 6516 4764 6644 4796
rect 6676 4764 6804 4796
rect 6836 4764 6964 4796
rect 6996 4764 7124 4796
rect 7156 4764 7284 4796
rect 7316 4764 7320 4796
rect 5520 4760 7320 4764
rect 7360 4796 7720 4800
rect 7360 4764 7364 4796
rect 7396 4764 7524 4796
rect 7556 4764 7684 4796
rect 7716 4764 7720 4796
rect 7360 4760 7720 4764
rect 6160 4716 7320 4720
rect 6160 4684 6164 4716
rect 6196 4684 6324 4716
rect 6356 4684 6484 4716
rect 6516 4684 6644 4716
rect 6676 4684 6804 4716
rect 6836 4684 6964 4716
rect 6996 4684 7124 4716
rect 7156 4684 7284 4716
rect 7316 4684 7320 4716
rect 6160 4680 7320 4684
rect 7360 4716 7720 4720
rect 7360 4684 7364 4716
rect 7396 4684 7524 4716
rect 7556 4684 7684 4716
rect 7716 4684 7720 4716
rect 7360 4680 7720 4684
rect 5520 4636 7320 4640
rect 5520 4604 5524 4636
rect 5556 4604 5684 4636
rect 5716 4604 5844 4636
rect 5876 4604 6004 4636
rect 6036 4604 6164 4636
rect 6196 4604 6324 4636
rect 6356 4604 6484 4636
rect 6516 4604 6644 4636
rect 6676 4604 6804 4636
rect 6836 4604 6964 4636
rect 6996 4604 7124 4636
rect 7156 4604 7284 4636
rect 7316 4604 7320 4636
rect 5520 4600 7320 4604
rect 7360 4636 7720 4640
rect 7360 4604 7364 4636
rect 7396 4604 7524 4636
rect 7556 4604 7684 4636
rect 7716 4604 7720 4636
rect 7360 4600 7720 4604
rect 5520 4556 7320 4560
rect 5520 4524 5524 4556
rect 5556 4524 5684 4556
rect 5716 4524 5844 4556
rect 5876 4524 6004 4556
rect 6036 4524 6164 4556
rect 6196 4524 6324 4556
rect 6356 4524 6484 4556
rect 6516 4524 6644 4556
rect 6676 4524 6804 4556
rect 6836 4524 6964 4556
rect 6996 4524 7124 4556
rect 7156 4524 7284 4556
rect 7316 4524 7320 4556
rect 5520 4520 7320 4524
rect 7360 4556 7720 4560
rect 7360 4524 7364 4556
rect 7396 4524 7524 4556
rect 7556 4524 7684 4556
rect 7716 4524 7720 4556
rect 7360 4520 7720 4524
rect 6320 4476 7320 4480
rect 6320 4444 6324 4476
rect 6356 4444 6484 4476
rect 6516 4444 6644 4476
rect 6676 4444 6804 4476
rect 6836 4444 6964 4476
rect 6996 4444 7124 4476
rect 7156 4444 7284 4476
rect 7316 4444 7320 4476
rect 6320 4440 7320 4444
rect 7360 4476 7720 4480
rect 7360 4444 7364 4476
rect 7396 4444 7524 4476
rect 7556 4444 7684 4476
rect 7716 4444 7720 4476
rect 7360 4440 7720 4444
rect 5520 4396 7320 4400
rect 5520 4364 5524 4396
rect 5556 4364 5684 4396
rect 5716 4364 5844 4396
rect 5876 4364 6004 4396
rect 6036 4364 6164 4396
rect 6196 4364 6324 4396
rect 6356 4364 6484 4396
rect 6516 4364 6644 4396
rect 6676 4364 6804 4396
rect 6836 4364 6964 4396
rect 6996 4364 7124 4396
rect 7156 4364 7284 4396
rect 7316 4364 7320 4396
rect 5520 4360 7320 4364
rect 7360 4396 7720 4400
rect 7360 4364 7364 4396
rect 7396 4364 7524 4396
rect 7556 4364 7684 4396
rect 7716 4364 7720 4396
rect 7360 4360 7720 4364
rect 5520 4316 7320 4320
rect 5520 4284 5524 4316
rect 5556 4284 5684 4316
rect 5716 4284 5844 4316
rect 5876 4284 6004 4316
rect 6036 4284 6164 4316
rect 6196 4284 6324 4316
rect 6356 4284 6484 4316
rect 6516 4284 6644 4316
rect 6676 4284 6804 4316
rect 6836 4284 6964 4316
rect 6996 4284 7124 4316
rect 7156 4284 7284 4316
rect 7316 4284 7320 4316
rect 5520 4280 7320 4284
rect 7360 4316 7720 4320
rect 7360 4284 7364 4316
rect 7396 4284 7524 4316
rect 7556 4284 7684 4316
rect 7716 4284 7720 4316
rect 7360 4280 7720 4284
rect 5520 4236 7320 4240
rect 5520 4204 5524 4236
rect 5556 4204 5684 4236
rect 5716 4204 5844 4236
rect 5876 4204 6004 4236
rect 6036 4204 6164 4236
rect 6196 4204 6324 4236
rect 6356 4204 6484 4236
rect 6516 4204 6644 4236
rect 6676 4204 6804 4236
rect 6836 4204 6964 4236
rect 6996 4204 7124 4236
rect 7156 4204 7284 4236
rect 7316 4204 7320 4236
rect 5520 4200 7320 4204
rect 7360 4236 7720 4240
rect 7360 4204 7364 4236
rect 7396 4204 7524 4236
rect 7556 4204 7684 4236
rect 7716 4204 7720 4236
rect 7360 4200 7720 4204
rect 5520 4156 7320 4160
rect 5520 4124 5524 4156
rect 5556 4124 5684 4156
rect 5716 4124 5844 4156
rect 5876 4124 6004 4156
rect 6036 4124 6164 4156
rect 6196 4124 6324 4156
rect 6356 4124 6484 4156
rect 6516 4124 6644 4156
rect 6676 4124 6804 4156
rect 6836 4124 6964 4156
rect 6996 4124 7124 4156
rect 7156 4124 7284 4156
rect 7316 4124 7320 4156
rect 5520 4120 7320 4124
rect 7360 4156 7720 4160
rect 7360 4124 7364 4156
rect 7396 4124 7524 4156
rect 7556 4124 7684 4156
rect 7716 4124 7720 4156
rect 7360 4120 7720 4124
rect 5520 4076 7320 4080
rect 5520 4044 5524 4076
rect 5556 4044 5684 4076
rect 5716 4044 5844 4076
rect 5876 4044 6004 4076
rect 6036 4044 6164 4076
rect 6196 4044 6324 4076
rect 6356 4044 6484 4076
rect 6516 4044 6644 4076
rect 6676 4044 6804 4076
rect 6836 4044 6964 4076
rect 6996 4044 7124 4076
rect 7156 4044 7284 4076
rect 7316 4044 7320 4076
rect 5520 4040 7320 4044
rect 7360 4076 7720 4080
rect 7360 4044 7364 4076
rect 7396 4044 7524 4076
rect 7556 4044 7684 4076
rect 7716 4044 7720 4076
rect 7360 4040 7720 4044
rect 6480 3996 7320 4000
rect 6480 3964 6484 3996
rect 6516 3964 6644 3996
rect 6676 3964 6804 3996
rect 6836 3964 6964 3996
rect 6996 3964 7124 3996
rect 7156 3964 7284 3996
rect 7316 3964 7320 3996
rect 6480 3960 7320 3964
rect 7360 3996 7720 4000
rect 7360 3964 7364 3996
rect 7396 3964 7524 3996
rect 7556 3964 7684 3996
rect 7716 3964 7720 3996
rect 7360 3960 7720 3964
rect 5520 3916 7320 3920
rect 5520 3884 5524 3916
rect 5556 3884 5684 3916
rect 5716 3884 5844 3916
rect 5876 3884 6004 3916
rect 6036 3884 6164 3916
rect 6196 3884 6324 3916
rect 6356 3884 6484 3916
rect 6516 3884 6644 3916
rect 6676 3884 6804 3916
rect 6836 3884 6964 3916
rect 6996 3884 7124 3916
rect 7156 3884 7284 3916
rect 7316 3884 7320 3916
rect 5520 3880 7320 3884
rect 7360 3916 7720 3920
rect 7360 3884 7364 3916
rect 7396 3884 7524 3916
rect 7556 3884 7684 3916
rect 7716 3884 7720 3916
rect 7360 3880 7720 3884
rect 5520 3836 7320 3840
rect 5520 3804 5524 3836
rect 5556 3804 5684 3836
rect 5716 3804 5844 3836
rect 5876 3804 6004 3836
rect 6036 3804 6164 3836
rect 6196 3804 6324 3836
rect 6356 3804 6484 3836
rect 6516 3804 6644 3836
rect 6676 3804 6804 3836
rect 6836 3804 6964 3836
rect 6996 3804 7124 3836
rect 7156 3804 7284 3836
rect 7316 3804 7320 3836
rect 5520 3800 7320 3804
rect 7360 3836 7720 3840
rect 7360 3804 7364 3836
rect 7396 3804 7524 3836
rect 7556 3804 7684 3836
rect 7716 3804 7720 3836
rect 7360 3800 7720 3804
rect 5520 3756 7320 3760
rect 5520 3724 5524 3756
rect 5556 3724 5684 3756
rect 5716 3724 5844 3756
rect 5876 3724 6004 3756
rect 6036 3724 6164 3756
rect 6196 3724 6324 3756
rect 6356 3724 6484 3756
rect 6516 3724 6644 3756
rect 6676 3724 6804 3756
rect 6836 3724 6964 3756
rect 6996 3724 7124 3756
rect 7156 3724 7284 3756
rect 7316 3724 7320 3756
rect 5520 3720 7320 3724
rect 7360 3756 7720 3760
rect 7360 3724 7364 3756
rect 7396 3724 7524 3756
rect 7556 3724 7684 3756
rect 7716 3724 7720 3756
rect 7360 3720 7720 3724
rect 7120 3676 7320 3680
rect 7120 3644 7124 3676
rect 7156 3644 7284 3676
rect 7316 3644 7320 3676
rect 7120 3640 7320 3644
rect 7360 3676 7720 3680
rect 7360 3644 7364 3676
rect 7396 3644 7524 3676
rect 7556 3644 7684 3676
rect 7716 3644 7720 3676
rect 7360 3640 7720 3644
rect 5520 3596 7320 3600
rect 5520 3564 5524 3596
rect 5556 3564 5684 3596
rect 5716 3564 5844 3596
rect 5876 3564 6004 3596
rect 6036 3564 6164 3596
rect 6196 3564 6324 3596
rect 6356 3564 6484 3596
rect 6516 3564 6644 3596
rect 6676 3564 6804 3596
rect 6836 3564 6964 3596
rect 6996 3564 7124 3596
rect 7156 3564 7284 3596
rect 7316 3564 7320 3596
rect 5520 3560 7320 3564
rect 7360 3596 7720 3600
rect 7360 3564 7364 3596
rect 7396 3564 7524 3596
rect 7556 3564 7684 3596
rect 7716 3564 7720 3596
rect 7360 3560 7720 3564
rect 6800 3516 7320 3520
rect 6800 3484 6804 3516
rect 6836 3484 6964 3516
rect 6996 3484 7124 3516
rect 7156 3484 7284 3516
rect 7316 3484 7320 3516
rect 6800 3480 7320 3484
rect 7360 3516 7720 3520
rect 7360 3484 7364 3516
rect 7396 3484 7524 3516
rect 7556 3484 7684 3516
rect 7716 3484 7720 3516
rect 7360 3480 7720 3484
rect 5520 3436 7320 3440
rect 5520 3404 5524 3436
rect 5556 3404 5684 3436
rect 5716 3404 5844 3436
rect 5876 3404 6004 3436
rect 6036 3404 6164 3436
rect 6196 3404 6324 3436
rect 6356 3404 6484 3436
rect 6516 3404 6644 3436
rect 6676 3404 6804 3436
rect 6836 3404 6964 3436
rect 6996 3404 7124 3436
rect 7156 3404 7284 3436
rect 7316 3404 7320 3436
rect 5520 3400 7320 3404
rect 7360 3436 7720 3440
rect 7360 3404 7364 3436
rect 7396 3404 7524 3436
rect 7556 3404 7684 3436
rect 7716 3404 7720 3436
rect 7360 3400 7720 3404
rect 5520 3356 7320 3360
rect 5520 3324 5524 3356
rect 5556 3324 5684 3356
rect 5716 3324 5844 3356
rect 5876 3324 6004 3356
rect 6036 3324 6164 3356
rect 6196 3324 6324 3356
rect 6356 3324 6484 3356
rect 6516 3324 6644 3356
rect 6676 3324 6804 3356
rect 6836 3324 6964 3356
rect 6996 3324 7124 3356
rect 7156 3324 7284 3356
rect 7316 3324 7320 3356
rect 5520 3320 7320 3324
rect 7360 3356 7720 3360
rect 7360 3324 7364 3356
rect 7396 3324 7524 3356
rect 7556 3324 7684 3356
rect 7716 3324 7720 3356
rect 7360 3320 7720 3324
rect 5520 3276 7320 3280
rect 5520 3244 5524 3276
rect 5556 3244 5684 3276
rect 5716 3244 5844 3276
rect 5876 3244 6004 3276
rect 6036 3244 6164 3276
rect 6196 3244 6324 3276
rect 6356 3244 6484 3276
rect 6516 3244 6644 3276
rect 6676 3244 6804 3276
rect 6836 3244 6964 3276
rect 6996 3244 7124 3276
rect 7156 3244 7284 3276
rect 7316 3244 7320 3276
rect 5520 3240 7320 3244
rect 7360 3276 7720 3280
rect 7360 3244 7364 3276
rect 7396 3244 7524 3276
rect 7556 3244 7684 3276
rect 7716 3244 7720 3276
rect 7360 3240 7720 3244
rect 5520 3196 7320 3200
rect 5520 3164 5524 3196
rect 5556 3164 5684 3196
rect 5716 3164 5844 3196
rect 5876 3164 6004 3196
rect 6036 3164 6164 3196
rect 6196 3164 6324 3196
rect 6356 3164 6484 3196
rect 6516 3164 6644 3196
rect 6676 3164 6804 3196
rect 6836 3164 6964 3196
rect 6996 3164 7124 3196
rect 7156 3164 7284 3196
rect 7316 3164 7320 3196
rect 5520 3160 7320 3164
rect 7360 3196 7720 3200
rect 7360 3164 7364 3196
rect 7396 3164 7524 3196
rect 7556 3164 7684 3196
rect 7716 3164 7720 3196
rect 7360 3160 7720 3164
rect 5520 3116 7320 3120
rect 5520 3084 5524 3116
rect 5556 3084 5684 3116
rect 5716 3084 5844 3116
rect 5876 3084 6004 3116
rect 6036 3084 6164 3116
rect 6196 3084 6324 3116
rect 6356 3084 6484 3116
rect 6516 3084 6644 3116
rect 6676 3084 6804 3116
rect 6836 3084 6964 3116
rect 6996 3084 7124 3116
rect 7156 3084 7284 3116
rect 7316 3084 7320 3116
rect 5520 3080 7320 3084
rect 7360 3116 7720 3120
rect 7360 3084 7364 3116
rect 7396 3084 7524 3116
rect 7556 3084 7684 3116
rect 7716 3084 7720 3116
rect 7360 3080 7720 3084
rect 5520 3036 7320 3040
rect 5520 3004 5524 3036
rect 5556 3004 5684 3036
rect 5716 3004 5844 3036
rect 5876 3004 6004 3036
rect 6036 3004 6164 3036
rect 6196 3004 6324 3036
rect 6356 3004 6484 3036
rect 6516 3004 6644 3036
rect 6676 3004 6804 3036
rect 6836 3004 6964 3036
rect 6996 3004 7124 3036
rect 7156 3004 7284 3036
rect 7316 3004 7320 3036
rect 5520 3000 7320 3004
rect 7360 3036 7720 3040
rect 7360 3004 7364 3036
rect 7396 3004 7524 3036
rect 7556 3004 7684 3036
rect 7716 3004 7720 3036
rect 7360 3000 7720 3004
rect 5520 2956 7320 2960
rect 5520 2924 5524 2956
rect 5556 2924 5684 2956
rect 5716 2924 5844 2956
rect 5876 2924 6004 2956
rect 6036 2924 6164 2956
rect 6196 2924 6324 2956
rect 6356 2924 6484 2956
rect 6516 2924 6644 2956
rect 6676 2924 6804 2956
rect 6836 2924 6964 2956
rect 6996 2924 7124 2956
rect 7156 2924 7284 2956
rect 7316 2924 7320 2956
rect 5520 2920 7320 2924
rect 7360 2956 7720 2960
rect 7360 2924 7364 2956
rect 7396 2924 7524 2956
rect 7556 2924 7684 2956
rect 7716 2924 7720 2956
rect 7360 2920 7720 2924
rect 5520 2876 7320 2880
rect 5520 2844 5524 2876
rect 5556 2844 5684 2876
rect 5716 2844 5844 2876
rect 5876 2844 6004 2876
rect 6036 2844 6164 2876
rect 6196 2844 6324 2876
rect 6356 2844 6484 2876
rect 6516 2844 6644 2876
rect 6676 2844 6804 2876
rect 6836 2844 6964 2876
rect 6996 2844 7124 2876
rect 7156 2844 7284 2876
rect 7316 2844 7320 2876
rect 5520 2840 7320 2844
rect 7360 2876 7720 2880
rect 7360 2844 7364 2876
rect 7396 2844 7524 2876
rect 7556 2844 7684 2876
rect 7716 2844 7720 2876
rect 7360 2840 7720 2844
rect 5520 2796 7320 2800
rect 5520 2764 5524 2796
rect 5556 2764 5684 2796
rect 5716 2764 5844 2796
rect 5876 2764 6004 2796
rect 6036 2764 6164 2796
rect 6196 2764 6324 2796
rect 6356 2764 6484 2796
rect 6516 2764 6644 2796
rect 6676 2764 6804 2796
rect 6836 2764 6964 2796
rect 6996 2764 7124 2796
rect 7156 2764 7284 2796
rect 7316 2764 7320 2796
rect 5520 2760 7320 2764
rect 7360 2796 7720 2800
rect 7360 2764 7364 2796
rect 7396 2764 7524 2796
rect 7556 2764 7684 2796
rect 7716 2764 7720 2796
rect 7360 2760 7720 2764
rect 5520 2716 7320 2720
rect 5520 2684 5524 2716
rect 5556 2684 5684 2716
rect 5716 2684 5844 2716
rect 5876 2684 6004 2716
rect 6036 2684 6164 2716
rect 6196 2684 6324 2716
rect 6356 2684 6484 2716
rect 6516 2684 6644 2716
rect 6676 2684 6804 2716
rect 6836 2684 6964 2716
rect 6996 2684 7124 2716
rect 7156 2684 7284 2716
rect 7316 2684 7320 2716
rect 5520 2680 7320 2684
rect 7360 2716 7720 2720
rect 7360 2684 7364 2716
rect 7396 2684 7524 2716
rect 7556 2684 7684 2716
rect 7716 2684 7720 2716
rect 7360 2680 7720 2684
rect 5520 2636 7320 2640
rect 5520 2604 5524 2636
rect 5556 2604 5684 2636
rect 5716 2604 5844 2636
rect 5876 2604 6004 2636
rect 6036 2604 6164 2636
rect 6196 2604 6324 2636
rect 6356 2604 6484 2636
rect 6516 2604 6644 2636
rect 6676 2604 6804 2636
rect 6836 2604 6964 2636
rect 6996 2604 7124 2636
rect 7156 2604 7284 2636
rect 7316 2604 7320 2636
rect 5520 2600 7320 2604
rect 7360 2636 7720 2640
rect 7360 2604 7364 2636
rect 7396 2604 7524 2636
rect 7556 2604 7684 2636
rect 7716 2604 7720 2636
rect 7360 2600 7720 2604
rect 5520 2556 7320 2560
rect 5520 2524 5524 2556
rect 5556 2524 5684 2556
rect 5716 2524 5844 2556
rect 5876 2524 6004 2556
rect 6036 2524 6164 2556
rect 6196 2524 6324 2556
rect 6356 2524 6484 2556
rect 6516 2524 6644 2556
rect 6676 2524 6804 2556
rect 6836 2524 6964 2556
rect 6996 2524 7124 2556
rect 7156 2524 7284 2556
rect 7316 2524 7320 2556
rect 5520 2520 7320 2524
rect 7360 2556 7720 2560
rect 7360 2524 7364 2556
rect 7396 2524 7524 2556
rect 7556 2524 7684 2556
rect 7716 2524 7720 2556
rect 7360 2520 7720 2524
rect 5520 2476 7320 2480
rect 5520 2444 5524 2476
rect 5556 2444 5684 2476
rect 5716 2444 5844 2476
rect 5876 2444 6004 2476
rect 6036 2444 6164 2476
rect 6196 2444 6324 2476
rect 6356 2444 6484 2476
rect 6516 2444 6644 2476
rect 6676 2444 6804 2476
rect 6836 2444 6964 2476
rect 6996 2444 7124 2476
rect 7156 2444 7284 2476
rect 7316 2444 7320 2476
rect 5520 2440 7320 2444
rect 7360 2476 7720 2480
rect 7360 2444 7364 2476
rect 7396 2444 7524 2476
rect 7556 2444 7684 2476
rect 7716 2444 7720 2476
rect 7360 2440 7720 2444
rect 5520 2396 7320 2400
rect 5520 2364 5524 2396
rect 5556 2364 5684 2396
rect 5716 2364 5844 2396
rect 5876 2364 6004 2396
rect 6036 2364 6164 2396
rect 6196 2364 6324 2396
rect 6356 2364 6484 2396
rect 6516 2364 6644 2396
rect 6676 2364 6804 2396
rect 6836 2364 6964 2396
rect 6996 2364 7124 2396
rect 7156 2364 7284 2396
rect 7316 2364 7320 2396
rect 5520 2360 7320 2364
rect 7360 2396 7720 2400
rect 7360 2364 7364 2396
rect 7396 2364 7524 2396
rect 7556 2364 7684 2396
rect 7716 2364 7720 2396
rect 7360 2360 7720 2364
rect 6160 2316 7320 2320
rect 6160 2284 6164 2316
rect 6196 2284 6324 2316
rect 6356 2284 6484 2316
rect 6516 2284 6644 2316
rect 6676 2284 6804 2316
rect 6836 2284 6964 2316
rect 6996 2284 7124 2316
rect 7156 2284 7284 2316
rect 7316 2284 7320 2316
rect 6160 2280 7320 2284
rect 7360 2316 7720 2320
rect 7360 2284 7364 2316
rect 7396 2284 7524 2316
rect 7556 2284 7684 2316
rect 7716 2284 7720 2316
rect 7360 2280 7720 2284
rect 5520 2236 7320 2240
rect 5520 2204 5524 2236
rect 5556 2204 5684 2236
rect 5716 2204 5844 2236
rect 5876 2204 6004 2236
rect 6036 2204 6164 2236
rect 6196 2204 6324 2236
rect 6356 2204 6484 2236
rect 6516 2204 6644 2236
rect 6676 2204 6804 2236
rect 6836 2204 6964 2236
rect 6996 2204 7124 2236
rect 7156 2204 7284 2236
rect 7316 2204 7320 2236
rect 5520 2200 7320 2204
rect 7360 2236 7720 2240
rect 7360 2204 7364 2236
rect 7396 2204 7524 2236
rect 7556 2204 7684 2236
rect 7716 2204 7720 2236
rect 7360 2200 7720 2204
rect 5520 2156 7320 2160
rect 5520 2124 5524 2156
rect 5556 2124 5684 2156
rect 5716 2124 5844 2156
rect 5876 2124 6004 2156
rect 6036 2124 6164 2156
rect 6196 2124 6324 2156
rect 6356 2124 6484 2156
rect 6516 2124 6644 2156
rect 6676 2124 6804 2156
rect 6836 2124 6964 2156
rect 6996 2124 7124 2156
rect 7156 2124 7284 2156
rect 7316 2124 7320 2156
rect 5520 2120 7320 2124
rect 7360 2156 7720 2160
rect 7360 2124 7364 2156
rect 7396 2124 7524 2156
rect 7556 2124 7684 2156
rect 7716 2124 7720 2156
rect 7360 2120 7720 2124
rect 5520 2076 7320 2080
rect 5520 2044 5524 2076
rect 5556 2044 5684 2076
rect 5716 2044 5844 2076
rect 5876 2044 6004 2076
rect 6036 2044 6164 2076
rect 6196 2044 6324 2076
rect 6356 2044 6484 2076
rect 6516 2044 6644 2076
rect 6676 2044 6804 2076
rect 6836 2044 6964 2076
rect 6996 2044 7124 2076
rect 7156 2044 7284 2076
rect 7316 2044 7320 2076
rect 5520 2040 7320 2044
rect 7360 2076 7720 2080
rect 7360 2044 7364 2076
rect 7396 2044 7524 2076
rect 7556 2044 7684 2076
rect 7716 2044 7720 2076
rect 7360 2040 7720 2044
rect 5520 1996 7320 2000
rect 5520 1964 5524 1996
rect 5556 1964 5684 1996
rect 5716 1964 5844 1996
rect 5876 1964 6004 1996
rect 6036 1964 6164 1996
rect 6196 1964 6324 1996
rect 6356 1964 6484 1996
rect 6516 1964 6644 1996
rect 6676 1964 6804 1996
rect 6836 1964 6964 1996
rect 6996 1964 7124 1996
rect 7156 1964 7284 1996
rect 7316 1964 7320 1996
rect 5520 1960 7320 1964
rect 7360 1996 7720 2000
rect 7360 1964 7364 1996
rect 7396 1964 7524 1996
rect 7556 1964 7684 1996
rect 7716 1964 7720 1996
rect 7360 1960 7720 1964
rect 5520 1916 7320 1920
rect 5520 1884 5524 1916
rect 5556 1884 5684 1916
rect 5716 1884 5844 1916
rect 5876 1884 6004 1916
rect 6036 1884 6164 1916
rect 6196 1884 6324 1916
rect 6356 1884 6484 1916
rect 6516 1884 6644 1916
rect 6676 1884 6804 1916
rect 6836 1884 6964 1916
rect 6996 1884 7124 1916
rect 7156 1884 7284 1916
rect 7316 1884 7320 1916
rect 5520 1880 7320 1884
rect 7360 1916 7720 1920
rect 7360 1884 7364 1916
rect 7396 1884 7524 1916
rect 7556 1884 7684 1916
rect 7716 1884 7720 1916
rect 7360 1880 7720 1884
rect 5520 1836 7320 1840
rect 5520 1804 5524 1836
rect 5556 1804 5684 1836
rect 5716 1804 5844 1836
rect 5876 1804 6004 1836
rect 6036 1804 6164 1836
rect 6196 1804 6324 1836
rect 6356 1804 6484 1836
rect 6516 1804 6644 1836
rect 6676 1804 6804 1836
rect 6836 1804 6964 1836
rect 6996 1804 7124 1836
rect 7156 1804 7284 1836
rect 7316 1804 7320 1836
rect 5520 1800 7320 1804
rect 7360 1836 7720 1840
rect 7360 1804 7364 1836
rect 7396 1804 7524 1836
rect 7556 1804 7684 1836
rect 7716 1804 7720 1836
rect 7360 1800 7720 1804
rect 5520 1756 7320 1760
rect 5520 1724 5524 1756
rect 5556 1724 5684 1756
rect 5716 1724 5844 1756
rect 5876 1724 6004 1756
rect 6036 1724 6164 1756
rect 6196 1724 6324 1756
rect 6356 1724 6484 1756
rect 6516 1724 6644 1756
rect 6676 1724 6804 1756
rect 6836 1724 6964 1756
rect 6996 1724 7124 1756
rect 7156 1724 7284 1756
rect 7316 1724 7320 1756
rect 5520 1720 7320 1724
rect 7360 1756 7720 1760
rect 7360 1724 7364 1756
rect 7396 1724 7524 1756
rect 7556 1724 7684 1756
rect 7716 1724 7720 1756
rect 7360 1720 7720 1724
rect 5520 1676 7320 1680
rect 5520 1644 5524 1676
rect 5556 1644 5684 1676
rect 5716 1644 5844 1676
rect 5876 1644 6004 1676
rect 6036 1644 6164 1676
rect 6196 1644 6324 1676
rect 6356 1644 6484 1676
rect 6516 1644 6644 1676
rect 6676 1644 6804 1676
rect 6836 1644 6964 1676
rect 6996 1644 7124 1676
rect 7156 1644 7284 1676
rect 7316 1644 7320 1676
rect 5520 1640 7320 1644
rect 7360 1676 7720 1680
rect 7360 1644 7364 1676
rect 7396 1644 7524 1676
rect 7556 1644 7684 1676
rect 7716 1644 7720 1676
rect 7360 1640 7720 1644
rect 6000 1596 7320 1600
rect 6000 1564 6004 1596
rect 6036 1564 6164 1596
rect 6196 1564 6324 1596
rect 6356 1564 6484 1596
rect 6516 1564 6644 1596
rect 6676 1564 6804 1596
rect 6836 1564 6964 1596
rect 6996 1564 7124 1596
rect 7156 1564 7284 1596
rect 7316 1564 7320 1596
rect 6000 1560 7320 1564
rect 7360 1596 7720 1600
rect 7360 1564 7364 1596
rect 7396 1564 7524 1596
rect 7556 1564 7684 1596
rect 7716 1564 7720 1596
rect 7360 1560 7720 1564
rect 5520 1516 7320 1520
rect 5520 1484 5524 1516
rect 5556 1484 5684 1516
rect 5716 1484 5844 1516
rect 5876 1484 6004 1516
rect 6036 1484 6164 1516
rect 6196 1484 6324 1516
rect 6356 1484 6484 1516
rect 6516 1484 6644 1516
rect 6676 1484 6804 1516
rect 6836 1484 6964 1516
rect 6996 1484 7124 1516
rect 7156 1484 7284 1516
rect 7316 1484 7320 1516
rect 5520 1480 7320 1484
rect 7360 1516 7720 1520
rect 7360 1484 7364 1516
rect 7396 1484 7524 1516
rect 7556 1484 7684 1516
rect 7716 1484 7720 1516
rect 7360 1480 7720 1484
rect 5520 1436 7320 1440
rect 5520 1404 5524 1436
rect 5556 1404 5684 1436
rect 5716 1404 5844 1436
rect 5876 1404 6004 1436
rect 6036 1404 6164 1436
rect 6196 1404 6324 1436
rect 6356 1404 6484 1436
rect 6516 1404 6644 1436
rect 6676 1404 6804 1436
rect 6836 1404 6964 1436
rect 6996 1404 7124 1436
rect 7156 1404 7284 1436
rect 7316 1404 7320 1436
rect 5520 1400 7320 1404
rect 7360 1436 7720 1440
rect 7360 1404 7364 1436
rect 7396 1404 7524 1436
rect 7556 1404 7684 1436
rect 7716 1404 7720 1436
rect 7360 1400 7720 1404
rect 5520 1356 7320 1360
rect 5520 1324 5524 1356
rect 5556 1324 5684 1356
rect 5716 1324 5844 1356
rect 5876 1324 6004 1356
rect 6036 1324 6164 1356
rect 6196 1324 6324 1356
rect 6356 1324 6484 1356
rect 6516 1324 6644 1356
rect 6676 1324 6804 1356
rect 6836 1324 6964 1356
rect 6996 1324 7124 1356
rect 7156 1324 7284 1356
rect 7316 1324 7320 1356
rect 5520 1320 7320 1324
rect 7360 1356 7720 1360
rect 7360 1324 7364 1356
rect 7396 1324 7524 1356
rect 7556 1324 7684 1356
rect 7716 1324 7720 1356
rect 7360 1320 7720 1324
rect 5680 1276 7320 1280
rect 5680 1244 5684 1276
rect 5716 1244 5844 1276
rect 5876 1244 6004 1276
rect 6036 1244 6164 1276
rect 6196 1244 6324 1276
rect 6356 1244 6484 1276
rect 6516 1244 6644 1276
rect 6676 1244 6804 1276
rect 6836 1244 6964 1276
rect 6996 1244 7124 1276
rect 7156 1244 7284 1276
rect 7316 1244 7320 1276
rect 5680 1240 7320 1244
rect 7360 1276 7720 1280
rect 7360 1244 7364 1276
rect 7396 1244 7524 1276
rect 7556 1244 7684 1276
rect 7716 1244 7720 1276
rect 7360 1240 7720 1244
rect 5520 1196 7320 1200
rect 5520 1164 5524 1196
rect 5556 1164 5684 1196
rect 5716 1164 5844 1196
rect 5876 1164 6004 1196
rect 6036 1164 6164 1196
rect 6196 1164 6324 1196
rect 6356 1164 6484 1196
rect 6516 1164 6644 1196
rect 6676 1164 6804 1196
rect 6836 1164 6964 1196
rect 6996 1164 7124 1196
rect 7156 1164 7284 1196
rect 7316 1164 7320 1196
rect 5520 1160 7320 1164
rect 7360 1196 7720 1200
rect 7360 1164 7364 1196
rect 7396 1164 7524 1196
rect 7556 1164 7684 1196
rect 7716 1164 7720 1196
rect 7360 1160 7720 1164
rect 5520 1116 7320 1120
rect 5520 1084 5524 1116
rect 5556 1084 5684 1116
rect 5716 1084 5844 1116
rect 5876 1084 6004 1116
rect 6036 1084 6164 1116
rect 6196 1084 6324 1116
rect 6356 1084 6484 1116
rect 6516 1084 6644 1116
rect 6676 1084 6804 1116
rect 6836 1084 6964 1116
rect 6996 1084 7124 1116
rect 7156 1084 7284 1116
rect 7316 1084 7320 1116
rect 5520 1080 7320 1084
rect 7360 1116 7720 1120
rect 7360 1084 7364 1116
rect 7396 1084 7524 1116
rect 7556 1084 7684 1116
rect 7716 1084 7720 1116
rect 7360 1080 7720 1084
rect 5520 1036 7320 1040
rect 5520 1004 5524 1036
rect 5556 1004 5684 1036
rect 5716 1004 5844 1036
rect 5876 1004 6004 1036
rect 6036 1004 6164 1036
rect 6196 1004 6324 1036
rect 6356 1004 6484 1036
rect 6516 1004 6644 1036
rect 6676 1004 6804 1036
rect 6836 1004 6964 1036
rect 6996 1004 7124 1036
rect 7156 1004 7284 1036
rect 7316 1004 7320 1036
rect 5520 1000 7320 1004
rect 7360 1036 7720 1040
rect 7360 1004 7364 1036
rect 7396 1004 7524 1036
rect 7556 1004 7684 1036
rect 7716 1004 7720 1036
rect 7360 1000 7720 1004
rect 5520 956 7320 960
rect 5520 924 5524 956
rect 5556 924 5684 956
rect 5716 924 5844 956
rect 5876 924 6004 956
rect 6036 924 6164 956
rect 6196 924 6324 956
rect 6356 924 6484 956
rect 6516 924 6644 956
rect 6676 924 6804 956
rect 6836 924 6964 956
rect 6996 924 7124 956
rect 7156 924 7284 956
rect 7316 924 7320 956
rect 5520 920 7320 924
rect 7360 956 7720 960
rect 7360 924 7364 956
rect 7396 924 7524 956
rect 7556 924 7684 956
rect 7716 924 7720 956
rect 7360 920 7720 924
rect 5520 876 7320 880
rect 5520 844 5524 876
rect 5556 844 5684 876
rect 5716 844 5844 876
rect 5876 844 6004 876
rect 6036 844 6164 876
rect 6196 844 6324 876
rect 6356 844 6484 876
rect 6516 844 6644 876
rect 6676 844 6804 876
rect 6836 844 6964 876
rect 6996 844 7124 876
rect 7156 844 7284 876
rect 7316 844 7320 876
rect 5520 840 7320 844
rect 7360 876 7720 880
rect 7360 844 7364 876
rect 7396 844 7524 876
rect 7556 844 7684 876
rect 7716 844 7720 876
rect 7360 840 7720 844
rect 5520 796 7320 800
rect 5520 764 5524 796
rect 5556 764 5684 796
rect 5716 764 5844 796
rect 5876 764 6004 796
rect 6036 764 6164 796
rect 6196 764 6324 796
rect 6356 764 6484 796
rect 6516 764 6644 796
rect 6676 764 6804 796
rect 6836 764 6964 796
rect 6996 764 7124 796
rect 7156 764 7284 796
rect 7316 764 7320 796
rect 5520 760 7320 764
rect 7360 796 7720 800
rect 7360 764 7364 796
rect 7396 764 7524 796
rect 7556 764 7684 796
rect 7716 764 7720 796
rect 7360 760 7720 764
rect 5840 716 7320 720
rect 5840 684 5844 716
rect 5876 684 6004 716
rect 6036 684 6164 716
rect 6196 684 6324 716
rect 6356 684 6484 716
rect 6516 684 6644 716
rect 6676 684 6804 716
rect 6836 684 6964 716
rect 6996 684 7124 716
rect 7156 684 7284 716
rect 7316 684 7320 716
rect 5840 680 7320 684
rect 7360 716 7720 720
rect 7360 684 7364 716
rect 7396 684 7524 716
rect 7556 684 7684 716
rect 7716 684 7720 716
rect 7360 680 7720 684
rect 5520 596 7320 600
rect 5520 564 5524 596
rect 5556 564 5684 596
rect 5716 564 5844 596
rect 5876 564 6004 596
rect 6036 564 6164 596
rect 6196 564 6324 596
rect 6356 564 6484 596
rect 6516 564 6644 596
rect 6676 564 6804 596
rect 6836 564 6964 596
rect 6996 564 7124 596
rect 7156 564 7284 596
rect 7316 564 7320 596
rect 5520 560 7320 564
rect 7360 596 7720 600
rect 7360 564 7364 596
rect 7396 564 7524 596
rect 7556 564 7684 596
rect 7716 564 7720 596
rect 7360 560 7720 564
rect 5520 516 7320 520
rect 5520 484 5524 516
rect 5556 484 5684 516
rect 5716 484 5844 516
rect 5876 484 6004 516
rect 6036 484 6164 516
rect 6196 484 6324 516
rect 6356 484 6484 516
rect 6516 484 6644 516
rect 6676 484 6804 516
rect 6836 484 6964 516
rect 6996 484 7124 516
rect 7156 484 7284 516
rect 7316 484 7320 516
rect 5520 480 7320 484
rect 7360 516 7720 520
rect 7360 484 7364 516
rect 7396 484 7524 516
rect 7556 484 7684 516
rect 7716 484 7720 516
rect 7360 480 7720 484
rect 5680 436 7320 440
rect 5680 404 5684 436
rect 5716 404 5844 436
rect 5876 404 6004 436
rect 6036 404 6164 436
rect 6196 404 6324 436
rect 6356 404 6484 436
rect 6516 404 6644 436
rect 6676 404 6804 436
rect 6836 404 6964 436
rect 6996 404 7124 436
rect 7156 404 7284 436
rect 7316 404 7320 436
rect 5680 400 7320 404
rect 7360 436 7720 440
rect 7360 404 7364 436
rect 7396 404 7524 436
rect 7556 404 7684 436
rect 7716 404 7720 436
rect 7360 400 7720 404
rect 5520 356 7320 360
rect 5520 324 5524 356
rect 5556 324 5684 356
rect 5716 324 5844 356
rect 5876 324 6004 356
rect 6036 324 6164 356
rect 6196 324 6324 356
rect 6356 324 6484 356
rect 6516 324 6644 356
rect 6676 324 6804 356
rect 6836 324 6964 356
rect 6996 324 7124 356
rect 7156 324 7284 356
rect 7316 324 7320 356
rect 5520 320 7320 324
rect 7360 356 7720 360
rect 7360 324 7364 356
rect 7396 324 7524 356
rect 7556 324 7684 356
rect 7716 324 7720 356
rect 7360 320 7720 324
rect 5520 276 7320 280
rect 5520 244 5524 276
rect 5556 244 5684 276
rect 5716 244 5844 276
rect 5876 244 6004 276
rect 6036 244 6164 276
rect 6196 244 6324 276
rect 6356 244 6484 276
rect 6516 244 6644 276
rect 6676 244 6804 276
rect 6836 244 6964 276
rect 6996 244 7124 276
rect 7156 244 7284 276
rect 7316 244 7320 276
rect 5520 240 7320 244
rect 7360 276 7720 280
rect 7360 244 7364 276
rect 7396 244 7524 276
rect 7556 244 7684 276
rect 7716 244 7720 276
rect 7360 240 7720 244
rect 5520 196 7320 200
rect 5520 164 5524 196
rect 5556 164 5684 196
rect 5716 164 5844 196
rect 5876 164 6004 196
rect 6036 164 6164 196
rect 6196 164 6324 196
rect 6356 164 6484 196
rect 6516 164 6644 196
rect 6676 164 6804 196
rect 6836 164 6964 196
rect 6996 164 7124 196
rect 7156 164 7284 196
rect 7316 164 7320 196
rect 5520 160 7320 164
rect 7360 196 7720 200
rect 7360 164 7364 196
rect 7396 164 7524 196
rect 7556 164 7684 196
rect 7716 164 7720 196
rect 7360 160 7720 164
rect 5520 116 7320 120
rect 5520 84 5524 116
rect 5556 84 5684 116
rect 5716 84 5844 116
rect 5876 84 6004 116
rect 6036 84 6164 116
rect 6196 84 6324 116
rect 6356 84 6484 116
rect 6516 84 6644 116
rect 6676 84 6804 116
rect 6836 84 6964 116
rect 6996 84 7124 116
rect 7156 84 7284 116
rect 7316 84 7320 116
rect 5520 80 7320 84
rect 7360 116 7720 120
rect 7360 84 7364 116
rect 7396 84 7524 116
rect 7556 84 7684 116
rect 7716 84 7720 116
rect 7360 80 7720 84
rect 5520 36 7320 40
rect 5520 4 5524 36
rect 5556 4 5684 36
rect 5716 4 5844 36
rect 5876 4 6004 36
rect 6036 4 6164 36
rect 6196 4 6324 36
rect 6356 4 6484 36
rect 6516 4 6644 36
rect 6676 4 6804 36
rect 6836 4 6964 36
rect 6996 4 7124 36
rect 7156 4 7284 36
rect 7316 4 7320 36
rect 5520 0 7320 4
rect 7360 36 7720 40
rect 7360 4 7364 36
rect 7396 4 7524 36
rect 7556 4 7684 36
rect 7716 4 7720 36
rect 7360 0 7720 4
<< via4 >>
rect 120 16920 240 17040
rect 760 16680 880 16800
<< metal5 >>
rect 80 17040 280 17080
rect 80 16920 120 17040
rect 240 16920 280 17040
rect 80 16600 280 16920
rect 720 16800 920 17080
rect 720 16680 760 16800
rect 880 16680 920 16800
rect 720 16600 920 16680
rect 80 15120 280 15160
rect 720 15120 920 15160
rect 1360 15120 1560 15160
rect 2000 15120 2200 15160
rect 2640 15120 2840 15160
rect 3280 15120 3480 15160
rect 3920 15120 4120 15160
rect 4560 15120 4760 15160
rect 5200 15120 5400 15160
rect 80 13640 280 13680
rect 720 13640 920 13680
rect 1360 13640 1560 13680
rect 2000 13640 2200 13680
rect 2640 13640 2840 13680
rect 3280 13640 3480 13680
rect 3920 13640 4120 13680
rect 4560 13640 4760 13680
rect 5200 13640 5400 13680
rect 80 12160 280 12200
rect 720 12160 920 12200
rect 1360 12160 1560 12200
rect 2000 12160 2200 12200
rect 2640 12160 2840 12200
rect 3280 12160 3480 12200
rect 3920 12160 4120 12200
rect 4560 12160 4760 12200
rect 5200 12160 5400 12200
rect 80 10080 280 10120
rect 720 10080 920 10120
rect 1360 10080 1560 10120
rect 2000 10080 2200 10120
rect 2640 10080 2840 10120
rect 3280 10080 3480 10120
rect 3920 10080 4120 10120
rect 4560 10080 4760 10120
rect 5200 10080 5400 10120
rect 80 8000 280 8040
rect 720 8000 920 8040
rect 1360 8000 1560 8040
rect 2000 8000 2200 8040
rect 2640 8000 2840 8040
rect 3280 8000 3480 8040
rect 3920 8000 4120 8040
rect 4560 8000 4760 8040
rect 5200 8000 5400 8040
rect 80 5600 280 5640
rect 720 5600 920 5640
rect 1360 5600 1560 5640
rect 2000 5600 2200 5640
rect 2640 5600 2840 5640
rect 3280 5600 3480 5640
rect 3920 5600 4120 5640
rect 4560 5600 4760 5640
rect 5200 5600 5400 5640
rect 80 3200 280 3240
rect 720 3200 920 3240
rect 1360 3200 1560 3240
rect 2000 3200 2200 3240
rect 2640 3200 2840 3240
rect 3280 3200 3480 3240
rect 3920 3200 4120 3240
rect 4560 3200 4760 3240
rect 5200 3200 5400 3240
rect 80 800 280 840
rect 720 800 920 840
rect 1360 800 1560 840
rect 2000 800 2200 840
rect 2640 800 2840 840
rect 3280 800 3480 840
rect 3920 800 4120 840
rect 4560 800 4760 840
rect 5200 800 5400 840
rect 80 -40 280 0
rect 720 -40 920 0
use opamp_coreb2  opamp_coreb2_1
timestamp 1637857574
transform 1 0 240 0 1 7160
box -240 -1520 5240 840
use opamp_coreb2  opamp_coreb2_0
timestamp 1637857574
transform 1 0 240 0 1 4760
box -240 -1520 5240 840
use opamp_corea2  a2
timestamp 1637779110
transform 1 0 240 0 1 2360
box -240 -1520 5240 840
use opamp_corec  cp
timestamp 1637779139
transform 1 0 240 0 1 9560
box -240 -1520 5240 520
use opamp_corec  cm
timestamp 1637779139
transform 1 0 240 0 1 11640
box -240 -1520 5240 520
use opamp_cored  dp
timestamp 1637789704
transform 1 0 240 0 1 13720
box -240 -1520 5240 -80
use opamp_cored  dm
timestamp 1637789704
transform 1 0 240 0 1 15200
box -240 -1520 5240 -80
use opamp_coree  e
timestamp 1637788580
transform 1 0 240 0 1 16680
box -240 -1520 5240 -80
use opamp_corea1  a1
timestamp 1637806411
transform 1 0 240 0 1 1520
box -240 -1520 5240 -720
<< labels >>
rlabel metal5 80 -40 280 0 0 vdda
port 15 nsew
rlabel metal5 720 -40 920 0 0 vssa
port 16 nsew
rlabel metal3 5600 -40 5640 0 0 gna
port 1 nsew
rlabel metal3 5760 -40 5800 0 0 gnb
port 2 nsew
rlabel metal3 5920 -40 5960 0 0 gpb
port 3 nsew
rlabel metal3 6080 -40 6120 0 0 gpa
port 4 nsew
rlabel metal3 6240 -40 6280 0 0 x
port 5 nsew
rlabel metal3 6400 -40 6440 0 0 ip
port 6 nsew
rlabel metal3 6560 -40 6600 0 0 im
port 7 nsew
rlabel metal3 6720 -40 6760 0 0 yp
port 8 nsew
rlabel metal3 6880 -40 6920 0 0 ym
port 9 nsew
rlabel metal3 7040 -40 7080 0 0 zn
port 10 nsew
rlabel metal3 7200 -40 7240 0 0 zp
port 11 nsew
rlabel metal3 7360 -40 7400 0 0 out
rlabel metal3 7440 -40 7480 0 0 dn
port 12 nsew
rlabel metal3 7520 -40 7560 0 0 out
rlabel metal3 7600 -40 7640 0 0 dp
port 13 nsew
rlabel metal3 7680 -40 7720 0 0 out
port 14 nsew
<< end >>
