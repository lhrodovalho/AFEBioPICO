* lna-ota buffer testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "lna_ota.spice"

vdd vdd 0 1.8
vss vss 0 0.0
ecm cm vss vdd vss 0.5

vin in cm dc 0 ac 1 SINE(0 0.9 0.5k 0 0 0)

* DUT
IB ib vss 10n
RIB vdd ib 100Meg
*VB ib vss 1.2
X0 out in out ib vdd vss lna_ota
CL out cm 1p

.save v(in) v(out) v(ib) v(x0.x) v(x0.y) i(vdd)
*.option gmin=1e-12
.option scale=1e-6
.control

	op
	print in out ib x0.x x0.y i(vdd)

	dc vin -0.9 0.9 10m
	let dc_vo = v(out)
	wrdata lna_ota_dc_vo.txt dc_vo
	plot dc_vo

	ac dec 10 1m 1Meg
	plot vdb(out)

	tran 10u 4m
	let tran_vi = v(in)
	let tran_vo = v(out)
	wrdata lna_ota_tran.txt tran_vi tran_vo
	plot tran_vi tran_vo
	plot ib x0.y
    
.endc

.end
