* NGSPICE file created from opamp.ext - technology: sky130A

.subckt p1_8 D G S B SUB
X0 D G a7 B sky130_fd_pr__pfet_01v8_lvt ad=3.75e+11p pd=3.5e+06u as=7.5e+11p ps=7e+06u w=3e+06u l=8e+06u
X1 a6 G a5 B sky130_fd_pr__pfet_01v8_lvt ad=7.5e+11p pd=7e+06u as=7.5e+11p ps=7e+06u w=3e+06u l=8e+06u
X2 S G a1 B sky130_fd_pr__pfet_01v8_lvt ad=3.75e+11p pd=3.5e+06u as=7.5e+11p ps=7e+06u w=3e+06u l=8e+06u
X3 a6 G a7 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X4 a2 G a3 B sky130_fd_pr__pfet_01v8_lvt ad=7.5e+11p pd=7e+06u as=7.5e+11p ps=7e+06u w=3e+06u l=8e+06u
X5 a2 G a1 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X6 a4 G a5 B sky130_fd_pr__pfet_01v8_lvt ad=7.5e+11p pd=7e+06u as=0p ps=0u w=3e+06u l=8e+06u
X7 a4 G a3 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
.ends

.subckt p8_1 D G S B SUB
X0 S G D B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=2.8e+07u as=3e+12p ps=2.8e+07u w=3e+06u l=8e+06u
X1 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X2 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X3 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X4 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X5 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X6 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X7 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
.ends

.subckt n8_1 D G S B
X0 D G S B sky130_fd_pr__nfet_01v8_lvt ad=1e+12p pd=1.2e+07u as=1e+12p ps=1.2e+07u w=1e+06u l=8e+06u
X1 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X2 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X3 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X4 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X5 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X6 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X7 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
.ends

.subckt n1_8 D G S B
X0 a5 G a6 B sky130_fd_pr__nfet_01v8_lvt ad=2.5e+11p pd=3e+06u as=2.5e+11p ps=3e+06u w=1e+06u l=8e+06u
X1 a1 G a2 B sky130_fd_pr__nfet_01v8_lvt ad=2.5e+11p pd=3e+06u as=2.5e+11p ps=3e+06u w=1e+06u l=8e+06u
X2 a1 G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.25e+11p ps=1.5e+06u w=1e+06u l=8e+06u
X3 a7 G D B sky130_fd_pr__nfet_01v8_lvt ad=2.5e+11p pd=3e+06u as=1.25e+11p ps=1.5e+06u w=1e+06u l=8e+06u
X4 a3 G a4 B sky130_fd_pr__nfet_01v8_lvt ad=2.5e+11p pd=3e+06u as=2.5e+11p ps=3e+06u w=1e+06u l=8e+06u
X5 a5 G a4 B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X6 a3 G a2 B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X7 a7 G a6 B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
.ends

.subckt opamp inm inp out ib vdda gnda vssa
Xp1_8_5 b p1 vdda vdda vssa p1_8
Xpa2_1 ib ib p1 vdda vssa p8_1
Xpd2_1 x inp xp vdda vssa p8_1
Xpd2_2 x inp xp vdda vssa p8_1
Xn8_1_0 n2 n2 n1 vssa n8_1
Xn8_1_1 a a xm vssa n8_1
Xn8_1_2 c a xp vssa n8_1
Xn8_1_3 c a xp vssa n8_1
Xn8_1_4 a a xm vssa n8_1
Xn8_1_5 c n2 b vssa n8_1
Xnf4_1 xp a vssa vssa n1_8
Xpc1_1 x p1 vdda vdda vssa p1_8
Xn8_1_6 out c vssa vssa n8_1
Xpf1_1 b p1 vdda vdda vssa p1_8
Xnf4_2 xp a vssa vssa n1_8
Xn8_1_7 vssa n1 vssa vssa n8_1
Xnf2_1 c n2 b vssa n8_1
Xn8_1_8 vssa n1 vssa vssa n8_1
Xnb3_1 n2 n2 n1 vssa n8_1
Xn1_8_0 n1 n1 vssa vssa n1_8
Xne3_1 a a xm vssa n8_1
Xn1_8_1 vssa n1 vssa vssa n1_8
Xp8_1_0 ib ib p1 vdda vssa p8_1
Xn1_8_2 xm a vssa vssa n1_8
Xne3_2 a a xm vssa n8_1
Xp8_1_1 x inm xm vdda vssa p8_1
Xn1_8_3 xp a vssa vssa n1_8
Xp8_1_2 x inp xp vdda vssa p8_1
Xn1_8_4 xp a vssa vssa n1_8
Xna4_1 vssa n1 vssa vssa n1_8
Xp8_1_3 x inp xp vdda vssa p8_1
Xn1_8_5 xm a vssa vssa n1_8
Xng4_1 out c vssa vssa n8_1
Xpd1_1 x p1 vdda vdda vssa p1_8
Xpa1_1 p1 p1 vdda vdda vssa p1_8
Xp8_1_4 x inm xm vdda vssa p8_1
Xpg1_1 out b vdda vdda vssa p8_1
Xp8_1_5 b ib c vdda vssa p8_1
Xp8_1_6 out b vdda vdda vssa p8_1
Xp8_1_7 vdda p1 vdda vdda vssa p8_1
Xp8_1_8 vdda p1 vdda vdda vssa p8_1
Xpc2_1 x inm xm vdda vssa p8_1
Xpf2_1 b ib c vdda vssa p8_1
Xpc2_2 x inm xm vdda vssa p8_1
Xnf3_1 c a xp vssa n8_1
Xp1_8_0 p1 p1 vdda vdda vssa p1_8
Xnf3_2 c a xp vssa n8_1
Xp1_8_1 n2 p1 vdda vdda vssa p1_8
Xp1_8_2 x p1 vdda vdda vssa p1_8
Xnb4_1 n1 n1 vssa vssa n1_8
Xp1_8_3 x p1 vdda vdda vssa p1_8
Xp1_8_4 a p1 vdda vdda vssa p1_8
Xne4_2 xm a vssa vssa n1_8
Xpe1_1 a p1 vdda vdda vssa p1_8
Xne4_1 xm a vssa vssa n1_8
Xpb1_1 n2 p1 vdda vdda vssa p1_8
.ends

