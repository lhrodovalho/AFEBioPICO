magic
tech sky130A
timestamp 1638148091
<< error_p >>
rect 10080 4927 10553 4930
rect 10080 3200 10596 3236
rect 10080 3180 10553 3193
rect 10080 3147 10520 3160
rect 10484 2676 10520 3147
rect 10080 2640 10520 2676
rect 10540 2620 10553 3180
rect 10560 3160 10596 3200
rect 10080 2607 10553 2620
rect 10080 2480 10596 2516
rect 10080 2460 10553 2473
rect 10080 2427 10520 2440
rect 10484 1956 10520 2427
rect 10080 1920 10520 1956
rect 10540 1900 10553 2460
rect 10560 2440 10596 2480
rect 10080 1887 10553 1900
rect 10080 1760 10596 1796
rect 10080 1740 10553 1753
rect 10080 1707 10520 1720
rect 10484 1236 10520 1707
rect 10080 1200 10520 1236
rect 10540 1180 10553 1740
rect 10560 1720 10596 1760
rect 10080 1167 10553 1180
<< error_s >>
rect 4 12640 4196 12676
rect 4 12600 40 12640
rect 47 12620 4153 12633
rect 47 12060 60 12620
rect 80 12587 4120 12600
rect 80 12116 116 12587
rect 4107 12116 4120 12587
rect 80 12080 4120 12116
rect 4140 12060 4153 12620
rect 4160 12080 4196 12640
rect 6404 12640 10596 12676
rect 6404 12600 6440 12640
rect 6447 12620 10553 12633
rect 47 12047 4153 12060
rect 6447 12060 6460 12620
rect 6480 12587 10520 12600
rect 6480 12116 6516 12587
rect 10507 12116 10520 12587
rect 6480 12080 10520 12116
rect 10540 12060 10553 12620
rect 10560 12080 10596 12640
rect 6447 12047 10553 12060
rect 4 11920 4196 11956
rect 4 11880 40 11920
rect 47 11900 4153 11913
rect 47 11340 60 11900
rect 80 11867 4120 11880
rect 80 11396 116 11867
rect 4107 11396 4120 11867
rect 80 11360 4120 11396
rect 4140 11340 4153 11900
rect 4160 11360 4196 11920
rect 6404 11920 10596 11956
rect 6404 11880 6440 11920
rect 6447 11900 10553 11913
rect 47 11327 4153 11340
rect 6447 11340 6460 11900
rect 6480 11867 10520 11880
rect 6480 11396 6516 11867
rect 10507 11396 10520 11867
rect 6480 11360 10520 11396
rect 10540 11340 10553 11900
rect 10560 11360 10596 11920
rect 6447 11327 10553 11340
rect 4 10600 4196 10636
rect 4 10560 40 10600
rect 47 10580 4153 10593
rect 47 9620 60 10580
rect 80 10547 4120 10560
rect 80 9676 116 10547
rect 4107 9676 4120 10547
rect 80 9640 4120 9676
rect 4140 9620 4153 10580
rect 4160 9640 4196 10600
rect 6404 10600 10596 10636
rect 6404 10560 6440 10600
rect 6447 10580 10553 10593
rect 47 9607 4153 9620
rect 6447 9620 6460 10580
rect 6480 10547 10520 10560
rect 6480 9676 6516 10547
rect 10507 9676 10520 10547
rect 6480 9640 10520 9676
rect 10540 9620 10553 10580
rect 10560 9640 10596 10600
rect 6447 9607 10553 9620
rect 4 9480 4196 9516
rect 4 9440 40 9480
rect 47 9460 4153 9473
rect 47 8500 60 9460
rect 80 9427 4120 9440
rect 80 8556 116 9427
rect 4107 8556 4120 9427
rect 80 8520 4120 8556
rect 4140 8500 4153 9460
rect 4160 8520 4196 9480
rect 6404 9480 10596 9516
rect 6404 9440 6440 9480
rect 6447 9460 10553 9473
rect 47 8487 4153 8500
rect 6447 8500 6460 9460
rect 6480 9427 10520 9440
rect 6480 8556 6516 9427
rect 10507 8556 10520 9427
rect 6480 8520 10520 8556
rect 10540 8500 10553 9460
rect 10560 8520 10596 9480
rect 6447 8487 10553 8500
rect 4 7560 4196 7596
rect 4 7520 40 7560
rect 47 7540 4153 7553
rect 47 6980 60 7540
rect 80 7507 4120 7520
rect 80 7036 116 7507
rect 4107 7036 4120 7507
rect 80 7000 4120 7036
rect 4140 6980 4153 7540
rect 4160 7000 4196 7560
rect 6404 7560 10596 7596
rect 6404 7520 6440 7560
rect 6447 7540 10553 7553
rect 47 6967 4153 6980
rect 6447 6980 6460 7540
rect 6480 7507 10520 7520
rect 6480 7036 6516 7507
rect 10507 7036 10520 7507
rect 6480 7000 10520 7036
rect 10540 6980 10553 7540
rect 10560 7000 10596 7560
rect 6447 6967 10553 6980
rect 4 6840 4196 6876
rect 4 6800 40 6840
rect 47 6820 4153 6833
rect 47 6260 60 6820
rect 80 6787 4120 6800
rect 80 6316 116 6787
rect 4107 6316 4120 6787
rect 80 6280 4120 6316
rect 4140 6260 4153 6820
rect 4160 6280 4196 6840
rect 6404 6840 10596 6876
rect 6404 6800 6440 6840
rect 6447 6820 10553 6833
rect 47 6247 4153 6260
rect 6447 6260 6460 6820
rect 6480 6787 10520 6800
rect 6480 6316 6516 6787
rect 10507 6316 10520 6787
rect 6480 6280 10520 6316
rect 10540 6260 10553 6820
rect 10560 6280 10596 6840
rect 6447 6247 10553 6260
rect 4 5520 4196 5556
rect 4 5480 40 5520
rect 47 5500 4153 5513
rect 47 4940 60 5500
rect 80 5467 4120 5480
rect 80 4996 116 5467
rect 4107 4996 4120 5467
rect 80 4960 4120 4996
rect 4140 4940 4153 5500
rect 4160 4960 4196 5520
rect 6404 5520 10596 5556
rect 6404 5480 6440 5520
rect 6447 5500 10553 5513
rect 47 4927 4153 4940
rect 6447 4940 6460 5500
rect 6480 5467 10520 5480
rect 6480 4996 6516 5467
rect 10507 4996 10520 5467
rect 6480 4960 10520 4996
rect 10540 4940 10553 5500
rect 10560 4960 10596 5520
rect 6447 4930 10553 4940
rect 6447 4927 10080 4930
rect 4 3200 4196 3236
rect 4 3160 40 3200
rect 47 3180 4153 3193
rect 47 2620 60 3180
rect 80 3147 4120 3160
rect 80 2676 116 3147
rect 4107 2676 4120 3147
rect 80 2640 4120 2676
rect 4140 2620 4153 3180
rect 4160 2640 4196 3200
rect 6404 3200 10080 3236
rect 6404 3160 6440 3200
rect 6447 3180 10080 3193
rect 47 2607 4153 2620
rect 6447 2620 6460 3180
rect 6480 3147 10080 3160
rect 6480 2676 6516 3147
rect 6480 2640 10080 2676
rect 6447 2607 10080 2620
rect 4 2480 4196 2516
rect 4 2440 40 2480
rect 47 2460 4153 2473
rect 47 1900 60 2460
rect 80 2427 4120 2440
rect 80 1956 116 2427
rect 4107 1956 4120 2427
rect 80 1920 4120 1956
rect 4140 1900 4153 2460
rect 4160 1920 4196 2480
rect 6404 2480 10080 2516
rect 6404 2440 6440 2480
rect 6447 2460 10080 2473
rect 47 1887 4153 1900
rect 6447 1900 6460 2460
rect 6480 2427 10080 2440
rect 6480 1956 6516 2427
rect 6480 1920 10080 1956
rect 6447 1887 10080 1900
rect 4 1760 4196 1796
rect 4 1720 40 1760
rect 47 1740 4153 1753
rect 47 1180 60 1740
rect 80 1707 4120 1720
rect 80 1236 116 1707
rect 4107 1236 4120 1707
rect 80 1200 4120 1236
rect 4140 1180 4153 1740
rect 4160 1200 4196 1760
rect 6404 1760 10080 1796
rect 6404 1720 6440 1760
rect 6447 1740 10080 1753
rect 47 1167 4153 1180
rect 6447 1180 6460 1740
rect 6480 1707 10080 1720
rect 6480 1236 6516 1707
rect 6480 1200 10080 1236
rect 6447 1167 10080 1180
<< metal2 >>
rect 4240 12634 4440 12640
rect 4240 12606 4246 12634
rect 4274 12606 4406 12634
rect 4434 12606 4440 12634
rect 4240 12600 4440 12606
rect 4480 12634 4680 12640
rect 4480 12606 4486 12634
rect 4514 12606 4646 12634
rect 4674 12606 4680 12634
rect 4480 12600 4680 12606
rect 4720 12634 5080 12640
rect 4720 12606 4726 12634
rect 4754 12606 4886 12634
rect 4914 12606 5046 12634
rect 5074 12606 5080 12634
rect 4720 12600 5080 12606
rect 5120 12634 5480 12640
rect 5120 12606 5126 12634
rect 5154 12606 5286 12634
rect 5314 12606 5446 12634
rect 5474 12606 5480 12634
rect 5120 12600 5480 12606
rect 5520 12634 5880 12640
rect 5520 12606 5526 12634
rect 5554 12606 5686 12634
rect 5714 12606 5846 12634
rect 5874 12606 5880 12634
rect 5520 12600 5880 12606
rect 5920 12634 6120 12640
rect 5920 12606 5926 12634
rect 5954 12606 6086 12634
rect 6114 12606 6120 12634
rect 5920 12600 6120 12606
rect 6160 12634 6360 12640
rect 6160 12606 6166 12634
rect 6194 12606 6326 12634
rect 6354 12606 6360 12634
rect 6160 12600 6360 12606
rect 4240 12554 4440 12560
rect 4240 12526 4246 12554
rect 4274 12526 4406 12554
rect 4434 12526 4440 12554
rect 4240 12520 4440 12526
rect 4480 12554 4680 12560
rect 4480 12526 4486 12554
rect 4514 12526 4646 12554
rect 4674 12526 4680 12554
rect 4480 12520 4680 12526
rect 4720 12554 5080 12560
rect 4720 12526 4726 12554
rect 4754 12526 4886 12554
rect 4914 12526 5046 12554
rect 5074 12526 5080 12554
rect 4720 12520 5080 12526
rect 5120 12554 5480 12560
rect 5120 12526 5126 12554
rect 5154 12526 5286 12554
rect 5314 12526 5446 12554
rect 5474 12526 5480 12554
rect 5120 12520 5480 12526
rect 5520 12554 5880 12560
rect 5520 12526 5526 12554
rect 5554 12526 5686 12554
rect 5714 12526 5846 12554
rect 5874 12526 5880 12554
rect 5520 12520 5880 12526
rect 5920 12554 6120 12560
rect 5920 12526 5926 12554
rect 5954 12526 6086 12554
rect 6114 12526 6120 12554
rect 5920 12520 6120 12526
rect 6160 12554 6360 12560
rect 6160 12526 6166 12554
rect 6194 12526 6326 12554
rect 6354 12526 6360 12554
rect 6160 12520 6360 12526
rect 4240 12474 4440 12480
rect 4240 12446 4246 12474
rect 4274 12446 4406 12474
rect 4434 12446 4440 12474
rect 4240 12440 4440 12446
rect 4480 12474 4680 12480
rect 4480 12446 4486 12474
rect 4514 12446 4646 12474
rect 4674 12446 4680 12474
rect 4480 12440 4680 12446
rect 4720 12474 5080 12480
rect 4720 12446 4726 12474
rect 4754 12446 4886 12474
rect 4914 12446 5046 12474
rect 5074 12446 5080 12474
rect 4720 12440 5080 12446
rect 5120 12474 5480 12480
rect 5120 12446 5126 12474
rect 5154 12446 5286 12474
rect 5314 12446 5446 12474
rect 5474 12446 5480 12474
rect 5120 12440 5480 12446
rect 5520 12474 5880 12480
rect 5520 12446 5526 12474
rect 5554 12446 5686 12474
rect 5714 12446 5846 12474
rect 5874 12446 5880 12474
rect 5520 12440 5880 12446
rect 5920 12474 6120 12480
rect 5920 12446 5926 12474
rect 5954 12446 6086 12474
rect 6114 12446 6120 12474
rect 5920 12440 6120 12446
rect 6160 12474 6360 12480
rect 6160 12446 6166 12474
rect 6194 12446 6326 12474
rect 6354 12446 6360 12474
rect 6160 12440 6360 12446
rect 4240 12394 4440 12400
rect 4240 12366 4246 12394
rect 4274 12366 4406 12394
rect 4434 12366 4440 12394
rect 4240 12360 4440 12366
rect 4480 12394 4680 12400
rect 4480 12366 4486 12394
rect 4514 12366 4646 12394
rect 4674 12366 4680 12394
rect 4480 12360 4680 12366
rect 4720 12394 5080 12400
rect 4720 12366 4726 12394
rect 4754 12366 4886 12394
rect 4914 12366 5046 12394
rect 5074 12366 5080 12394
rect 4720 12360 5080 12366
rect 5120 12394 5480 12400
rect 5120 12366 5126 12394
rect 5154 12366 5286 12394
rect 5314 12366 5446 12394
rect 5474 12366 5480 12394
rect 5120 12360 5480 12366
rect 5520 12394 5880 12400
rect 5520 12366 5526 12394
rect 5554 12366 5686 12394
rect 5714 12366 5846 12394
rect 5874 12366 5880 12394
rect 5520 12360 5880 12366
rect 5920 12394 6120 12400
rect 5920 12366 5926 12394
rect 5954 12366 6086 12394
rect 6114 12366 6120 12394
rect 5920 12360 6120 12366
rect 6160 12394 6360 12400
rect 6160 12366 6166 12394
rect 6194 12366 6326 12394
rect 6354 12366 6360 12394
rect 6160 12360 6360 12366
rect 4240 12314 4440 12320
rect 4240 12286 4246 12314
rect 4274 12286 4406 12314
rect 4434 12286 4440 12314
rect 4240 12280 4440 12286
rect 4480 12314 4680 12320
rect 4480 12286 4486 12314
rect 4514 12286 4646 12314
rect 4674 12286 4680 12314
rect 4480 12280 4680 12286
rect 4720 12314 5080 12320
rect 4720 12286 4726 12314
rect 4754 12286 4886 12314
rect 4914 12286 5046 12314
rect 5074 12286 5080 12314
rect 4720 12280 5080 12286
rect 5120 12314 5480 12320
rect 5120 12286 5126 12314
rect 5154 12286 5286 12314
rect 5314 12286 5446 12314
rect 5474 12286 5480 12314
rect 5120 12280 5480 12286
rect 5520 12314 5880 12320
rect 5520 12286 5526 12314
rect 5554 12286 5686 12314
rect 5714 12286 5846 12314
rect 5874 12286 5880 12314
rect 5520 12280 5880 12286
rect 5920 12314 6120 12320
rect 5920 12286 5926 12314
rect 5954 12286 6086 12314
rect 6114 12286 6120 12314
rect 5920 12280 6120 12286
rect 6160 12314 6360 12320
rect 6160 12286 6166 12314
rect 6194 12286 6326 12314
rect 6354 12286 6360 12314
rect 6160 12280 6360 12286
rect 4240 12234 4440 12240
rect 4240 12206 4246 12234
rect 4274 12206 4406 12234
rect 4434 12206 4440 12234
rect 4240 12200 4440 12206
rect 4480 12234 4680 12240
rect 4480 12206 4486 12234
rect 4514 12206 4646 12234
rect 4674 12206 4680 12234
rect 4480 12200 4680 12206
rect 4720 12234 5080 12240
rect 4720 12206 4726 12234
rect 4754 12206 4886 12234
rect 4914 12206 5046 12234
rect 5074 12206 5080 12234
rect 4720 12200 5080 12206
rect 5120 12234 5480 12240
rect 5120 12206 5126 12234
rect 5154 12206 5286 12234
rect 5314 12206 5446 12234
rect 5474 12206 5480 12234
rect 5120 12200 5480 12206
rect 5520 12234 5880 12240
rect 5520 12206 5526 12234
rect 5554 12206 5686 12234
rect 5714 12206 5846 12234
rect 5874 12206 5880 12234
rect 5520 12200 5880 12206
rect 5920 12234 6120 12240
rect 5920 12206 5926 12234
rect 5954 12206 6086 12234
rect 6114 12206 6120 12234
rect 5920 12200 6120 12206
rect 6160 12234 6360 12240
rect 6160 12206 6166 12234
rect 6194 12206 6326 12234
rect 6354 12206 6360 12234
rect 6160 12200 6360 12206
rect 4240 12154 4440 12160
rect 4240 12126 4246 12154
rect 4274 12126 4406 12154
rect 4434 12126 4440 12154
rect 4240 12120 4440 12126
rect 4480 12154 4680 12160
rect 4480 12126 4486 12154
rect 4514 12126 4646 12154
rect 4674 12126 4680 12154
rect 4480 12120 4680 12126
rect 4720 12154 5080 12160
rect 4720 12126 4726 12154
rect 4754 12126 4886 12154
rect 4914 12126 5046 12154
rect 5074 12126 5080 12154
rect 4720 12120 5080 12126
rect 5120 12154 5480 12160
rect 5120 12126 5126 12154
rect 5154 12126 5286 12154
rect 5314 12126 5446 12154
rect 5474 12126 5480 12154
rect 5120 12120 5480 12126
rect 5520 12154 5880 12160
rect 5520 12126 5526 12154
rect 5554 12126 5686 12154
rect 5714 12126 5846 12154
rect 5874 12126 5880 12154
rect 5520 12120 5880 12126
rect 5920 12154 6120 12160
rect 5920 12126 5926 12154
rect 5954 12126 6086 12154
rect 6114 12126 6120 12154
rect 5920 12120 6120 12126
rect 6160 12154 6360 12160
rect 6160 12126 6166 12154
rect 6194 12126 6326 12154
rect 6354 12126 6360 12154
rect 6160 12120 6360 12126
rect 4200 12074 6400 12080
rect 4200 12046 4486 12074
rect 4514 12046 4646 12074
rect 4674 12046 6400 12074
rect 4200 12040 6400 12046
rect 4200 11994 6400 12000
rect 4200 11966 4566 11994
rect 4594 11966 6400 11994
rect 4200 11960 6400 11966
rect 4200 11914 6400 11920
rect 4200 11886 4486 11914
rect 4514 11886 4646 11914
rect 4674 11886 6400 11914
rect 4200 11880 6400 11886
rect 4240 11834 4440 11840
rect 4240 11806 4246 11834
rect 4274 11806 4406 11834
rect 4434 11806 4440 11834
rect 4240 11800 4440 11806
rect 4480 11834 4680 11840
rect 4480 11806 4486 11834
rect 4514 11806 4646 11834
rect 4674 11806 4680 11834
rect 4480 11800 4680 11806
rect 4720 11834 5080 11840
rect 4720 11806 4726 11834
rect 4754 11806 4886 11834
rect 4914 11806 5046 11834
rect 5074 11806 5080 11834
rect 4720 11800 5080 11806
rect 5120 11834 5480 11840
rect 5120 11806 5126 11834
rect 5154 11806 5286 11834
rect 5314 11806 5446 11834
rect 5474 11806 5480 11834
rect 5120 11800 5480 11806
rect 5520 11834 5880 11840
rect 5520 11806 5526 11834
rect 5554 11806 5686 11834
rect 5714 11806 5846 11834
rect 5874 11806 5880 11834
rect 5520 11800 5880 11806
rect 5920 11834 6120 11840
rect 5920 11806 5926 11834
rect 5954 11806 6086 11834
rect 6114 11806 6120 11834
rect 5920 11800 6120 11806
rect 6160 11834 6360 11840
rect 6160 11806 6166 11834
rect 6194 11806 6326 11834
rect 6354 11806 6360 11834
rect 6160 11800 6360 11806
rect 4240 11754 4440 11760
rect 4240 11726 4246 11754
rect 4274 11726 4406 11754
rect 4434 11726 4440 11754
rect 4240 11720 4440 11726
rect 4480 11754 4680 11760
rect 4480 11726 4486 11754
rect 4514 11726 4646 11754
rect 4674 11726 4680 11754
rect 4480 11720 4680 11726
rect 4720 11754 5080 11760
rect 4720 11726 4726 11754
rect 4754 11726 4886 11754
rect 4914 11726 5046 11754
rect 5074 11726 5080 11754
rect 4720 11720 5080 11726
rect 5120 11754 5480 11760
rect 5120 11726 5126 11754
rect 5154 11726 5286 11754
rect 5314 11726 5446 11754
rect 5474 11726 5480 11754
rect 5120 11720 5480 11726
rect 5520 11754 5880 11760
rect 5520 11726 5526 11754
rect 5554 11726 5686 11754
rect 5714 11726 5846 11754
rect 5874 11726 5880 11754
rect 5520 11720 5880 11726
rect 5920 11754 6120 11760
rect 5920 11726 5926 11754
rect 5954 11726 6086 11754
rect 6114 11726 6120 11754
rect 5920 11720 6120 11726
rect 6160 11754 6360 11760
rect 6160 11726 6166 11754
rect 6194 11726 6326 11754
rect 6354 11726 6360 11754
rect 6160 11720 6360 11726
rect 4240 11674 4440 11680
rect 4240 11646 4246 11674
rect 4274 11646 4406 11674
rect 4434 11646 4440 11674
rect 4240 11640 4440 11646
rect 4480 11674 4680 11680
rect 4480 11646 4486 11674
rect 4514 11646 4646 11674
rect 4674 11646 4680 11674
rect 4480 11640 4680 11646
rect 4720 11674 5080 11680
rect 4720 11646 4726 11674
rect 4754 11646 4886 11674
rect 4914 11646 5046 11674
rect 5074 11646 5080 11674
rect 4720 11640 5080 11646
rect 5120 11674 5480 11680
rect 5120 11646 5126 11674
rect 5154 11646 5286 11674
rect 5314 11646 5446 11674
rect 5474 11646 5480 11674
rect 5120 11640 5480 11646
rect 5520 11674 5880 11680
rect 5520 11646 5526 11674
rect 5554 11646 5686 11674
rect 5714 11646 5846 11674
rect 5874 11646 5880 11674
rect 5520 11640 5880 11646
rect 5920 11674 6120 11680
rect 5920 11646 5926 11674
rect 5954 11646 6086 11674
rect 6114 11646 6120 11674
rect 5920 11640 6120 11646
rect 6160 11674 6360 11680
rect 6160 11646 6166 11674
rect 6194 11646 6326 11674
rect 6354 11646 6360 11674
rect 6160 11640 6360 11646
rect 4240 11594 4440 11600
rect 4240 11566 4246 11594
rect 4274 11566 4406 11594
rect 4434 11566 4440 11594
rect 4240 11560 4440 11566
rect 4480 11594 4680 11600
rect 4480 11566 4486 11594
rect 4514 11566 4646 11594
rect 4674 11566 4680 11594
rect 4480 11560 4680 11566
rect 4720 11594 5080 11600
rect 4720 11566 4726 11594
rect 4754 11566 4886 11594
rect 4914 11566 5046 11594
rect 5074 11566 5080 11594
rect 4720 11560 5080 11566
rect 5120 11594 5480 11600
rect 5120 11566 5126 11594
rect 5154 11566 5286 11594
rect 5314 11566 5446 11594
rect 5474 11566 5480 11594
rect 5120 11560 5480 11566
rect 5520 11594 5880 11600
rect 5520 11566 5526 11594
rect 5554 11566 5686 11594
rect 5714 11566 5846 11594
rect 5874 11566 5880 11594
rect 5520 11560 5880 11566
rect 5920 11594 6120 11600
rect 5920 11566 5926 11594
rect 5954 11566 6086 11594
rect 6114 11566 6120 11594
rect 5920 11560 6120 11566
rect 6160 11594 6360 11600
rect 6160 11566 6166 11594
rect 6194 11566 6326 11594
rect 6354 11566 6360 11594
rect 6160 11560 6360 11566
rect 4240 11514 4440 11520
rect 4240 11486 4246 11514
rect 4274 11486 4406 11514
rect 4434 11486 4440 11514
rect 4240 11480 4440 11486
rect 4480 11514 4680 11520
rect 4480 11486 4486 11514
rect 4514 11486 4646 11514
rect 4674 11486 4680 11514
rect 4480 11480 4680 11486
rect 4720 11514 5080 11520
rect 4720 11486 4726 11514
rect 4754 11486 4886 11514
rect 4914 11486 5046 11514
rect 5074 11486 5080 11514
rect 4720 11480 5080 11486
rect 5120 11514 5480 11520
rect 5120 11486 5126 11514
rect 5154 11486 5286 11514
rect 5314 11486 5446 11514
rect 5474 11486 5480 11514
rect 5120 11480 5480 11486
rect 5520 11514 5880 11520
rect 5520 11486 5526 11514
rect 5554 11486 5686 11514
rect 5714 11486 5846 11514
rect 5874 11486 5880 11514
rect 5520 11480 5880 11486
rect 5920 11514 6120 11520
rect 5920 11486 5926 11514
rect 5954 11486 6086 11514
rect 6114 11486 6120 11514
rect 5920 11480 6120 11486
rect 6160 11514 6360 11520
rect 6160 11486 6166 11514
rect 6194 11486 6326 11514
rect 6354 11486 6360 11514
rect 6160 11480 6360 11486
rect 4240 11434 4440 11440
rect 4240 11406 4246 11434
rect 4274 11406 4406 11434
rect 4434 11406 4440 11434
rect 4240 11400 4440 11406
rect 4480 11434 4680 11440
rect 4480 11406 4486 11434
rect 4514 11406 4646 11434
rect 4674 11406 4680 11434
rect 4480 11400 4680 11406
rect 4720 11434 5080 11440
rect 4720 11406 4726 11434
rect 4754 11406 4886 11434
rect 4914 11406 5046 11434
rect 5074 11406 5080 11434
rect 4720 11400 5080 11406
rect 5120 11434 5480 11440
rect 5120 11406 5126 11434
rect 5154 11406 5286 11434
rect 5314 11406 5446 11434
rect 5474 11406 5480 11434
rect 5120 11400 5480 11406
rect 5520 11434 5880 11440
rect 5520 11406 5526 11434
rect 5554 11406 5686 11434
rect 5714 11406 5846 11434
rect 5874 11406 5880 11434
rect 5520 11400 5880 11406
rect 5920 11434 6120 11440
rect 5920 11406 5926 11434
rect 5954 11406 6086 11434
rect 6114 11406 6120 11434
rect 5920 11400 6120 11406
rect 6160 11434 6360 11440
rect 6160 11406 6166 11434
rect 6194 11406 6326 11434
rect 6354 11406 6360 11434
rect 6160 11400 6360 11406
rect 4200 11314 6400 11320
rect 4200 11286 5526 11314
rect 5554 11286 5686 11314
rect 5714 11286 6400 11314
rect 4200 11280 6400 11286
rect 4200 11234 6400 11240
rect 4200 11206 5606 11234
rect 5634 11206 6400 11234
rect 4200 11200 6400 11206
rect 4200 11154 6400 11160
rect 4200 11126 5046 11154
rect 5074 11126 5526 11154
rect 5554 11126 5686 11154
rect 5714 11126 6400 11154
rect 4200 11120 6400 11126
rect 4200 11074 6400 11080
rect 4200 11046 5126 11074
rect 5154 11046 5286 11074
rect 5314 11046 5446 11074
rect 5474 11046 6400 11074
rect 4200 11040 6400 11046
rect 4200 10994 6400 11000
rect 4200 10966 5046 10994
rect 5074 10966 5526 10994
rect 5554 10966 6400 10994
rect 4200 10960 6400 10966
rect 4240 10874 4440 10880
rect 4240 10846 4246 10874
rect 4274 10846 4406 10874
rect 4434 10846 4440 10874
rect 4240 10840 4440 10846
rect 4480 10874 4680 10880
rect 4480 10846 4486 10874
rect 4514 10846 4646 10874
rect 4674 10846 4680 10874
rect 4480 10840 4680 10846
rect 4720 10874 5080 10880
rect 4720 10846 4726 10874
rect 4754 10846 4886 10874
rect 4914 10846 5046 10874
rect 5074 10846 5080 10874
rect 4720 10840 5080 10846
rect 5120 10874 5480 10880
rect 5120 10846 5126 10874
rect 5154 10846 5286 10874
rect 5314 10846 5446 10874
rect 5474 10846 5480 10874
rect 5120 10840 5480 10846
rect 5520 10874 5880 10880
rect 5520 10846 5526 10874
rect 5554 10846 5686 10874
rect 5714 10846 5846 10874
rect 5874 10846 5880 10874
rect 5520 10840 5880 10846
rect 5920 10874 6120 10880
rect 5920 10846 5926 10874
rect 5954 10846 6086 10874
rect 6114 10846 6120 10874
rect 5920 10840 6120 10846
rect 6160 10874 6360 10880
rect 6160 10846 6166 10874
rect 6194 10846 6326 10874
rect 6354 10846 6360 10874
rect 6160 10840 6360 10846
rect 4240 10794 4440 10800
rect 4240 10766 4246 10794
rect 4274 10766 4406 10794
rect 4434 10766 4440 10794
rect 4240 10760 4440 10766
rect 4480 10794 4680 10800
rect 4480 10766 4486 10794
rect 4514 10766 4646 10794
rect 4674 10766 4680 10794
rect 4480 10760 4680 10766
rect 4720 10794 5080 10800
rect 4720 10766 4726 10794
rect 4754 10766 4886 10794
rect 4914 10766 5046 10794
rect 5074 10766 5080 10794
rect 4720 10760 5080 10766
rect 5120 10794 5480 10800
rect 5120 10766 5126 10794
rect 5154 10766 5286 10794
rect 5314 10766 5446 10794
rect 5474 10766 5480 10794
rect 5120 10760 5480 10766
rect 5520 10794 5880 10800
rect 5520 10766 5526 10794
rect 5554 10766 5686 10794
rect 5714 10766 5846 10794
rect 5874 10766 5880 10794
rect 5520 10760 5880 10766
rect 5920 10794 6120 10800
rect 5920 10766 5926 10794
rect 5954 10766 6086 10794
rect 6114 10766 6120 10794
rect 5920 10760 6120 10766
rect 6160 10794 6360 10800
rect 6160 10766 6166 10794
rect 6194 10766 6326 10794
rect 6354 10766 6360 10794
rect 6160 10760 6360 10766
rect 4240 10714 4440 10720
rect 4240 10686 4246 10714
rect 4274 10686 4406 10714
rect 4434 10686 4440 10714
rect 4240 10680 4440 10686
rect 4480 10714 4680 10720
rect 4480 10686 4486 10714
rect 4514 10686 4646 10714
rect 4674 10686 4680 10714
rect 4480 10680 4680 10686
rect 4720 10714 5080 10720
rect 4720 10686 4726 10714
rect 4754 10686 4886 10714
rect 4914 10686 5046 10714
rect 5074 10686 5080 10714
rect 4720 10680 5080 10686
rect 5120 10714 5480 10720
rect 5120 10686 5126 10714
rect 5154 10686 5286 10714
rect 5314 10686 5446 10714
rect 5474 10686 5480 10714
rect 5120 10680 5480 10686
rect 5520 10714 5880 10720
rect 5520 10686 5526 10714
rect 5554 10686 5686 10714
rect 5714 10686 5846 10714
rect 5874 10686 5880 10714
rect 5520 10680 5880 10686
rect 5920 10714 6120 10720
rect 5920 10686 5926 10714
rect 5954 10686 6086 10714
rect 6114 10686 6120 10714
rect 5920 10680 6120 10686
rect 6160 10714 6360 10720
rect 6160 10686 6166 10714
rect 6194 10686 6326 10714
rect 6354 10686 6360 10714
rect 6160 10680 6360 10686
rect 4240 10634 4440 10640
rect 4240 10606 4246 10634
rect 4274 10606 4406 10634
rect 4434 10606 4440 10634
rect 4240 10600 4440 10606
rect 4480 10634 4680 10640
rect 4480 10606 4486 10634
rect 4514 10606 4646 10634
rect 4674 10606 4680 10634
rect 4480 10600 4680 10606
rect 4720 10634 5080 10640
rect 4720 10606 4726 10634
rect 4754 10606 4886 10634
rect 4914 10606 5046 10634
rect 5074 10606 5080 10634
rect 4720 10600 5080 10606
rect 5120 10634 5480 10640
rect 5120 10606 5126 10634
rect 5154 10606 5286 10634
rect 5314 10606 5446 10634
rect 5474 10606 5480 10634
rect 5120 10600 5480 10606
rect 5520 10634 5880 10640
rect 5520 10606 5526 10634
rect 5554 10606 5686 10634
rect 5714 10606 5846 10634
rect 5874 10606 5880 10634
rect 5520 10600 5880 10606
rect 5920 10634 6120 10640
rect 5920 10606 5926 10634
rect 5954 10606 6086 10634
rect 6114 10606 6120 10634
rect 5920 10600 6120 10606
rect 6160 10634 6360 10640
rect 6160 10606 6166 10634
rect 6194 10606 6326 10634
rect 6354 10606 6360 10634
rect 6160 10600 6360 10606
rect 4240 10554 4440 10560
rect 4240 10526 4246 10554
rect 4274 10526 4406 10554
rect 4434 10526 4440 10554
rect 4240 10520 4440 10526
rect 4480 10554 4680 10560
rect 4480 10526 4486 10554
rect 4514 10526 4646 10554
rect 4674 10526 4680 10554
rect 4480 10520 4680 10526
rect 4720 10554 5080 10560
rect 4720 10526 4726 10554
rect 4754 10526 4886 10554
rect 4914 10526 5046 10554
rect 5074 10526 5080 10554
rect 4720 10520 5080 10526
rect 5120 10554 5480 10560
rect 5120 10526 5126 10554
rect 5154 10526 5286 10554
rect 5314 10526 5446 10554
rect 5474 10526 5480 10554
rect 5120 10520 5480 10526
rect 5520 10554 5880 10560
rect 5520 10526 5526 10554
rect 5554 10526 5686 10554
rect 5714 10526 5846 10554
rect 5874 10526 5880 10554
rect 5520 10520 5880 10526
rect 5920 10554 6120 10560
rect 5920 10526 5926 10554
rect 5954 10526 6086 10554
rect 6114 10526 6120 10554
rect 5920 10520 6120 10526
rect 6160 10554 6360 10560
rect 6160 10526 6166 10554
rect 6194 10526 6326 10554
rect 6354 10526 6360 10554
rect 6160 10520 6360 10526
rect 4240 10474 4440 10480
rect 4240 10446 4246 10474
rect 4274 10446 4406 10474
rect 4434 10446 4440 10474
rect 4240 10440 4440 10446
rect 4480 10474 4680 10480
rect 4480 10446 4486 10474
rect 4514 10446 4646 10474
rect 4674 10446 4680 10474
rect 4480 10440 4680 10446
rect 4720 10474 5080 10480
rect 4720 10446 4726 10474
rect 4754 10446 4886 10474
rect 4914 10446 5046 10474
rect 5074 10446 5080 10474
rect 4720 10440 5080 10446
rect 5120 10474 5480 10480
rect 5120 10446 5126 10474
rect 5154 10446 5286 10474
rect 5314 10446 5446 10474
rect 5474 10446 5480 10474
rect 5120 10440 5480 10446
rect 5520 10474 5880 10480
rect 5520 10446 5526 10474
rect 5554 10446 5686 10474
rect 5714 10446 5846 10474
rect 5874 10446 5880 10474
rect 5520 10440 5880 10446
rect 5920 10474 6120 10480
rect 5920 10446 5926 10474
rect 5954 10446 6086 10474
rect 6114 10446 6120 10474
rect 5920 10440 6120 10446
rect 6160 10474 6360 10480
rect 6160 10446 6166 10474
rect 6194 10446 6326 10474
rect 6354 10446 6360 10474
rect 6160 10440 6360 10446
rect 4240 10394 4440 10400
rect 4240 10366 4246 10394
rect 4274 10366 4406 10394
rect 4434 10366 4440 10394
rect 4240 10360 4440 10366
rect 4480 10394 4680 10400
rect 4480 10366 4486 10394
rect 4514 10366 4646 10394
rect 4674 10366 4680 10394
rect 4480 10360 4680 10366
rect 4720 10394 5080 10400
rect 4720 10366 4726 10394
rect 4754 10366 4886 10394
rect 4914 10366 5046 10394
rect 5074 10366 5080 10394
rect 4720 10360 5080 10366
rect 5120 10394 5480 10400
rect 5120 10366 5126 10394
rect 5154 10366 5286 10394
rect 5314 10366 5446 10394
rect 5474 10366 5480 10394
rect 5120 10360 5480 10366
rect 5520 10394 5880 10400
rect 5520 10366 5526 10394
rect 5554 10366 5686 10394
rect 5714 10366 5846 10394
rect 5874 10366 5880 10394
rect 5520 10360 5880 10366
rect 5920 10394 6120 10400
rect 5920 10366 5926 10394
rect 5954 10366 6086 10394
rect 6114 10366 6120 10394
rect 5920 10360 6120 10366
rect 6160 10394 6360 10400
rect 6160 10366 6166 10394
rect 6194 10366 6326 10394
rect 6354 10366 6360 10394
rect 6160 10360 6360 10366
rect 4240 10314 4440 10320
rect 4240 10286 4246 10314
rect 4274 10286 4406 10314
rect 4434 10286 4440 10314
rect 4240 10280 4440 10286
rect 4480 10314 4680 10320
rect 4480 10286 4486 10314
rect 4514 10286 4646 10314
rect 4674 10286 4680 10314
rect 4480 10280 4680 10286
rect 4720 10314 5080 10320
rect 4720 10286 4726 10314
rect 4754 10286 4886 10314
rect 4914 10286 5046 10314
rect 5074 10286 5080 10314
rect 4720 10280 5080 10286
rect 5120 10314 5480 10320
rect 5120 10286 5126 10314
rect 5154 10286 5286 10314
rect 5314 10286 5446 10314
rect 5474 10286 5480 10314
rect 5120 10280 5480 10286
rect 5520 10314 5880 10320
rect 5520 10286 5526 10314
rect 5554 10286 5686 10314
rect 5714 10286 5846 10314
rect 5874 10286 5880 10314
rect 5520 10280 5880 10286
rect 5920 10314 6120 10320
rect 5920 10286 5926 10314
rect 5954 10286 6086 10314
rect 6114 10286 6120 10314
rect 5920 10280 6120 10286
rect 6160 10314 6360 10320
rect 6160 10286 6166 10314
rect 6194 10286 6326 10314
rect 6354 10286 6360 10314
rect 6160 10280 6360 10286
rect 4240 10234 4440 10240
rect 4240 10206 4246 10234
rect 4274 10206 4406 10234
rect 4434 10206 4440 10234
rect 4240 10200 4440 10206
rect 4480 10234 4680 10240
rect 4480 10206 4486 10234
rect 4514 10206 4646 10234
rect 4674 10206 4680 10234
rect 4480 10200 4680 10206
rect 4720 10234 5080 10240
rect 4720 10206 4726 10234
rect 4754 10206 4886 10234
rect 4914 10206 5046 10234
rect 5074 10206 5080 10234
rect 4720 10200 5080 10206
rect 5120 10234 5480 10240
rect 5120 10206 5126 10234
rect 5154 10206 5286 10234
rect 5314 10206 5446 10234
rect 5474 10206 5480 10234
rect 5120 10200 5480 10206
rect 5520 10234 5880 10240
rect 5520 10206 5526 10234
rect 5554 10206 5686 10234
rect 5714 10206 5846 10234
rect 5874 10206 5880 10234
rect 5520 10200 5880 10206
rect 5920 10234 6120 10240
rect 5920 10206 5926 10234
rect 5954 10206 6086 10234
rect 6114 10206 6120 10234
rect 5920 10200 6120 10206
rect 6160 10234 6360 10240
rect 6160 10206 6166 10234
rect 6194 10206 6326 10234
rect 6354 10206 6360 10234
rect 6160 10200 6360 10206
rect 4240 10154 4440 10160
rect 4240 10126 4246 10154
rect 4274 10126 4406 10154
rect 4434 10126 4440 10154
rect 4240 10120 4440 10126
rect 4480 10154 4680 10160
rect 4480 10126 4486 10154
rect 4514 10126 4646 10154
rect 4674 10126 4680 10154
rect 4480 10120 4680 10126
rect 4720 10154 5080 10160
rect 4720 10126 4726 10154
rect 4754 10126 4886 10154
rect 4914 10126 5046 10154
rect 5074 10126 5080 10154
rect 4720 10120 5080 10126
rect 5120 10154 5480 10160
rect 5120 10126 5126 10154
rect 5154 10126 5286 10154
rect 5314 10126 5446 10154
rect 5474 10126 5480 10154
rect 5120 10120 5480 10126
rect 5520 10154 5880 10160
rect 5520 10126 5526 10154
rect 5554 10126 5686 10154
rect 5714 10126 5846 10154
rect 5874 10126 5880 10154
rect 5520 10120 5880 10126
rect 5920 10154 6120 10160
rect 5920 10126 5926 10154
rect 5954 10126 6086 10154
rect 6114 10126 6120 10154
rect 5920 10120 6120 10126
rect 6160 10154 6360 10160
rect 6160 10126 6166 10154
rect 6194 10126 6326 10154
rect 6354 10126 6360 10154
rect 6160 10120 6360 10126
rect 4240 10074 4440 10080
rect 4240 10046 4246 10074
rect 4274 10046 4406 10074
rect 4434 10046 4440 10074
rect 4240 10040 4440 10046
rect 4480 10074 4680 10080
rect 4480 10046 4486 10074
rect 4514 10046 4646 10074
rect 4674 10046 4680 10074
rect 4480 10040 4680 10046
rect 4720 10074 5080 10080
rect 4720 10046 4726 10074
rect 4754 10046 4886 10074
rect 4914 10046 5046 10074
rect 5074 10046 5080 10074
rect 4720 10040 5080 10046
rect 5120 10074 5480 10080
rect 5120 10046 5126 10074
rect 5154 10046 5286 10074
rect 5314 10046 5446 10074
rect 5474 10046 5480 10074
rect 5120 10040 5480 10046
rect 5520 10074 5880 10080
rect 5520 10046 5526 10074
rect 5554 10046 5686 10074
rect 5714 10046 5846 10074
rect 5874 10046 5880 10074
rect 5520 10040 5880 10046
rect 5920 10074 6120 10080
rect 5920 10046 5926 10074
rect 5954 10046 6086 10074
rect 6114 10046 6120 10074
rect 5920 10040 6120 10046
rect 6160 10074 6360 10080
rect 6160 10046 6166 10074
rect 6194 10046 6326 10074
rect 6354 10046 6360 10074
rect 6160 10040 6360 10046
rect 4240 9994 4440 10000
rect 4240 9966 4246 9994
rect 4274 9966 4406 9994
rect 4434 9966 4440 9994
rect 4240 9960 4440 9966
rect 4480 9994 4680 10000
rect 4480 9966 4486 9994
rect 4514 9966 4646 9994
rect 4674 9966 4680 9994
rect 4480 9960 4680 9966
rect 4720 9994 5080 10000
rect 4720 9966 4726 9994
rect 4754 9966 4886 9994
rect 4914 9966 5046 9994
rect 5074 9966 5080 9994
rect 4720 9960 5080 9966
rect 5120 9994 5480 10000
rect 5120 9966 5126 9994
rect 5154 9966 5286 9994
rect 5314 9966 5446 9994
rect 5474 9966 5480 9994
rect 5120 9960 5480 9966
rect 5520 9994 5880 10000
rect 5520 9966 5526 9994
rect 5554 9966 5686 9994
rect 5714 9966 5846 9994
rect 5874 9966 5880 9994
rect 5520 9960 5880 9966
rect 5920 9994 6120 10000
rect 5920 9966 5926 9994
rect 5954 9966 6086 9994
rect 6114 9966 6120 9994
rect 5920 9960 6120 9966
rect 6160 9994 6360 10000
rect 6160 9966 6166 9994
rect 6194 9966 6326 9994
rect 6354 9966 6360 9994
rect 6160 9960 6360 9966
rect 4240 9914 4440 9920
rect 4240 9886 4246 9914
rect 4274 9886 4406 9914
rect 4434 9886 4440 9914
rect 4240 9880 4440 9886
rect 4480 9914 4680 9920
rect 4480 9886 4486 9914
rect 4514 9886 4646 9914
rect 4674 9886 4680 9914
rect 4480 9880 4680 9886
rect 4720 9914 5080 9920
rect 4720 9886 4726 9914
rect 4754 9886 4886 9914
rect 4914 9886 5046 9914
rect 5074 9886 5080 9914
rect 4720 9880 5080 9886
rect 5120 9914 5480 9920
rect 5120 9886 5126 9914
rect 5154 9886 5286 9914
rect 5314 9886 5446 9914
rect 5474 9886 5480 9914
rect 5120 9880 5480 9886
rect 5520 9914 5880 9920
rect 5520 9886 5526 9914
rect 5554 9886 5686 9914
rect 5714 9886 5846 9914
rect 5874 9886 5880 9914
rect 5520 9880 5880 9886
rect 5920 9914 6120 9920
rect 5920 9886 5926 9914
rect 5954 9886 6086 9914
rect 6114 9886 6120 9914
rect 5920 9880 6120 9886
rect 6160 9914 6360 9920
rect 6160 9886 6166 9914
rect 6194 9886 6326 9914
rect 6354 9886 6360 9914
rect 6160 9880 6360 9886
rect 4240 9834 4440 9840
rect 4240 9806 4246 9834
rect 4274 9806 4406 9834
rect 4434 9806 4440 9834
rect 4240 9800 4440 9806
rect 4480 9834 4680 9840
rect 4480 9806 4486 9834
rect 4514 9806 4646 9834
rect 4674 9806 4680 9834
rect 4480 9800 4680 9806
rect 4720 9834 5080 9840
rect 4720 9806 4726 9834
rect 4754 9806 4886 9834
rect 4914 9806 5046 9834
rect 5074 9806 5080 9834
rect 4720 9800 5080 9806
rect 5120 9834 5480 9840
rect 5120 9806 5126 9834
rect 5154 9806 5286 9834
rect 5314 9806 5446 9834
rect 5474 9806 5480 9834
rect 5120 9800 5480 9806
rect 5520 9834 5880 9840
rect 5520 9806 5526 9834
rect 5554 9806 5686 9834
rect 5714 9806 5846 9834
rect 5874 9806 5880 9834
rect 5520 9800 5880 9806
rect 5920 9834 6120 9840
rect 5920 9806 5926 9834
rect 5954 9806 6086 9834
rect 6114 9806 6120 9834
rect 5920 9800 6120 9806
rect 6160 9834 6360 9840
rect 6160 9806 6166 9834
rect 6194 9806 6326 9834
rect 6354 9806 6360 9834
rect 6160 9800 6360 9806
rect 4240 9754 4440 9760
rect 4240 9726 4246 9754
rect 4274 9726 4406 9754
rect 4434 9726 4440 9754
rect 4240 9720 4440 9726
rect 4480 9754 4680 9760
rect 4480 9726 4486 9754
rect 4514 9726 4646 9754
rect 4674 9726 4680 9754
rect 4480 9720 4680 9726
rect 4720 9754 5080 9760
rect 4720 9726 4726 9754
rect 4754 9726 4886 9754
rect 4914 9726 5046 9754
rect 5074 9726 5080 9754
rect 4720 9720 5080 9726
rect 5120 9754 5480 9760
rect 5120 9726 5126 9754
rect 5154 9726 5286 9754
rect 5314 9726 5446 9754
rect 5474 9726 5480 9754
rect 5120 9720 5480 9726
rect 5520 9754 5880 9760
rect 5520 9726 5526 9754
rect 5554 9726 5686 9754
rect 5714 9726 5846 9754
rect 5874 9726 5880 9754
rect 5520 9720 5880 9726
rect 5920 9754 6120 9760
rect 5920 9726 5926 9754
rect 5954 9726 6086 9754
rect 6114 9726 6120 9754
rect 5920 9720 6120 9726
rect 6160 9754 6360 9760
rect 6160 9726 6166 9754
rect 6194 9726 6326 9754
rect 6354 9726 6360 9754
rect 6160 9720 6360 9726
rect 4240 9634 6360 9640
rect 4240 9606 4486 9634
rect 4514 9606 4646 9634
rect 4674 9606 6360 9634
rect 4240 9600 6360 9606
rect 4200 9554 6400 9560
rect 4200 9526 4566 9554
rect 4594 9526 6400 9554
rect 4200 9520 6400 9526
rect 4240 9474 6360 9480
rect 4240 9446 4486 9474
rect 4514 9446 4646 9474
rect 4674 9446 6360 9474
rect 4240 9440 6360 9446
rect 4240 9354 4440 9360
rect 4240 9326 4246 9354
rect 4274 9326 4406 9354
rect 4434 9326 4440 9354
rect 4240 9320 4440 9326
rect 4480 9354 4680 9360
rect 4480 9326 4486 9354
rect 4514 9326 4646 9354
rect 4674 9326 4680 9354
rect 4480 9320 4680 9326
rect 4720 9354 5080 9360
rect 4720 9326 4726 9354
rect 4754 9326 4886 9354
rect 4914 9326 5046 9354
rect 5074 9326 5080 9354
rect 4720 9320 5080 9326
rect 5120 9354 5480 9360
rect 5120 9326 5126 9354
rect 5154 9326 5286 9354
rect 5314 9326 5446 9354
rect 5474 9326 5480 9354
rect 5120 9320 5480 9326
rect 5520 9354 5880 9360
rect 5520 9326 5526 9354
rect 5554 9326 5686 9354
rect 5714 9326 5846 9354
rect 5874 9326 5880 9354
rect 5520 9320 5880 9326
rect 5920 9354 6120 9360
rect 5920 9326 5926 9354
rect 5954 9326 6086 9354
rect 6114 9326 6120 9354
rect 5920 9320 6120 9326
rect 6160 9354 6360 9360
rect 6160 9326 6166 9354
rect 6194 9326 6326 9354
rect 6354 9326 6360 9354
rect 6160 9320 6360 9326
rect 4240 9274 4440 9280
rect 4240 9246 4246 9274
rect 4274 9246 4406 9274
rect 4434 9246 4440 9274
rect 4240 9240 4440 9246
rect 4480 9274 4680 9280
rect 4480 9246 4486 9274
rect 4514 9246 4646 9274
rect 4674 9246 4680 9274
rect 4480 9240 4680 9246
rect 4720 9274 5080 9280
rect 4720 9246 4726 9274
rect 4754 9246 4886 9274
rect 4914 9246 5046 9274
rect 5074 9246 5080 9274
rect 4720 9240 5080 9246
rect 5120 9274 5480 9280
rect 5120 9246 5126 9274
rect 5154 9246 5286 9274
rect 5314 9246 5446 9274
rect 5474 9246 5480 9274
rect 5120 9240 5480 9246
rect 5520 9274 5880 9280
rect 5520 9246 5526 9274
rect 5554 9246 5686 9274
rect 5714 9246 5846 9274
rect 5874 9246 5880 9274
rect 5520 9240 5880 9246
rect 5920 9274 6120 9280
rect 5920 9246 5926 9274
rect 5954 9246 6086 9274
rect 6114 9246 6120 9274
rect 5920 9240 6120 9246
rect 6160 9274 6360 9280
rect 6160 9246 6166 9274
rect 6194 9246 6326 9274
rect 6354 9246 6360 9274
rect 6160 9240 6360 9246
rect 4240 9194 4440 9200
rect 4240 9166 4246 9194
rect 4274 9166 4406 9194
rect 4434 9166 4440 9194
rect 4240 9160 4440 9166
rect 4480 9194 4680 9200
rect 4480 9166 4486 9194
rect 4514 9166 4646 9194
rect 4674 9166 4680 9194
rect 4480 9160 4680 9166
rect 4720 9194 5080 9200
rect 4720 9166 4726 9194
rect 4754 9166 4886 9194
rect 4914 9166 5046 9194
rect 5074 9166 5080 9194
rect 4720 9160 5080 9166
rect 5120 9194 5480 9200
rect 5120 9166 5126 9194
rect 5154 9166 5286 9194
rect 5314 9166 5446 9194
rect 5474 9166 5480 9194
rect 5120 9160 5480 9166
rect 5520 9194 5880 9200
rect 5520 9166 5526 9194
rect 5554 9166 5686 9194
rect 5714 9166 5846 9194
rect 5874 9166 5880 9194
rect 5520 9160 5880 9166
rect 5920 9194 6120 9200
rect 5920 9166 5926 9194
rect 5954 9166 6086 9194
rect 6114 9166 6120 9194
rect 5920 9160 6120 9166
rect 6160 9194 6360 9200
rect 6160 9166 6166 9194
rect 6194 9166 6326 9194
rect 6354 9166 6360 9194
rect 6160 9160 6360 9166
rect 4240 9114 6360 9120
rect 4240 9086 5126 9114
rect 5154 9086 5286 9114
rect 5314 9086 5446 9114
rect 5474 9086 6360 9114
rect 4240 9080 6360 9086
rect 4200 9034 6400 9040
rect 4200 9006 5366 9034
rect 5394 9006 6400 9034
rect 4200 9000 6400 9006
rect 4240 8954 6360 8960
rect 4240 8926 5126 8954
rect 5154 8926 5286 8954
rect 5314 8926 5446 8954
rect 5474 8926 6360 8954
rect 4240 8920 6360 8926
rect 4240 8874 4440 8880
rect 4240 8846 4246 8874
rect 4274 8846 4406 8874
rect 4434 8846 4440 8874
rect 4240 8840 4440 8846
rect 4480 8874 4680 8880
rect 4480 8846 4486 8874
rect 4514 8846 4646 8874
rect 4674 8846 4680 8874
rect 4480 8840 4680 8846
rect 4720 8874 5080 8880
rect 4720 8846 4726 8874
rect 4754 8846 4886 8874
rect 4914 8846 5046 8874
rect 5074 8846 5080 8874
rect 4720 8840 5080 8846
rect 5120 8874 5480 8880
rect 5120 8846 5126 8874
rect 5154 8846 5286 8874
rect 5314 8846 5446 8874
rect 5474 8846 5480 8874
rect 5120 8840 5480 8846
rect 5520 8874 5880 8880
rect 5520 8846 5526 8874
rect 5554 8846 5686 8874
rect 5714 8846 5846 8874
rect 5874 8846 5880 8874
rect 5520 8840 5880 8846
rect 5920 8874 6120 8880
rect 5920 8846 5926 8874
rect 5954 8846 6086 8874
rect 6114 8846 6120 8874
rect 5920 8840 6120 8846
rect 6160 8874 6360 8880
rect 6160 8846 6166 8874
rect 6194 8846 6326 8874
rect 6354 8846 6360 8874
rect 6160 8840 6360 8846
rect 4240 8794 4440 8800
rect 4240 8766 4246 8794
rect 4274 8766 4406 8794
rect 4434 8766 4440 8794
rect 4240 8760 4440 8766
rect 4480 8794 4680 8800
rect 4480 8766 4486 8794
rect 4514 8766 4646 8794
rect 4674 8766 4680 8794
rect 4480 8760 4680 8766
rect 4720 8794 5080 8800
rect 4720 8766 4726 8794
rect 4754 8766 4886 8794
rect 4914 8766 5046 8794
rect 5074 8766 5080 8794
rect 4720 8760 5080 8766
rect 5120 8794 5480 8800
rect 5120 8766 5126 8794
rect 5154 8766 5286 8794
rect 5314 8766 5446 8794
rect 5474 8766 5480 8794
rect 5120 8760 5480 8766
rect 5520 8794 5880 8800
rect 5520 8766 5526 8794
rect 5554 8766 5686 8794
rect 5714 8766 5846 8794
rect 5874 8766 5880 8794
rect 5520 8760 5880 8766
rect 5920 8794 6120 8800
rect 5920 8766 5926 8794
rect 5954 8766 6086 8794
rect 6114 8766 6120 8794
rect 5920 8760 6120 8766
rect 6160 8794 6360 8800
rect 6160 8766 6166 8794
rect 6194 8766 6326 8794
rect 6354 8766 6360 8794
rect 6160 8760 6360 8766
rect 4240 8714 4440 8720
rect 4240 8686 4246 8714
rect 4274 8686 4406 8714
rect 4434 8686 4440 8714
rect 4240 8680 4440 8686
rect 4480 8714 4680 8720
rect 4480 8686 4486 8714
rect 4514 8686 4646 8714
rect 4674 8686 4680 8714
rect 4480 8680 4680 8686
rect 4720 8714 5080 8720
rect 4720 8686 4726 8714
rect 4754 8686 4886 8714
rect 4914 8686 5046 8714
rect 5074 8686 5080 8714
rect 4720 8680 5080 8686
rect 5120 8714 5480 8720
rect 5120 8686 5126 8714
rect 5154 8686 5286 8714
rect 5314 8686 5446 8714
rect 5474 8686 5480 8714
rect 5120 8680 5480 8686
rect 5520 8714 5880 8720
rect 5520 8686 5526 8714
rect 5554 8686 5686 8714
rect 5714 8686 5846 8714
rect 5874 8686 5880 8714
rect 5520 8680 5880 8686
rect 5920 8714 6120 8720
rect 5920 8686 5926 8714
rect 5954 8686 6086 8714
rect 6114 8686 6120 8714
rect 5920 8680 6120 8686
rect 6160 8714 6360 8720
rect 6160 8686 6166 8714
rect 6194 8686 6326 8714
rect 6354 8686 6360 8714
rect 6160 8680 6360 8686
rect 4240 8634 4440 8640
rect 4240 8606 4246 8634
rect 4274 8606 4406 8634
rect 4434 8606 4440 8634
rect 4240 8600 4440 8606
rect 4480 8634 4680 8640
rect 4480 8606 4486 8634
rect 4514 8606 4646 8634
rect 4674 8606 4680 8634
rect 4480 8600 4680 8606
rect 4720 8634 5080 8640
rect 4720 8606 4726 8634
rect 4754 8606 4886 8634
rect 4914 8606 5046 8634
rect 5074 8606 5080 8634
rect 4720 8600 5080 8606
rect 5120 8634 5480 8640
rect 5120 8606 5126 8634
rect 5154 8606 5286 8634
rect 5314 8606 5446 8634
rect 5474 8606 5480 8634
rect 5120 8600 5480 8606
rect 5520 8634 5880 8640
rect 5520 8606 5526 8634
rect 5554 8606 5686 8634
rect 5714 8606 5846 8634
rect 5874 8606 5880 8634
rect 5520 8600 5880 8606
rect 5920 8634 6120 8640
rect 5920 8606 5926 8634
rect 5954 8606 6086 8634
rect 6114 8606 6120 8634
rect 5920 8600 6120 8606
rect 6160 8634 6360 8640
rect 6160 8606 6166 8634
rect 6194 8606 6326 8634
rect 6354 8606 6360 8634
rect 6160 8600 6360 8606
rect 4240 8554 4440 8560
rect 4240 8526 4246 8554
rect 4274 8526 4406 8554
rect 4434 8526 4440 8554
rect 4240 8520 4440 8526
rect 4480 8554 4680 8560
rect 4480 8526 4486 8554
rect 4514 8526 4646 8554
rect 4674 8526 4680 8554
rect 4480 8520 4680 8526
rect 4720 8554 5080 8560
rect 4720 8526 4726 8554
rect 4754 8526 4886 8554
rect 4914 8526 5046 8554
rect 5074 8526 5080 8554
rect 4720 8520 5080 8526
rect 5120 8554 5480 8560
rect 5120 8526 5126 8554
rect 5154 8526 5286 8554
rect 5314 8526 5446 8554
rect 5474 8526 5480 8554
rect 5120 8520 5480 8526
rect 5520 8554 5880 8560
rect 5520 8526 5526 8554
rect 5554 8526 5686 8554
rect 5714 8526 5846 8554
rect 5874 8526 5880 8554
rect 5520 8520 5880 8526
rect 5920 8554 6120 8560
rect 5920 8526 5926 8554
rect 5954 8526 6086 8554
rect 6114 8526 6120 8554
rect 5920 8520 6120 8526
rect 6160 8554 6360 8560
rect 6160 8526 6166 8554
rect 6194 8526 6326 8554
rect 6354 8526 6360 8554
rect 6160 8520 6360 8526
rect 4240 8474 6360 8480
rect 4240 8446 4886 8474
rect 4914 8446 5046 8474
rect 5074 8446 5686 8474
rect 5714 8446 5846 8474
rect 5874 8446 6360 8474
rect 4240 8440 6360 8446
rect 4200 8394 5000 8400
rect 4200 8366 4966 8394
rect 4994 8366 5000 8394
rect 4200 8360 5000 8366
rect 5760 8394 6400 8400
rect 5760 8366 5766 8394
rect 5794 8366 6400 8394
rect 5760 8360 6400 8366
rect 4240 8314 6360 8320
rect 4240 8286 4886 8314
rect 4914 8286 5046 8314
rect 5074 8286 5526 8314
rect 5554 8286 5686 8314
rect 5714 8286 5846 8314
rect 5874 8286 6360 8314
rect 4240 8280 6360 8286
rect 4200 8234 6400 8240
rect 4200 8206 5606 8234
rect 5634 8206 6400 8234
rect 4200 8200 6400 8206
rect 4240 8154 6360 8160
rect 4240 8126 5526 8154
rect 5554 8126 5686 8154
rect 5714 8126 6360 8154
rect 4240 8120 6360 8126
rect 4240 8074 6360 8080
rect 4240 8046 5046 8074
rect 5074 8046 5526 8074
rect 5554 8046 6360 8074
rect 4240 8040 6360 8046
rect 4240 7994 6360 8000
rect 4240 7966 5126 7994
rect 5154 7966 5286 7994
rect 5314 7966 5446 7994
rect 5474 7966 6360 7994
rect 4240 7960 6360 7966
rect 4200 7914 6400 7920
rect 4200 7886 5206 7914
rect 5234 7886 6400 7914
rect 4200 7880 6400 7886
rect 4240 7834 6360 7840
rect 4240 7806 5126 7834
rect 5154 7806 5286 7834
rect 5314 7806 5446 7834
rect 5474 7806 6360 7834
rect 4240 7800 6360 7806
rect 4240 7754 6360 7760
rect 4240 7726 5046 7754
rect 5074 7726 5526 7754
rect 5554 7726 6360 7754
rect 4240 7720 6360 7726
rect 4240 7634 4440 7640
rect 4240 7606 4246 7634
rect 4274 7606 4406 7634
rect 4434 7606 4440 7634
rect 4240 7600 4440 7606
rect 4480 7634 4680 7640
rect 4480 7606 4486 7634
rect 4514 7606 4646 7634
rect 4674 7606 4680 7634
rect 4480 7600 4680 7606
rect 4720 7634 5080 7640
rect 4720 7606 4726 7634
rect 4754 7606 4886 7634
rect 4914 7606 5046 7634
rect 5074 7606 5080 7634
rect 4720 7600 5080 7606
rect 5120 7634 5480 7640
rect 5120 7606 5126 7634
rect 5154 7606 5286 7634
rect 5314 7606 5446 7634
rect 5474 7606 5480 7634
rect 5120 7600 5480 7606
rect 5520 7634 5880 7640
rect 5520 7606 5526 7634
rect 5554 7606 5686 7634
rect 5714 7606 5846 7634
rect 5874 7606 5880 7634
rect 5520 7600 5880 7606
rect 5920 7634 6120 7640
rect 5920 7606 5926 7634
rect 5954 7606 6086 7634
rect 6114 7606 6120 7634
rect 5920 7600 6120 7606
rect 6160 7634 6360 7640
rect 6160 7606 6166 7634
rect 6194 7606 6326 7634
rect 6354 7606 6360 7634
rect 6160 7600 6360 7606
rect 4240 7554 4440 7560
rect 4240 7526 4246 7554
rect 4274 7526 4406 7554
rect 4434 7526 4440 7554
rect 4240 7520 4440 7526
rect 4480 7554 4680 7560
rect 4480 7526 4486 7554
rect 4514 7526 4646 7554
rect 4674 7526 4680 7554
rect 4480 7520 4680 7526
rect 4720 7554 5080 7560
rect 4720 7526 4726 7554
rect 4754 7526 4886 7554
rect 4914 7526 5046 7554
rect 5074 7526 5080 7554
rect 4720 7520 5080 7526
rect 5120 7554 5480 7560
rect 5120 7526 5126 7554
rect 5154 7526 5286 7554
rect 5314 7526 5446 7554
rect 5474 7526 5480 7554
rect 5120 7520 5480 7526
rect 5520 7554 5880 7560
rect 5520 7526 5526 7554
rect 5554 7526 5686 7554
rect 5714 7526 5846 7554
rect 5874 7526 5880 7554
rect 5520 7520 5880 7526
rect 5920 7554 6120 7560
rect 5920 7526 5926 7554
rect 5954 7526 6086 7554
rect 6114 7526 6120 7554
rect 5920 7520 6120 7526
rect 6160 7554 6360 7560
rect 6160 7526 6166 7554
rect 6194 7526 6326 7554
rect 6354 7526 6360 7554
rect 6160 7520 6360 7526
rect 4240 7474 4440 7480
rect 4240 7446 4246 7474
rect 4274 7446 4406 7474
rect 4434 7446 4440 7474
rect 4240 7440 4440 7446
rect 4480 7474 4680 7480
rect 4480 7446 4486 7474
rect 4514 7446 4646 7474
rect 4674 7446 4680 7474
rect 4480 7440 4680 7446
rect 4720 7474 5080 7480
rect 4720 7446 4726 7474
rect 4754 7446 4886 7474
rect 4914 7446 5046 7474
rect 5074 7446 5080 7474
rect 4720 7440 5080 7446
rect 5120 7474 5480 7480
rect 5120 7446 5126 7474
rect 5154 7446 5286 7474
rect 5314 7446 5446 7474
rect 5474 7446 5480 7474
rect 5120 7440 5480 7446
rect 5520 7474 5880 7480
rect 5520 7446 5526 7474
rect 5554 7446 5686 7474
rect 5714 7446 5846 7474
rect 5874 7446 5880 7474
rect 5520 7440 5880 7446
rect 5920 7474 6120 7480
rect 5920 7446 5926 7474
rect 5954 7446 6086 7474
rect 6114 7446 6120 7474
rect 5920 7440 6120 7446
rect 6160 7474 6360 7480
rect 6160 7446 6166 7474
rect 6194 7446 6326 7474
rect 6354 7446 6360 7474
rect 6160 7440 6360 7446
rect 4240 7394 4440 7400
rect 4240 7366 4246 7394
rect 4274 7366 4406 7394
rect 4434 7366 4440 7394
rect 4240 7360 4440 7366
rect 4480 7394 4680 7400
rect 4480 7366 4486 7394
rect 4514 7366 4646 7394
rect 4674 7366 4680 7394
rect 4480 7360 4680 7366
rect 4720 7394 5080 7400
rect 4720 7366 4726 7394
rect 4754 7366 4886 7394
rect 4914 7366 5046 7394
rect 5074 7366 5080 7394
rect 4720 7360 5080 7366
rect 5120 7394 5480 7400
rect 5120 7366 5126 7394
rect 5154 7366 5286 7394
rect 5314 7366 5446 7394
rect 5474 7366 5480 7394
rect 5120 7360 5480 7366
rect 5520 7394 5880 7400
rect 5520 7366 5526 7394
rect 5554 7366 5686 7394
rect 5714 7366 5846 7394
rect 5874 7366 5880 7394
rect 5520 7360 5880 7366
rect 5920 7394 6120 7400
rect 5920 7366 5926 7394
rect 5954 7366 6086 7394
rect 6114 7366 6120 7394
rect 5920 7360 6120 7366
rect 6160 7394 6360 7400
rect 6160 7366 6166 7394
rect 6194 7366 6326 7394
rect 6354 7366 6360 7394
rect 6160 7360 6360 7366
rect 4240 7314 4440 7320
rect 4240 7286 4246 7314
rect 4274 7286 4406 7314
rect 4434 7286 4440 7314
rect 4240 7280 4440 7286
rect 4480 7314 4680 7320
rect 4480 7286 4486 7314
rect 4514 7286 4646 7314
rect 4674 7286 4680 7314
rect 4480 7280 4680 7286
rect 4720 7314 5080 7320
rect 4720 7286 4726 7314
rect 4754 7286 4886 7314
rect 4914 7286 5046 7314
rect 5074 7286 5080 7314
rect 4720 7280 5080 7286
rect 5120 7314 5480 7320
rect 5120 7286 5126 7314
rect 5154 7286 5286 7314
rect 5314 7286 5446 7314
rect 5474 7286 5480 7314
rect 5120 7280 5480 7286
rect 5520 7314 5880 7320
rect 5520 7286 5526 7314
rect 5554 7286 5686 7314
rect 5714 7286 5846 7314
rect 5874 7286 5880 7314
rect 5520 7280 5880 7286
rect 5920 7314 6120 7320
rect 5920 7286 5926 7314
rect 5954 7286 6086 7314
rect 6114 7286 6120 7314
rect 5920 7280 6120 7286
rect 6160 7314 6360 7320
rect 6160 7286 6166 7314
rect 6194 7286 6326 7314
rect 6354 7286 6360 7314
rect 6160 7280 6360 7286
rect 4240 7234 4440 7240
rect 4240 7206 4246 7234
rect 4274 7206 4406 7234
rect 4434 7206 4440 7234
rect 4240 7200 4440 7206
rect 4480 7234 4680 7240
rect 4480 7206 4486 7234
rect 4514 7206 4646 7234
rect 4674 7206 4680 7234
rect 4480 7200 4680 7206
rect 4720 7234 5080 7240
rect 4720 7206 4726 7234
rect 4754 7206 4886 7234
rect 4914 7206 5046 7234
rect 5074 7206 5080 7234
rect 4720 7200 5080 7206
rect 5120 7234 5480 7240
rect 5120 7206 5126 7234
rect 5154 7206 5286 7234
rect 5314 7206 5446 7234
rect 5474 7206 5480 7234
rect 5120 7200 5480 7206
rect 5520 7234 5880 7240
rect 5520 7206 5526 7234
rect 5554 7206 5686 7234
rect 5714 7206 5846 7234
rect 5874 7206 5880 7234
rect 5520 7200 5880 7206
rect 5920 7234 6120 7240
rect 5920 7206 5926 7234
rect 5954 7206 6086 7234
rect 6114 7206 6120 7234
rect 5920 7200 6120 7206
rect 6160 7234 6360 7240
rect 6160 7206 6166 7234
rect 6194 7206 6326 7234
rect 6354 7206 6360 7234
rect 6160 7200 6360 7206
rect 4240 7154 4440 7160
rect 4240 7126 4246 7154
rect 4274 7126 4406 7154
rect 4434 7126 4440 7154
rect 4240 7120 4440 7126
rect 4480 7154 4680 7160
rect 4480 7126 4486 7154
rect 4514 7126 4646 7154
rect 4674 7126 4680 7154
rect 4480 7120 4680 7126
rect 4720 7154 5080 7160
rect 4720 7126 4726 7154
rect 4754 7126 4886 7154
rect 4914 7126 5046 7154
rect 5074 7126 5080 7154
rect 4720 7120 5080 7126
rect 5120 7154 5480 7160
rect 5120 7126 5126 7154
rect 5154 7126 5286 7154
rect 5314 7126 5446 7154
rect 5474 7126 5480 7154
rect 5120 7120 5480 7126
rect 5520 7154 5880 7160
rect 5520 7126 5526 7154
rect 5554 7126 5686 7154
rect 5714 7126 5846 7154
rect 5874 7126 5880 7154
rect 5520 7120 5880 7126
rect 5920 7154 6120 7160
rect 5920 7126 5926 7154
rect 5954 7126 6086 7154
rect 6114 7126 6120 7154
rect 5920 7120 6120 7126
rect 6160 7154 6360 7160
rect 6160 7126 6166 7154
rect 6194 7126 6326 7154
rect 6354 7126 6360 7154
rect 6160 7120 6360 7126
rect 4240 7074 4440 7080
rect 4240 7046 4246 7074
rect 4274 7046 4406 7074
rect 4434 7046 4440 7074
rect 4240 7040 4440 7046
rect 4480 7074 4680 7080
rect 4480 7046 4486 7074
rect 4514 7046 4646 7074
rect 4674 7046 4680 7074
rect 4480 7040 4680 7046
rect 4720 7074 5080 7080
rect 4720 7046 4726 7074
rect 4754 7046 4886 7074
rect 4914 7046 5046 7074
rect 5074 7046 5080 7074
rect 4720 7040 5080 7046
rect 5120 7074 5480 7080
rect 5120 7046 5126 7074
rect 5154 7046 5286 7074
rect 5314 7046 5446 7074
rect 5474 7046 5480 7074
rect 5120 7040 5480 7046
rect 5520 7074 5880 7080
rect 5520 7046 5526 7074
rect 5554 7046 5686 7074
rect 5714 7046 5846 7074
rect 5874 7046 5880 7074
rect 5520 7040 5880 7046
rect 5920 7074 6120 7080
rect 5920 7046 5926 7074
rect 5954 7046 6086 7074
rect 6114 7046 6120 7074
rect 5920 7040 6120 7046
rect 6160 7074 6360 7080
rect 6160 7046 6166 7074
rect 6194 7046 6326 7074
rect 6354 7046 6360 7074
rect 6160 7040 6360 7046
rect 4200 6994 6400 7000
rect 4200 6966 4486 6994
rect 4514 6966 4646 6994
rect 4674 6966 6400 6994
rect 4200 6960 6400 6966
rect 4200 6914 6400 6920
rect 4200 6886 4566 6914
rect 4594 6886 6400 6914
rect 4200 6880 6400 6886
rect 4200 6834 6400 6840
rect 4200 6806 4486 6834
rect 4514 6806 4646 6834
rect 4674 6806 6400 6834
rect 4200 6800 6400 6806
rect 4240 6754 4440 6760
rect 4240 6726 4246 6754
rect 4274 6726 4406 6754
rect 4434 6726 4440 6754
rect 4240 6720 4440 6726
rect 4480 6754 4680 6760
rect 4480 6726 4486 6754
rect 4514 6726 4646 6754
rect 4674 6726 4680 6754
rect 4480 6720 4680 6726
rect 4720 6754 5080 6760
rect 4720 6726 4726 6754
rect 4754 6726 4886 6754
rect 4914 6726 5046 6754
rect 5074 6726 5080 6754
rect 4720 6720 5080 6726
rect 5120 6754 5480 6760
rect 5120 6726 5126 6754
rect 5154 6726 5286 6754
rect 5314 6726 5446 6754
rect 5474 6726 5480 6754
rect 5120 6720 5480 6726
rect 5520 6754 5880 6760
rect 5520 6726 5526 6754
rect 5554 6726 5686 6754
rect 5714 6726 5846 6754
rect 5874 6726 5880 6754
rect 5520 6720 5880 6726
rect 5920 6754 6120 6760
rect 5920 6726 5926 6754
rect 5954 6726 6086 6754
rect 6114 6726 6120 6754
rect 5920 6720 6120 6726
rect 6160 6754 6360 6760
rect 6160 6726 6166 6754
rect 6194 6726 6326 6754
rect 6354 6726 6360 6754
rect 6160 6720 6360 6726
rect 4240 6674 4440 6680
rect 4240 6646 4246 6674
rect 4274 6646 4406 6674
rect 4434 6646 4440 6674
rect 4240 6640 4440 6646
rect 4480 6674 4680 6680
rect 4480 6646 4486 6674
rect 4514 6646 4646 6674
rect 4674 6646 4680 6674
rect 4480 6640 4680 6646
rect 4720 6674 5080 6680
rect 4720 6646 4726 6674
rect 4754 6646 4886 6674
rect 4914 6646 5046 6674
rect 5074 6646 5080 6674
rect 4720 6640 5080 6646
rect 5120 6674 5480 6680
rect 5120 6646 5126 6674
rect 5154 6646 5286 6674
rect 5314 6646 5446 6674
rect 5474 6646 5480 6674
rect 5120 6640 5480 6646
rect 5520 6674 5880 6680
rect 5520 6646 5526 6674
rect 5554 6646 5686 6674
rect 5714 6646 5846 6674
rect 5874 6646 5880 6674
rect 5520 6640 5880 6646
rect 5920 6674 6120 6680
rect 5920 6646 5926 6674
rect 5954 6646 6086 6674
rect 6114 6646 6120 6674
rect 5920 6640 6120 6646
rect 6160 6674 6360 6680
rect 6160 6646 6166 6674
rect 6194 6646 6326 6674
rect 6354 6646 6360 6674
rect 6160 6640 6360 6646
rect 4240 6594 4440 6600
rect 4240 6566 4246 6594
rect 4274 6566 4406 6594
rect 4434 6566 4440 6594
rect 4240 6560 4440 6566
rect 4480 6594 4680 6600
rect 4480 6566 4486 6594
rect 4514 6566 4646 6594
rect 4674 6566 4680 6594
rect 4480 6560 4680 6566
rect 4720 6594 5080 6600
rect 4720 6566 4726 6594
rect 4754 6566 4886 6594
rect 4914 6566 5046 6594
rect 5074 6566 5080 6594
rect 4720 6560 5080 6566
rect 5120 6594 5480 6600
rect 5120 6566 5126 6594
rect 5154 6566 5286 6594
rect 5314 6566 5446 6594
rect 5474 6566 5480 6594
rect 5120 6560 5480 6566
rect 5520 6594 5880 6600
rect 5520 6566 5526 6594
rect 5554 6566 5686 6594
rect 5714 6566 5846 6594
rect 5874 6566 5880 6594
rect 5520 6560 5880 6566
rect 5920 6594 6120 6600
rect 5920 6566 5926 6594
rect 5954 6566 6086 6594
rect 6114 6566 6120 6594
rect 5920 6560 6120 6566
rect 6160 6594 6360 6600
rect 6160 6566 6166 6594
rect 6194 6566 6326 6594
rect 6354 6566 6360 6594
rect 6160 6560 6360 6566
rect 4240 6514 4440 6520
rect 4240 6486 4246 6514
rect 4274 6486 4406 6514
rect 4434 6486 4440 6514
rect 4240 6480 4440 6486
rect 4480 6514 4680 6520
rect 4480 6486 4486 6514
rect 4514 6486 4646 6514
rect 4674 6486 4680 6514
rect 4480 6480 4680 6486
rect 4720 6514 5080 6520
rect 4720 6486 4726 6514
rect 4754 6486 4886 6514
rect 4914 6486 5046 6514
rect 5074 6486 5080 6514
rect 4720 6480 5080 6486
rect 5120 6514 5480 6520
rect 5120 6486 5126 6514
rect 5154 6486 5286 6514
rect 5314 6486 5446 6514
rect 5474 6486 5480 6514
rect 5120 6480 5480 6486
rect 5520 6514 5880 6520
rect 5520 6486 5526 6514
rect 5554 6486 5686 6514
rect 5714 6486 5846 6514
rect 5874 6486 5880 6514
rect 5520 6480 5880 6486
rect 5920 6514 6120 6520
rect 5920 6486 5926 6514
rect 5954 6486 6086 6514
rect 6114 6486 6120 6514
rect 5920 6480 6120 6486
rect 6160 6514 6360 6520
rect 6160 6486 6166 6514
rect 6194 6486 6326 6514
rect 6354 6486 6360 6514
rect 6160 6480 6360 6486
rect 4240 6434 4440 6440
rect 4240 6406 4246 6434
rect 4274 6406 4406 6434
rect 4434 6406 4440 6434
rect 4240 6400 4440 6406
rect 4480 6434 4680 6440
rect 4480 6406 4486 6434
rect 4514 6406 4646 6434
rect 4674 6406 4680 6434
rect 4480 6400 4680 6406
rect 4720 6434 5080 6440
rect 4720 6406 4726 6434
rect 4754 6406 4886 6434
rect 4914 6406 5046 6434
rect 5074 6406 5080 6434
rect 4720 6400 5080 6406
rect 5120 6434 5480 6440
rect 5120 6406 5126 6434
rect 5154 6406 5286 6434
rect 5314 6406 5446 6434
rect 5474 6406 5480 6434
rect 5120 6400 5480 6406
rect 5520 6434 5880 6440
rect 5520 6406 5526 6434
rect 5554 6406 5686 6434
rect 5714 6406 5846 6434
rect 5874 6406 5880 6434
rect 5520 6400 5880 6406
rect 5920 6434 6120 6440
rect 5920 6406 5926 6434
rect 5954 6406 6086 6434
rect 6114 6406 6120 6434
rect 5920 6400 6120 6406
rect 6160 6434 6360 6440
rect 6160 6406 6166 6434
rect 6194 6406 6326 6434
rect 6354 6406 6360 6434
rect 6160 6400 6360 6406
rect 4240 6354 4440 6360
rect 4240 6326 4246 6354
rect 4274 6326 4406 6354
rect 4434 6326 4440 6354
rect 4240 6320 4440 6326
rect 4480 6354 4680 6360
rect 4480 6326 4486 6354
rect 4514 6326 4646 6354
rect 4674 6326 4680 6354
rect 4480 6320 4680 6326
rect 4720 6354 5080 6360
rect 4720 6326 4726 6354
rect 4754 6326 4886 6354
rect 4914 6326 5046 6354
rect 5074 6326 5080 6354
rect 4720 6320 5080 6326
rect 5120 6354 5480 6360
rect 5120 6326 5126 6354
rect 5154 6326 5286 6354
rect 5314 6326 5446 6354
rect 5474 6326 5480 6354
rect 5120 6320 5480 6326
rect 5520 6354 5880 6360
rect 5520 6326 5526 6354
rect 5554 6326 5686 6354
rect 5714 6326 5846 6354
rect 5874 6326 5880 6354
rect 5520 6320 5880 6326
rect 5920 6354 6120 6360
rect 5920 6326 5926 6354
rect 5954 6326 6086 6354
rect 6114 6326 6120 6354
rect 5920 6320 6120 6326
rect 6160 6354 6360 6360
rect 6160 6326 6166 6354
rect 6194 6326 6326 6354
rect 6354 6326 6360 6354
rect 6160 6320 6360 6326
rect 4240 6234 6360 6240
rect 4240 6206 4726 6234
rect 4754 6206 4886 6234
rect 4914 6206 5046 6234
rect 5074 6206 6360 6234
rect 4240 6200 6360 6206
rect 4200 6154 4840 6160
rect 4200 6126 4806 6154
rect 4834 6126 4840 6154
rect 4200 6120 4840 6126
rect 4960 6154 6400 6160
rect 4960 6126 4966 6154
rect 4994 6126 6400 6154
rect 4960 6120 6400 6126
rect 4240 6074 6360 6080
rect 4240 6046 4726 6074
rect 4754 6046 4886 6074
rect 4914 6046 5046 6074
rect 5074 6046 6360 6074
rect 4240 6040 6360 6046
rect 4200 5994 6400 6000
rect 4200 5966 4966 5994
rect 4994 5966 6400 5994
rect 4200 5960 6400 5966
rect 4240 5914 6360 5920
rect 4240 5886 4726 5914
rect 4754 5886 4886 5914
rect 4914 5886 5046 5914
rect 5074 5886 6360 5914
rect 4240 5880 6360 5886
rect 4240 5794 4440 5800
rect 4240 5766 4246 5794
rect 4274 5766 4406 5794
rect 4434 5766 4440 5794
rect 4240 5760 4440 5766
rect 4480 5794 4680 5800
rect 4480 5766 4486 5794
rect 4514 5766 4646 5794
rect 4674 5766 4680 5794
rect 4480 5760 4680 5766
rect 4720 5794 5080 5800
rect 4720 5766 4726 5794
rect 4754 5766 4886 5794
rect 4914 5766 5046 5794
rect 5074 5766 5080 5794
rect 4720 5760 5080 5766
rect 5120 5794 5480 5800
rect 5120 5766 5126 5794
rect 5154 5766 5286 5794
rect 5314 5766 5446 5794
rect 5474 5766 5480 5794
rect 5120 5760 5480 5766
rect 5520 5794 5880 5800
rect 5520 5766 5526 5794
rect 5554 5766 5686 5794
rect 5714 5766 5846 5794
rect 5874 5766 5880 5794
rect 5520 5760 5880 5766
rect 5920 5794 6120 5800
rect 5920 5766 5926 5794
rect 5954 5766 6086 5794
rect 6114 5766 6120 5794
rect 5920 5760 6120 5766
rect 6160 5794 6360 5800
rect 6160 5766 6166 5794
rect 6194 5766 6326 5794
rect 6354 5766 6360 5794
rect 6160 5760 6360 5766
rect 4240 5714 4440 5720
rect 4240 5686 4246 5714
rect 4274 5686 4406 5714
rect 4434 5686 4440 5714
rect 4240 5680 4440 5686
rect 4480 5714 4680 5720
rect 4480 5686 4486 5714
rect 4514 5686 4646 5714
rect 4674 5686 4680 5714
rect 4480 5680 4680 5686
rect 4720 5714 5080 5720
rect 4720 5686 4726 5714
rect 4754 5686 4886 5714
rect 4914 5686 5046 5714
rect 5074 5686 5080 5714
rect 4720 5680 5080 5686
rect 5120 5714 5480 5720
rect 5120 5686 5126 5714
rect 5154 5686 5286 5714
rect 5314 5686 5446 5714
rect 5474 5686 5480 5714
rect 5120 5680 5480 5686
rect 5520 5714 5880 5720
rect 5520 5686 5526 5714
rect 5554 5686 5686 5714
rect 5714 5686 5846 5714
rect 5874 5686 5880 5714
rect 5520 5680 5880 5686
rect 5920 5714 6120 5720
rect 5920 5686 5926 5714
rect 5954 5686 6086 5714
rect 6114 5686 6120 5714
rect 5920 5680 6120 5686
rect 6160 5714 6360 5720
rect 6160 5686 6166 5714
rect 6194 5686 6326 5714
rect 6354 5686 6360 5714
rect 6160 5680 6360 5686
rect 4240 5634 4440 5640
rect 4240 5606 4246 5634
rect 4274 5606 4406 5634
rect 4434 5606 4440 5634
rect 4240 5600 4440 5606
rect 4480 5634 4680 5640
rect 4480 5606 4486 5634
rect 4514 5606 4646 5634
rect 4674 5606 4680 5634
rect 4480 5600 4680 5606
rect 4720 5634 5080 5640
rect 4720 5606 4726 5634
rect 4754 5606 4886 5634
rect 4914 5606 5046 5634
rect 5074 5606 5080 5634
rect 4720 5600 5080 5606
rect 5120 5634 5480 5640
rect 5120 5606 5126 5634
rect 5154 5606 5286 5634
rect 5314 5606 5446 5634
rect 5474 5606 5480 5634
rect 5120 5600 5480 5606
rect 5520 5634 5880 5640
rect 5520 5606 5526 5634
rect 5554 5606 5686 5634
rect 5714 5606 5846 5634
rect 5874 5606 5880 5634
rect 5520 5600 5880 5606
rect 5920 5634 6120 5640
rect 5920 5606 5926 5634
rect 5954 5606 6086 5634
rect 6114 5606 6120 5634
rect 5920 5600 6120 5606
rect 6160 5634 6360 5640
rect 6160 5606 6166 5634
rect 6194 5606 6326 5634
rect 6354 5606 6360 5634
rect 6160 5600 6360 5606
rect 4240 5554 4440 5560
rect 4240 5526 4246 5554
rect 4274 5526 4406 5554
rect 4434 5526 4440 5554
rect 4240 5520 4440 5526
rect 4480 5554 4680 5560
rect 4480 5526 4486 5554
rect 4514 5526 4646 5554
rect 4674 5526 4680 5554
rect 4480 5520 4680 5526
rect 4720 5554 5080 5560
rect 4720 5526 4726 5554
rect 4754 5526 4886 5554
rect 4914 5526 5046 5554
rect 5074 5526 5080 5554
rect 4720 5520 5080 5526
rect 5120 5554 5480 5560
rect 5120 5526 5126 5554
rect 5154 5526 5286 5554
rect 5314 5526 5446 5554
rect 5474 5526 5480 5554
rect 5120 5520 5480 5526
rect 5520 5554 5880 5560
rect 5520 5526 5526 5554
rect 5554 5526 5686 5554
rect 5714 5526 5846 5554
rect 5874 5526 5880 5554
rect 5520 5520 5880 5526
rect 5920 5554 6120 5560
rect 5920 5526 5926 5554
rect 5954 5526 6086 5554
rect 6114 5526 6120 5554
rect 5920 5520 6120 5526
rect 6160 5554 6360 5560
rect 6160 5526 6166 5554
rect 6194 5526 6326 5554
rect 6354 5526 6360 5554
rect 6160 5520 6360 5526
rect 4240 5474 4440 5480
rect 4240 5446 4246 5474
rect 4274 5446 4406 5474
rect 4434 5446 4440 5474
rect 4240 5440 4440 5446
rect 4480 5474 4680 5480
rect 4480 5446 4486 5474
rect 4514 5446 4646 5474
rect 4674 5446 4680 5474
rect 4480 5440 4680 5446
rect 4720 5474 5080 5480
rect 4720 5446 4726 5474
rect 4754 5446 4886 5474
rect 4914 5446 5046 5474
rect 5074 5446 5080 5474
rect 4720 5440 5080 5446
rect 5120 5474 5480 5480
rect 5120 5446 5126 5474
rect 5154 5446 5286 5474
rect 5314 5446 5446 5474
rect 5474 5446 5480 5474
rect 5120 5440 5480 5446
rect 5520 5474 5880 5480
rect 5520 5446 5526 5474
rect 5554 5446 5686 5474
rect 5714 5446 5846 5474
rect 5874 5446 5880 5474
rect 5520 5440 5880 5446
rect 5920 5474 6120 5480
rect 5920 5446 5926 5474
rect 5954 5446 6086 5474
rect 6114 5446 6120 5474
rect 5920 5440 6120 5446
rect 6160 5474 6360 5480
rect 6160 5446 6166 5474
rect 6194 5446 6326 5474
rect 6354 5446 6360 5474
rect 6160 5440 6360 5446
rect 4240 5394 4440 5400
rect 4240 5366 4246 5394
rect 4274 5366 4406 5394
rect 4434 5366 4440 5394
rect 4240 5360 4440 5366
rect 4480 5394 4680 5400
rect 4480 5366 4486 5394
rect 4514 5366 4646 5394
rect 4674 5366 4680 5394
rect 4480 5360 4680 5366
rect 4720 5394 5080 5400
rect 4720 5366 4726 5394
rect 4754 5366 4886 5394
rect 4914 5366 5046 5394
rect 5074 5366 5080 5394
rect 4720 5360 5080 5366
rect 5120 5394 5480 5400
rect 5120 5366 5126 5394
rect 5154 5366 5286 5394
rect 5314 5366 5446 5394
rect 5474 5366 5480 5394
rect 5120 5360 5480 5366
rect 5520 5394 5880 5400
rect 5520 5366 5526 5394
rect 5554 5366 5686 5394
rect 5714 5366 5846 5394
rect 5874 5366 5880 5394
rect 5520 5360 5880 5366
rect 5920 5394 6120 5400
rect 5920 5366 5926 5394
rect 5954 5366 6086 5394
rect 6114 5366 6120 5394
rect 5920 5360 6120 5366
rect 6160 5394 6360 5400
rect 6160 5366 6166 5394
rect 6194 5366 6326 5394
rect 6354 5366 6360 5394
rect 6160 5360 6360 5366
rect 4240 5314 4440 5320
rect 4240 5286 4246 5314
rect 4274 5286 4406 5314
rect 4434 5286 4440 5314
rect 4240 5280 4440 5286
rect 4480 5314 4680 5320
rect 4480 5286 4486 5314
rect 4514 5286 4646 5314
rect 4674 5286 4680 5314
rect 4480 5280 4680 5286
rect 4720 5314 5080 5320
rect 4720 5286 4726 5314
rect 4754 5286 4886 5314
rect 4914 5286 5046 5314
rect 5074 5286 5080 5314
rect 4720 5280 5080 5286
rect 5120 5314 5480 5320
rect 5120 5286 5126 5314
rect 5154 5286 5286 5314
rect 5314 5286 5446 5314
rect 5474 5286 5480 5314
rect 5120 5280 5480 5286
rect 5520 5314 5880 5320
rect 5520 5286 5526 5314
rect 5554 5286 5686 5314
rect 5714 5286 5846 5314
rect 5874 5286 5880 5314
rect 5520 5280 5880 5286
rect 5920 5314 6120 5320
rect 5920 5286 5926 5314
rect 5954 5286 6086 5314
rect 6114 5286 6120 5314
rect 5920 5280 6120 5286
rect 6160 5314 6360 5320
rect 6160 5286 6166 5314
rect 6194 5286 6326 5314
rect 6354 5286 6360 5314
rect 6160 5280 6360 5286
rect 4240 5234 4440 5240
rect 4240 5206 4246 5234
rect 4274 5206 4406 5234
rect 4434 5206 4440 5234
rect 4240 5200 4440 5206
rect 4480 5234 4680 5240
rect 4480 5206 4486 5234
rect 4514 5206 4646 5234
rect 4674 5206 4680 5234
rect 4480 5200 4680 5206
rect 4720 5234 5080 5240
rect 4720 5206 4726 5234
rect 4754 5206 4886 5234
rect 4914 5206 5046 5234
rect 5074 5206 5080 5234
rect 4720 5200 5080 5206
rect 5120 5234 5480 5240
rect 5120 5206 5126 5234
rect 5154 5206 5286 5234
rect 5314 5206 5446 5234
rect 5474 5206 5480 5234
rect 5120 5200 5480 5206
rect 5520 5234 5880 5240
rect 5520 5206 5526 5234
rect 5554 5206 5686 5234
rect 5714 5206 5846 5234
rect 5874 5206 5880 5234
rect 5520 5200 5880 5206
rect 5920 5234 6120 5240
rect 5920 5206 5926 5234
rect 5954 5206 6086 5234
rect 6114 5206 6120 5234
rect 5920 5200 6120 5206
rect 6160 5234 6360 5240
rect 6160 5206 6166 5234
rect 6194 5206 6326 5234
rect 6354 5206 6360 5234
rect 6160 5200 6360 5206
rect 4240 5154 4440 5160
rect 4240 5126 4246 5154
rect 4274 5126 4406 5154
rect 4434 5126 4440 5154
rect 4240 5120 4440 5126
rect 4480 5154 4680 5160
rect 4480 5126 4486 5154
rect 4514 5126 4646 5154
rect 4674 5126 4680 5154
rect 4480 5120 4680 5126
rect 4720 5154 5080 5160
rect 4720 5126 4726 5154
rect 4754 5126 4886 5154
rect 4914 5126 5046 5154
rect 5074 5126 5080 5154
rect 4720 5120 5080 5126
rect 5120 5154 5480 5160
rect 5120 5126 5126 5154
rect 5154 5126 5286 5154
rect 5314 5126 5446 5154
rect 5474 5126 5480 5154
rect 5120 5120 5480 5126
rect 5520 5154 5880 5160
rect 5520 5126 5526 5154
rect 5554 5126 5686 5154
rect 5714 5126 5846 5154
rect 5874 5126 5880 5154
rect 5520 5120 5880 5126
rect 5920 5154 6120 5160
rect 5920 5126 5926 5154
rect 5954 5126 6086 5154
rect 6114 5126 6120 5154
rect 5920 5120 6120 5126
rect 6160 5154 6360 5160
rect 6160 5126 6166 5154
rect 6194 5126 6326 5154
rect 6354 5126 6360 5154
rect 6160 5120 6360 5126
rect 4240 5074 4440 5080
rect 4240 5046 4246 5074
rect 4274 5046 4406 5074
rect 4434 5046 4440 5074
rect 4240 5040 4440 5046
rect 4480 5074 4680 5080
rect 4480 5046 4486 5074
rect 4514 5046 4646 5074
rect 4674 5046 4680 5074
rect 4480 5040 4680 5046
rect 4720 5074 5080 5080
rect 4720 5046 4726 5074
rect 4754 5046 4886 5074
rect 4914 5046 5046 5074
rect 5074 5046 5080 5074
rect 4720 5040 5080 5046
rect 5120 5074 5480 5080
rect 5120 5046 5126 5074
rect 5154 5046 5286 5074
rect 5314 5046 5446 5074
rect 5474 5046 5480 5074
rect 5120 5040 5480 5046
rect 5520 5074 5880 5080
rect 5520 5046 5526 5074
rect 5554 5046 5686 5074
rect 5714 5046 5846 5074
rect 5874 5046 5880 5074
rect 5520 5040 5880 5046
rect 5920 5074 6120 5080
rect 5920 5046 5926 5074
rect 5954 5046 6086 5074
rect 6114 5046 6120 5074
rect 5920 5040 6120 5046
rect 6160 5074 6360 5080
rect 6160 5046 6166 5074
rect 6194 5046 6326 5074
rect 6354 5046 6360 5074
rect 6160 5040 6360 5046
rect 4240 4994 4440 5000
rect 4240 4966 4246 4994
rect 4274 4966 4406 4994
rect 4434 4966 4440 4994
rect 4240 4960 4440 4966
rect 4480 4994 4680 5000
rect 4480 4966 4486 4994
rect 4514 4966 4646 4994
rect 4674 4966 4680 4994
rect 4480 4960 4680 4966
rect 4720 4994 5080 5000
rect 4720 4966 4726 4994
rect 4754 4966 4886 4994
rect 4914 4966 5046 4994
rect 5074 4966 5080 4994
rect 4720 4960 5080 4966
rect 5120 4994 5480 5000
rect 5120 4966 5126 4994
rect 5154 4966 5286 4994
rect 5314 4966 5446 4994
rect 5474 4966 5480 4994
rect 5120 4960 5480 4966
rect 5520 4994 5880 5000
rect 5520 4966 5526 4994
rect 5554 4966 5686 4994
rect 5714 4966 5846 4994
rect 5874 4966 5880 4994
rect 5520 4960 5880 4966
rect 5920 4994 6120 5000
rect 5920 4966 5926 4994
rect 5954 4966 6086 4994
rect 6114 4966 6120 4994
rect 5920 4960 6120 4966
rect 6160 4994 6360 5000
rect 6160 4966 6166 4994
rect 6194 4966 6326 4994
rect 6354 4966 6360 4994
rect 6160 4960 6360 4966
rect 4240 4914 6360 4920
rect 4240 4886 5926 4914
rect 5954 4886 6086 4914
rect 6114 4886 6360 4914
rect 4240 4880 6360 4886
rect 4200 4834 6400 4840
rect 4200 4806 6006 4834
rect 6034 4806 6400 4834
rect 4200 4800 6400 4806
rect 4240 4754 6360 4760
rect 4240 4726 5926 4754
rect 5954 4726 6086 4754
rect 6114 4726 6360 4754
rect 4240 4720 6360 4726
rect 4240 4674 6360 4680
rect 4240 4646 6166 4674
rect 6194 4646 6326 4674
rect 6354 4646 6360 4674
rect 4240 4640 6360 4646
rect 4200 4594 6400 4600
rect 4200 4566 6246 4594
rect 6274 4566 6400 4594
rect 4200 4560 6400 4566
rect 4240 4514 6360 4520
rect 4240 4486 6166 4514
rect 6194 4486 6326 4514
rect 6354 4486 6360 4514
rect 4240 4480 6360 4486
rect 4240 4434 4440 4440
rect 4240 4406 4246 4434
rect 4274 4406 4406 4434
rect 4434 4406 4440 4434
rect 4240 4400 4440 4406
rect 4480 4434 4680 4440
rect 4480 4406 4486 4434
rect 4514 4406 4646 4434
rect 4674 4406 4680 4434
rect 4480 4400 4680 4406
rect 4720 4434 5080 4440
rect 4720 4406 4726 4434
rect 4754 4406 4886 4434
rect 4914 4406 5046 4434
rect 5074 4406 5080 4434
rect 4720 4400 5080 4406
rect 5120 4434 5480 4440
rect 5120 4406 5126 4434
rect 5154 4406 5286 4434
rect 5314 4406 5446 4434
rect 5474 4406 5480 4434
rect 5120 4400 5480 4406
rect 5520 4434 5880 4440
rect 5520 4406 5526 4434
rect 5554 4406 5686 4434
rect 5714 4406 5846 4434
rect 5874 4406 5880 4434
rect 5520 4400 5880 4406
rect 5920 4434 6120 4440
rect 5920 4406 5926 4434
rect 5954 4406 6086 4434
rect 6114 4406 6120 4434
rect 5920 4400 6120 4406
rect 6160 4434 6360 4440
rect 6160 4406 6166 4434
rect 6194 4406 6326 4434
rect 6354 4406 6360 4434
rect 6160 4400 6360 4406
rect 4240 4354 4440 4360
rect 4240 4326 4246 4354
rect 4274 4326 4406 4354
rect 4434 4326 4440 4354
rect 4240 4320 4440 4326
rect 4480 4354 4680 4360
rect 4480 4326 4486 4354
rect 4514 4326 4646 4354
rect 4674 4326 4680 4354
rect 4480 4320 4680 4326
rect 4720 4354 5080 4360
rect 4720 4326 4726 4354
rect 4754 4326 4886 4354
rect 4914 4326 5046 4354
rect 5074 4326 5080 4354
rect 4720 4320 5080 4326
rect 5120 4354 5480 4360
rect 5120 4326 5126 4354
rect 5154 4326 5286 4354
rect 5314 4326 5446 4354
rect 5474 4326 5480 4354
rect 5120 4320 5480 4326
rect 5520 4354 5880 4360
rect 5520 4326 5526 4354
rect 5554 4326 5686 4354
rect 5714 4326 5846 4354
rect 5874 4326 5880 4354
rect 5520 4320 5880 4326
rect 5920 4354 6120 4360
rect 5920 4326 5926 4354
rect 5954 4326 6086 4354
rect 6114 4326 6120 4354
rect 5920 4320 6120 4326
rect 6160 4354 6360 4360
rect 6160 4326 6166 4354
rect 6194 4326 6326 4354
rect 6354 4326 6360 4354
rect 6160 4320 6360 4326
rect 4240 4274 4440 4280
rect 4240 4246 4246 4274
rect 4274 4246 4406 4274
rect 4434 4246 4440 4274
rect 4240 4240 4440 4246
rect 4480 4274 4680 4280
rect 4480 4246 4486 4274
rect 4514 4246 4646 4274
rect 4674 4246 4680 4274
rect 4480 4240 4680 4246
rect 4720 4274 5080 4280
rect 4720 4246 4726 4274
rect 4754 4246 4886 4274
rect 4914 4246 5046 4274
rect 5074 4246 5080 4274
rect 4720 4240 5080 4246
rect 5120 4274 5480 4280
rect 5120 4246 5126 4274
rect 5154 4246 5286 4274
rect 5314 4246 5446 4274
rect 5474 4246 5480 4274
rect 5120 4240 5480 4246
rect 5520 4274 5880 4280
rect 5520 4246 5526 4274
rect 5554 4246 5686 4274
rect 5714 4246 5846 4274
rect 5874 4246 5880 4274
rect 5520 4240 5880 4246
rect 5920 4274 6120 4280
rect 5920 4246 5926 4274
rect 5954 4246 6086 4274
rect 6114 4246 6120 4274
rect 5920 4240 6120 4246
rect 6160 4274 6360 4280
rect 6160 4246 6166 4274
rect 6194 4246 6326 4274
rect 6354 4246 6360 4274
rect 6160 4240 6360 4246
rect 4240 4194 4440 4200
rect 4240 4166 4246 4194
rect 4274 4166 4406 4194
rect 4434 4166 4440 4194
rect 4240 4160 4440 4166
rect 4480 4194 4680 4200
rect 4480 4166 4486 4194
rect 4514 4166 4646 4194
rect 4674 4166 4680 4194
rect 4480 4160 4680 4166
rect 4720 4194 5080 4200
rect 4720 4166 4726 4194
rect 4754 4166 4886 4194
rect 4914 4166 5046 4194
rect 5074 4166 5080 4194
rect 4720 4160 5080 4166
rect 5120 4194 5480 4200
rect 5120 4166 5126 4194
rect 5154 4166 5286 4194
rect 5314 4166 5446 4194
rect 5474 4166 5480 4194
rect 5120 4160 5480 4166
rect 5520 4194 5880 4200
rect 5520 4166 5526 4194
rect 5554 4166 5686 4194
rect 5714 4166 5846 4194
rect 5874 4166 5880 4194
rect 5520 4160 5880 4166
rect 5920 4194 6120 4200
rect 5920 4166 5926 4194
rect 5954 4166 6086 4194
rect 6114 4166 6120 4194
rect 5920 4160 6120 4166
rect 6160 4194 6360 4200
rect 6160 4166 6166 4194
rect 6194 4166 6326 4194
rect 6354 4166 6360 4194
rect 6160 4160 6360 4166
rect 4240 4114 4440 4120
rect 4240 4086 4246 4114
rect 4274 4086 4406 4114
rect 4434 4086 4440 4114
rect 4240 4080 4440 4086
rect 4480 4114 4680 4120
rect 4480 4086 4486 4114
rect 4514 4086 4646 4114
rect 4674 4086 4680 4114
rect 4480 4080 4680 4086
rect 4720 4114 5080 4120
rect 4720 4086 4726 4114
rect 4754 4086 4886 4114
rect 4914 4086 5046 4114
rect 5074 4086 5080 4114
rect 4720 4080 5080 4086
rect 5120 4114 5480 4120
rect 5120 4086 5126 4114
rect 5154 4086 5286 4114
rect 5314 4086 5446 4114
rect 5474 4086 5480 4114
rect 5120 4080 5480 4086
rect 5520 4114 5880 4120
rect 5520 4086 5526 4114
rect 5554 4086 5686 4114
rect 5714 4086 5846 4114
rect 5874 4086 5880 4114
rect 5520 4080 5880 4086
rect 5920 4114 6120 4120
rect 5920 4086 5926 4114
rect 5954 4086 6086 4114
rect 6114 4086 6120 4114
rect 5920 4080 6120 4086
rect 6160 4114 6360 4120
rect 6160 4086 6166 4114
rect 6194 4086 6326 4114
rect 6354 4086 6360 4114
rect 6160 4080 6360 4086
rect 4240 4034 4440 4040
rect 4240 4006 4246 4034
rect 4274 4006 4406 4034
rect 4434 4006 4440 4034
rect 4240 4000 4440 4006
rect 4480 4034 4680 4040
rect 4480 4006 4486 4034
rect 4514 4006 4646 4034
rect 4674 4006 4680 4034
rect 4480 4000 4680 4006
rect 4720 4034 5080 4040
rect 4720 4006 4726 4034
rect 4754 4006 4886 4034
rect 4914 4006 5046 4034
rect 5074 4006 5080 4034
rect 4720 4000 5080 4006
rect 5120 4034 5480 4040
rect 5120 4006 5126 4034
rect 5154 4006 5286 4034
rect 5314 4006 5446 4034
rect 5474 4006 5480 4034
rect 5120 4000 5480 4006
rect 5520 4034 5880 4040
rect 5520 4006 5526 4034
rect 5554 4006 5686 4034
rect 5714 4006 5846 4034
rect 5874 4006 5880 4034
rect 5520 4000 5880 4006
rect 5920 4034 6120 4040
rect 5920 4006 5926 4034
rect 5954 4006 6086 4034
rect 6114 4006 6120 4034
rect 5920 4000 6120 4006
rect 6160 4034 6360 4040
rect 6160 4006 6166 4034
rect 6194 4006 6326 4034
rect 6354 4006 6360 4034
rect 6160 4000 6360 4006
rect 4240 3954 4440 3960
rect 4240 3926 4246 3954
rect 4274 3926 4406 3954
rect 4434 3926 4440 3954
rect 4240 3920 4440 3926
rect 4480 3954 4680 3960
rect 4480 3926 4486 3954
rect 4514 3926 4646 3954
rect 4674 3926 4680 3954
rect 4480 3920 4680 3926
rect 4720 3954 5080 3960
rect 4720 3926 4726 3954
rect 4754 3926 4886 3954
rect 4914 3926 5046 3954
rect 5074 3926 5080 3954
rect 4720 3920 5080 3926
rect 5120 3954 5480 3960
rect 5120 3926 5126 3954
rect 5154 3926 5286 3954
rect 5314 3926 5446 3954
rect 5474 3926 5480 3954
rect 5120 3920 5480 3926
rect 5520 3954 5880 3960
rect 5520 3926 5526 3954
rect 5554 3926 5686 3954
rect 5714 3926 5846 3954
rect 5874 3926 5880 3954
rect 5520 3920 5880 3926
rect 5920 3954 6120 3960
rect 5920 3926 5926 3954
rect 5954 3926 6086 3954
rect 6114 3926 6120 3954
rect 5920 3920 6120 3926
rect 6160 3954 6360 3960
rect 6160 3926 6166 3954
rect 6194 3926 6326 3954
rect 6354 3926 6360 3954
rect 6160 3920 6360 3926
rect 4240 3874 6360 3880
rect 4240 3846 4246 3874
rect 4274 3846 4406 3874
rect 4434 3846 6360 3874
rect 4240 3840 6360 3846
rect 4200 3794 6400 3800
rect 4200 3766 4326 3794
rect 4354 3766 6400 3794
rect 4200 3760 6400 3766
rect 4240 3714 6360 3720
rect 4240 3686 4246 3714
rect 4274 3686 4406 3714
rect 4434 3686 6360 3714
rect 4240 3680 6360 3686
rect 4240 3634 6360 3640
rect 4240 3606 4486 3634
rect 4514 3606 4646 3634
rect 4674 3606 6360 3634
rect 4240 3600 6360 3606
rect 4200 3554 6400 3560
rect 4200 3526 4566 3554
rect 4594 3526 6400 3554
rect 4200 3520 6400 3526
rect 4240 3474 6360 3480
rect 4240 3446 4486 3474
rect 4514 3446 4646 3474
rect 4674 3446 6360 3474
rect 4240 3440 6360 3446
rect 4240 3394 6360 3400
rect 4240 3366 5926 3394
rect 5954 3366 6086 3394
rect 6114 3366 6360 3394
rect 4240 3360 6360 3366
rect 4200 3314 6400 3320
rect 4200 3286 6006 3314
rect 6034 3286 6400 3314
rect 4200 3280 6400 3286
rect 4240 3234 6360 3240
rect 4240 3206 5926 3234
rect 5954 3206 6086 3234
rect 6114 3206 6360 3234
rect 4240 3200 6360 3206
rect 4240 3154 4440 3160
rect 4240 3126 4246 3154
rect 4274 3126 4406 3154
rect 4434 3126 4440 3154
rect 4240 3120 4440 3126
rect 4480 3154 4680 3160
rect 4480 3126 4486 3154
rect 4514 3126 4646 3154
rect 4674 3126 4680 3154
rect 4480 3120 4680 3126
rect 4720 3154 5080 3160
rect 4720 3126 4726 3154
rect 4754 3126 4886 3154
rect 4914 3126 5046 3154
rect 5074 3126 5080 3154
rect 4720 3120 5080 3126
rect 5120 3154 5480 3160
rect 5120 3126 5126 3154
rect 5154 3126 5286 3154
rect 5314 3126 5446 3154
rect 5474 3126 5480 3154
rect 5120 3120 5480 3126
rect 5520 3154 5880 3160
rect 5520 3126 5526 3154
rect 5554 3126 5686 3154
rect 5714 3126 5846 3154
rect 5874 3126 5880 3154
rect 5520 3120 5880 3126
rect 5920 3154 6120 3160
rect 5920 3126 5926 3154
rect 5954 3126 6086 3154
rect 6114 3126 6120 3154
rect 5920 3120 6120 3126
rect 6160 3154 6360 3160
rect 6160 3126 6166 3154
rect 6194 3126 6326 3154
rect 6354 3126 6360 3154
rect 6160 3120 6360 3126
rect 4240 3074 4440 3080
rect 4240 3046 4246 3074
rect 4274 3046 4406 3074
rect 4434 3046 4440 3074
rect 4240 3040 4440 3046
rect 4480 3074 4680 3080
rect 4480 3046 4486 3074
rect 4514 3046 4646 3074
rect 4674 3046 4680 3074
rect 4480 3040 4680 3046
rect 4720 3074 5080 3080
rect 4720 3046 4726 3074
rect 4754 3046 4886 3074
rect 4914 3046 5046 3074
rect 5074 3046 5080 3074
rect 4720 3040 5080 3046
rect 5120 3074 5480 3080
rect 5120 3046 5126 3074
rect 5154 3046 5286 3074
rect 5314 3046 5446 3074
rect 5474 3046 5480 3074
rect 5120 3040 5480 3046
rect 5520 3074 5880 3080
rect 5520 3046 5526 3074
rect 5554 3046 5686 3074
rect 5714 3046 5846 3074
rect 5874 3046 5880 3074
rect 5520 3040 5880 3046
rect 5920 3074 6120 3080
rect 5920 3046 5926 3074
rect 5954 3046 6086 3074
rect 6114 3046 6120 3074
rect 5920 3040 6120 3046
rect 6160 3074 6360 3080
rect 6160 3046 6166 3074
rect 6194 3046 6326 3074
rect 6354 3046 6360 3074
rect 6160 3040 6360 3046
rect 4240 2994 4440 3000
rect 4240 2966 4246 2994
rect 4274 2966 4406 2994
rect 4434 2966 4440 2994
rect 4240 2960 4440 2966
rect 4480 2994 4680 3000
rect 4480 2966 4486 2994
rect 4514 2966 4646 2994
rect 4674 2966 4680 2994
rect 4480 2960 4680 2966
rect 4720 2994 5080 3000
rect 4720 2966 4726 2994
rect 4754 2966 4886 2994
rect 4914 2966 5046 2994
rect 5074 2966 5080 2994
rect 4720 2960 5080 2966
rect 5120 2994 5480 3000
rect 5120 2966 5126 2994
rect 5154 2966 5286 2994
rect 5314 2966 5446 2994
rect 5474 2966 5480 2994
rect 5120 2960 5480 2966
rect 5520 2994 5880 3000
rect 5520 2966 5526 2994
rect 5554 2966 5686 2994
rect 5714 2966 5846 2994
rect 5874 2966 5880 2994
rect 5520 2960 5880 2966
rect 5920 2994 6120 3000
rect 5920 2966 5926 2994
rect 5954 2966 6086 2994
rect 6114 2966 6120 2994
rect 5920 2960 6120 2966
rect 6160 2994 6360 3000
rect 6160 2966 6166 2994
rect 6194 2966 6326 2994
rect 6354 2966 6360 2994
rect 6160 2960 6360 2966
rect 4240 2914 4440 2920
rect 4240 2886 4246 2914
rect 4274 2886 4406 2914
rect 4434 2886 4440 2914
rect 4240 2880 4440 2886
rect 4480 2914 4680 2920
rect 4480 2886 4486 2914
rect 4514 2886 4646 2914
rect 4674 2886 4680 2914
rect 4480 2880 4680 2886
rect 4720 2914 5080 2920
rect 4720 2886 4726 2914
rect 4754 2886 4886 2914
rect 4914 2886 5046 2914
rect 5074 2886 5080 2914
rect 4720 2880 5080 2886
rect 5120 2914 5480 2920
rect 5120 2886 5126 2914
rect 5154 2886 5286 2914
rect 5314 2886 5446 2914
rect 5474 2886 5480 2914
rect 5120 2880 5480 2886
rect 5520 2914 5880 2920
rect 5520 2886 5526 2914
rect 5554 2886 5686 2914
rect 5714 2886 5846 2914
rect 5874 2886 5880 2914
rect 5520 2880 5880 2886
rect 5920 2914 6120 2920
rect 5920 2886 5926 2914
rect 5954 2886 6086 2914
rect 6114 2886 6120 2914
rect 5920 2880 6120 2886
rect 6160 2914 6360 2920
rect 6160 2886 6166 2914
rect 6194 2886 6326 2914
rect 6354 2886 6360 2914
rect 6160 2880 6360 2886
rect 4240 2834 4440 2840
rect 4240 2806 4246 2834
rect 4274 2806 4406 2834
rect 4434 2806 4440 2834
rect 4240 2800 4440 2806
rect 4480 2834 4680 2840
rect 4480 2806 4486 2834
rect 4514 2806 4646 2834
rect 4674 2806 4680 2834
rect 4480 2800 4680 2806
rect 4720 2834 5080 2840
rect 4720 2806 4726 2834
rect 4754 2806 4886 2834
rect 4914 2806 5046 2834
rect 5074 2806 5080 2834
rect 4720 2800 5080 2806
rect 5120 2834 5480 2840
rect 5120 2806 5126 2834
rect 5154 2806 5286 2834
rect 5314 2806 5446 2834
rect 5474 2806 5480 2834
rect 5120 2800 5480 2806
rect 5520 2834 5880 2840
rect 5520 2806 5526 2834
rect 5554 2806 5686 2834
rect 5714 2806 5846 2834
rect 5874 2806 5880 2834
rect 5520 2800 5880 2806
rect 5920 2834 6120 2840
rect 5920 2806 5926 2834
rect 5954 2806 6086 2834
rect 6114 2806 6120 2834
rect 5920 2800 6120 2806
rect 6160 2834 6360 2840
rect 6160 2806 6166 2834
rect 6194 2806 6326 2834
rect 6354 2806 6360 2834
rect 6160 2800 6360 2806
rect 4240 2754 4440 2760
rect 4240 2726 4246 2754
rect 4274 2726 4406 2754
rect 4434 2726 4440 2754
rect 4240 2720 4440 2726
rect 4480 2754 4680 2760
rect 4480 2726 4486 2754
rect 4514 2726 4646 2754
rect 4674 2726 4680 2754
rect 4480 2720 4680 2726
rect 4720 2754 5080 2760
rect 4720 2726 4726 2754
rect 4754 2726 4886 2754
rect 4914 2726 5046 2754
rect 5074 2726 5080 2754
rect 4720 2720 5080 2726
rect 5120 2754 5480 2760
rect 5120 2726 5126 2754
rect 5154 2726 5286 2754
rect 5314 2726 5446 2754
rect 5474 2726 5480 2754
rect 5120 2720 5480 2726
rect 5520 2754 5880 2760
rect 5520 2726 5526 2754
rect 5554 2726 5686 2754
rect 5714 2726 5846 2754
rect 5874 2726 5880 2754
rect 5520 2720 5880 2726
rect 5920 2754 6120 2760
rect 5920 2726 5926 2754
rect 5954 2726 6086 2754
rect 6114 2726 6120 2754
rect 5920 2720 6120 2726
rect 6160 2754 6360 2760
rect 6160 2726 6166 2754
rect 6194 2726 6326 2754
rect 6354 2726 6360 2754
rect 6160 2720 6360 2726
rect 4240 2674 4440 2680
rect 4240 2646 4246 2674
rect 4274 2646 4406 2674
rect 4434 2646 4440 2674
rect 4240 2640 4440 2646
rect 4480 2674 4680 2680
rect 4480 2646 4486 2674
rect 4514 2646 4646 2674
rect 4674 2646 4680 2674
rect 4480 2640 4680 2646
rect 4720 2674 5080 2680
rect 4720 2646 4726 2674
rect 4754 2646 4886 2674
rect 4914 2646 5046 2674
rect 5074 2646 5080 2674
rect 4720 2640 5080 2646
rect 5120 2674 5480 2680
rect 5120 2646 5126 2674
rect 5154 2646 5286 2674
rect 5314 2646 5446 2674
rect 5474 2646 5480 2674
rect 5120 2640 5480 2646
rect 5520 2674 5880 2680
rect 5520 2646 5526 2674
rect 5554 2646 5686 2674
rect 5714 2646 5846 2674
rect 5874 2646 5880 2674
rect 5520 2640 5880 2646
rect 5920 2674 6120 2680
rect 5920 2646 5926 2674
rect 5954 2646 6086 2674
rect 6114 2646 6120 2674
rect 5920 2640 6120 2646
rect 6160 2674 6360 2680
rect 6160 2646 6166 2674
rect 6194 2646 6326 2674
rect 6354 2646 6360 2674
rect 6160 2640 6360 2646
rect 4240 2594 4440 2600
rect 4240 2566 4246 2594
rect 4274 2566 4406 2594
rect 4434 2566 4440 2594
rect 4240 2560 4440 2566
rect 4480 2594 4680 2600
rect 4480 2566 4486 2594
rect 4514 2566 4646 2594
rect 4674 2566 4680 2594
rect 4480 2560 4680 2566
rect 4720 2594 5080 2600
rect 4720 2566 4726 2594
rect 4754 2566 4886 2594
rect 4914 2566 5046 2594
rect 5074 2566 5080 2594
rect 4720 2560 5080 2566
rect 5120 2594 5480 2600
rect 5120 2566 5126 2594
rect 5154 2566 5286 2594
rect 5314 2566 5446 2594
rect 5474 2566 5480 2594
rect 5120 2560 5480 2566
rect 5520 2594 5880 2600
rect 5520 2566 5526 2594
rect 5554 2566 5686 2594
rect 5714 2566 5846 2594
rect 5874 2566 5880 2594
rect 5520 2560 5880 2566
rect 5920 2594 6120 2600
rect 5920 2566 5926 2594
rect 5954 2566 6086 2594
rect 6114 2566 6120 2594
rect 5920 2560 6120 2566
rect 6160 2594 6360 2600
rect 6160 2566 6166 2594
rect 6194 2566 6326 2594
rect 6354 2566 6360 2594
rect 6160 2560 6360 2566
rect 4240 2514 4440 2520
rect 4240 2486 4246 2514
rect 4274 2486 4406 2514
rect 4434 2486 4440 2514
rect 4240 2480 4440 2486
rect 4480 2514 4680 2520
rect 4480 2486 4486 2514
rect 4514 2486 4646 2514
rect 4674 2486 4680 2514
rect 4480 2480 4680 2486
rect 4720 2514 5080 2520
rect 4720 2486 4726 2514
rect 4754 2486 4886 2514
rect 4914 2486 5046 2514
rect 5074 2486 5080 2514
rect 4720 2480 5080 2486
rect 5120 2514 5480 2520
rect 5120 2486 5126 2514
rect 5154 2486 5286 2514
rect 5314 2486 5446 2514
rect 5474 2486 5480 2514
rect 5120 2480 5480 2486
rect 5520 2514 5880 2520
rect 5520 2486 5526 2514
rect 5554 2486 5686 2514
rect 5714 2486 5846 2514
rect 5874 2486 5880 2514
rect 5520 2480 5880 2486
rect 5920 2514 6120 2520
rect 5920 2486 5926 2514
rect 5954 2486 6086 2514
rect 6114 2486 6120 2514
rect 5920 2480 6120 2486
rect 6160 2514 6360 2520
rect 6160 2486 6166 2514
rect 6194 2486 6326 2514
rect 6354 2486 6360 2514
rect 6160 2480 6360 2486
rect 4240 2434 4440 2440
rect 4240 2406 4246 2434
rect 4274 2406 4406 2434
rect 4434 2406 4440 2434
rect 4240 2400 4440 2406
rect 4480 2434 4680 2440
rect 4480 2406 4486 2434
rect 4514 2406 4646 2434
rect 4674 2406 4680 2434
rect 4480 2400 4680 2406
rect 4720 2434 5080 2440
rect 4720 2406 4726 2434
rect 4754 2406 4886 2434
rect 4914 2406 5046 2434
rect 5074 2406 5080 2434
rect 4720 2400 5080 2406
rect 5120 2434 5480 2440
rect 5120 2406 5126 2434
rect 5154 2406 5286 2434
rect 5314 2406 5446 2434
rect 5474 2406 5480 2434
rect 5120 2400 5480 2406
rect 5520 2434 5880 2440
rect 5520 2406 5526 2434
rect 5554 2406 5686 2434
rect 5714 2406 5846 2434
rect 5874 2406 5880 2434
rect 5520 2400 5880 2406
rect 5920 2434 6120 2440
rect 5920 2406 5926 2434
rect 5954 2406 6086 2434
rect 6114 2406 6120 2434
rect 5920 2400 6120 2406
rect 6160 2434 6360 2440
rect 6160 2406 6166 2434
rect 6194 2406 6326 2434
rect 6354 2406 6360 2434
rect 6160 2400 6360 2406
rect 4240 2354 4440 2360
rect 4240 2326 4246 2354
rect 4274 2326 4406 2354
rect 4434 2326 4440 2354
rect 4240 2320 4440 2326
rect 4480 2354 4680 2360
rect 4480 2326 4486 2354
rect 4514 2326 4646 2354
rect 4674 2326 4680 2354
rect 4480 2320 4680 2326
rect 4720 2354 5080 2360
rect 4720 2326 4726 2354
rect 4754 2326 4886 2354
rect 4914 2326 5046 2354
rect 5074 2326 5080 2354
rect 4720 2320 5080 2326
rect 5120 2354 5480 2360
rect 5120 2326 5126 2354
rect 5154 2326 5286 2354
rect 5314 2326 5446 2354
rect 5474 2326 5480 2354
rect 5120 2320 5480 2326
rect 5520 2354 5880 2360
rect 5520 2326 5526 2354
rect 5554 2326 5686 2354
rect 5714 2326 5846 2354
rect 5874 2326 5880 2354
rect 5520 2320 5880 2326
rect 5920 2354 6120 2360
rect 5920 2326 5926 2354
rect 5954 2326 6086 2354
rect 6114 2326 6120 2354
rect 5920 2320 6120 2326
rect 6160 2354 6360 2360
rect 6160 2326 6166 2354
rect 6194 2326 6326 2354
rect 6354 2326 6360 2354
rect 6160 2320 6360 2326
rect 4240 2274 4440 2280
rect 4240 2246 4246 2274
rect 4274 2246 4406 2274
rect 4434 2246 4440 2274
rect 4240 2240 4440 2246
rect 4480 2274 4680 2280
rect 4480 2246 4486 2274
rect 4514 2246 4646 2274
rect 4674 2246 4680 2274
rect 4480 2240 4680 2246
rect 4720 2274 5080 2280
rect 4720 2246 4726 2274
rect 4754 2246 4886 2274
rect 4914 2246 5046 2274
rect 5074 2246 5080 2274
rect 4720 2240 5080 2246
rect 5120 2274 5480 2280
rect 5120 2246 5126 2274
rect 5154 2246 5286 2274
rect 5314 2246 5446 2274
rect 5474 2246 5480 2274
rect 5120 2240 5480 2246
rect 5520 2274 5880 2280
rect 5520 2246 5526 2274
rect 5554 2246 5686 2274
rect 5714 2246 5846 2274
rect 5874 2246 5880 2274
rect 5520 2240 5880 2246
rect 5920 2274 6120 2280
rect 5920 2246 5926 2274
rect 5954 2246 6086 2274
rect 6114 2246 6120 2274
rect 5920 2240 6120 2246
rect 6160 2274 6360 2280
rect 6160 2246 6166 2274
rect 6194 2246 6326 2274
rect 6354 2246 6360 2274
rect 6160 2240 6360 2246
rect 4240 2194 4440 2200
rect 4240 2166 4246 2194
rect 4274 2166 4406 2194
rect 4434 2166 4440 2194
rect 4240 2160 4440 2166
rect 4480 2194 4680 2200
rect 4480 2166 4486 2194
rect 4514 2166 4646 2194
rect 4674 2166 4680 2194
rect 4480 2160 4680 2166
rect 4720 2194 5080 2200
rect 4720 2166 4726 2194
rect 4754 2166 4886 2194
rect 4914 2166 5046 2194
rect 5074 2166 5080 2194
rect 4720 2160 5080 2166
rect 5120 2194 5480 2200
rect 5120 2166 5126 2194
rect 5154 2166 5286 2194
rect 5314 2166 5446 2194
rect 5474 2166 5480 2194
rect 5120 2160 5480 2166
rect 5520 2194 5880 2200
rect 5520 2166 5526 2194
rect 5554 2166 5686 2194
rect 5714 2166 5846 2194
rect 5874 2166 5880 2194
rect 5520 2160 5880 2166
rect 5920 2194 6120 2200
rect 5920 2166 5926 2194
rect 5954 2166 6086 2194
rect 6114 2166 6120 2194
rect 5920 2160 6120 2166
rect 6160 2194 6360 2200
rect 6160 2166 6166 2194
rect 6194 2166 6326 2194
rect 6354 2166 6360 2194
rect 6160 2160 6360 2166
rect 4240 2114 4440 2120
rect 4240 2086 4246 2114
rect 4274 2086 4406 2114
rect 4434 2086 4440 2114
rect 4240 2080 4440 2086
rect 4480 2114 4680 2120
rect 4480 2086 4486 2114
rect 4514 2086 4646 2114
rect 4674 2086 4680 2114
rect 4480 2080 4680 2086
rect 4720 2114 5080 2120
rect 4720 2086 4726 2114
rect 4754 2086 4886 2114
rect 4914 2086 5046 2114
rect 5074 2086 5080 2114
rect 4720 2080 5080 2086
rect 5120 2114 5480 2120
rect 5120 2086 5126 2114
rect 5154 2086 5286 2114
rect 5314 2086 5446 2114
rect 5474 2086 5480 2114
rect 5120 2080 5480 2086
rect 5520 2114 5880 2120
rect 5520 2086 5526 2114
rect 5554 2086 5686 2114
rect 5714 2086 5846 2114
rect 5874 2086 5880 2114
rect 5520 2080 5880 2086
rect 5920 2114 6120 2120
rect 5920 2086 5926 2114
rect 5954 2086 6086 2114
rect 6114 2086 6120 2114
rect 5920 2080 6120 2086
rect 6160 2114 6360 2120
rect 6160 2086 6166 2114
rect 6194 2086 6326 2114
rect 6354 2086 6360 2114
rect 6160 2080 6360 2086
rect 4240 2034 4440 2040
rect 4240 2006 4246 2034
rect 4274 2006 4406 2034
rect 4434 2006 4440 2034
rect 4240 2000 4440 2006
rect 4480 2034 4680 2040
rect 4480 2006 4486 2034
rect 4514 2006 4646 2034
rect 4674 2006 4680 2034
rect 4480 2000 4680 2006
rect 4720 2034 5080 2040
rect 4720 2006 4726 2034
rect 4754 2006 4886 2034
rect 4914 2006 5046 2034
rect 5074 2006 5080 2034
rect 4720 2000 5080 2006
rect 5120 2034 5480 2040
rect 5120 2006 5126 2034
rect 5154 2006 5286 2034
rect 5314 2006 5446 2034
rect 5474 2006 5480 2034
rect 5120 2000 5480 2006
rect 5520 2034 5880 2040
rect 5520 2006 5526 2034
rect 5554 2006 5686 2034
rect 5714 2006 5846 2034
rect 5874 2006 5880 2034
rect 5520 2000 5880 2006
rect 5920 2034 6120 2040
rect 5920 2006 5926 2034
rect 5954 2006 6086 2034
rect 6114 2006 6120 2034
rect 5920 2000 6120 2006
rect 6160 2034 6360 2040
rect 6160 2006 6166 2034
rect 6194 2006 6326 2034
rect 6354 2006 6360 2034
rect 6160 2000 6360 2006
rect 4240 1914 6360 1920
rect 4240 1886 4486 1914
rect 4514 1886 4646 1914
rect 4674 1886 6360 1914
rect 4240 1880 6360 1886
rect 4200 1834 6400 1840
rect 4200 1806 4566 1834
rect 4594 1806 6400 1834
rect 4200 1800 6400 1806
rect 4240 1754 6360 1760
rect 4240 1726 4486 1754
rect 4514 1726 4646 1754
rect 4674 1726 6360 1754
rect 4240 1720 6360 1726
rect 4240 1634 4440 1640
rect 4240 1606 4246 1634
rect 4274 1606 4406 1634
rect 4434 1606 4440 1634
rect 4240 1600 4440 1606
rect 4480 1634 4680 1640
rect 4480 1606 4486 1634
rect 4514 1606 4646 1634
rect 4674 1606 4680 1634
rect 4480 1600 4680 1606
rect 4720 1634 5080 1640
rect 4720 1606 4726 1634
rect 4754 1606 4886 1634
rect 4914 1606 5046 1634
rect 5074 1606 5080 1634
rect 4720 1600 5080 1606
rect 5120 1634 5480 1640
rect 5120 1606 5126 1634
rect 5154 1606 5286 1634
rect 5314 1606 5446 1634
rect 5474 1606 5480 1634
rect 5120 1600 5480 1606
rect 5520 1634 5880 1640
rect 5520 1606 5526 1634
rect 5554 1606 5686 1634
rect 5714 1606 5846 1634
rect 5874 1606 5880 1634
rect 5520 1600 5880 1606
rect 5920 1634 6120 1640
rect 5920 1606 5926 1634
rect 5954 1606 6086 1634
rect 6114 1606 6120 1634
rect 5920 1600 6120 1606
rect 6160 1634 6360 1640
rect 6160 1606 6166 1634
rect 6194 1606 6326 1634
rect 6354 1606 6360 1634
rect 6160 1600 6360 1606
rect 4240 1554 4440 1560
rect 4240 1526 4246 1554
rect 4274 1526 4406 1554
rect 4434 1526 4440 1554
rect 4240 1520 4440 1526
rect 4480 1554 4680 1560
rect 4480 1526 4486 1554
rect 4514 1526 4646 1554
rect 4674 1526 4680 1554
rect 4480 1520 4680 1526
rect 4720 1554 5080 1560
rect 4720 1526 4726 1554
rect 4754 1526 4886 1554
rect 4914 1526 5046 1554
rect 5074 1526 5080 1554
rect 4720 1520 5080 1526
rect 5120 1554 5480 1560
rect 5120 1526 5126 1554
rect 5154 1526 5286 1554
rect 5314 1526 5446 1554
rect 5474 1526 5480 1554
rect 5120 1520 5480 1526
rect 5520 1554 5880 1560
rect 5520 1526 5526 1554
rect 5554 1526 5686 1554
rect 5714 1526 5846 1554
rect 5874 1526 5880 1554
rect 5520 1520 5880 1526
rect 5920 1554 6120 1560
rect 5920 1526 5926 1554
rect 5954 1526 6086 1554
rect 6114 1526 6120 1554
rect 5920 1520 6120 1526
rect 6160 1554 6360 1560
rect 6160 1526 6166 1554
rect 6194 1526 6326 1554
rect 6354 1526 6360 1554
rect 6160 1520 6360 1526
rect 4240 1474 4440 1480
rect 4240 1446 4246 1474
rect 4274 1446 4406 1474
rect 4434 1446 4440 1474
rect 4240 1440 4440 1446
rect 4480 1474 4680 1480
rect 4480 1446 4486 1474
rect 4514 1446 4646 1474
rect 4674 1446 4680 1474
rect 4480 1440 4680 1446
rect 4720 1474 5080 1480
rect 4720 1446 4726 1474
rect 4754 1446 4886 1474
rect 4914 1446 5046 1474
rect 5074 1446 5080 1474
rect 4720 1440 5080 1446
rect 5120 1474 5480 1480
rect 5120 1446 5126 1474
rect 5154 1446 5286 1474
rect 5314 1446 5446 1474
rect 5474 1446 5480 1474
rect 5120 1440 5480 1446
rect 5520 1474 5880 1480
rect 5520 1446 5526 1474
rect 5554 1446 5686 1474
rect 5714 1446 5846 1474
rect 5874 1446 5880 1474
rect 5520 1440 5880 1446
rect 5920 1474 6120 1480
rect 5920 1446 5926 1474
rect 5954 1446 6086 1474
rect 6114 1446 6120 1474
rect 5920 1440 6120 1446
rect 6160 1474 6360 1480
rect 6160 1446 6166 1474
rect 6194 1446 6326 1474
rect 6354 1446 6360 1474
rect 6160 1440 6360 1446
rect 4240 1394 4440 1400
rect 4240 1366 4246 1394
rect 4274 1366 4406 1394
rect 4434 1366 4440 1394
rect 4240 1360 4440 1366
rect 4480 1394 4680 1400
rect 4480 1366 4486 1394
rect 4514 1366 4646 1394
rect 4674 1366 4680 1394
rect 4480 1360 4680 1366
rect 4720 1394 5080 1400
rect 4720 1366 4726 1394
rect 4754 1366 4886 1394
rect 4914 1366 5046 1394
rect 5074 1366 5080 1394
rect 4720 1360 5080 1366
rect 5120 1394 5480 1400
rect 5120 1366 5126 1394
rect 5154 1366 5286 1394
rect 5314 1366 5446 1394
rect 5474 1366 5480 1394
rect 5120 1360 5480 1366
rect 5520 1394 5880 1400
rect 5520 1366 5526 1394
rect 5554 1366 5686 1394
rect 5714 1366 5846 1394
rect 5874 1366 5880 1394
rect 5520 1360 5880 1366
rect 5920 1394 6120 1400
rect 5920 1366 5926 1394
rect 5954 1366 6086 1394
rect 6114 1366 6120 1394
rect 5920 1360 6120 1366
rect 6160 1394 6360 1400
rect 6160 1366 6166 1394
rect 6194 1366 6326 1394
rect 6354 1366 6360 1394
rect 6160 1360 6360 1366
rect 4240 1314 4440 1320
rect 4240 1286 4246 1314
rect 4274 1286 4406 1314
rect 4434 1286 4440 1314
rect 4240 1280 4440 1286
rect 4480 1314 4680 1320
rect 4480 1286 4486 1314
rect 4514 1286 4646 1314
rect 4674 1286 4680 1314
rect 4480 1280 4680 1286
rect 4720 1314 5080 1320
rect 4720 1286 4726 1314
rect 4754 1286 4886 1314
rect 4914 1286 5046 1314
rect 5074 1286 5080 1314
rect 4720 1280 5080 1286
rect 5120 1314 5480 1320
rect 5120 1286 5126 1314
rect 5154 1286 5286 1314
rect 5314 1286 5446 1314
rect 5474 1286 5480 1314
rect 5120 1280 5480 1286
rect 5520 1314 5880 1320
rect 5520 1286 5526 1314
rect 5554 1286 5686 1314
rect 5714 1286 5846 1314
rect 5874 1286 5880 1314
rect 5520 1280 5880 1286
rect 5920 1314 6120 1320
rect 5920 1286 5926 1314
rect 5954 1286 6086 1314
rect 6114 1286 6120 1314
rect 5920 1280 6120 1286
rect 6160 1314 6360 1320
rect 6160 1286 6166 1314
rect 6194 1286 6326 1314
rect 6354 1286 6360 1314
rect 6160 1280 6360 1286
rect 4240 1234 4440 1240
rect 4240 1206 4246 1234
rect 4274 1206 4406 1234
rect 4434 1206 4440 1234
rect 4240 1200 4440 1206
rect 4480 1234 4680 1240
rect 4480 1206 4486 1234
rect 4514 1206 4646 1234
rect 4674 1206 4680 1234
rect 4480 1200 4680 1206
rect 4720 1234 5080 1240
rect 4720 1206 4726 1234
rect 4754 1206 4886 1234
rect 4914 1206 5046 1234
rect 5074 1206 5080 1234
rect 4720 1200 5080 1206
rect 5120 1234 5480 1240
rect 5120 1206 5126 1234
rect 5154 1206 5286 1234
rect 5314 1206 5446 1234
rect 5474 1206 5480 1234
rect 5120 1200 5480 1206
rect 5520 1234 5880 1240
rect 5520 1206 5526 1234
rect 5554 1206 5686 1234
rect 5714 1206 5846 1234
rect 5874 1206 5880 1234
rect 5520 1200 5880 1206
rect 5920 1234 6120 1240
rect 5920 1206 5926 1234
rect 5954 1206 6086 1234
rect 6114 1206 6120 1234
rect 5920 1200 6120 1206
rect 6160 1234 6360 1240
rect 6160 1206 6166 1234
rect 6194 1206 6326 1234
rect 6354 1206 6360 1234
rect 6160 1200 6360 1206
rect 4240 1154 4440 1160
rect 4240 1126 4246 1154
rect 4274 1126 4406 1154
rect 4434 1126 4440 1154
rect 4240 1120 4440 1126
rect 4480 1154 4680 1160
rect 4480 1126 4486 1154
rect 4514 1126 4646 1154
rect 4674 1126 4680 1154
rect 4480 1120 4680 1126
rect 4720 1154 5080 1160
rect 4720 1126 4726 1154
rect 4754 1126 4886 1154
rect 4914 1126 5046 1154
rect 5074 1126 5080 1154
rect 4720 1120 5080 1126
rect 5120 1154 5480 1160
rect 5120 1126 5126 1154
rect 5154 1126 5286 1154
rect 5314 1126 5446 1154
rect 5474 1126 5480 1154
rect 5120 1120 5480 1126
rect 5520 1154 5880 1160
rect 5520 1126 5526 1154
rect 5554 1126 5686 1154
rect 5714 1126 5846 1154
rect 5874 1126 5880 1154
rect 5520 1120 5880 1126
rect 5920 1154 6120 1160
rect 5920 1126 5926 1154
rect 5954 1126 6086 1154
rect 6114 1126 6120 1154
rect 5920 1120 6120 1126
rect 6160 1154 6360 1160
rect 6160 1126 6166 1154
rect 6194 1126 6326 1154
rect 6354 1126 6360 1154
rect 6160 1120 6360 1126
rect 4240 1074 4440 1080
rect 4240 1046 4246 1074
rect 4274 1046 4406 1074
rect 4434 1046 4440 1074
rect 4240 1040 4440 1046
rect 4480 1074 4680 1080
rect 4480 1046 4486 1074
rect 4514 1046 4646 1074
rect 4674 1046 4680 1074
rect 4480 1040 4680 1046
rect 4720 1074 5080 1080
rect 4720 1046 4726 1074
rect 4754 1046 4886 1074
rect 4914 1046 5046 1074
rect 5074 1046 5080 1074
rect 4720 1040 5080 1046
rect 5120 1074 5480 1080
rect 5120 1046 5126 1074
rect 5154 1046 5286 1074
rect 5314 1046 5446 1074
rect 5474 1046 5480 1074
rect 5120 1040 5480 1046
rect 5520 1074 5880 1080
rect 5520 1046 5526 1074
rect 5554 1046 5686 1074
rect 5714 1046 5846 1074
rect 5874 1046 5880 1074
rect 5520 1040 5880 1046
rect 5920 1074 6120 1080
rect 5920 1046 5926 1074
rect 5954 1046 6086 1074
rect 6114 1046 6120 1074
rect 5920 1040 6120 1046
rect 6160 1074 6360 1080
rect 6160 1046 6166 1074
rect 6194 1046 6326 1074
rect 6354 1046 6360 1074
rect 6160 1040 6360 1046
rect 4240 994 6360 1000
rect 4240 966 6166 994
rect 6194 966 6326 994
rect 6354 966 6360 994
rect 4240 960 6360 966
rect 4200 914 6400 920
rect 4200 886 6246 914
rect 6274 886 6400 914
rect 4200 880 6400 886
rect 4240 834 6360 840
rect 4240 806 6166 834
rect 6194 806 6326 834
rect 6354 806 6360 834
rect 4240 800 6360 806
rect 4240 754 4440 760
rect 4240 726 4246 754
rect 4274 726 4406 754
rect 4434 726 4440 754
rect 4240 720 4440 726
rect 4480 754 4680 760
rect 4480 726 4486 754
rect 4514 726 4646 754
rect 4674 726 4680 754
rect 4480 720 4680 726
rect 4720 754 5080 760
rect 4720 726 4726 754
rect 4754 726 4886 754
rect 4914 726 5046 754
rect 5074 726 5080 754
rect 4720 720 5080 726
rect 5120 754 5480 760
rect 5120 726 5126 754
rect 5154 726 5286 754
rect 5314 726 5446 754
rect 5474 726 5480 754
rect 5120 720 5480 726
rect 5520 754 5880 760
rect 5520 726 5526 754
rect 5554 726 5686 754
rect 5714 726 5846 754
rect 5874 726 5880 754
rect 5520 720 5880 726
rect 5920 754 6120 760
rect 5920 726 5926 754
rect 5954 726 6086 754
rect 6114 726 6120 754
rect 5920 720 6120 726
rect 6160 754 6360 760
rect 6160 726 6166 754
rect 6194 726 6326 754
rect 6354 726 6360 754
rect 6160 720 6360 726
rect 4240 674 4440 680
rect 4240 646 4246 674
rect 4274 646 4406 674
rect 4434 646 4440 674
rect 4240 640 4440 646
rect 4480 674 4680 680
rect 4480 646 4486 674
rect 4514 646 4646 674
rect 4674 646 4680 674
rect 4480 640 4680 646
rect 4720 674 5080 680
rect 4720 646 4726 674
rect 4754 646 4886 674
rect 4914 646 5046 674
rect 5074 646 5080 674
rect 4720 640 5080 646
rect 5120 674 5480 680
rect 5120 646 5126 674
rect 5154 646 5286 674
rect 5314 646 5446 674
rect 5474 646 5480 674
rect 5120 640 5480 646
rect 5520 674 5880 680
rect 5520 646 5526 674
rect 5554 646 5686 674
rect 5714 646 5846 674
rect 5874 646 5880 674
rect 5520 640 5880 646
rect 5920 674 6120 680
rect 5920 646 5926 674
rect 5954 646 6086 674
rect 6114 646 6120 674
rect 5920 640 6120 646
rect 6160 674 6360 680
rect 6160 646 6166 674
rect 6194 646 6326 674
rect 6354 646 6360 674
rect 6160 640 6360 646
rect 4240 594 4440 600
rect 4240 566 4246 594
rect 4274 566 4406 594
rect 4434 566 4440 594
rect 4240 560 4440 566
rect 4480 594 4680 600
rect 4480 566 4486 594
rect 4514 566 4646 594
rect 4674 566 4680 594
rect 4480 560 4680 566
rect 4720 594 5080 600
rect 4720 566 4726 594
rect 4754 566 4886 594
rect 4914 566 5046 594
rect 5074 566 5080 594
rect 4720 560 5080 566
rect 5120 594 5480 600
rect 5120 566 5126 594
rect 5154 566 5286 594
rect 5314 566 5446 594
rect 5474 566 5480 594
rect 5120 560 5480 566
rect 5520 594 5880 600
rect 5520 566 5526 594
rect 5554 566 5686 594
rect 5714 566 5846 594
rect 5874 566 5880 594
rect 5520 560 5880 566
rect 5920 594 6120 600
rect 5920 566 5926 594
rect 5954 566 6086 594
rect 6114 566 6120 594
rect 5920 560 6120 566
rect 6160 594 6360 600
rect 6160 566 6166 594
rect 6194 566 6326 594
rect 6354 566 6360 594
rect 6160 560 6360 566
rect 4240 474 6360 480
rect 4240 446 4246 474
rect 4274 446 4406 474
rect 4434 446 6360 474
rect 4240 440 6360 446
rect 4200 394 6400 400
rect 4200 366 4326 394
rect 4354 366 6400 394
rect 4200 360 6400 366
rect 4240 314 6360 320
rect 4240 286 4246 314
rect 4274 286 4406 314
rect 4434 286 6360 314
rect 4240 280 6360 286
rect 4240 194 4440 200
rect 4240 166 4246 194
rect 4274 166 4406 194
rect 4434 166 4440 194
rect 4240 160 4440 166
rect 4480 194 4680 200
rect 4480 166 4486 194
rect 4514 166 4646 194
rect 4674 166 4680 194
rect 4480 160 4680 166
rect 4720 194 5080 200
rect 4720 166 4726 194
rect 4754 166 4886 194
rect 4914 166 5046 194
rect 5074 166 5080 194
rect 4720 160 5080 166
rect 5120 194 5480 200
rect 5120 166 5126 194
rect 5154 166 5286 194
rect 5314 166 5446 194
rect 5474 166 5480 194
rect 5120 160 5480 166
rect 5520 194 5880 200
rect 5520 166 5526 194
rect 5554 166 5686 194
rect 5714 166 5846 194
rect 5874 166 5880 194
rect 5520 160 5880 166
rect 5920 194 6120 200
rect 5920 166 5926 194
rect 5954 166 6086 194
rect 6114 166 6120 194
rect 5920 160 6120 166
rect 6160 194 6360 200
rect 6160 166 6166 194
rect 6194 166 6326 194
rect 6354 166 6360 194
rect 6160 160 6360 166
rect 4240 114 4440 120
rect 4240 86 4246 114
rect 4274 86 4406 114
rect 4434 86 4440 114
rect 4240 80 4440 86
rect 4480 114 4680 120
rect 4480 86 4486 114
rect 4514 86 4646 114
rect 4674 86 4680 114
rect 4480 80 4680 86
rect 4720 114 5080 120
rect 4720 86 4726 114
rect 4754 86 4886 114
rect 4914 86 5046 114
rect 5074 86 5080 114
rect 4720 80 5080 86
rect 5120 114 5480 120
rect 5120 86 5126 114
rect 5154 86 5286 114
rect 5314 86 5446 114
rect 5474 86 5480 114
rect 5120 80 5480 86
rect 5520 114 5880 120
rect 5520 86 5526 114
rect 5554 86 5686 114
rect 5714 86 5846 114
rect 5874 86 5880 114
rect 5520 80 5880 86
rect 5920 114 6120 120
rect 5920 86 5926 114
rect 5954 86 6086 114
rect 6114 86 6120 114
rect 5920 80 6120 86
rect 6160 114 6360 120
rect 6160 86 6166 114
rect 6194 86 6326 114
rect 6354 86 6360 114
rect 6160 80 6360 86
rect 4240 34 4440 40
rect 4240 6 4246 34
rect 4274 6 4406 34
rect 4434 6 4440 34
rect 4240 0 4440 6
rect 4480 34 4680 40
rect 4480 6 4486 34
rect 4514 6 4646 34
rect 4674 6 4680 34
rect 4480 0 4680 6
rect 4720 34 5080 40
rect 4720 6 4726 34
rect 4754 6 4886 34
rect 4914 6 5046 34
rect 5074 6 5080 34
rect 4720 0 5080 6
rect 5120 34 5480 40
rect 5120 6 5126 34
rect 5154 6 5286 34
rect 5314 6 5446 34
rect 5474 6 5480 34
rect 5120 0 5480 6
rect 5520 34 5880 40
rect 5520 6 5526 34
rect 5554 6 5686 34
rect 5714 6 5846 34
rect 5874 6 5880 34
rect 5520 0 5880 6
rect 5920 34 6120 40
rect 5920 6 5926 34
rect 5954 6 6086 34
rect 6114 6 6120 34
rect 5920 0 6120 6
rect 6160 34 6360 40
rect 6160 6 6166 34
rect 6194 6 6326 34
rect 6354 6 6360 34
rect 6160 0 6360 6
<< via2 >>
rect 4246 12606 4274 12634
rect 4406 12606 4434 12634
rect 4486 12606 4514 12634
rect 4646 12606 4674 12634
rect 4726 12606 4754 12634
rect 4886 12606 4914 12634
rect 5046 12606 5074 12634
rect 5126 12606 5154 12634
rect 5286 12606 5314 12634
rect 5446 12606 5474 12634
rect 5526 12606 5554 12634
rect 5686 12606 5714 12634
rect 5846 12606 5874 12634
rect 5926 12606 5954 12634
rect 6086 12606 6114 12634
rect 6166 12606 6194 12634
rect 6326 12606 6354 12634
rect 4246 12526 4274 12554
rect 4406 12526 4434 12554
rect 4486 12526 4514 12554
rect 4646 12526 4674 12554
rect 4726 12526 4754 12554
rect 4886 12526 4914 12554
rect 5046 12526 5074 12554
rect 5126 12526 5154 12554
rect 5286 12526 5314 12554
rect 5446 12526 5474 12554
rect 5526 12526 5554 12554
rect 5686 12526 5714 12554
rect 5846 12526 5874 12554
rect 5926 12526 5954 12554
rect 6086 12526 6114 12554
rect 6166 12526 6194 12554
rect 6326 12526 6354 12554
rect 4246 12446 4274 12474
rect 4406 12446 4434 12474
rect 4486 12446 4514 12474
rect 4646 12446 4674 12474
rect 4726 12446 4754 12474
rect 4886 12446 4914 12474
rect 5046 12446 5074 12474
rect 5126 12446 5154 12474
rect 5286 12446 5314 12474
rect 5446 12446 5474 12474
rect 5526 12446 5554 12474
rect 5686 12446 5714 12474
rect 5846 12446 5874 12474
rect 5926 12446 5954 12474
rect 6086 12446 6114 12474
rect 6166 12446 6194 12474
rect 6326 12446 6354 12474
rect 4246 12366 4274 12394
rect 4406 12366 4434 12394
rect 4486 12366 4514 12394
rect 4646 12366 4674 12394
rect 4726 12366 4754 12394
rect 4886 12366 4914 12394
rect 5046 12366 5074 12394
rect 5126 12366 5154 12394
rect 5286 12366 5314 12394
rect 5446 12366 5474 12394
rect 5526 12366 5554 12394
rect 5686 12366 5714 12394
rect 5846 12366 5874 12394
rect 5926 12366 5954 12394
rect 6086 12366 6114 12394
rect 6166 12366 6194 12394
rect 6326 12366 6354 12394
rect 4246 12286 4274 12314
rect 4406 12286 4434 12314
rect 4486 12286 4514 12314
rect 4646 12286 4674 12314
rect 4726 12286 4754 12314
rect 4886 12286 4914 12314
rect 5046 12286 5074 12314
rect 5126 12286 5154 12314
rect 5286 12286 5314 12314
rect 5446 12286 5474 12314
rect 5526 12286 5554 12314
rect 5686 12286 5714 12314
rect 5846 12286 5874 12314
rect 5926 12286 5954 12314
rect 6086 12286 6114 12314
rect 6166 12286 6194 12314
rect 6326 12286 6354 12314
rect 4246 12206 4274 12234
rect 4406 12206 4434 12234
rect 4486 12206 4514 12234
rect 4646 12206 4674 12234
rect 4726 12206 4754 12234
rect 4886 12206 4914 12234
rect 5046 12206 5074 12234
rect 5126 12206 5154 12234
rect 5286 12206 5314 12234
rect 5446 12206 5474 12234
rect 5526 12206 5554 12234
rect 5686 12206 5714 12234
rect 5846 12206 5874 12234
rect 5926 12206 5954 12234
rect 6086 12206 6114 12234
rect 6166 12206 6194 12234
rect 6326 12206 6354 12234
rect 4246 12126 4274 12154
rect 4406 12126 4434 12154
rect 4486 12126 4514 12154
rect 4646 12126 4674 12154
rect 4726 12126 4754 12154
rect 4886 12126 4914 12154
rect 5046 12126 5074 12154
rect 5126 12126 5154 12154
rect 5286 12126 5314 12154
rect 5446 12126 5474 12154
rect 5526 12126 5554 12154
rect 5686 12126 5714 12154
rect 5846 12126 5874 12154
rect 5926 12126 5954 12154
rect 6086 12126 6114 12154
rect 6166 12126 6194 12154
rect 6326 12126 6354 12154
rect 4486 12046 4514 12074
rect 4646 12046 4674 12074
rect 4566 11966 4594 11994
rect 4486 11886 4514 11914
rect 4646 11886 4674 11914
rect 4246 11806 4274 11834
rect 4406 11806 4434 11834
rect 4486 11806 4514 11834
rect 4646 11806 4674 11834
rect 4726 11806 4754 11834
rect 4886 11806 4914 11834
rect 5046 11806 5074 11834
rect 5126 11806 5154 11834
rect 5286 11806 5314 11834
rect 5446 11806 5474 11834
rect 5526 11806 5554 11834
rect 5686 11806 5714 11834
rect 5846 11806 5874 11834
rect 5926 11806 5954 11834
rect 6086 11806 6114 11834
rect 6166 11806 6194 11834
rect 6326 11806 6354 11834
rect 4246 11726 4274 11754
rect 4406 11726 4434 11754
rect 4486 11726 4514 11754
rect 4646 11726 4674 11754
rect 4726 11726 4754 11754
rect 4886 11726 4914 11754
rect 5046 11726 5074 11754
rect 5126 11726 5154 11754
rect 5286 11726 5314 11754
rect 5446 11726 5474 11754
rect 5526 11726 5554 11754
rect 5686 11726 5714 11754
rect 5846 11726 5874 11754
rect 5926 11726 5954 11754
rect 6086 11726 6114 11754
rect 6166 11726 6194 11754
rect 6326 11726 6354 11754
rect 4246 11646 4274 11674
rect 4406 11646 4434 11674
rect 4486 11646 4514 11674
rect 4646 11646 4674 11674
rect 4726 11646 4754 11674
rect 4886 11646 4914 11674
rect 5046 11646 5074 11674
rect 5126 11646 5154 11674
rect 5286 11646 5314 11674
rect 5446 11646 5474 11674
rect 5526 11646 5554 11674
rect 5686 11646 5714 11674
rect 5846 11646 5874 11674
rect 5926 11646 5954 11674
rect 6086 11646 6114 11674
rect 6166 11646 6194 11674
rect 6326 11646 6354 11674
rect 4246 11566 4274 11594
rect 4406 11566 4434 11594
rect 4486 11566 4514 11594
rect 4646 11566 4674 11594
rect 4726 11566 4754 11594
rect 4886 11566 4914 11594
rect 5046 11566 5074 11594
rect 5126 11566 5154 11594
rect 5286 11566 5314 11594
rect 5446 11566 5474 11594
rect 5526 11566 5554 11594
rect 5686 11566 5714 11594
rect 5846 11566 5874 11594
rect 5926 11566 5954 11594
rect 6086 11566 6114 11594
rect 6166 11566 6194 11594
rect 6326 11566 6354 11594
rect 4246 11486 4274 11514
rect 4406 11486 4434 11514
rect 4486 11486 4514 11514
rect 4646 11486 4674 11514
rect 4726 11486 4754 11514
rect 4886 11486 4914 11514
rect 5046 11486 5074 11514
rect 5126 11486 5154 11514
rect 5286 11486 5314 11514
rect 5446 11486 5474 11514
rect 5526 11486 5554 11514
rect 5686 11486 5714 11514
rect 5846 11486 5874 11514
rect 5926 11486 5954 11514
rect 6086 11486 6114 11514
rect 6166 11486 6194 11514
rect 6326 11486 6354 11514
rect 4246 11406 4274 11434
rect 4406 11406 4434 11434
rect 4486 11406 4514 11434
rect 4646 11406 4674 11434
rect 4726 11406 4754 11434
rect 4886 11406 4914 11434
rect 5046 11406 5074 11434
rect 5126 11406 5154 11434
rect 5286 11406 5314 11434
rect 5446 11406 5474 11434
rect 5526 11406 5554 11434
rect 5686 11406 5714 11434
rect 5846 11406 5874 11434
rect 5926 11406 5954 11434
rect 6086 11406 6114 11434
rect 6166 11406 6194 11434
rect 6326 11406 6354 11434
rect 5526 11286 5554 11314
rect 5686 11286 5714 11314
rect 5606 11206 5634 11234
rect 5046 11126 5074 11154
rect 5526 11126 5554 11154
rect 5686 11126 5714 11154
rect 5126 11046 5154 11074
rect 5286 11046 5314 11074
rect 5446 11046 5474 11074
rect 5046 10966 5074 10994
rect 5526 10966 5554 10994
rect 4246 10846 4274 10874
rect 4406 10846 4434 10874
rect 4486 10846 4514 10874
rect 4646 10846 4674 10874
rect 4726 10846 4754 10874
rect 4886 10846 4914 10874
rect 5046 10846 5074 10874
rect 5126 10846 5154 10874
rect 5286 10846 5314 10874
rect 5446 10846 5474 10874
rect 5526 10846 5554 10874
rect 5686 10846 5714 10874
rect 5846 10846 5874 10874
rect 5926 10846 5954 10874
rect 6086 10846 6114 10874
rect 6166 10846 6194 10874
rect 6326 10846 6354 10874
rect 4246 10766 4274 10794
rect 4406 10766 4434 10794
rect 4486 10766 4514 10794
rect 4646 10766 4674 10794
rect 4726 10766 4754 10794
rect 4886 10766 4914 10794
rect 5046 10766 5074 10794
rect 5126 10766 5154 10794
rect 5286 10766 5314 10794
rect 5446 10766 5474 10794
rect 5526 10766 5554 10794
rect 5686 10766 5714 10794
rect 5846 10766 5874 10794
rect 5926 10766 5954 10794
rect 6086 10766 6114 10794
rect 6166 10766 6194 10794
rect 6326 10766 6354 10794
rect 4246 10686 4274 10714
rect 4406 10686 4434 10714
rect 4486 10686 4514 10714
rect 4646 10686 4674 10714
rect 4726 10686 4754 10714
rect 4886 10686 4914 10714
rect 5046 10686 5074 10714
rect 5126 10686 5154 10714
rect 5286 10686 5314 10714
rect 5446 10686 5474 10714
rect 5526 10686 5554 10714
rect 5686 10686 5714 10714
rect 5846 10686 5874 10714
rect 5926 10686 5954 10714
rect 6086 10686 6114 10714
rect 6166 10686 6194 10714
rect 6326 10686 6354 10714
rect 4246 10606 4274 10634
rect 4406 10606 4434 10634
rect 4486 10606 4514 10634
rect 4646 10606 4674 10634
rect 4726 10606 4754 10634
rect 4886 10606 4914 10634
rect 5046 10606 5074 10634
rect 5126 10606 5154 10634
rect 5286 10606 5314 10634
rect 5446 10606 5474 10634
rect 5526 10606 5554 10634
rect 5686 10606 5714 10634
rect 5846 10606 5874 10634
rect 5926 10606 5954 10634
rect 6086 10606 6114 10634
rect 6166 10606 6194 10634
rect 6326 10606 6354 10634
rect 4246 10526 4274 10554
rect 4406 10526 4434 10554
rect 4486 10526 4514 10554
rect 4646 10526 4674 10554
rect 4726 10526 4754 10554
rect 4886 10526 4914 10554
rect 5046 10526 5074 10554
rect 5126 10526 5154 10554
rect 5286 10526 5314 10554
rect 5446 10526 5474 10554
rect 5526 10526 5554 10554
rect 5686 10526 5714 10554
rect 5846 10526 5874 10554
rect 5926 10526 5954 10554
rect 6086 10526 6114 10554
rect 6166 10526 6194 10554
rect 6326 10526 6354 10554
rect 4246 10446 4274 10474
rect 4406 10446 4434 10474
rect 4486 10446 4514 10474
rect 4646 10446 4674 10474
rect 4726 10446 4754 10474
rect 4886 10446 4914 10474
rect 5046 10446 5074 10474
rect 5126 10446 5154 10474
rect 5286 10446 5314 10474
rect 5446 10446 5474 10474
rect 5526 10446 5554 10474
rect 5686 10446 5714 10474
rect 5846 10446 5874 10474
rect 5926 10446 5954 10474
rect 6086 10446 6114 10474
rect 6166 10446 6194 10474
rect 6326 10446 6354 10474
rect 4246 10366 4274 10394
rect 4406 10366 4434 10394
rect 4486 10366 4514 10394
rect 4646 10366 4674 10394
rect 4726 10366 4754 10394
rect 4886 10366 4914 10394
rect 5046 10366 5074 10394
rect 5126 10366 5154 10394
rect 5286 10366 5314 10394
rect 5446 10366 5474 10394
rect 5526 10366 5554 10394
rect 5686 10366 5714 10394
rect 5846 10366 5874 10394
rect 5926 10366 5954 10394
rect 6086 10366 6114 10394
rect 6166 10366 6194 10394
rect 6326 10366 6354 10394
rect 4246 10286 4274 10314
rect 4406 10286 4434 10314
rect 4486 10286 4514 10314
rect 4646 10286 4674 10314
rect 4726 10286 4754 10314
rect 4886 10286 4914 10314
rect 5046 10286 5074 10314
rect 5126 10286 5154 10314
rect 5286 10286 5314 10314
rect 5446 10286 5474 10314
rect 5526 10286 5554 10314
rect 5686 10286 5714 10314
rect 5846 10286 5874 10314
rect 5926 10286 5954 10314
rect 6086 10286 6114 10314
rect 6166 10286 6194 10314
rect 6326 10286 6354 10314
rect 4246 10206 4274 10234
rect 4406 10206 4434 10234
rect 4486 10206 4514 10234
rect 4646 10206 4674 10234
rect 4726 10206 4754 10234
rect 4886 10206 4914 10234
rect 5046 10206 5074 10234
rect 5126 10206 5154 10234
rect 5286 10206 5314 10234
rect 5446 10206 5474 10234
rect 5526 10206 5554 10234
rect 5686 10206 5714 10234
rect 5846 10206 5874 10234
rect 5926 10206 5954 10234
rect 6086 10206 6114 10234
rect 6166 10206 6194 10234
rect 6326 10206 6354 10234
rect 4246 10126 4274 10154
rect 4406 10126 4434 10154
rect 4486 10126 4514 10154
rect 4646 10126 4674 10154
rect 4726 10126 4754 10154
rect 4886 10126 4914 10154
rect 5046 10126 5074 10154
rect 5126 10126 5154 10154
rect 5286 10126 5314 10154
rect 5446 10126 5474 10154
rect 5526 10126 5554 10154
rect 5686 10126 5714 10154
rect 5846 10126 5874 10154
rect 5926 10126 5954 10154
rect 6086 10126 6114 10154
rect 6166 10126 6194 10154
rect 6326 10126 6354 10154
rect 4246 10046 4274 10074
rect 4406 10046 4434 10074
rect 4486 10046 4514 10074
rect 4646 10046 4674 10074
rect 4726 10046 4754 10074
rect 4886 10046 4914 10074
rect 5046 10046 5074 10074
rect 5126 10046 5154 10074
rect 5286 10046 5314 10074
rect 5446 10046 5474 10074
rect 5526 10046 5554 10074
rect 5686 10046 5714 10074
rect 5846 10046 5874 10074
rect 5926 10046 5954 10074
rect 6086 10046 6114 10074
rect 6166 10046 6194 10074
rect 6326 10046 6354 10074
rect 4246 9966 4274 9994
rect 4406 9966 4434 9994
rect 4486 9966 4514 9994
rect 4646 9966 4674 9994
rect 4726 9966 4754 9994
rect 4886 9966 4914 9994
rect 5046 9966 5074 9994
rect 5126 9966 5154 9994
rect 5286 9966 5314 9994
rect 5446 9966 5474 9994
rect 5526 9966 5554 9994
rect 5686 9966 5714 9994
rect 5846 9966 5874 9994
rect 5926 9966 5954 9994
rect 6086 9966 6114 9994
rect 6166 9966 6194 9994
rect 6326 9966 6354 9994
rect 4246 9886 4274 9914
rect 4406 9886 4434 9914
rect 4486 9886 4514 9914
rect 4646 9886 4674 9914
rect 4726 9886 4754 9914
rect 4886 9886 4914 9914
rect 5046 9886 5074 9914
rect 5126 9886 5154 9914
rect 5286 9886 5314 9914
rect 5446 9886 5474 9914
rect 5526 9886 5554 9914
rect 5686 9886 5714 9914
rect 5846 9886 5874 9914
rect 5926 9886 5954 9914
rect 6086 9886 6114 9914
rect 6166 9886 6194 9914
rect 6326 9886 6354 9914
rect 4246 9806 4274 9834
rect 4406 9806 4434 9834
rect 4486 9806 4514 9834
rect 4646 9806 4674 9834
rect 4726 9806 4754 9834
rect 4886 9806 4914 9834
rect 5046 9806 5074 9834
rect 5126 9806 5154 9834
rect 5286 9806 5314 9834
rect 5446 9806 5474 9834
rect 5526 9806 5554 9834
rect 5686 9806 5714 9834
rect 5846 9806 5874 9834
rect 5926 9806 5954 9834
rect 6086 9806 6114 9834
rect 6166 9806 6194 9834
rect 6326 9806 6354 9834
rect 4246 9726 4274 9754
rect 4406 9726 4434 9754
rect 4486 9726 4514 9754
rect 4646 9726 4674 9754
rect 4726 9726 4754 9754
rect 4886 9726 4914 9754
rect 5046 9726 5074 9754
rect 5126 9726 5154 9754
rect 5286 9726 5314 9754
rect 5446 9726 5474 9754
rect 5526 9726 5554 9754
rect 5686 9726 5714 9754
rect 5846 9726 5874 9754
rect 5926 9726 5954 9754
rect 6086 9726 6114 9754
rect 6166 9726 6194 9754
rect 6326 9726 6354 9754
rect 4486 9606 4514 9634
rect 4646 9606 4674 9634
rect 4566 9526 4594 9554
rect 4486 9446 4514 9474
rect 4646 9446 4674 9474
rect 4246 9326 4274 9354
rect 4406 9326 4434 9354
rect 4486 9326 4514 9354
rect 4646 9326 4674 9354
rect 4726 9326 4754 9354
rect 4886 9326 4914 9354
rect 5046 9326 5074 9354
rect 5126 9326 5154 9354
rect 5286 9326 5314 9354
rect 5446 9326 5474 9354
rect 5526 9326 5554 9354
rect 5686 9326 5714 9354
rect 5846 9326 5874 9354
rect 5926 9326 5954 9354
rect 6086 9326 6114 9354
rect 6166 9326 6194 9354
rect 6326 9326 6354 9354
rect 4246 9246 4274 9274
rect 4406 9246 4434 9274
rect 4486 9246 4514 9274
rect 4646 9246 4674 9274
rect 4726 9246 4754 9274
rect 4886 9246 4914 9274
rect 5046 9246 5074 9274
rect 5126 9246 5154 9274
rect 5286 9246 5314 9274
rect 5446 9246 5474 9274
rect 5526 9246 5554 9274
rect 5686 9246 5714 9274
rect 5846 9246 5874 9274
rect 5926 9246 5954 9274
rect 6086 9246 6114 9274
rect 6166 9246 6194 9274
rect 6326 9246 6354 9274
rect 4246 9166 4274 9194
rect 4406 9166 4434 9194
rect 4486 9166 4514 9194
rect 4646 9166 4674 9194
rect 4726 9166 4754 9194
rect 4886 9166 4914 9194
rect 5046 9166 5074 9194
rect 5126 9166 5154 9194
rect 5286 9166 5314 9194
rect 5446 9166 5474 9194
rect 5526 9166 5554 9194
rect 5686 9166 5714 9194
rect 5846 9166 5874 9194
rect 5926 9166 5954 9194
rect 6086 9166 6114 9194
rect 6166 9166 6194 9194
rect 6326 9166 6354 9194
rect 5126 9086 5154 9114
rect 5286 9086 5314 9114
rect 5446 9086 5474 9114
rect 5366 9006 5394 9034
rect 5126 8926 5154 8954
rect 5286 8926 5314 8954
rect 5446 8926 5474 8954
rect 4246 8846 4274 8874
rect 4406 8846 4434 8874
rect 4486 8846 4514 8874
rect 4646 8846 4674 8874
rect 4726 8846 4754 8874
rect 4886 8846 4914 8874
rect 5046 8846 5074 8874
rect 5126 8846 5154 8874
rect 5286 8846 5314 8874
rect 5446 8846 5474 8874
rect 5526 8846 5554 8874
rect 5686 8846 5714 8874
rect 5846 8846 5874 8874
rect 5926 8846 5954 8874
rect 6086 8846 6114 8874
rect 6166 8846 6194 8874
rect 6326 8846 6354 8874
rect 4246 8766 4274 8794
rect 4406 8766 4434 8794
rect 4486 8766 4514 8794
rect 4646 8766 4674 8794
rect 4726 8766 4754 8794
rect 4886 8766 4914 8794
rect 5046 8766 5074 8794
rect 5126 8766 5154 8794
rect 5286 8766 5314 8794
rect 5446 8766 5474 8794
rect 5526 8766 5554 8794
rect 5686 8766 5714 8794
rect 5846 8766 5874 8794
rect 5926 8766 5954 8794
rect 6086 8766 6114 8794
rect 6166 8766 6194 8794
rect 6326 8766 6354 8794
rect 4246 8686 4274 8714
rect 4406 8686 4434 8714
rect 4486 8686 4514 8714
rect 4646 8686 4674 8714
rect 4726 8686 4754 8714
rect 4886 8686 4914 8714
rect 5046 8686 5074 8714
rect 5126 8686 5154 8714
rect 5286 8686 5314 8714
rect 5446 8686 5474 8714
rect 5526 8686 5554 8714
rect 5686 8686 5714 8714
rect 5846 8686 5874 8714
rect 5926 8686 5954 8714
rect 6086 8686 6114 8714
rect 6166 8686 6194 8714
rect 6326 8686 6354 8714
rect 4246 8606 4274 8634
rect 4406 8606 4434 8634
rect 4486 8606 4514 8634
rect 4646 8606 4674 8634
rect 4726 8606 4754 8634
rect 4886 8606 4914 8634
rect 5046 8606 5074 8634
rect 5126 8606 5154 8634
rect 5286 8606 5314 8634
rect 5446 8606 5474 8634
rect 5526 8606 5554 8634
rect 5686 8606 5714 8634
rect 5846 8606 5874 8634
rect 5926 8606 5954 8634
rect 6086 8606 6114 8634
rect 6166 8606 6194 8634
rect 6326 8606 6354 8634
rect 4246 8526 4274 8554
rect 4406 8526 4434 8554
rect 4486 8526 4514 8554
rect 4646 8526 4674 8554
rect 4726 8526 4754 8554
rect 4886 8526 4914 8554
rect 5046 8526 5074 8554
rect 5126 8526 5154 8554
rect 5286 8526 5314 8554
rect 5446 8526 5474 8554
rect 5526 8526 5554 8554
rect 5686 8526 5714 8554
rect 5846 8526 5874 8554
rect 5926 8526 5954 8554
rect 6086 8526 6114 8554
rect 6166 8526 6194 8554
rect 6326 8526 6354 8554
rect 4886 8446 4914 8474
rect 5046 8446 5074 8474
rect 5686 8446 5714 8474
rect 5846 8446 5874 8474
rect 4966 8366 4994 8394
rect 5766 8366 5794 8394
rect 4886 8286 4914 8314
rect 5046 8286 5074 8314
rect 5526 8286 5554 8314
rect 5686 8286 5714 8314
rect 5846 8286 5874 8314
rect 5606 8206 5634 8234
rect 5526 8126 5554 8154
rect 5686 8126 5714 8154
rect 5046 8046 5074 8074
rect 5526 8046 5554 8074
rect 5126 7966 5154 7994
rect 5286 7966 5314 7994
rect 5446 7966 5474 7994
rect 5206 7886 5234 7914
rect 5126 7806 5154 7834
rect 5286 7806 5314 7834
rect 5446 7806 5474 7834
rect 5046 7726 5074 7754
rect 5526 7726 5554 7754
rect 4246 7606 4274 7634
rect 4406 7606 4434 7634
rect 4486 7606 4514 7634
rect 4646 7606 4674 7634
rect 4726 7606 4754 7634
rect 4886 7606 4914 7634
rect 5046 7606 5074 7634
rect 5126 7606 5154 7634
rect 5286 7606 5314 7634
rect 5446 7606 5474 7634
rect 5526 7606 5554 7634
rect 5686 7606 5714 7634
rect 5846 7606 5874 7634
rect 5926 7606 5954 7634
rect 6086 7606 6114 7634
rect 6166 7606 6194 7634
rect 6326 7606 6354 7634
rect 4246 7526 4274 7554
rect 4406 7526 4434 7554
rect 4486 7526 4514 7554
rect 4646 7526 4674 7554
rect 4726 7526 4754 7554
rect 4886 7526 4914 7554
rect 5046 7526 5074 7554
rect 5126 7526 5154 7554
rect 5286 7526 5314 7554
rect 5446 7526 5474 7554
rect 5526 7526 5554 7554
rect 5686 7526 5714 7554
rect 5846 7526 5874 7554
rect 5926 7526 5954 7554
rect 6086 7526 6114 7554
rect 6166 7526 6194 7554
rect 6326 7526 6354 7554
rect 4246 7446 4274 7474
rect 4406 7446 4434 7474
rect 4486 7446 4514 7474
rect 4646 7446 4674 7474
rect 4726 7446 4754 7474
rect 4886 7446 4914 7474
rect 5046 7446 5074 7474
rect 5126 7446 5154 7474
rect 5286 7446 5314 7474
rect 5446 7446 5474 7474
rect 5526 7446 5554 7474
rect 5686 7446 5714 7474
rect 5846 7446 5874 7474
rect 5926 7446 5954 7474
rect 6086 7446 6114 7474
rect 6166 7446 6194 7474
rect 6326 7446 6354 7474
rect 4246 7366 4274 7394
rect 4406 7366 4434 7394
rect 4486 7366 4514 7394
rect 4646 7366 4674 7394
rect 4726 7366 4754 7394
rect 4886 7366 4914 7394
rect 5046 7366 5074 7394
rect 5126 7366 5154 7394
rect 5286 7366 5314 7394
rect 5446 7366 5474 7394
rect 5526 7366 5554 7394
rect 5686 7366 5714 7394
rect 5846 7366 5874 7394
rect 5926 7366 5954 7394
rect 6086 7366 6114 7394
rect 6166 7366 6194 7394
rect 6326 7366 6354 7394
rect 4246 7286 4274 7314
rect 4406 7286 4434 7314
rect 4486 7286 4514 7314
rect 4646 7286 4674 7314
rect 4726 7286 4754 7314
rect 4886 7286 4914 7314
rect 5046 7286 5074 7314
rect 5126 7286 5154 7314
rect 5286 7286 5314 7314
rect 5446 7286 5474 7314
rect 5526 7286 5554 7314
rect 5686 7286 5714 7314
rect 5846 7286 5874 7314
rect 5926 7286 5954 7314
rect 6086 7286 6114 7314
rect 6166 7286 6194 7314
rect 6326 7286 6354 7314
rect 4246 7206 4274 7234
rect 4406 7206 4434 7234
rect 4486 7206 4514 7234
rect 4646 7206 4674 7234
rect 4726 7206 4754 7234
rect 4886 7206 4914 7234
rect 5046 7206 5074 7234
rect 5126 7206 5154 7234
rect 5286 7206 5314 7234
rect 5446 7206 5474 7234
rect 5526 7206 5554 7234
rect 5686 7206 5714 7234
rect 5846 7206 5874 7234
rect 5926 7206 5954 7234
rect 6086 7206 6114 7234
rect 6166 7206 6194 7234
rect 6326 7206 6354 7234
rect 4246 7126 4274 7154
rect 4406 7126 4434 7154
rect 4486 7126 4514 7154
rect 4646 7126 4674 7154
rect 4726 7126 4754 7154
rect 4886 7126 4914 7154
rect 5046 7126 5074 7154
rect 5126 7126 5154 7154
rect 5286 7126 5314 7154
rect 5446 7126 5474 7154
rect 5526 7126 5554 7154
rect 5686 7126 5714 7154
rect 5846 7126 5874 7154
rect 5926 7126 5954 7154
rect 6086 7126 6114 7154
rect 6166 7126 6194 7154
rect 6326 7126 6354 7154
rect 4246 7046 4274 7074
rect 4406 7046 4434 7074
rect 4486 7046 4514 7074
rect 4646 7046 4674 7074
rect 4726 7046 4754 7074
rect 4886 7046 4914 7074
rect 5046 7046 5074 7074
rect 5126 7046 5154 7074
rect 5286 7046 5314 7074
rect 5446 7046 5474 7074
rect 5526 7046 5554 7074
rect 5686 7046 5714 7074
rect 5846 7046 5874 7074
rect 5926 7046 5954 7074
rect 6086 7046 6114 7074
rect 6166 7046 6194 7074
rect 6326 7046 6354 7074
rect 4486 6966 4514 6994
rect 4646 6966 4674 6994
rect 4566 6886 4594 6914
rect 4486 6806 4514 6834
rect 4646 6806 4674 6834
rect 4246 6726 4274 6754
rect 4406 6726 4434 6754
rect 4486 6726 4514 6754
rect 4646 6726 4674 6754
rect 4726 6726 4754 6754
rect 4886 6726 4914 6754
rect 5046 6726 5074 6754
rect 5126 6726 5154 6754
rect 5286 6726 5314 6754
rect 5446 6726 5474 6754
rect 5526 6726 5554 6754
rect 5686 6726 5714 6754
rect 5846 6726 5874 6754
rect 5926 6726 5954 6754
rect 6086 6726 6114 6754
rect 6166 6726 6194 6754
rect 6326 6726 6354 6754
rect 4246 6646 4274 6674
rect 4406 6646 4434 6674
rect 4486 6646 4514 6674
rect 4646 6646 4674 6674
rect 4726 6646 4754 6674
rect 4886 6646 4914 6674
rect 5046 6646 5074 6674
rect 5126 6646 5154 6674
rect 5286 6646 5314 6674
rect 5446 6646 5474 6674
rect 5526 6646 5554 6674
rect 5686 6646 5714 6674
rect 5846 6646 5874 6674
rect 5926 6646 5954 6674
rect 6086 6646 6114 6674
rect 6166 6646 6194 6674
rect 6326 6646 6354 6674
rect 4246 6566 4274 6594
rect 4406 6566 4434 6594
rect 4486 6566 4514 6594
rect 4646 6566 4674 6594
rect 4726 6566 4754 6594
rect 4886 6566 4914 6594
rect 5046 6566 5074 6594
rect 5126 6566 5154 6594
rect 5286 6566 5314 6594
rect 5446 6566 5474 6594
rect 5526 6566 5554 6594
rect 5686 6566 5714 6594
rect 5846 6566 5874 6594
rect 5926 6566 5954 6594
rect 6086 6566 6114 6594
rect 6166 6566 6194 6594
rect 6326 6566 6354 6594
rect 4246 6486 4274 6514
rect 4406 6486 4434 6514
rect 4486 6486 4514 6514
rect 4646 6486 4674 6514
rect 4726 6486 4754 6514
rect 4886 6486 4914 6514
rect 5046 6486 5074 6514
rect 5126 6486 5154 6514
rect 5286 6486 5314 6514
rect 5446 6486 5474 6514
rect 5526 6486 5554 6514
rect 5686 6486 5714 6514
rect 5846 6486 5874 6514
rect 5926 6486 5954 6514
rect 6086 6486 6114 6514
rect 6166 6486 6194 6514
rect 6326 6486 6354 6514
rect 4246 6406 4274 6434
rect 4406 6406 4434 6434
rect 4486 6406 4514 6434
rect 4646 6406 4674 6434
rect 4726 6406 4754 6434
rect 4886 6406 4914 6434
rect 5046 6406 5074 6434
rect 5126 6406 5154 6434
rect 5286 6406 5314 6434
rect 5446 6406 5474 6434
rect 5526 6406 5554 6434
rect 5686 6406 5714 6434
rect 5846 6406 5874 6434
rect 5926 6406 5954 6434
rect 6086 6406 6114 6434
rect 6166 6406 6194 6434
rect 6326 6406 6354 6434
rect 4246 6326 4274 6354
rect 4406 6326 4434 6354
rect 4486 6326 4514 6354
rect 4646 6326 4674 6354
rect 4726 6326 4754 6354
rect 4886 6326 4914 6354
rect 5046 6326 5074 6354
rect 5126 6326 5154 6354
rect 5286 6326 5314 6354
rect 5446 6326 5474 6354
rect 5526 6326 5554 6354
rect 5686 6326 5714 6354
rect 5846 6326 5874 6354
rect 5926 6326 5954 6354
rect 6086 6326 6114 6354
rect 6166 6326 6194 6354
rect 6326 6326 6354 6354
rect 4726 6206 4754 6234
rect 4886 6206 4914 6234
rect 5046 6206 5074 6234
rect 4806 6126 4834 6154
rect 4966 6126 4994 6154
rect 4726 6046 4754 6074
rect 4886 6046 4914 6074
rect 5046 6046 5074 6074
rect 4966 5966 4994 5994
rect 4726 5886 4754 5914
rect 4886 5886 4914 5914
rect 5046 5886 5074 5914
rect 4246 5766 4274 5794
rect 4406 5766 4434 5794
rect 4486 5766 4514 5794
rect 4646 5766 4674 5794
rect 4726 5766 4754 5794
rect 4886 5766 4914 5794
rect 5046 5766 5074 5794
rect 5126 5766 5154 5794
rect 5286 5766 5314 5794
rect 5446 5766 5474 5794
rect 5526 5766 5554 5794
rect 5686 5766 5714 5794
rect 5846 5766 5874 5794
rect 5926 5766 5954 5794
rect 6086 5766 6114 5794
rect 6166 5766 6194 5794
rect 6326 5766 6354 5794
rect 4246 5686 4274 5714
rect 4406 5686 4434 5714
rect 4486 5686 4514 5714
rect 4646 5686 4674 5714
rect 4726 5686 4754 5714
rect 4886 5686 4914 5714
rect 5046 5686 5074 5714
rect 5126 5686 5154 5714
rect 5286 5686 5314 5714
rect 5446 5686 5474 5714
rect 5526 5686 5554 5714
rect 5686 5686 5714 5714
rect 5846 5686 5874 5714
rect 5926 5686 5954 5714
rect 6086 5686 6114 5714
rect 6166 5686 6194 5714
rect 6326 5686 6354 5714
rect 4246 5606 4274 5634
rect 4406 5606 4434 5634
rect 4486 5606 4514 5634
rect 4646 5606 4674 5634
rect 4726 5606 4754 5634
rect 4886 5606 4914 5634
rect 5046 5606 5074 5634
rect 5126 5606 5154 5634
rect 5286 5606 5314 5634
rect 5446 5606 5474 5634
rect 5526 5606 5554 5634
rect 5686 5606 5714 5634
rect 5846 5606 5874 5634
rect 5926 5606 5954 5634
rect 6086 5606 6114 5634
rect 6166 5606 6194 5634
rect 6326 5606 6354 5634
rect 4246 5526 4274 5554
rect 4406 5526 4434 5554
rect 4486 5526 4514 5554
rect 4646 5526 4674 5554
rect 4726 5526 4754 5554
rect 4886 5526 4914 5554
rect 5046 5526 5074 5554
rect 5126 5526 5154 5554
rect 5286 5526 5314 5554
rect 5446 5526 5474 5554
rect 5526 5526 5554 5554
rect 5686 5526 5714 5554
rect 5846 5526 5874 5554
rect 5926 5526 5954 5554
rect 6086 5526 6114 5554
rect 6166 5526 6194 5554
rect 6326 5526 6354 5554
rect 4246 5446 4274 5474
rect 4406 5446 4434 5474
rect 4486 5446 4514 5474
rect 4646 5446 4674 5474
rect 4726 5446 4754 5474
rect 4886 5446 4914 5474
rect 5046 5446 5074 5474
rect 5126 5446 5154 5474
rect 5286 5446 5314 5474
rect 5446 5446 5474 5474
rect 5526 5446 5554 5474
rect 5686 5446 5714 5474
rect 5846 5446 5874 5474
rect 5926 5446 5954 5474
rect 6086 5446 6114 5474
rect 6166 5446 6194 5474
rect 6326 5446 6354 5474
rect 4246 5366 4274 5394
rect 4406 5366 4434 5394
rect 4486 5366 4514 5394
rect 4646 5366 4674 5394
rect 4726 5366 4754 5394
rect 4886 5366 4914 5394
rect 5046 5366 5074 5394
rect 5126 5366 5154 5394
rect 5286 5366 5314 5394
rect 5446 5366 5474 5394
rect 5526 5366 5554 5394
rect 5686 5366 5714 5394
rect 5846 5366 5874 5394
rect 5926 5366 5954 5394
rect 6086 5366 6114 5394
rect 6166 5366 6194 5394
rect 6326 5366 6354 5394
rect 4246 5286 4274 5314
rect 4406 5286 4434 5314
rect 4486 5286 4514 5314
rect 4646 5286 4674 5314
rect 4726 5286 4754 5314
rect 4886 5286 4914 5314
rect 5046 5286 5074 5314
rect 5126 5286 5154 5314
rect 5286 5286 5314 5314
rect 5446 5286 5474 5314
rect 5526 5286 5554 5314
rect 5686 5286 5714 5314
rect 5846 5286 5874 5314
rect 5926 5286 5954 5314
rect 6086 5286 6114 5314
rect 6166 5286 6194 5314
rect 6326 5286 6354 5314
rect 4246 5206 4274 5234
rect 4406 5206 4434 5234
rect 4486 5206 4514 5234
rect 4646 5206 4674 5234
rect 4726 5206 4754 5234
rect 4886 5206 4914 5234
rect 5046 5206 5074 5234
rect 5126 5206 5154 5234
rect 5286 5206 5314 5234
rect 5446 5206 5474 5234
rect 5526 5206 5554 5234
rect 5686 5206 5714 5234
rect 5846 5206 5874 5234
rect 5926 5206 5954 5234
rect 6086 5206 6114 5234
rect 6166 5206 6194 5234
rect 6326 5206 6354 5234
rect 4246 5126 4274 5154
rect 4406 5126 4434 5154
rect 4486 5126 4514 5154
rect 4646 5126 4674 5154
rect 4726 5126 4754 5154
rect 4886 5126 4914 5154
rect 5046 5126 5074 5154
rect 5126 5126 5154 5154
rect 5286 5126 5314 5154
rect 5446 5126 5474 5154
rect 5526 5126 5554 5154
rect 5686 5126 5714 5154
rect 5846 5126 5874 5154
rect 5926 5126 5954 5154
rect 6086 5126 6114 5154
rect 6166 5126 6194 5154
rect 6326 5126 6354 5154
rect 4246 5046 4274 5074
rect 4406 5046 4434 5074
rect 4486 5046 4514 5074
rect 4646 5046 4674 5074
rect 4726 5046 4754 5074
rect 4886 5046 4914 5074
rect 5046 5046 5074 5074
rect 5126 5046 5154 5074
rect 5286 5046 5314 5074
rect 5446 5046 5474 5074
rect 5526 5046 5554 5074
rect 5686 5046 5714 5074
rect 5846 5046 5874 5074
rect 5926 5046 5954 5074
rect 6086 5046 6114 5074
rect 6166 5046 6194 5074
rect 6326 5046 6354 5074
rect 4246 4966 4274 4994
rect 4406 4966 4434 4994
rect 4486 4966 4514 4994
rect 4646 4966 4674 4994
rect 4726 4966 4754 4994
rect 4886 4966 4914 4994
rect 5046 4966 5074 4994
rect 5126 4966 5154 4994
rect 5286 4966 5314 4994
rect 5446 4966 5474 4994
rect 5526 4966 5554 4994
rect 5686 4966 5714 4994
rect 5846 4966 5874 4994
rect 5926 4966 5954 4994
rect 6086 4966 6114 4994
rect 6166 4966 6194 4994
rect 6326 4966 6354 4994
rect 5926 4886 5954 4914
rect 6086 4886 6114 4914
rect 6006 4806 6034 4834
rect 5926 4726 5954 4754
rect 6086 4726 6114 4754
rect 6166 4646 6194 4674
rect 6326 4646 6354 4674
rect 6246 4566 6274 4594
rect 6166 4486 6194 4514
rect 6326 4486 6354 4514
rect 4246 4406 4274 4434
rect 4406 4406 4434 4434
rect 4486 4406 4514 4434
rect 4646 4406 4674 4434
rect 4726 4406 4754 4434
rect 4886 4406 4914 4434
rect 5046 4406 5074 4434
rect 5126 4406 5154 4434
rect 5286 4406 5314 4434
rect 5446 4406 5474 4434
rect 5526 4406 5554 4434
rect 5686 4406 5714 4434
rect 5846 4406 5874 4434
rect 5926 4406 5954 4434
rect 6086 4406 6114 4434
rect 6166 4406 6194 4434
rect 6326 4406 6354 4434
rect 4246 4326 4274 4354
rect 4406 4326 4434 4354
rect 4486 4326 4514 4354
rect 4646 4326 4674 4354
rect 4726 4326 4754 4354
rect 4886 4326 4914 4354
rect 5046 4326 5074 4354
rect 5126 4326 5154 4354
rect 5286 4326 5314 4354
rect 5446 4326 5474 4354
rect 5526 4326 5554 4354
rect 5686 4326 5714 4354
rect 5846 4326 5874 4354
rect 5926 4326 5954 4354
rect 6086 4326 6114 4354
rect 6166 4326 6194 4354
rect 6326 4326 6354 4354
rect 4246 4246 4274 4274
rect 4406 4246 4434 4274
rect 4486 4246 4514 4274
rect 4646 4246 4674 4274
rect 4726 4246 4754 4274
rect 4886 4246 4914 4274
rect 5046 4246 5074 4274
rect 5126 4246 5154 4274
rect 5286 4246 5314 4274
rect 5446 4246 5474 4274
rect 5526 4246 5554 4274
rect 5686 4246 5714 4274
rect 5846 4246 5874 4274
rect 5926 4246 5954 4274
rect 6086 4246 6114 4274
rect 6166 4246 6194 4274
rect 6326 4246 6354 4274
rect 4246 4166 4274 4194
rect 4406 4166 4434 4194
rect 4486 4166 4514 4194
rect 4646 4166 4674 4194
rect 4726 4166 4754 4194
rect 4886 4166 4914 4194
rect 5046 4166 5074 4194
rect 5126 4166 5154 4194
rect 5286 4166 5314 4194
rect 5446 4166 5474 4194
rect 5526 4166 5554 4194
rect 5686 4166 5714 4194
rect 5846 4166 5874 4194
rect 5926 4166 5954 4194
rect 6086 4166 6114 4194
rect 6166 4166 6194 4194
rect 6326 4166 6354 4194
rect 4246 4086 4274 4114
rect 4406 4086 4434 4114
rect 4486 4086 4514 4114
rect 4646 4086 4674 4114
rect 4726 4086 4754 4114
rect 4886 4086 4914 4114
rect 5046 4086 5074 4114
rect 5126 4086 5154 4114
rect 5286 4086 5314 4114
rect 5446 4086 5474 4114
rect 5526 4086 5554 4114
rect 5686 4086 5714 4114
rect 5846 4086 5874 4114
rect 5926 4086 5954 4114
rect 6086 4086 6114 4114
rect 6166 4086 6194 4114
rect 6326 4086 6354 4114
rect 4246 4006 4274 4034
rect 4406 4006 4434 4034
rect 4486 4006 4514 4034
rect 4646 4006 4674 4034
rect 4726 4006 4754 4034
rect 4886 4006 4914 4034
rect 5046 4006 5074 4034
rect 5126 4006 5154 4034
rect 5286 4006 5314 4034
rect 5446 4006 5474 4034
rect 5526 4006 5554 4034
rect 5686 4006 5714 4034
rect 5846 4006 5874 4034
rect 5926 4006 5954 4034
rect 6086 4006 6114 4034
rect 6166 4006 6194 4034
rect 6326 4006 6354 4034
rect 4246 3926 4274 3954
rect 4406 3926 4434 3954
rect 4486 3926 4514 3954
rect 4646 3926 4674 3954
rect 4726 3926 4754 3954
rect 4886 3926 4914 3954
rect 5046 3926 5074 3954
rect 5126 3926 5154 3954
rect 5286 3926 5314 3954
rect 5446 3926 5474 3954
rect 5526 3926 5554 3954
rect 5686 3926 5714 3954
rect 5846 3926 5874 3954
rect 5926 3926 5954 3954
rect 6086 3926 6114 3954
rect 6166 3926 6194 3954
rect 6326 3926 6354 3954
rect 4246 3846 4274 3874
rect 4406 3846 4434 3874
rect 4326 3766 4354 3794
rect 4246 3686 4274 3714
rect 4406 3686 4434 3714
rect 4486 3606 4514 3634
rect 4646 3606 4674 3634
rect 4566 3526 4594 3554
rect 4486 3446 4514 3474
rect 4646 3446 4674 3474
rect 5926 3366 5954 3394
rect 6086 3366 6114 3394
rect 6006 3286 6034 3314
rect 5926 3206 5954 3234
rect 6086 3206 6114 3234
rect 4246 3126 4274 3154
rect 4406 3126 4434 3154
rect 4486 3126 4514 3154
rect 4646 3126 4674 3154
rect 4726 3126 4754 3154
rect 4886 3126 4914 3154
rect 5046 3126 5074 3154
rect 5126 3126 5154 3154
rect 5286 3126 5314 3154
rect 5446 3126 5474 3154
rect 5526 3126 5554 3154
rect 5686 3126 5714 3154
rect 5846 3126 5874 3154
rect 5926 3126 5954 3154
rect 6086 3126 6114 3154
rect 6166 3126 6194 3154
rect 6326 3126 6354 3154
rect 4246 3046 4274 3074
rect 4406 3046 4434 3074
rect 4486 3046 4514 3074
rect 4646 3046 4674 3074
rect 4726 3046 4754 3074
rect 4886 3046 4914 3074
rect 5046 3046 5074 3074
rect 5126 3046 5154 3074
rect 5286 3046 5314 3074
rect 5446 3046 5474 3074
rect 5526 3046 5554 3074
rect 5686 3046 5714 3074
rect 5846 3046 5874 3074
rect 5926 3046 5954 3074
rect 6086 3046 6114 3074
rect 6166 3046 6194 3074
rect 6326 3046 6354 3074
rect 4246 2966 4274 2994
rect 4406 2966 4434 2994
rect 4486 2966 4514 2994
rect 4646 2966 4674 2994
rect 4726 2966 4754 2994
rect 4886 2966 4914 2994
rect 5046 2966 5074 2994
rect 5126 2966 5154 2994
rect 5286 2966 5314 2994
rect 5446 2966 5474 2994
rect 5526 2966 5554 2994
rect 5686 2966 5714 2994
rect 5846 2966 5874 2994
rect 5926 2966 5954 2994
rect 6086 2966 6114 2994
rect 6166 2966 6194 2994
rect 6326 2966 6354 2994
rect 4246 2886 4274 2914
rect 4406 2886 4434 2914
rect 4486 2886 4514 2914
rect 4646 2886 4674 2914
rect 4726 2886 4754 2914
rect 4886 2886 4914 2914
rect 5046 2886 5074 2914
rect 5126 2886 5154 2914
rect 5286 2886 5314 2914
rect 5446 2886 5474 2914
rect 5526 2886 5554 2914
rect 5686 2886 5714 2914
rect 5846 2886 5874 2914
rect 5926 2886 5954 2914
rect 6086 2886 6114 2914
rect 6166 2886 6194 2914
rect 6326 2886 6354 2914
rect 4246 2806 4274 2834
rect 4406 2806 4434 2834
rect 4486 2806 4514 2834
rect 4646 2806 4674 2834
rect 4726 2806 4754 2834
rect 4886 2806 4914 2834
rect 5046 2806 5074 2834
rect 5126 2806 5154 2834
rect 5286 2806 5314 2834
rect 5446 2806 5474 2834
rect 5526 2806 5554 2834
rect 5686 2806 5714 2834
rect 5846 2806 5874 2834
rect 5926 2806 5954 2834
rect 6086 2806 6114 2834
rect 6166 2806 6194 2834
rect 6326 2806 6354 2834
rect 4246 2726 4274 2754
rect 4406 2726 4434 2754
rect 4486 2726 4514 2754
rect 4646 2726 4674 2754
rect 4726 2726 4754 2754
rect 4886 2726 4914 2754
rect 5046 2726 5074 2754
rect 5126 2726 5154 2754
rect 5286 2726 5314 2754
rect 5446 2726 5474 2754
rect 5526 2726 5554 2754
rect 5686 2726 5714 2754
rect 5846 2726 5874 2754
rect 5926 2726 5954 2754
rect 6086 2726 6114 2754
rect 6166 2726 6194 2754
rect 6326 2726 6354 2754
rect 4246 2646 4274 2674
rect 4406 2646 4434 2674
rect 4486 2646 4514 2674
rect 4646 2646 4674 2674
rect 4726 2646 4754 2674
rect 4886 2646 4914 2674
rect 5046 2646 5074 2674
rect 5126 2646 5154 2674
rect 5286 2646 5314 2674
rect 5446 2646 5474 2674
rect 5526 2646 5554 2674
rect 5686 2646 5714 2674
rect 5846 2646 5874 2674
rect 5926 2646 5954 2674
rect 6086 2646 6114 2674
rect 6166 2646 6194 2674
rect 6326 2646 6354 2674
rect 4246 2566 4274 2594
rect 4406 2566 4434 2594
rect 4486 2566 4514 2594
rect 4646 2566 4674 2594
rect 4726 2566 4754 2594
rect 4886 2566 4914 2594
rect 5046 2566 5074 2594
rect 5126 2566 5154 2594
rect 5286 2566 5314 2594
rect 5446 2566 5474 2594
rect 5526 2566 5554 2594
rect 5686 2566 5714 2594
rect 5846 2566 5874 2594
rect 5926 2566 5954 2594
rect 6086 2566 6114 2594
rect 6166 2566 6194 2594
rect 6326 2566 6354 2594
rect 4246 2486 4274 2514
rect 4406 2486 4434 2514
rect 4486 2486 4514 2514
rect 4646 2486 4674 2514
rect 4726 2486 4754 2514
rect 4886 2486 4914 2514
rect 5046 2486 5074 2514
rect 5126 2486 5154 2514
rect 5286 2486 5314 2514
rect 5446 2486 5474 2514
rect 5526 2486 5554 2514
rect 5686 2486 5714 2514
rect 5846 2486 5874 2514
rect 5926 2486 5954 2514
rect 6086 2486 6114 2514
rect 6166 2486 6194 2514
rect 6326 2486 6354 2514
rect 4246 2406 4274 2434
rect 4406 2406 4434 2434
rect 4486 2406 4514 2434
rect 4646 2406 4674 2434
rect 4726 2406 4754 2434
rect 4886 2406 4914 2434
rect 5046 2406 5074 2434
rect 5126 2406 5154 2434
rect 5286 2406 5314 2434
rect 5446 2406 5474 2434
rect 5526 2406 5554 2434
rect 5686 2406 5714 2434
rect 5846 2406 5874 2434
rect 5926 2406 5954 2434
rect 6086 2406 6114 2434
rect 6166 2406 6194 2434
rect 6326 2406 6354 2434
rect 4246 2326 4274 2354
rect 4406 2326 4434 2354
rect 4486 2326 4514 2354
rect 4646 2326 4674 2354
rect 4726 2326 4754 2354
rect 4886 2326 4914 2354
rect 5046 2326 5074 2354
rect 5126 2326 5154 2354
rect 5286 2326 5314 2354
rect 5446 2326 5474 2354
rect 5526 2326 5554 2354
rect 5686 2326 5714 2354
rect 5846 2326 5874 2354
rect 5926 2326 5954 2354
rect 6086 2326 6114 2354
rect 6166 2326 6194 2354
rect 6326 2326 6354 2354
rect 4246 2246 4274 2274
rect 4406 2246 4434 2274
rect 4486 2246 4514 2274
rect 4646 2246 4674 2274
rect 4726 2246 4754 2274
rect 4886 2246 4914 2274
rect 5046 2246 5074 2274
rect 5126 2246 5154 2274
rect 5286 2246 5314 2274
rect 5446 2246 5474 2274
rect 5526 2246 5554 2274
rect 5686 2246 5714 2274
rect 5846 2246 5874 2274
rect 5926 2246 5954 2274
rect 6086 2246 6114 2274
rect 6166 2246 6194 2274
rect 6326 2246 6354 2274
rect 4246 2166 4274 2194
rect 4406 2166 4434 2194
rect 4486 2166 4514 2194
rect 4646 2166 4674 2194
rect 4726 2166 4754 2194
rect 4886 2166 4914 2194
rect 5046 2166 5074 2194
rect 5126 2166 5154 2194
rect 5286 2166 5314 2194
rect 5446 2166 5474 2194
rect 5526 2166 5554 2194
rect 5686 2166 5714 2194
rect 5846 2166 5874 2194
rect 5926 2166 5954 2194
rect 6086 2166 6114 2194
rect 6166 2166 6194 2194
rect 6326 2166 6354 2194
rect 4246 2086 4274 2114
rect 4406 2086 4434 2114
rect 4486 2086 4514 2114
rect 4646 2086 4674 2114
rect 4726 2086 4754 2114
rect 4886 2086 4914 2114
rect 5046 2086 5074 2114
rect 5126 2086 5154 2114
rect 5286 2086 5314 2114
rect 5446 2086 5474 2114
rect 5526 2086 5554 2114
rect 5686 2086 5714 2114
rect 5846 2086 5874 2114
rect 5926 2086 5954 2114
rect 6086 2086 6114 2114
rect 6166 2086 6194 2114
rect 6326 2086 6354 2114
rect 4246 2006 4274 2034
rect 4406 2006 4434 2034
rect 4486 2006 4514 2034
rect 4646 2006 4674 2034
rect 4726 2006 4754 2034
rect 4886 2006 4914 2034
rect 5046 2006 5074 2034
rect 5126 2006 5154 2034
rect 5286 2006 5314 2034
rect 5446 2006 5474 2034
rect 5526 2006 5554 2034
rect 5686 2006 5714 2034
rect 5846 2006 5874 2034
rect 5926 2006 5954 2034
rect 6086 2006 6114 2034
rect 6166 2006 6194 2034
rect 6326 2006 6354 2034
rect 4486 1886 4514 1914
rect 4646 1886 4674 1914
rect 4566 1806 4594 1834
rect 4486 1726 4514 1754
rect 4646 1726 4674 1754
rect 4246 1606 4274 1634
rect 4406 1606 4434 1634
rect 4486 1606 4514 1634
rect 4646 1606 4674 1634
rect 4726 1606 4754 1634
rect 4886 1606 4914 1634
rect 5046 1606 5074 1634
rect 5126 1606 5154 1634
rect 5286 1606 5314 1634
rect 5446 1606 5474 1634
rect 5526 1606 5554 1634
rect 5686 1606 5714 1634
rect 5846 1606 5874 1634
rect 5926 1606 5954 1634
rect 6086 1606 6114 1634
rect 6166 1606 6194 1634
rect 6326 1606 6354 1634
rect 4246 1526 4274 1554
rect 4406 1526 4434 1554
rect 4486 1526 4514 1554
rect 4646 1526 4674 1554
rect 4726 1526 4754 1554
rect 4886 1526 4914 1554
rect 5046 1526 5074 1554
rect 5126 1526 5154 1554
rect 5286 1526 5314 1554
rect 5446 1526 5474 1554
rect 5526 1526 5554 1554
rect 5686 1526 5714 1554
rect 5846 1526 5874 1554
rect 5926 1526 5954 1554
rect 6086 1526 6114 1554
rect 6166 1526 6194 1554
rect 6326 1526 6354 1554
rect 4246 1446 4274 1474
rect 4406 1446 4434 1474
rect 4486 1446 4514 1474
rect 4646 1446 4674 1474
rect 4726 1446 4754 1474
rect 4886 1446 4914 1474
rect 5046 1446 5074 1474
rect 5126 1446 5154 1474
rect 5286 1446 5314 1474
rect 5446 1446 5474 1474
rect 5526 1446 5554 1474
rect 5686 1446 5714 1474
rect 5846 1446 5874 1474
rect 5926 1446 5954 1474
rect 6086 1446 6114 1474
rect 6166 1446 6194 1474
rect 6326 1446 6354 1474
rect 4246 1366 4274 1394
rect 4406 1366 4434 1394
rect 4486 1366 4514 1394
rect 4646 1366 4674 1394
rect 4726 1366 4754 1394
rect 4886 1366 4914 1394
rect 5046 1366 5074 1394
rect 5126 1366 5154 1394
rect 5286 1366 5314 1394
rect 5446 1366 5474 1394
rect 5526 1366 5554 1394
rect 5686 1366 5714 1394
rect 5846 1366 5874 1394
rect 5926 1366 5954 1394
rect 6086 1366 6114 1394
rect 6166 1366 6194 1394
rect 6326 1366 6354 1394
rect 4246 1286 4274 1314
rect 4406 1286 4434 1314
rect 4486 1286 4514 1314
rect 4646 1286 4674 1314
rect 4726 1286 4754 1314
rect 4886 1286 4914 1314
rect 5046 1286 5074 1314
rect 5126 1286 5154 1314
rect 5286 1286 5314 1314
rect 5446 1286 5474 1314
rect 5526 1286 5554 1314
rect 5686 1286 5714 1314
rect 5846 1286 5874 1314
rect 5926 1286 5954 1314
rect 6086 1286 6114 1314
rect 6166 1286 6194 1314
rect 6326 1286 6354 1314
rect 4246 1206 4274 1234
rect 4406 1206 4434 1234
rect 4486 1206 4514 1234
rect 4646 1206 4674 1234
rect 4726 1206 4754 1234
rect 4886 1206 4914 1234
rect 5046 1206 5074 1234
rect 5126 1206 5154 1234
rect 5286 1206 5314 1234
rect 5446 1206 5474 1234
rect 5526 1206 5554 1234
rect 5686 1206 5714 1234
rect 5846 1206 5874 1234
rect 5926 1206 5954 1234
rect 6086 1206 6114 1234
rect 6166 1206 6194 1234
rect 6326 1206 6354 1234
rect 4246 1126 4274 1154
rect 4406 1126 4434 1154
rect 4486 1126 4514 1154
rect 4646 1126 4674 1154
rect 4726 1126 4754 1154
rect 4886 1126 4914 1154
rect 5046 1126 5074 1154
rect 5126 1126 5154 1154
rect 5286 1126 5314 1154
rect 5446 1126 5474 1154
rect 5526 1126 5554 1154
rect 5686 1126 5714 1154
rect 5846 1126 5874 1154
rect 5926 1126 5954 1154
rect 6086 1126 6114 1154
rect 6166 1126 6194 1154
rect 6326 1126 6354 1154
rect 4246 1046 4274 1074
rect 4406 1046 4434 1074
rect 4486 1046 4514 1074
rect 4646 1046 4674 1074
rect 4726 1046 4754 1074
rect 4886 1046 4914 1074
rect 5046 1046 5074 1074
rect 5126 1046 5154 1074
rect 5286 1046 5314 1074
rect 5446 1046 5474 1074
rect 5526 1046 5554 1074
rect 5686 1046 5714 1074
rect 5846 1046 5874 1074
rect 5926 1046 5954 1074
rect 6086 1046 6114 1074
rect 6166 1046 6194 1074
rect 6326 1046 6354 1074
rect 6166 966 6194 994
rect 6326 966 6354 994
rect 6246 886 6274 914
rect 6166 806 6194 834
rect 6326 806 6354 834
rect 4246 726 4274 754
rect 4406 726 4434 754
rect 4486 726 4514 754
rect 4646 726 4674 754
rect 4726 726 4754 754
rect 4886 726 4914 754
rect 5046 726 5074 754
rect 5126 726 5154 754
rect 5286 726 5314 754
rect 5446 726 5474 754
rect 5526 726 5554 754
rect 5686 726 5714 754
rect 5846 726 5874 754
rect 5926 726 5954 754
rect 6086 726 6114 754
rect 6166 726 6194 754
rect 6326 726 6354 754
rect 4246 646 4274 674
rect 4406 646 4434 674
rect 4486 646 4514 674
rect 4646 646 4674 674
rect 4726 646 4754 674
rect 4886 646 4914 674
rect 5046 646 5074 674
rect 5126 646 5154 674
rect 5286 646 5314 674
rect 5446 646 5474 674
rect 5526 646 5554 674
rect 5686 646 5714 674
rect 5846 646 5874 674
rect 5926 646 5954 674
rect 6086 646 6114 674
rect 6166 646 6194 674
rect 6326 646 6354 674
rect 4246 566 4274 594
rect 4406 566 4434 594
rect 4486 566 4514 594
rect 4646 566 4674 594
rect 4726 566 4754 594
rect 4886 566 4914 594
rect 5046 566 5074 594
rect 5126 566 5154 594
rect 5286 566 5314 594
rect 5446 566 5474 594
rect 5526 566 5554 594
rect 5686 566 5714 594
rect 5846 566 5874 594
rect 5926 566 5954 594
rect 6086 566 6114 594
rect 6166 566 6194 594
rect 6326 566 6354 594
rect 4246 446 4274 474
rect 4406 446 4434 474
rect 4326 366 4354 394
rect 4246 286 4274 314
rect 4406 286 4434 314
rect 4246 166 4274 194
rect 4406 166 4434 194
rect 4486 166 4514 194
rect 4646 166 4674 194
rect 4726 166 4754 194
rect 4886 166 4914 194
rect 5046 166 5074 194
rect 5126 166 5154 194
rect 5286 166 5314 194
rect 5446 166 5474 194
rect 5526 166 5554 194
rect 5686 166 5714 194
rect 5846 166 5874 194
rect 5926 166 5954 194
rect 6086 166 6114 194
rect 6166 166 6194 194
rect 6326 166 6354 194
rect 4246 86 4274 114
rect 4406 86 4434 114
rect 4486 86 4514 114
rect 4646 86 4674 114
rect 4726 86 4754 114
rect 4886 86 4914 114
rect 5046 86 5074 114
rect 5126 86 5154 114
rect 5286 86 5314 114
rect 5446 86 5474 114
rect 5526 86 5554 114
rect 5686 86 5714 114
rect 5846 86 5874 114
rect 5926 86 5954 114
rect 6086 86 6114 114
rect 6166 86 6194 114
rect 6326 86 6354 114
rect 4246 6 4274 34
rect 4406 6 4434 34
rect 4486 6 4514 34
rect 4646 6 4674 34
rect 4726 6 4754 34
rect 4886 6 4914 34
rect 5046 6 5074 34
rect 5126 6 5154 34
rect 5286 6 5314 34
rect 5446 6 5474 34
rect 5526 6 5554 34
rect 5686 6 5714 34
rect 5846 6 5874 34
rect 5926 6 5954 34
rect 6086 6 6114 34
rect 6166 6 6194 34
rect 6326 6 6354 34
<< metal3 >>
rect 0 16916 40 16920
rect 0 16884 4 16916
rect 36 16884 40 16916
rect 0 15476 40 16884
rect 0 15444 4 15476
rect 36 15444 40 15476
rect 0 14036 40 15444
rect 0 14004 4 14036
rect 36 14004 40 14036
rect 0 13716 40 14004
rect 80 16836 120 16920
rect 80 16804 84 16836
rect 116 16804 120 16836
rect 80 15556 120 16804
rect 80 15524 84 15556
rect 116 15524 120 15556
rect 80 13956 120 15524
rect 80 13924 84 13956
rect 116 13924 120 13956
rect 80 13796 120 13924
rect 80 13764 84 13796
rect 116 13764 120 13796
rect 80 13760 120 13764
rect 160 16756 200 16920
rect 160 16724 164 16756
rect 196 16724 200 16756
rect 160 13876 200 16724
rect 160 13844 164 13876
rect 196 13844 200 13876
rect 160 13760 200 13844
rect 240 16836 280 16920
rect 240 16804 244 16836
rect 276 16804 280 16836
rect 240 15556 280 16804
rect 240 15524 244 15556
rect 276 15524 280 15556
rect 240 13956 280 15524
rect 240 13924 244 13956
rect 276 13924 280 13956
rect 240 13796 280 13924
rect 240 13764 244 13796
rect 276 13764 280 13796
rect 240 13760 280 13764
rect 320 16916 360 16920
rect 320 16884 324 16916
rect 356 16884 360 16916
rect 320 15476 360 16884
rect 10240 16916 10280 16920
rect 10240 16884 10244 16916
rect 10276 16884 10280 16916
rect 400 16836 440 16840
rect 400 16804 404 16836
rect 436 16804 440 16836
rect 400 15556 440 16804
rect 10160 16836 10200 16840
rect 10160 16804 10164 16836
rect 10196 16804 10200 16836
rect 480 16756 520 16760
rect 480 16724 484 16756
rect 516 16724 520 16756
rect 480 16680 520 16724
rect 1520 16756 1560 16760
rect 1520 16724 1524 16756
rect 1556 16724 1560 16756
rect 1520 16680 1560 16724
rect 480 15600 1560 16680
rect 1600 16756 1640 16760
rect 1600 16724 1604 16756
rect 1636 16724 1640 16756
rect 1600 16680 1640 16724
rect 2640 16756 2680 16760
rect 2640 16724 2644 16756
rect 2676 16724 2680 16756
rect 2640 16680 2680 16724
rect 1600 15600 2680 16680
rect 2720 16756 2760 16760
rect 2720 16724 2724 16756
rect 2756 16724 2760 16756
rect 2720 16680 2760 16724
rect 3760 16756 3800 16760
rect 3760 16724 3764 16756
rect 3796 16724 3800 16756
rect 3760 16680 3800 16724
rect 2720 15600 3800 16680
rect 3840 16756 3880 16760
rect 3840 16724 3844 16756
rect 3876 16724 3880 16756
rect 3840 16680 3880 16724
rect 4880 16756 4920 16760
rect 4880 16724 4884 16756
rect 4916 16724 4920 16756
rect 4880 16680 4920 16724
rect 3840 15600 4920 16680
rect 5680 16756 5720 16760
rect 5680 16724 5684 16756
rect 5716 16724 5720 16756
rect 5680 16680 5720 16724
rect 6720 16756 6760 16760
rect 6720 16724 6724 16756
rect 6756 16724 6760 16756
rect 6720 16680 6760 16724
rect 5680 15600 6760 16680
rect 6800 16756 6840 16760
rect 6800 16724 6804 16756
rect 6836 16724 6840 16756
rect 6800 16680 6840 16724
rect 7840 16756 7880 16760
rect 7840 16724 7844 16756
rect 7876 16724 7880 16756
rect 7840 16680 7880 16724
rect 6800 15600 7880 16680
rect 7920 16756 7960 16760
rect 7920 16724 7924 16756
rect 7956 16724 7960 16756
rect 7920 16680 7960 16724
rect 8960 16756 9000 16760
rect 8960 16724 8964 16756
rect 8996 16724 9000 16756
rect 8960 16680 9000 16724
rect 7920 15600 9000 16680
rect 9040 16756 9080 16760
rect 9040 16724 9044 16756
rect 9076 16724 9080 16756
rect 9040 16680 9080 16724
rect 10080 16756 10120 16760
rect 10080 16724 10084 16756
rect 10116 16724 10120 16756
rect 10080 16680 10120 16724
rect 9040 15600 10120 16680
rect 400 15524 404 15556
rect 436 15524 440 15556
rect 400 15520 440 15524
rect 10160 15556 10200 16804
rect 10160 15524 10164 15556
rect 10196 15524 10200 15556
rect 10160 15520 10200 15524
rect 320 15444 324 15476
rect 356 15444 360 15476
rect 320 14036 360 15444
rect 10240 15476 10280 16884
rect 10240 15444 10244 15476
rect 10276 15444 10280 15476
rect 400 15396 440 15400
rect 400 15364 404 15396
rect 436 15364 440 15396
rect 400 14116 440 15364
rect 4960 15396 5000 15400
rect 4960 15364 4964 15396
rect 4996 15364 5000 15396
rect 480 15316 520 15320
rect 480 15284 484 15316
rect 516 15284 520 15316
rect 480 15240 520 15284
rect 1520 15316 1560 15320
rect 1520 15284 1524 15316
rect 1556 15284 1560 15316
rect 1520 15240 1560 15284
rect 480 14160 1560 15240
rect 1600 15316 1640 15320
rect 1600 15284 1604 15316
rect 1636 15284 1640 15316
rect 1600 15240 1640 15284
rect 2640 15316 2680 15320
rect 2640 15284 2644 15316
rect 2676 15284 2680 15316
rect 2640 15240 2680 15284
rect 1600 14160 2680 15240
rect 2720 15316 2760 15320
rect 2720 15284 2724 15316
rect 2756 15284 2760 15316
rect 2720 15240 2760 15284
rect 3760 15316 3800 15320
rect 3760 15284 3764 15316
rect 3796 15284 3800 15316
rect 3760 15240 3800 15284
rect 2720 14160 3800 15240
rect 3840 15316 3880 15320
rect 3840 15284 3844 15316
rect 3876 15284 3880 15316
rect 3840 15240 3880 15284
rect 4880 15316 4920 15320
rect 4880 15284 4884 15316
rect 4916 15284 4920 15316
rect 4880 15240 4920 15284
rect 3840 14160 4920 15240
rect 400 14084 404 14116
rect 436 14084 440 14116
rect 400 14080 440 14084
rect 4960 14116 5000 15364
rect 4960 14084 4964 14116
rect 4996 14084 5000 14116
rect 4960 14080 5000 14084
rect 320 14004 324 14036
rect 356 14004 360 14036
rect 0 13684 4 13716
rect 36 13684 40 13716
rect 0 13680 40 13684
rect 320 13716 360 14004
rect 5040 14036 5080 15400
rect 5040 14004 5044 14036
rect 5076 14004 5080 14036
rect 320 13684 324 13716
rect 356 13684 360 13716
rect 320 13680 360 13684
rect 4480 13956 4520 13960
rect 4480 13924 4484 13956
rect 4516 13924 4520 13956
rect 4480 13796 4520 13924
rect 4480 13764 4484 13796
rect 4516 13764 4520 13796
rect 4240 13636 4280 13640
rect 4240 13604 4244 13636
rect 4276 13604 4280 13636
rect 4240 13596 4280 13604
rect 4240 13564 4244 13596
rect 4276 13564 4280 13596
rect 4240 13556 4280 13564
rect 4240 13524 4244 13556
rect 4276 13524 4280 13556
rect 4240 13516 4280 13524
rect 4240 13484 4244 13516
rect 4276 13484 4280 13516
rect 4240 13476 4280 13484
rect 4240 13444 4244 13476
rect 4276 13444 4280 13476
rect 4240 12636 4280 13444
rect 4400 13636 4440 13640
rect 4400 13604 4404 13636
rect 4436 13604 4440 13636
rect 4400 13596 4440 13604
rect 4400 13564 4404 13596
rect 4436 13564 4440 13596
rect 4400 13556 4440 13564
rect 4400 13524 4404 13556
rect 4436 13524 4440 13556
rect 4400 13516 4440 13524
rect 4400 13484 4404 13516
rect 4436 13484 4440 13516
rect 4400 13476 4440 13484
rect 4400 13444 4404 13476
rect 4436 13444 4440 13476
rect 4240 12604 4244 12636
rect 4276 12604 4280 12636
rect 4240 12556 4280 12604
rect 4240 12524 4244 12556
rect 4276 12524 4280 12556
rect 4240 12476 4280 12524
rect 4240 12444 4244 12476
rect 4276 12444 4280 12476
rect 4240 12396 4280 12444
rect 4240 12364 4244 12396
rect 4276 12364 4280 12396
rect 4240 12316 4280 12364
rect 4240 12284 4244 12316
rect 4276 12284 4280 12316
rect 4240 12236 4280 12284
rect 4240 12204 4244 12236
rect 4276 12204 4280 12236
rect 4240 12156 4280 12204
rect 4240 12124 4244 12156
rect 4276 12124 4280 12156
rect 4240 11836 4280 12124
rect 4240 11804 4244 11836
rect 4276 11804 4280 11836
rect 4240 11756 4280 11804
rect 4240 11724 4244 11756
rect 4276 11724 4280 11756
rect 4240 11676 4280 11724
rect 4240 11644 4244 11676
rect 4276 11644 4280 11676
rect 4240 11596 4280 11644
rect 4240 11564 4244 11596
rect 4276 11564 4280 11596
rect 4240 11516 4280 11564
rect 4240 11484 4244 11516
rect 4276 11484 4280 11516
rect 4240 11436 4280 11484
rect 4240 11404 4244 11436
rect 4276 11404 4280 11436
rect 4240 10876 4280 11404
rect 4240 10844 4244 10876
rect 4276 10844 4280 10876
rect 4240 10796 4280 10844
rect 4240 10764 4244 10796
rect 4276 10764 4280 10796
rect 4240 10716 4280 10764
rect 4240 10684 4244 10716
rect 4276 10684 4280 10716
rect 4240 10636 4280 10684
rect 4240 10604 4244 10636
rect 4276 10604 4280 10636
rect 4240 10556 4280 10604
rect 4240 10524 4244 10556
rect 4276 10524 4280 10556
rect 4240 10476 4280 10524
rect 4240 10444 4244 10476
rect 4276 10444 4280 10476
rect 4240 10396 4280 10444
rect 4240 10364 4244 10396
rect 4276 10364 4280 10396
rect 4240 10316 4280 10364
rect 4240 10284 4244 10316
rect 4276 10284 4280 10316
rect 4240 10236 4280 10284
rect 4240 10204 4244 10236
rect 4276 10204 4280 10236
rect 4240 10156 4280 10204
rect 4240 10124 4244 10156
rect 4276 10124 4280 10156
rect 4240 10076 4280 10124
rect 4240 10044 4244 10076
rect 4276 10044 4280 10076
rect 4240 9996 4280 10044
rect 4240 9964 4244 9996
rect 4276 9964 4280 9996
rect 4240 9916 4280 9964
rect 4240 9884 4244 9916
rect 4276 9884 4280 9916
rect 4240 9836 4280 9884
rect 4240 9804 4244 9836
rect 4276 9804 4280 9836
rect 4240 9756 4280 9804
rect 4240 9724 4244 9756
rect 4276 9724 4280 9756
rect 4240 9356 4280 9724
rect 4240 9324 4244 9356
rect 4276 9324 4280 9356
rect 4240 9276 4280 9324
rect 4240 9244 4244 9276
rect 4276 9244 4280 9276
rect 4240 9196 4280 9244
rect 4240 9164 4244 9196
rect 4276 9164 4280 9196
rect 4240 8876 4280 9164
rect 4240 8844 4244 8876
rect 4276 8844 4280 8876
rect 4240 8796 4280 8844
rect 4240 8764 4244 8796
rect 4276 8764 4280 8796
rect 4240 8716 4280 8764
rect 4240 8684 4244 8716
rect 4276 8684 4280 8716
rect 4240 8636 4280 8684
rect 4240 8604 4244 8636
rect 4276 8604 4280 8636
rect 4240 8556 4280 8604
rect 4240 8524 4244 8556
rect 4276 8524 4280 8556
rect 4240 7636 4280 8524
rect 4240 7604 4244 7636
rect 4276 7604 4280 7636
rect 4240 7556 4280 7604
rect 4240 7524 4244 7556
rect 4276 7524 4280 7556
rect 4240 7476 4280 7524
rect 4240 7444 4244 7476
rect 4276 7444 4280 7476
rect 4240 7396 4280 7444
rect 4240 7364 4244 7396
rect 4276 7364 4280 7396
rect 4240 7316 4280 7364
rect 4240 7284 4244 7316
rect 4276 7284 4280 7316
rect 4240 7236 4280 7284
rect 4240 7204 4244 7236
rect 4276 7204 4280 7236
rect 4240 7156 4280 7204
rect 4240 7124 4244 7156
rect 4276 7124 4280 7156
rect 4240 7076 4280 7124
rect 4240 7044 4244 7076
rect 4276 7044 4280 7076
rect 4240 6756 4280 7044
rect 4240 6724 4244 6756
rect 4276 6724 4280 6756
rect 4240 6676 4280 6724
rect 4240 6644 4244 6676
rect 4276 6644 4280 6676
rect 4240 6596 4280 6644
rect 4240 6564 4244 6596
rect 4276 6564 4280 6596
rect 4240 6516 4280 6564
rect 4240 6484 4244 6516
rect 4276 6484 4280 6516
rect 4240 6436 4280 6484
rect 4240 6404 4244 6436
rect 4276 6404 4280 6436
rect 4240 6356 4280 6404
rect 4240 6324 4244 6356
rect 4276 6324 4280 6356
rect 4240 5796 4280 6324
rect 4240 5764 4244 5796
rect 4276 5764 4280 5796
rect 4240 5716 4280 5764
rect 4240 5684 4244 5716
rect 4276 5684 4280 5716
rect 4240 5636 4280 5684
rect 4240 5604 4244 5636
rect 4276 5604 4280 5636
rect 4240 5556 4280 5604
rect 4240 5524 4244 5556
rect 4276 5524 4280 5556
rect 4240 5476 4280 5524
rect 4240 5444 4244 5476
rect 4276 5444 4280 5476
rect 4240 5396 4280 5444
rect 4240 5364 4244 5396
rect 4276 5364 4280 5396
rect 4240 5316 4280 5364
rect 4240 5284 4244 5316
rect 4276 5284 4280 5316
rect 4240 5236 4280 5284
rect 4240 5204 4244 5236
rect 4276 5204 4280 5236
rect 4240 5156 4280 5204
rect 4240 5124 4244 5156
rect 4276 5124 4280 5156
rect 4240 5076 4280 5124
rect 4240 5044 4244 5076
rect 4276 5044 4280 5076
rect 4240 4996 4280 5044
rect 4240 4964 4244 4996
rect 4276 4964 4280 4996
rect 4240 4436 4280 4964
rect 4240 4404 4244 4436
rect 4276 4404 4280 4436
rect 4240 4356 4280 4404
rect 4240 4324 4244 4356
rect 4276 4324 4280 4356
rect 4240 4276 4280 4324
rect 4240 4244 4244 4276
rect 4276 4244 4280 4276
rect 4240 4196 4280 4244
rect 4240 4164 4244 4196
rect 4276 4164 4280 4196
rect 4240 4116 4280 4164
rect 4240 4084 4244 4116
rect 4276 4084 4280 4116
rect 4240 4036 4280 4084
rect 4240 4004 4244 4036
rect 4276 4004 4280 4036
rect 4240 3956 4280 4004
rect 4240 3924 4244 3956
rect 4276 3924 4280 3956
rect 4240 3874 4280 3924
rect 4240 3846 4246 3874
rect 4274 3846 4280 3874
rect 4240 3714 4280 3846
rect 4240 3686 4246 3714
rect 4274 3686 4280 3714
rect 4240 3156 4280 3686
rect 4240 3124 4244 3156
rect 4276 3124 4280 3156
rect 4240 3076 4280 3124
rect 4240 3044 4244 3076
rect 4276 3044 4280 3076
rect 4240 2996 4280 3044
rect 4240 2964 4244 2996
rect 4276 2964 4280 2996
rect 4240 2916 4280 2964
rect 4240 2884 4244 2916
rect 4276 2884 4280 2916
rect 4240 2836 4280 2884
rect 4240 2804 4244 2836
rect 4276 2804 4280 2836
rect 4240 2756 4280 2804
rect 4240 2724 4244 2756
rect 4276 2724 4280 2756
rect 4240 2676 4280 2724
rect 4240 2644 4244 2676
rect 4276 2644 4280 2676
rect 4240 2596 4280 2644
rect 4240 2564 4244 2596
rect 4276 2564 4280 2596
rect 4240 2516 4280 2564
rect 4240 2484 4244 2516
rect 4276 2484 4280 2516
rect 4240 2436 4280 2484
rect 4240 2404 4244 2436
rect 4276 2404 4280 2436
rect 4240 2356 4280 2404
rect 4240 2324 4244 2356
rect 4276 2324 4280 2356
rect 4240 2276 4280 2324
rect 4240 2244 4244 2276
rect 4276 2244 4280 2276
rect 4240 2196 4280 2244
rect 4240 2164 4244 2196
rect 4276 2164 4280 2196
rect 4240 2116 4280 2164
rect 4240 2084 4244 2116
rect 4276 2084 4280 2116
rect 4240 2036 4280 2084
rect 4240 2004 4244 2036
rect 4276 2004 4280 2036
rect 4240 1636 4280 2004
rect 4240 1604 4244 1636
rect 4276 1604 4280 1636
rect 4240 1556 4280 1604
rect 4240 1524 4244 1556
rect 4276 1524 4280 1556
rect 4240 1476 4280 1524
rect 4240 1444 4244 1476
rect 4276 1444 4280 1476
rect 4240 1396 4280 1444
rect 4240 1364 4244 1396
rect 4276 1364 4280 1396
rect 4240 1316 4280 1364
rect 4240 1284 4244 1316
rect 4276 1284 4280 1316
rect 4240 1236 4280 1284
rect 4240 1204 4244 1236
rect 4276 1204 4280 1236
rect 4240 1156 4280 1204
rect 4240 1124 4244 1156
rect 4276 1124 4280 1156
rect 4240 1076 4280 1124
rect 4240 1044 4244 1076
rect 4276 1044 4280 1076
rect 4240 756 4280 1044
rect 4240 724 4244 756
rect 4276 724 4280 756
rect 4240 676 4280 724
rect 4240 644 4244 676
rect 4276 644 4280 676
rect 4240 596 4280 644
rect 4240 564 4244 596
rect 4276 564 4280 596
rect 4240 474 4280 564
rect 4240 446 4246 474
rect 4274 446 4280 474
rect 4240 314 4280 446
rect 4240 286 4246 314
rect 4274 286 4280 314
rect 4240 196 4280 286
rect 4240 164 4244 196
rect 4276 164 4280 196
rect 4240 116 4280 164
rect 4240 84 4244 116
rect 4276 84 4280 116
rect 4240 36 4280 84
rect 4240 4 4244 36
rect 4276 4 4280 36
rect 4240 -40 4280 4
rect 4320 3794 4360 12680
rect 4320 3766 4326 3794
rect 4354 3766 4360 3794
rect 4320 394 4360 3766
rect 4320 366 4326 394
rect 4354 366 4360 394
rect 4320 -40 4360 366
rect 4400 12636 4440 13444
rect 4400 12604 4404 12636
rect 4436 12604 4440 12636
rect 4400 12556 4440 12604
rect 4400 12524 4404 12556
rect 4436 12524 4440 12556
rect 4400 12476 4440 12524
rect 4400 12444 4404 12476
rect 4436 12444 4440 12476
rect 4400 12396 4440 12444
rect 4400 12364 4404 12396
rect 4436 12364 4440 12396
rect 4400 12316 4440 12364
rect 4400 12284 4404 12316
rect 4436 12284 4440 12316
rect 4400 12236 4440 12284
rect 4400 12204 4404 12236
rect 4436 12204 4440 12236
rect 4400 12156 4440 12204
rect 4400 12124 4404 12156
rect 4436 12124 4440 12156
rect 4400 11836 4440 12124
rect 4400 11804 4404 11836
rect 4436 11804 4440 11836
rect 4400 11756 4440 11804
rect 4400 11724 4404 11756
rect 4436 11724 4440 11756
rect 4400 11676 4440 11724
rect 4400 11644 4404 11676
rect 4436 11644 4440 11676
rect 4400 11596 4440 11644
rect 4400 11564 4404 11596
rect 4436 11564 4440 11596
rect 4400 11516 4440 11564
rect 4400 11484 4404 11516
rect 4436 11484 4440 11516
rect 4400 11436 4440 11484
rect 4400 11404 4404 11436
rect 4436 11404 4440 11436
rect 4400 10876 4440 11404
rect 4400 10844 4404 10876
rect 4436 10844 4440 10876
rect 4400 10796 4440 10844
rect 4400 10764 4404 10796
rect 4436 10764 4440 10796
rect 4400 10716 4440 10764
rect 4400 10684 4404 10716
rect 4436 10684 4440 10716
rect 4400 10636 4440 10684
rect 4400 10604 4404 10636
rect 4436 10604 4440 10636
rect 4400 10556 4440 10604
rect 4400 10524 4404 10556
rect 4436 10524 4440 10556
rect 4400 10476 4440 10524
rect 4400 10444 4404 10476
rect 4436 10444 4440 10476
rect 4400 10396 4440 10444
rect 4400 10364 4404 10396
rect 4436 10364 4440 10396
rect 4400 10316 4440 10364
rect 4400 10284 4404 10316
rect 4436 10284 4440 10316
rect 4400 10236 4440 10284
rect 4400 10204 4404 10236
rect 4436 10204 4440 10236
rect 4400 10156 4440 10204
rect 4400 10124 4404 10156
rect 4436 10124 4440 10156
rect 4400 10076 4440 10124
rect 4400 10044 4404 10076
rect 4436 10044 4440 10076
rect 4400 9996 4440 10044
rect 4400 9964 4404 9996
rect 4436 9964 4440 9996
rect 4400 9916 4440 9964
rect 4400 9884 4404 9916
rect 4436 9884 4440 9916
rect 4400 9836 4440 9884
rect 4400 9804 4404 9836
rect 4436 9804 4440 9836
rect 4400 9756 4440 9804
rect 4400 9724 4404 9756
rect 4436 9724 4440 9756
rect 4400 9356 4440 9724
rect 4400 9324 4404 9356
rect 4436 9324 4440 9356
rect 4400 9276 4440 9324
rect 4400 9244 4404 9276
rect 4436 9244 4440 9276
rect 4400 9196 4440 9244
rect 4400 9164 4404 9196
rect 4436 9164 4440 9196
rect 4400 8876 4440 9164
rect 4400 8844 4404 8876
rect 4436 8844 4440 8876
rect 4400 8796 4440 8844
rect 4400 8764 4404 8796
rect 4436 8764 4440 8796
rect 4400 8716 4440 8764
rect 4400 8684 4404 8716
rect 4436 8684 4440 8716
rect 4400 8636 4440 8684
rect 4400 8604 4404 8636
rect 4436 8604 4440 8636
rect 4400 8556 4440 8604
rect 4400 8524 4404 8556
rect 4436 8524 4440 8556
rect 4400 7636 4440 8524
rect 4400 7604 4404 7636
rect 4436 7604 4440 7636
rect 4400 7556 4440 7604
rect 4400 7524 4404 7556
rect 4436 7524 4440 7556
rect 4400 7476 4440 7524
rect 4400 7444 4404 7476
rect 4436 7444 4440 7476
rect 4400 7396 4440 7444
rect 4400 7364 4404 7396
rect 4436 7364 4440 7396
rect 4400 7316 4440 7364
rect 4400 7284 4404 7316
rect 4436 7284 4440 7316
rect 4400 7236 4440 7284
rect 4400 7204 4404 7236
rect 4436 7204 4440 7236
rect 4400 7156 4440 7204
rect 4400 7124 4404 7156
rect 4436 7124 4440 7156
rect 4400 7076 4440 7124
rect 4400 7044 4404 7076
rect 4436 7044 4440 7076
rect 4400 6756 4440 7044
rect 4400 6724 4404 6756
rect 4436 6724 4440 6756
rect 4400 6676 4440 6724
rect 4400 6644 4404 6676
rect 4436 6644 4440 6676
rect 4400 6596 4440 6644
rect 4400 6564 4404 6596
rect 4436 6564 4440 6596
rect 4400 6516 4440 6564
rect 4400 6484 4404 6516
rect 4436 6484 4440 6516
rect 4400 6436 4440 6484
rect 4400 6404 4404 6436
rect 4436 6404 4440 6436
rect 4400 6356 4440 6404
rect 4400 6324 4404 6356
rect 4436 6324 4440 6356
rect 4400 5796 4440 6324
rect 4400 5764 4404 5796
rect 4436 5764 4440 5796
rect 4400 5716 4440 5764
rect 4400 5684 4404 5716
rect 4436 5684 4440 5716
rect 4400 5636 4440 5684
rect 4400 5604 4404 5636
rect 4436 5604 4440 5636
rect 4400 5556 4440 5604
rect 4400 5524 4404 5556
rect 4436 5524 4440 5556
rect 4400 5476 4440 5524
rect 4400 5444 4404 5476
rect 4436 5444 4440 5476
rect 4400 5396 4440 5444
rect 4400 5364 4404 5396
rect 4436 5364 4440 5396
rect 4400 5316 4440 5364
rect 4400 5284 4404 5316
rect 4436 5284 4440 5316
rect 4400 5236 4440 5284
rect 4400 5204 4404 5236
rect 4436 5204 4440 5236
rect 4400 5156 4440 5204
rect 4400 5124 4404 5156
rect 4436 5124 4440 5156
rect 4400 5076 4440 5124
rect 4400 5044 4404 5076
rect 4436 5044 4440 5076
rect 4400 4996 4440 5044
rect 4400 4964 4404 4996
rect 4436 4964 4440 4996
rect 4400 4436 4440 4964
rect 4400 4404 4404 4436
rect 4436 4404 4440 4436
rect 4400 4356 4440 4404
rect 4400 4324 4404 4356
rect 4436 4324 4440 4356
rect 4400 4276 4440 4324
rect 4400 4244 4404 4276
rect 4436 4244 4440 4276
rect 4400 4196 4440 4244
rect 4400 4164 4404 4196
rect 4436 4164 4440 4196
rect 4400 4116 4440 4164
rect 4400 4084 4404 4116
rect 4436 4084 4440 4116
rect 4400 4036 4440 4084
rect 4400 4004 4404 4036
rect 4436 4004 4440 4036
rect 4400 3956 4440 4004
rect 4400 3924 4404 3956
rect 4436 3924 4440 3956
rect 4400 3874 4440 3924
rect 4400 3846 4406 3874
rect 4434 3846 4440 3874
rect 4400 3714 4440 3846
rect 4400 3686 4406 3714
rect 4434 3686 4440 3714
rect 4400 3156 4440 3686
rect 4400 3124 4404 3156
rect 4436 3124 4440 3156
rect 4400 3076 4440 3124
rect 4400 3044 4404 3076
rect 4436 3044 4440 3076
rect 4400 2996 4440 3044
rect 4400 2964 4404 2996
rect 4436 2964 4440 2996
rect 4400 2916 4440 2964
rect 4400 2884 4404 2916
rect 4436 2884 4440 2916
rect 4400 2836 4440 2884
rect 4400 2804 4404 2836
rect 4436 2804 4440 2836
rect 4400 2756 4440 2804
rect 4400 2724 4404 2756
rect 4436 2724 4440 2756
rect 4400 2676 4440 2724
rect 4400 2644 4404 2676
rect 4436 2644 4440 2676
rect 4400 2596 4440 2644
rect 4400 2564 4404 2596
rect 4436 2564 4440 2596
rect 4400 2516 4440 2564
rect 4400 2484 4404 2516
rect 4436 2484 4440 2516
rect 4400 2436 4440 2484
rect 4400 2404 4404 2436
rect 4436 2404 4440 2436
rect 4400 2356 4440 2404
rect 4400 2324 4404 2356
rect 4436 2324 4440 2356
rect 4400 2276 4440 2324
rect 4400 2244 4404 2276
rect 4436 2244 4440 2276
rect 4400 2196 4440 2244
rect 4400 2164 4404 2196
rect 4436 2164 4440 2196
rect 4400 2116 4440 2164
rect 4400 2084 4404 2116
rect 4436 2084 4440 2116
rect 4400 2036 4440 2084
rect 4400 2004 4404 2036
rect 4436 2004 4440 2036
rect 4400 1636 4440 2004
rect 4400 1604 4404 1636
rect 4436 1604 4440 1636
rect 4400 1556 4440 1604
rect 4400 1524 4404 1556
rect 4436 1524 4440 1556
rect 4400 1476 4440 1524
rect 4400 1444 4404 1476
rect 4436 1444 4440 1476
rect 4400 1396 4440 1444
rect 4400 1364 4404 1396
rect 4436 1364 4440 1396
rect 4400 1316 4440 1364
rect 4400 1284 4404 1316
rect 4436 1284 4440 1316
rect 4400 1236 4440 1284
rect 4400 1204 4404 1236
rect 4436 1204 4440 1236
rect 4400 1156 4440 1204
rect 4400 1124 4404 1156
rect 4436 1124 4440 1156
rect 4400 1076 4440 1124
rect 4400 1044 4404 1076
rect 4436 1044 4440 1076
rect 4400 756 4440 1044
rect 4400 724 4404 756
rect 4436 724 4440 756
rect 4400 676 4440 724
rect 4400 644 4404 676
rect 4436 644 4440 676
rect 4400 596 4440 644
rect 4400 564 4404 596
rect 4436 564 4440 596
rect 4400 474 4440 564
rect 4400 446 4406 474
rect 4434 446 4440 474
rect 4400 314 4440 446
rect 4400 286 4406 314
rect 4434 286 4440 314
rect 4400 196 4440 286
rect 4400 164 4404 196
rect 4436 164 4440 196
rect 4400 116 4440 164
rect 4400 84 4404 116
rect 4436 84 4440 116
rect 4400 36 4440 84
rect 4400 4 4404 36
rect 4436 4 4440 36
rect 4400 -40 4440 4
rect 4480 13156 4520 13764
rect 4480 13124 4484 13156
rect 4516 13124 4520 13156
rect 4480 13116 4520 13124
rect 4480 13084 4484 13116
rect 4516 13084 4520 13116
rect 4480 13076 4520 13084
rect 4480 13044 4484 13076
rect 4516 13044 4520 13076
rect 4480 13036 4520 13044
rect 4480 13004 4484 13036
rect 4516 13004 4520 13036
rect 4480 12996 4520 13004
rect 4480 12964 4484 12996
rect 4516 12964 4520 12996
rect 4480 12636 4520 12964
rect 4480 12604 4484 12636
rect 4516 12604 4520 12636
rect 4480 12556 4520 12604
rect 4480 12524 4484 12556
rect 4516 12524 4520 12556
rect 4480 12476 4520 12524
rect 4480 12444 4484 12476
rect 4516 12444 4520 12476
rect 4480 12396 4520 12444
rect 4480 12364 4484 12396
rect 4516 12364 4520 12396
rect 4480 12316 4520 12364
rect 4480 12284 4484 12316
rect 4516 12284 4520 12316
rect 4480 12236 4520 12284
rect 4480 12204 4484 12236
rect 4516 12204 4520 12236
rect 4480 12156 4520 12204
rect 4480 12124 4484 12156
rect 4516 12124 4520 12156
rect 4480 12074 4520 12124
rect 4480 12046 4486 12074
rect 4514 12046 4520 12074
rect 4480 11914 4520 12046
rect 4480 11886 4486 11914
rect 4514 11886 4520 11914
rect 4480 11836 4520 11886
rect 4480 11804 4484 11836
rect 4516 11804 4520 11836
rect 4480 11756 4520 11804
rect 4480 11724 4484 11756
rect 4516 11724 4520 11756
rect 4480 11676 4520 11724
rect 4480 11644 4484 11676
rect 4516 11644 4520 11676
rect 4480 11596 4520 11644
rect 4480 11564 4484 11596
rect 4516 11564 4520 11596
rect 4480 11516 4520 11564
rect 4480 11484 4484 11516
rect 4516 11484 4520 11516
rect 4480 11436 4520 11484
rect 4480 11404 4484 11436
rect 4516 11404 4520 11436
rect 4480 10876 4520 11404
rect 4480 10844 4484 10876
rect 4516 10844 4520 10876
rect 4480 10796 4520 10844
rect 4480 10764 4484 10796
rect 4516 10764 4520 10796
rect 4480 10716 4520 10764
rect 4480 10684 4484 10716
rect 4516 10684 4520 10716
rect 4480 10636 4520 10684
rect 4480 10604 4484 10636
rect 4516 10604 4520 10636
rect 4480 10556 4520 10604
rect 4480 10524 4484 10556
rect 4516 10524 4520 10556
rect 4480 10476 4520 10524
rect 4480 10444 4484 10476
rect 4516 10444 4520 10476
rect 4480 10396 4520 10444
rect 4480 10364 4484 10396
rect 4516 10364 4520 10396
rect 4480 10316 4520 10364
rect 4480 10284 4484 10316
rect 4516 10284 4520 10316
rect 4480 10236 4520 10284
rect 4480 10204 4484 10236
rect 4516 10204 4520 10236
rect 4480 10156 4520 10204
rect 4480 10124 4484 10156
rect 4516 10124 4520 10156
rect 4480 10076 4520 10124
rect 4480 10044 4484 10076
rect 4516 10044 4520 10076
rect 4480 9996 4520 10044
rect 4480 9964 4484 9996
rect 4516 9964 4520 9996
rect 4480 9916 4520 9964
rect 4480 9884 4484 9916
rect 4516 9884 4520 9916
rect 4480 9836 4520 9884
rect 4480 9804 4484 9836
rect 4516 9804 4520 9836
rect 4480 9756 4520 9804
rect 4480 9724 4484 9756
rect 4516 9724 4520 9756
rect 4480 9634 4520 9724
rect 4480 9606 4486 9634
rect 4514 9606 4520 9634
rect 4480 9474 4520 9606
rect 4480 9446 4486 9474
rect 4514 9446 4520 9474
rect 4480 9356 4520 9446
rect 4480 9324 4484 9356
rect 4516 9324 4520 9356
rect 4480 9276 4520 9324
rect 4480 9244 4484 9276
rect 4516 9244 4520 9276
rect 4480 9196 4520 9244
rect 4480 9164 4484 9196
rect 4516 9164 4520 9196
rect 4480 8876 4520 9164
rect 4480 8844 4484 8876
rect 4516 8844 4520 8876
rect 4480 8796 4520 8844
rect 4480 8764 4484 8796
rect 4516 8764 4520 8796
rect 4480 8716 4520 8764
rect 4480 8684 4484 8716
rect 4516 8684 4520 8716
rect 4480 8636 4520 8684
rect 4480 8604 4484 8636
rect 4516 8604 4520 8636
rect 4480 8556 4520 8604
rect 4480 8524 4484 8556
rect 4516 8524 4520 8556
rect 4480 7636 4520 8524
rect 4480 7604 4484 7636
rect 4516 7604 4520 7636
rect 4480 7556 4520 7604
rect 4480 7524 4484 7556
rect 4516 7524 4520 7556
rect 4480 7476 4520 7524
rect 4480 7444 4484 7476
rect 4516 7444 4520 7476
rect 4480 7396 4520 7444
rect 4480 7364 4484 7396
rect 4516 7364 4520 7396
rect 4480 7316 4520 7364
rect 4480 7284 4484 7316
rect 4516 7284 4520 7316
rect 4480 7236 4520 7284
rect 4480 7204 4484 7236
rect 4516 7204 4520 7236
rect 4480 7156 4520 7204
rect 4480 7124 4484 7156
rect 4516 7124 4520 7156
rect 4480 7076 4520 7124
rect 4480 7044 4484 7076
rect 4516 7044 4520 7076
rect 4480 6994 4520 7044
rect 4480 6966 4486 6994
rect 4514 6966 4520 6994
rect 4480 6834 4520 6966
rect 4480 6806 4486 6834
rect 4514 6806 4520 6834
rect 4480 6756 4520 6806
rect 4480 6724 4484 6756
rect 4516 6724 4520 6756
rect 4480 6676 4520 6724
rect 4480 6644 4484 6676
rect 4516 6644 4520 6676
rect 4480 6596 4520 6644
rect 4480 6564 4484 6596
rect 4516 6564 4520 6596
rect 4480 6516 4520 6564
rect 4480 6484 4484 6516
rect 4516 6484 4520 6516
rect 4480 6436 4520 6484
rect 4480 6404 4484 6436
rect 4516 6404 4520 6436
rect 4480 6356 4520 6404
rect 4480 6324 4484 6356
rect 4516 6324 4520 6356
rect 4480 5796 4520 6324
rect 4480 5764 4484 5796
rect 4516 5764 4520 5796
rect 4480 5716 4520 5764
rect 4480 5684 4484 5716
rect 4516 5684 4520 5716
rect 4480 5636 4520 5684
rect 4480 5604 4484 5636
rect 4516 5604 4520 5636
rect 4480 5556 4520 5604
rect 4480 5524 4484 5556
rect 4516 5524 4520 5556
rect 4480 5476 4520 5524
rect 4480 5444 4484 5476
rect 4516 5444 4520 5476
rect 4480 5396 4520 5444
rect 4480 5364 4484 5396
rect 4516 5364 4520 5396
rect 4480 5316 4520 5364
rect 4480 5284 4484 5316
rect 4516 5284 4520 5316
rect 4480 5236 4520 5284
rect 4480 5204 4484 5236
rect 4516 5204 4520 5236
rect 4480 5156 4520 5204
rect 4480 5124 4484 5156
rect 4516 5124 4520 5156
rect 4480 5076 4520 5124
rect 4480 5044 4484 5076
rect 4516 5044 4520 5076
rect 4480 4996 4520 5044
rect 4480 4964 4484 4996
rect 4516 4964 4520 4996
rect 4480 4436 4520 4964
rect 4480 4404 4484 4436
rect 4516 4404 4520 4436
rect 4480 4356 4520 4404
rect 4480 4324 4484 4356
rect 4516 4324 4520 4356
rect 4480 4276 4520 4324
rect 4480 4244 4484 4276
rect 4516 4244 4520 4276
rect 4480 4196 4520 4244
rect 4480 4164 4484 4196
rect 4516 4164 4520 4196
rect 4480 4116 4520 4164
rect 4480 4084 4484 4116
rect 4516 4084 4520 4116
rect 4480 4036 4520 4084
rect 4480 4004 4484 4036
rect 4516 4004 4520 4036
rect 4480 3956 4520 4004
rect 4480 3924 4484 3956
rect 4516 3924 4520 3956
rect 4480 3634 4520 3924
rect 4480 3606 4486 3634
rect 4514 3606 4520 3634
rect 4480 3474 4520 3606
rect 4480 3446 4486 3474
rect 4514 3446 4520 3474
rect 4480 3156 4520 3446
rect 4480 3124 4484 3156
rect 4516 3124 4520 3156
rect 4480 3076 4520 3124
rect 4480 3044 4484 3076
rect 4516 3044 4520 3076
rect 4480 2996 4520 3044
rect 4480 2964 4484 2996
rect 4516 2964 4520 2996
rect 4480 2916 4520 2964
rect 4480 2884 4484 2916
rect 4516 2884 4520 2916
rect 4480 2836 4520 2884
rect 4480 2804 4484 2836
rect 4516 2804 4520 2836
rect 4480 2756 4520 2804
rect 4480 2724 4484 2756
rect 4516 2724 4520 2756
rect 4480 2676 4520 2724
rect 4480 2644 4484 2676
rect 4516 2644 4520 2676
rect 4480 2596 4520 2644
rect 4480 2564 4484 2596
rect 4516 2564 4520 2596
rect 4480 2516 4520 2564
rect 4480 2484 4484 2516
rect 4516 2484 4520 2516
rect 4480 2436 4520 2484
rect 4480 2404 4484 2436
rect 4516 2404 4520 2436
rect 4480 2356 4520 2404
rect 4480 2324 4484 2356
rect 4516 2324 4520 2356
rect 4480 2276 4520 2324
rect 4480 2244 4484 2276
rect 4516 2244 4520 2276
rect 4480 2196 4520 2244
rect 4480 2164 4484 2196
rect 4516 2164 4520 2196
rect 4480 2116 4520 2164
rect 4480 2084 4484 2116
rect 4516 2084 4520 2116
rect 4480 2036 4520 2084
rect 4480 2004 4484 2036
rect 4516 2004 4520 2036
rect 4480 1914 4520 2004
rect 4480 1886 4486 1914
rect 4514 1886 4520 1914
rect 4480 1754 4520 1886
rect 4480 1726 4486 1754
rect 4514 1726 4520 1754
rect 4480 1636 4520 1726
rect 4480 1604 4484 1636
rect 4516 1604 4520 1636
rect 4480 1556 4520 1604
rect 4480 1524 4484 1556
rect 4516 1524 4520 1556
rect 4480 1476 4520 1524
rect 4480 1444 4484 1476
rect 4516 1444 4520 1476
rect 4480 1396 4520 1444
rect 4480 1364 4484 1396
rect 4516 1364 4520 1396
rect 4480 1316 4520 1364
rect 4480 1284 4484 1316
rect 4516 1284 4520 1316
rect 4480 1236 4520 1284
rect 4480 1204 4484 1236
rect 4516 1204 4520 1236
rect 4480 1156 4520 1204
rect 4480 1124 4484 1156
rect 4516 1124 4520 1156
rect 4480 1076 4520 1124
rect 4480 1044 4484 1076
rect 4516 1044 4520 1076
rect 4480 756 4520 1044
rect 4480 724 4484 756
rect 4516 724 4520 756
rect 4480 676 4520 724
rect 4480 644 4484 676
rect 4516 644 4520 676
rect 4480 596 4520 644
rect 4480 564 4484 596
rect 4516 564 4520 596
rect 4480 196 4520 564
rect 4480 164 4484 196
rect 4516 164 4520 196
rect 4480 116 4520 164
rect 4480 84 4484 116
rect 4516 84 4520 116
rect 4480 36 4520 84
rect 4480 4 4484 36
rect 4516 4 4520 36
rect 4480 -40 4520 4
rect 4560 13876 4600 13960
rect 4560 13844 4564 13876
rect 4596 13844 4600 13876
rect 4560 11994 4600 13844
rect 4560 11966 4566 11994
rect 4594 11966 4600 11994
rect 4560 9554 4600 11966
rect 4560 9526 4566 9554
rect 4594 9526 4600 9554
rect 4560 6914 4600 9526
rect 4560 6886 4566 6914
rect 4594 6886 4600 6914
rect 4560 3554 4600 6886
rect 4560 3526 4566 3554
rect 4594 3526 4600 3554
rect 4560 1834 4600 3526
rect 4560 1806 4566 1834
rect 4594 1806 4600 1834
rect 4560 -40 4600 1806
rect 4640 13956 4680 13960
rect 4640 13924 4644 13956
rect 4676 13924 4680 13956
rect 4640 13796 4680 13924
rect 4640 13764 4644 13796
rect 4676 13764 4680 13796
rect 4640 13156 4680 13764
rect 5040 13716 5080 14004
rect 5040 13684 5044 13716
rect 5076 13684 5080 13716
rect 4640 13124 4644 13156
rect 4676 13124 4680 13156
rect 4640 13116 4680 13124
rect 4640 13084 4644 13116
rect 4676 13084 4680 13116
rect 4640 13076 4680 13084
rect 4640 13044 4644 13076
rect 4676 13044 4680 13076
rect 4640 13036 4680 13044
rect 4640 13004 4644 13036
rect 4676 13004 4680 13036
rect 4640 12996 4680 13004
rect 4640 12964 4644 12996
rect 4676 12964 4680 12996
rect 4640 12636 4680 12964
rect 4640 12604 4644 12636
rect 4676 12604 4680 12636
rect 4640 12556 4680 12604
rect 4640 12524 4644 12556
rect 4676 12524 4680 12556
rect 4640 12476 4680 12524
rect 4640 12444 4644 12476
rect 4676 12444 4680 12476
rect 4640 12396 4680 12444
rect 4640 12364 4644 12396
rect 4676 12364 4680 12396
rect 4640 12316 4680 12364
rect 4640 12284 4644 12316
rect 4676 12284 4680 12316
rect 4640 12236 4680 12284
rect 4640 12204 4644 12236
rect 4676 12204 4680 12236
rect 4640 12156 4680 12204
rect 4640 12124 4644 12156
rect 4676 12124 4680 12156
rect 4640 12074 4680 12124
rect 4640 12046 4646 12074
rect 4674 12046 4680 12074
rect 4640 11914 4680 12046
rect 4640 11886 4646 11914
rect 4674 11886 4680 11914
rect 4640 11836 4680 11886
rect 4640 11804 4644 11836
rect 4676 11804 4680 11836
rect 4640 11756 4680 11804
rect 4640 11724 4644 11756
rect 4676 11724 4680 11756
rect 4640 11676 4680 11724
rect 4640 11644 4644 11676
rect 4676 11644 4680 11676
rect 4640 11596 4680 11644
rect 4640 11564 4644 11596
rect 4676 11564 4680 11596
rect 4640 11516 4680 11564
rect 4640 11484 4644 11516
rect 4676 11484 4680 11516
rect 4640 11436 4680 11484
rect 4640 11404 4644 11436
rect 4676 11404 4680 11436
rect 4640 10876 4680 11404
rect 4640 10844 4644 10876
rect 4676 10844 4680 10876
rect 4640 10796 4680 10844
rect 4640 10764 4644 10796
rect 4676 10764 4680 10796
rect 4640 10716 4680 10764
rect 4640 10684 4644 10716
rect 4676 10684 4680 10716
rect 4640 10636 4680 10684
rect 4640 10604 4644 10636
rect 4676 10604 4680 10636
rect 4640 10556 4680 10604
rect 4640 10524 4644 10556
rect 4676 10524 4680 10556
rect 4640 10476 4680 10524
rect 4640 10444 4644 10476
rect 4676 10444 4680 10476
rect 4640 10396 4680 10444
rect 4640 10364 4644 10396
rect 4676 10364 4680 10396
rect 4640 10316 4680 10364
rect 4640 10284 4644 10316
rect 4676 10284 4680 10316
rect 4640 10236 4680 10284
rect 4640 10204 4644 10236
rect 4676 10204 4680 10236
rect 4640 10156 4680 10204
rect 4640 10124 4644 10156
rect 4676 10124 4680 10156
rect 4640 10076 4680 10124
rect 4640 10044 4644 10076
rect 4676 10044 4680 10076
rect 4640 9996 4680 10044
rect 4640 9964 4644 9996
rect 4676 9964 4680 9996
rect 4640 9916 4680 9964
rect 4640 9884 4644 9916
rect 4676 9884 4680 9916
rect 4640 9836 4680 9884
rect 4640 9804 4644 9836
rect 4676 9804 4680 9836
rect 4640 9756 4680 9804
rect 4640 9724 4644 9756
rect 4676 9724 4680 9756
rect 4640 9634 4680 9724
rect 4640 9606 4646 9634
rect 4674 9606 4680 9634
rect 4640 9474 4680 9606
rect 4640 9446 4646 9474
rect 4674 9446 4680 9474
rect 4640 9356 4680 9446
rect 4640 9324 4644 9356
rect 4676 9324 4680 9356
rect 4640 9276 4680 9324
rect 4640 9244 4644 9276
rect 4676 9244 4680 9276
rect 4640 9196 4680 9244
rect 4640 9164 4644 9196
rect 4676 9164 4680 9196
rect 4640 8876 4680 9164
rect 4640 8844 4644 8876
rect 4676 8844 4680 8876
rect 4640 8796 4680 8844
rect 4640 8764 4644 8796
rect 4676 8764 4680 8796
rect 4640 8716 4680 8764
rect 4640 8684 4644 8716
rect 4676 8684 4680 8716
rect 4640 8636 4680 8684
rect 4640 8604 4644 8636
rect 4676 8604 4680 8636
rect 4640 8556 4680 8604
rect 4640 8524 4644 8556
rect 4676 8524 4680 8556
rect 4640 7636 4680 8524
rect 4640 7604 4644 7636
rect 4676 7604 4680 7636
rect 4640 7556 4680 7604
rect 4640 7524 4644 7556
rect 4676 7524 4680 7556
rect 4640 7476 4680 7524
rect 4640 7444 4644 7476
rect 4676 7444 4680 7476
rect 4640 7396 4680 7444
rect 4640 7364 4644 7396
rect 4676 7364 4680 7396
rect 4640 7316 4680 7364
rect 4640 7284 4644 7316
rect 4676 7284 4680 7316
rect 4640 7236 4680 7284
rect 4640 7204 4644 7236
rect 4676 7204 4680 7236
rect 4640 7156 4680 7204
rect 4640 7124 4644 7156
rect 4676 7124 4680 7156
rect 4640 7076 4680 7124
rect 4640 7044 4644 7076
rect 4676 7044 4680 7076
rect 4640 6994 4680 7044
rect 4640 6966 4646 6994
rect 4674 6966 4680 6994
rect 4640 6834 4680 6966
rect 4640 6806 4646 6834
rect 4674 6806 4680 6834
rect 4640 6756 4680 6806
rect 4640 6724 4644 6756
rect 4676 6724 4680 6756
rect 4640 6676 4680 6724
rect 4640 6644 4644 6676
rect 4676 6644 4680 6676
rect 4640 6596 4680 6644
rect 4640 6564 4644 6596
rect 4676 6564 4680 6596
rect 4640 6516 4680 6564
rect 4640 6484 4644 6516
rect 4676 6484 4680 6516
rect 4640 6436 4680 6484
rect 4640 6404 4644 6436
rect 4676 6404 4680 6436
rect 4640 6356 4680 6404
rect 4640 6324 4644 6356
rect 4676 6324 4680 6356
rect 4640 5796 4680 6324
rect 4640 5764 4644 5796
rect 4676 5764 4680 5796
rect 4640 5716 4680 5764
rect 4640 5684 4644 5716
rect 4676 5684 4680 5716
rect 4640 5636 4680 5684
rect 4640 5604 4644 5636
rect 4676 5604 4680 5636
rect 4640 5556 4680 5604
rect 4640 5524 4644 5556
rect 4676 5524 4680 5556
rect 4640 5476 4680 5524
rect 4640 5444 4644 5476
rect 4676 5444 4680 5476
rect 4640 5396 4680 5444
rect 4640 5364 4644 5396
rect 4676 5364 4680 5396
rect 4640 5316 4680 5364
rect 4640 5284 4644 5316
rect 4676 5284 4680 5316
rect 4640 5236 4680 5284
rect 4640 5204 4644 5236
rect 4676 5204 4680 5236
rect 4640 5156 4680 5204
rect 4640 5124 4644 5156
rect 4676 5124 4680 5156
rect 4640 5076 4680 5124
rect 4640 5044 4644 5076
rect 4676 5044 4680 5076
rect 4640 4996 4680 5044
rect 4640 4964 4644 4996
rect 4676 4964 4680 4996
rect 4640 4436 4680 4964
rect 4640 4404 4644 4436
rect 4676 4404 4680 4436
rect 4640 4356 4680 4404
rect 4640 4324 4644 4356
rect 4676 4324 4680 4356
rect 4640 4276 4680 4324
rect 4640 4244 4644 4276
rect 4676 4244 4680 4276
rect 4640 4196 4680 4244
rect 4640 4164 4644 4196
rect 4676 4164 4680 4196
rect 4640 4116 4680 4164
rect 4640 4084 4644 4116
rect 4676 4084 4680 4116
rect 4640 4036 4680 4084
rect 4640 4004 4644 4036
rect 4676 4004 4680 4036
rect 4640 3956 4680 4004
rect 4640 3924 4644 3956
rect 4676 3924 4680 3956
rect 4640 3634 4680 3924
rect 4640 3606 4646 3634
rect 4674 3606 4680 3634
rect 4640 3474 4680 3606
rect 4640 3446 4646 3474
rect 4674 3446 4680 3474
rect 4640 3156 4680 3446
rect 4640 3124 4644 3156
rect 4676 3124 4680 3156
rect 4640 3076 4680 3124
rect 4640 3044 4644 3076
rect 4676 3044 4680 3076
rect 4640 2996 4680 3044
rect 4640 2964 4644 2996
rect 4676 2964 4680 2996
rect 4640 2916 4680 2964
rect 4640 2884 4644 2916
rect 4676 2884 4680 2916
rect 4640 2836 4680 2884
rect 4640 2804 4644 2836
rect 4676 2804 4680 2836
rect 4640 2756 4680 2804
rect 4640 2724 4644 2756
rect 4676 2724 4680 2756
rect 4640 2676 4680 2724
rect 4640 2644 4644 2676
rect 4676 2644 4680 2676
rect 4640 2596 4680 2644
rect 4640 2564 4644 2596
rect 4676 2564 4680 2596
rect 4640 2516 4680 2564
rect 4640 2484 4644 2516
rect 4676 2484 4680 2516
rect 4640 2436 4680 2484
rect 4640 2404 4644 2436
rect 4676 2404 4680 2436
rect 4640 2356 4680 2404
rect 4640 2324 4644 2356
rect 4676 2324 4680 2356
rect 4640 2276 4680 2324
rect 4640 2244 4644 2276
rect 4676 2244 4680 2276
rect 4640 2196 4680 2244
rect 4640 2164 4644 2196
rect 4676 2164 4680 2196
rect 4640 2116 4680 2164
rect 4640 2084 4644 2116
rect 4676 2084 4680 2116
rect 4640 2036 4680 2084
rect 4640 2004 4644 2036
rect 4676 2004 4680 2036
rect 4640 1914 4680 2004
rect 4640 1886 4646 1914
rect 4674 1886 4680 1914
rect 4640 1754 4680 1886
rect 4640 1726 4646 1754
rect 4674 1726 4680 1754
rect 4640 1636 4680 1726
rect 4640 1604 4644 1636
rect 4676 1604 4680 1636
rect 4640 1556 4680 1604
rect 4640 1524 4644 1556
rect 4676 1524 4680 1556
rect 4640 1476 4680 1524
rect 4640 1444 4644 1476
rect 4676 1444 4680 1476
rect 4640 1396 4680 1444
rect 4640 1364 4644 1396
rect 4676 1364 4680 1396
rect 4640 1316 4680 1364
rect 4640 1284 4644 1316
rect 4676 1284 4680 1316
rect 4640 1236 4680 1284
rect 4640 1204 4644 1236
rect 4676 1204 4680 1236
rect 4640 1156 4680 1204
rect 4640 1124 4644 1156
rect 4676 1124 4680 1156
rect 4640 1076 4680 1124
rect 4640 1044 4644 1076
rect 4676 1044 4680 1076
rect 4640 756 4680 1044
rect 4640 724 4644 756
rect 4676 724 4680 756
rect 4640 676 4680 724
rect 4640 644 4644 676
rect 4676 644 4680 676
rect 4640 596 4680 644
rect 4640 564 4644 596
rect 4676 564 4680 596
rect 4640 196 4680 564
rect 4640 164 4644 196
rect 4676 164 4680 196
rect 4640 116 4680 164
rect 4640 84 4644 116
rect 4676 84 4680 116
rect 4640 36 4680 84
rect 4640 4 4644 36
rect 4676 4 4680 36
rect 4640 -40 4680 4
rect 4720 13396 4760 13400
rect 4720 13364 4724 13396
rect 4756 13364 4760 13396
rect 4720 13356 4760 13364
rect 4720 13324 4724 13356
rect 4756 13324 4760 13356
rect 4720 13316 4760 13324
rect 4720 13284 4724 13316
rect 4756 13284 4760 13316
rect 4720 13276 4760 13284
rect 4720 13244 4724 13276
rect 4756 13244 4760 13276
rect 4720 13236 4760 13244
rect 4720 13204 4724 13236
rect 4756 13204 4760 13236
rect 4720 12636 4760 13204
rect 4880 13396 4920 13400
rect 4880 13364 4884 13396
rect 4916 13364 4920 13396
rect 4880 13356 4920 13364
rect 4880 13324 4884 13356
rect 4916 13324 4920 13356
rect 4880 13316 4920 13324
rect 4880 13284 4884 13316
rect 4916 13284 4920 13316
rect 4880 13276 4920 13284
rect 4880 13244 4884 13276
rect 4916 13244 4920 13276
rect 4880 13236 4920 13244
rect 4880 13204 4884 13236
rect 4916 13204 4920 13236
rect 4720 12604 4724 12636
rect 4756 12604 4760 12636
rect 4720 12556 4760 12604
rect 4720 12524 4724 12556
rect 4756 12524 4760 12556
rect 4720 12476 4760 12524
rect 4720 12444 4724 12476
rect 4756 12444 4760 12476
rect 4720 12396 4760 12444
rect 4720 12364 4724 12396
rect 4756 12364 4760 12396
rect 4720 12316 4760 12364
rect 4720 12284 4724 12316
rect 4756 12284 4760 12316
rect 4720 12236 4760 12284
rect 4720 12204 4724 12236
rect 4756 12204 4760 12236
rect 4720 12156 4760 12204
rect 4720 12124 4724 12156
rect 4756 12124 4760 12156
rect 4720 11836 4760 12124
rect 4720 11804 4724 11836
rect 4756 11804 4760 11836
rect 4720 11756 4760 11804
rect 4720 11724 4724 11756
rect 4756 11724 4760 11756
rect 4720 11676 4760 11724
rect 4720 11644 4724 11676
rect 4756 11644 4760 11676
rect 4720 11596 4760 11644
rect 4720 11564 4724 11596
rect 4756 11564 4760 11596
rect 4720 11516 4760 11564
rect 4720 11484 4724 11516
rect 4756 11484 4760 11516
rect 4720 11436 4760 11484
rect 4720 11404 4724 11436
rect 4756 11404 4760 11436
rect 4720 10876 4760 11404
rect 4720 10844 4724 10876
rect 4756 10844 4760 10876
rect 4720 10796 4760 10844
rect 4720 10764 4724 10796
rect 4756 10764 4760 10796
rect 4720 10716 4760 10764
rect 4720 10684 4724 10716
rect 4756 10684 4760 10716
rect 4720 10636 4760 10684
rect 4720 10604 4724 10636
rect 4756 10604 4760 10636
rect 4720 10556 4760 10604
rect 4720 10524 4724 10556
rect 4756 10524 4760 10556
rect 4720 10476 4760 10524
rect 4720 10444 4724 10476
rect 4756 10444 4760 10476
rect 4720 10396 4760 10444
rect 4720 10364 4724 10396
rect 4756 10364 4760 10396
rect 4720 10316 4760 10364
rect 4720 10284 4724 10316
rect 4756 10284 4760 10316
rect 4720 10236 4760 10284
rect 4720 10204 4724 10236
rect 4756 10204 4760 10236
rect 4720 10156 4760 10204
rect 4720 10124 4724 10156
rect 4756 10124 4760 10156
rect 4720 10076 4760 10124
rect 4720 10044 4724 10076
rect 4756 10044 4760 10076
rect 4720 9996 4760 10044
rect 4720 9964 4724 9996
rect 4756 9964 4760 9996
rect 4720 9916 4760 9964
rect 4720 9884 4724 9916
rect 4756 9884 4760 9916
rect 4720 9836 4760 9884
rect 4720 9804 4724 9836
rect 4756 9804 4760 9836
rect 4720 9756 4760 9804
rect 4720 9724 4724 9756
rect 4756 9724 4760 9756
rect 4720 9356 4760 9724
rect 4720 9324 4724 9356
rect 4756 9324 4760 9356
rect 4720 9276 4760 9324
rect 4720 9244 4724 9276
rect 4756 9244 4760 9276
rect 4720 9196 4760 9244
rect 4720 9164 4724 9196
rect 4756 9164 4760 9196
rect 4720 8876 4760 9164
rect 4720 8844 4724 8876
rect 4756 8844 4760 8876
rect 4720 8796 4760 8844
rect 4720 8764 4724 8796
rect 4756 8764 4760 8796
rect 4720 8716 4760 8764
rect 4720 8684 4724 8716
rect 4756 8684 4760 8716
rect 4720 8636 4760 8684
rect 4720 8604 4724 8636
rect 4756 8604 4760 8636
rect 4720 8556 4760 8604
rect 4720 8524 4724 8556
rect 4756 8524 4760 8556
rect 4720 7636 4760 8524
rect 4720 7604 4724 7636
rect 4756 7604 4760 7636
rect 4720 7556 4760 7604
rect 4720 7524 4724 7556
rect 4756 7524 4760 7556
rect 4720 7476 4760 7524
rect 4720 7444 4724 7476
rect 4756 7444 4760 7476
rect 4720 7396 4760 7444
rect 4720 7364 4724 7396
rect 4756 7364 4760 7396
rect 4720 7316 4760 7364
rect 4720 7284 4724 7316
rect 4756 7284 4760 7316
rect 4720 7236 4760 7284
rect 4720 7204 4724 7236
rect 4756 7204 4760 7236
rect 4720 7156 4760 7204
rect 4720 7124 4724 7156
rect 4756 7124 4760 7156
rect 4720 7076 4760 7124
rect 4720 7044 4724 7076
rect 4756 7044 4760 7076
rect 4720 6756 4760 7044
rect 4720 6724 4724 6756
rect 4756 6724 4760 6756
rect 4720 6676 4760 6724
rect 4720 6644 4724 6676
rect 4756 6644 4760 6676
rect 4720 6596 4760 6644
rect 4720 6564 4724 6596
rect 4756 6564 4760 6596
rect 4720 6516 4760 6564
rect 4720 6484 4724 6516
rect 4756 6484 4760 6516
rect 4720 6436 4760 6484
rect 4720 6404 4724 6436
rect 4756 6404 4760 6436
rect 4720 6356 4760 6404
rect 4720 6324 4724 6356
rect 4756 6324 4760 6356
rect 4720 6234 4760 6324
rect 4720 6206 4726 6234
rect 4754 6206 4760 6234
rect 4720 6074 4760 6206
rect 4720 6046 4726 6074
rect 4754 6046 4760 6074
rect 4720 5914 4760 6046
rect 4720 5886 4726 5914
rect 4754 5886 4760 5914
rect 4720 5796 4760 5886
rect 4720 5764 4724 5796
rect 4756 5764 4760 5796
rect 4720 5716 4760 5764
rect 4720 5684 4724 5716
rect 4756 5684 4760 5716
rect 4720 5636 4760 5684
rect 4720 5604 4724 5636
rect 4756 5604 4760 5636
rect 4720 5556 4760 5604
rect 4720 5524 4724 5556
rect 4756 5524 4760 5556
rect 4720 5476 4760 5524
rect 4720 5444 4724 5476
rect 4756 5444 4760 5476
rect 4720 5396 4760 5444
rect 4720 5364 4724 5396
rect 4756 5364 4760 5396
rect 4720 5316 4760 5364
rect 4720 5284 4724 5316
rect 4756 5284 4760 5316
rect 4720 5236 4760 5284
rect 4720 5204 4724 5236
rect 4756 5204 4760 5236
rect 4720 5156 4760 5204
rect 4720 5124 4724 5156
rect 4756 5124 4760 5156
rect 4720 5076 4760 5124
rect 4720 5044 4724 5076
rect 4756 5044 4760 5076
rect 4720 4996 4760 5044
rect 4720 4964 4724 4996
rect 4756 4964 4760 4996
rect 4720 4436 4760 4964
rect 4720 4404 4724 4436
rect 4756 4404 4760 4436
rect 4720 4356 4760 4404
rect 4720 4324 4724 4356
rect 4756 4324 4760 4356
rect 4720 4276 4760 4324
rect 4720 4244 4724 4276
rect 4756 4244 4760 4276
rect 4720 4196 4760 4244
rect 4720 4164 4724 4196
rect 4756 4164 4760 4196
rect 4720 4116 4760 4164
rect 4720 4084 4724 4116
rect 4756 4084 4760 4116
rect 4720 4036 4760 4084
rect 4720 4004 4724 4036
rect 4756 4004 4760 4036
rect 4720 3956 4760 4004
rect 4720 3924 4724 3956
rect 4756 3924 4760 3956
rect 4720 3156 4760 3924
rect 4720 3124 4724 3156
rect 4756 3124 4760 3156
rect 4720 3076 4760 3124
rect 4720 3044 4724 3076
rect 4756 3044 4760 3076
rect 4720 2996 4760 3044
rect 4720 2964 4724 2996
rect 4756 2964 4760 2996
rect 4720 2916 4760 2964
rect 4720 2884 4724 2916
rect 4756 2884 4760 2916
rect 4720 2836 4760 2884
rect 4720 2804 4724 2836
rect 4756 2804 4760 2836
rect 4720 2756 4760 2804
rect 4720 2724 4724 2756
rect 4756 2724 4760 2756
rect 4720 2676 4760 2724
rect 4720 2644 4724 2676
rect 4756 2644 4760 2676
rect 4720 2596 4760 2644
rect 4720 2564 4724 2596
rect 4756 2564 4760 2596
rect 4720 2516 4760 2564
rect 4720 2484 4724 2516
rect 4756 2484 4760 2516
rect 4720 2436 4760 2484
rect 4720 2404 4724 2436
rect 4756 2404 4760 2436
rect 4720 2356 4760 2404
rect 4720 2324 4724 2356
rect 4756 2324 4760 2356
rect 4720 2276 4760 2324
rect 4720 2244 4724 2276
rect 4756 2244 4760 2276
rect 4720 2196 4760 2244
rect 4720 2164 4724 2196
rect 4756 2164 4760 2196
rect 4720 2116 4760 2164
rect 4720 2084 4724 2116
rect 4756 2084 4760 2116
rect 4720 2036 4760 2084
rect 4720 2004 4724 2036
rect 4756 2004 4760 2036
rect 4720 1636 4760 2004
rect 4720 1604 4724 1636
rect 4756 1604 4760 1636
rect 4720 1556 4760 1604
rect 4720 1524 4724 1556
rect 4756 1524 4760 1556
rect 4720 1476 4760 1524
rect 4720 1444 4724 1476
rect 4756 1444 4760 1476
rect 4720 1396 4760 1444
rect 4720 1364 4724 1396
rect 4756 1364 4760 1396
rect 4720 1316 4760 1364
rect 4720 1284 4724 1316
rect 4756 1284 4760 1316
rect 4720 1236 4760 1284
rect 4720 1204 4724 1236
rect 4756 1204 4760 1236
rect 4720 1156 4760 1204
rect 4720 1124 4724 1156
rect 4756 1124 4760 1156
rect 4720 1076 4760 1124
rect 4720 1044 4724 1076
rect 4756 1044 4760 1076
rect 4720 756 4760 1044
rect 4720 724 4724 756
rect 4756 724 4760 756
rect 4720 676 4760 724
rect 4720 644 4724 676
rect 4756 644 4760 676
rect 4720 596 4760 644
rect 4720 564 4724 596
rect 4756 564 4760 596
rect 4720 196 4760 564
rect 4720 164 4724 196
rect 4756 164 4760 196
rect 4720 116 4760 164
rect 4720 84 4724 116
rect 4756 84 4760 116
rect 4720 36 4760 84
rect 4720 4 4724 36
rect 4756 4 4760 36
rect 4720 -40 4760 4
rect 4800 6154 4840 12680
rect 4800 6126 4806 6154
rect 4834 6126 4840 6154
rect 4800 -40 4840 6126
rect 4880 12636 4920 13204
rect 5040 13396 5080 13684
rect 5040 13364 5044 13396
rect 5076 13364 5080 13396
rect 5040 13356 5080 13364
rect 5040 13324 5044 13356
rect 5076 13324 5080 13356
rect 5040 13316 5080 13324
rect 5040 13284 5044 13316
rect 5076 13284 5080 13316
rect 5040 13276 5080 13284
rect 5040 13244 5044 13276
rect 5076 13244 5080 13276
rect 5040 13236 5080 13244
rect 5040 13204 5044 13236
rect 5076 13204 5080 13236
rect 4880 12604 4884 12636
rect 4916 12604 4920 12636
rect 4880 12556 4920 12604
rect 4880 12524 4884 12556
rect 4916 12524 4920 12556
rect 4880 12476 4920 12524
rect 4880 12444 4884 12476
rect 4916 12444 4920 12476
rect 4880 12396 4920 12444
rect 4880 12364 4884 12396
rect 4916 12364 4920 12396
rect 4880 12316 4920 12364
rect 4880 12284 4884 12316
rect 4916 12284 4920 12316
rect 4880 12236 4920 12284
rect 4880 12204 4884 12236
rect 4916 12204 4920 12236
rect 4880 12156 4920 12204
rect 4880 12124 4884 12156
rect 4916 12124 4920 12156
rect 4880 11836 4920 12124
rect 4880 11804 4884 11836
rect 4916 11804 4920 11836
rect 4880 11756 4920 11804
rect 4880 11724 4884 11756
rect 4916 11724 4920 11756
rect 4880 11676 4920 11724
rect 4880 11644 4884 11676
rect 4916 11644 4920 11676
rect 4880 11596 4920 11644
rect 4880 11564 4884 11596
rect 4916 11564 4920 11596
rect 4880 11516 4920 11564
rect 4880 11484 4884 11516
rect 4916 11484 4920 11516
rect 4880 11436 4920 11484
rect 4880 11404 4884 11436
rect 4916 11404 4920 11436
rect 4880 10876 4920 11404
rect 4880 10844 4884 10876
rect 4916 10844 4920 10876
rect 4880 10796 4920 10844
rect 4880 10764 4884 10796
rect 4916 10764 4920 10796
rect 4880 10716 4920 10764
rect 4880 10684 4884 10716
rect 4916 10684 4920 10716
rect 4880 10636 4920 10684
rect 4880 10604 4884 10636
rect 4916 10604 4920 10636
rect 4880 10556 4920 10604
rect 4880 10524 4884 10556
rect 4916 10524 4920 10556
rect 4880 10476 4920 10524
rect 4880 10444 4884 10476
rect 4916 10444 4920 10476
rect 4880 10396 4920 10444
rect 4880 10364 4884 10396
rect 4916 10364 4920 10396
rect 4880 10316 4920 10364
rect 4880 10284 4884 10316
rect 4916 10284 4920 10316
rect 4880 10236 4920 10284
rect 4880 10204 4884 10236
rect 4916 10204 4920 10236
rect 4880 10156 4920 10204
rect 4880 10124 4884 10156
rect 4916 10124 4920 10156
rect 4880 10076 4920 10124
rect 4880 10044 4884 10076
rect 4916 10044 4920 10076
rect 4880 9996 4920 10044
rect 4880 9964 4884 9996
rect 4916 9964 4920 9996
rect 4880 9916 4920 9964
rect 4880 9884 4884 9916
rect 4916 9884 4920 9916
rect 4880 9836 4920 9884
rect 4880 9804 4884 9836
rect 4916 9804 4920 9836
rect 4880 9756 4920 9804
rect 4880 9724 4884 9756
rect 4916 9724 4920 9756
rect 4880 9356 4920 9724
rect 4880 9324 4884 9356
rect 4916 9324 4920 9356
rect 4880 9276 4920 9324
rect 4880 9244 4884 9276
rect 4916 9244 4920 9276
rect 4880 9196 4920 9244
rect 4880 9164 4884 9196
rect 4916 9164 4920 9196
rect 4880 8876 4920 9164
rect 4880 8844 4884 8876
rect 4916 8844 4920 8876
rect 4880 8796 4920 8844
rect 4880 8764 4884 8796
rect 4916 8764 4920 8796
rect 4880 8716 4920 8764
rect 4880 8684 4884 8716
rect 4916 8684 4920 8716
rect 4880 8636 4920 8684
rect 4880 8604 4884 8636
rect 4916 8604 4920 8636
rect 4880 8556 4920 8604
rect 4880 8524 4884 8556
rect 4916 8524 4920 8556
rect 4880 8474 4920 8524
rect 4880 8446 4886 8474
rect 4914 8446 4920 8474
rect 4880 8314 4920 8446
rect 4880 8286 4886 8314
rect 4914 8286 4920 8314
rect 4880 7636 4920 8286
rect 4880 7604 4884 7636
rect 4916 7604 4920 7636
rect 4880 7556 4920 7604
rect 4880 7524 4884 7556
rect 4916 7524 4920 7556
rect 4880 7476 4920 7524
rect 4880 7444 4884 7476
rect 4916 7444 4920 7476
rect 4880 7396 4920 7444
rect 4880 7364 4884 7396
rect 4916 7364 4920 7396
rect 4880 7316 4920 7364
rect 4880 7284 4884 7316
rect 4916 7284 4920 7316
rect 4880 7236 4920 7284
rect 4880 7204 4884 7236
rect 4916 7204 4920 7236
rect 4880 7156 4920 7204
rect 4880 7124 4884 7156
rect 4916 7124 4920 7156
rect 4880 7076 4920 7124
rect 4880 7044 4884 7076
rect 4916 7044 4920 7076
rect 4880 6756 4920 7044
rect 4880 6724 4884 6756
rect 4916 6724 4920 6756
rect 4880 6676 4920 6724
rect 4880 6644 4884 6676
rect 4916 6644 4920 6676
rect 4880 6596 4920 6644
rect 4880 6564 4884 6596
rect 4916 6564 4920 6596
rect 4880 6516 4920 6564
rect 4880 6484 4884 6516
rect 4916 6484 4920 6516
rect 4880 6436 4920 6484
rect 4880 6404 4884 6436
rect 4916 6404 4920 6436
rect 4880 6356 4920 6404
rect 4880 6324 4884 6356
rect 4916 6324 4920 6356
rect 4880 6234 4920 6324
rect 4880 6206 4886 6234
rect 4914 6206 4920 6234
rect 4880 6074 4920 6206
rect 4880 6046 4886 6074
rect 4914 6046 4920 6074
rect 4880 5914 4920 6046
rect 4880 5886 4886 5914
rect 4914 5886 4920 5914
rect 4880 5796 4920 5886
rect 4880 5764 4884 5796
rect 4916 5764 4920 5796
rect 4880 5716 4920 5764
rect 4880 5684 4884 5716
rect 4916 5684 4920 5716
rect 4880 5636 4920 5684
rect 4880 5604 4884 5636
rect 4916 5604 4920 5636
rect 4880 5556 4920 5604
rect 4880 5524 4884 5556
rect 4916 5524 4920 5556
rect 4880 5476 4920 5524
rect 4880 5444 4884 5476
rect 4916 5444 4920 5476
rect 4880 5396 4920 5444
rect 4880 5364 4884 5396
rect 4916 5364 4920 5396
rect 4880 5316 4920 5364
rect 4880 5284 4884 5316
rect 4916 5284 4920 5316
rect 4880 5236 4920 5284
rect 4880 5204 4884 5236
rect 4916 5204 4920 5236
rect 4880 5156 4920 5204
rect 4880 5124 4884 5156
rect 4916 5124 4920 5156
rect 4880 5076 4920 5124
rect 4880 5044 4884 5076
rect 4916 5044 4920 5076
rect 4880 4996 4920 5044
rect 4880 4964 4884 4996
rect 4916 4964 4920 4996
rect 4880 4436 4920 4964
rect 4880 4404 4884 4436
rect 4916 4404 4920 4436
rect 4880 4356 4920 4404
rect 4880 4324 4884 4356
rect 4916 4324 4920 4356
rect 4880 4276 4920 4324
rect 4880 4244 4884 4276
rect 4916 4244 4920 4276
rect 4880 4196 4920 4244
rect 4880 4164 4884 4196
rect 4916 4164 4920 4196
rect 4880 4116 4920 4164
rect 4880 4084 4884 4116
rect 4916 4084 4920 4116
rect 4880 4036 4920 4084
rect 4880 4004 4884 4036
rect 4916 4004 4920 4036
rect 4880 3956 4920 4004
rect 4880 3924 4884 3956
rect 4916 3924 4920 3956
rect 4880 3156 4920 3924
rect 4880 3124 4884 3156
rect 4916 3124 4920 3156
rect 4880 3076 4920 3124
rect 4880 3044 4884 3076
rect 4916 3044 4920 3076
rect 4880 2996 4920 3044
rect 4880 2964 4884 2996
rect 4916 2964 4920 2996
rect 4880 2916 4920 2964
rect 4880 2884 4884 2916
rect 4916 2884 4920 2916
rect 4880 2836 4920 2884
rect 4880 2804 4884 2836
rect 4916 2804 4920 2836
rect 4880 2756 4920 2804
rect 4880 2724 4884 2756
rect 4916 2724 4920 2756
rect 4880 2676 4920 2724
rect 4880 2644 4884 2676
rect 4916 2644 4920 2676
rect 4880 2596 4920 2644
rect 4880 2564 4884 2596
rect 4916 2564 4920 2596
rect 4880 2516 4920 2564
rect 4880 2484 4884 2516
rect 4916 2484 4920 2516
rect 4880 2436 4920 2484
rect 4880 2404 4884 2436
rect 4916 2404 4920 2436
rect 4880 2356 4920 2404
rect 4880 2324 4884 2356
rect 4916 2324 4920 2356
rect 4880 2276 4920 2324
rect 4880 2244 4884 2276
rect 4916 2244 4920 2276
rect 4880 2196 4920 2244
rect 4880 2164 4884 2196
rect 4916 2164 4920 2196
rect 4880 2116 4920 2164
rect 4880 2084 4884 2116
rect 4916 2084 4920 2116
rect 4880 2036 4920 2084
rect 4880 2004 4884 2036
rect 4916 2004 4920 2036
rect 4880 1636 4920 2004
rect 4880 1604 4884 1636
rect 4916 1604 4920 1636
rect 4880 1556 4920 1604
rect 4880 1524 4884 1556
rect 4916 1524 4920 1556
rect 4880 1476 4920 1524
rect 4880 1444 4884 1476
rect 4916 1444 4920 1476
rect 4880 1396 4920 1444
rect 4880 1364 4884 1396
rect 4916 1364 4920 1396
rect 4880 1316 4920 1364
rect 4880 1284 4884 1316
rect 4916 1284 4920 1316
rect 4880 1236 4920 1284
rect 4880 1204 4884 1236
rect 4916 1204 4920 1236
rect 4880 1156 4920 1204
rect 4880 1124 4884 1156
rect 4916 1124 4920 1156
rect 4880 1076 4920 1124
rect 4880 1044 4884 1076
rect 4916 1044 4920 1076
rect 4880 756 4920 1044
rect 4880 724 4884 756
rect 4916 724 4920 756
rect 4880 676 4920 724
rect 4880 644 4884 676
rect 4916 644 4920 676
rect 4880 596 4920 644
rect 4880 564 4884 596
rect 4916 564 4920 596
rect 4880 196 4920 564
rect 4880 164 4884 196
rect 4916 164 4920 196
rect 4880 116 4920 164
rect 4880 84 4884 116
rect 4916 84 4920 116
rect 4880 36 4920 84
rect 4880 4 4884 36
rect 4916 4 4920 36
rect 4880 -40 4920 4
rect 4960 8394 5000 12680
rect 4960 8366 4966 8394
rect 4994 8366 5000 8394
rect 4960 6154 5000 8366
rect 4960 6126 4966 6154
rect 4994 6126 5000 6154
rect 4960 5994 5000 6126
rect 4960 5966 4966 5994
rect 4994 5966 5000 5994
rect 4960 -40 5000 5966
rect 5040 12636 5080 13204
rect 5040 12604 5044 12636
rect 5076 12604 5080 12636
rect 5040 12556 5080 12604
rect 5040 12524 5044 12556
rect 5076 12524 5080 12556
rect 5040 12476 5080 12524
rect 5040 12444 5044 12476
rect 5076 12444 5080 12476
rect 5040 12396 5080 12444
rect 5040 12364 5044 12396
rect 5076 12364 5080 12396
rect 5040 12316 5080 12364
rect 5040 12284 5044 12316
rect 5076 12284 5080 12316
rect 5040 12236 5080 12284
rect 5040 12204 5044 12236
rect 5076 12204 5080 12236
rect 5040 12156 5080 12204
rect 5040 12124 5044 12156
rect 5076 12124 5080 12156
rect 5040 11836 5080 12124
rect 5040 11804 5044 11836
rect 5076 11804 5080 11836
rect 5040 11756 5080 11804
rect 5040 11724 5044 11756
rect 5076 11724 5080 11756
rect 5040 11676 5080 11724
rect 5040 11644 5044 11676
rect 5076 11644 5080 11676
rect 5040 11596 5080 11644
rect 5040 11564 5044 11596
rect 5076 11564 5080 11596
rect 5040 11516 5080 11564
rect 5040 11484 5044 11516
rect 5076 11484 5080 11516
rect 5040 11436 5080 11484
rect 5040 11404 5044 11436
rect 5076 11404 5080 11436
rect 5040 11154 5080 11404
rect 5040 11126 5046 11154
rect 5074 11126 5080 11154
rect 5040 10994 5080 11126
rect 5040 10966 5046 10994
rect 5074 10966 5080 10994
rect 5040 10876 5080 10966
rect 5040 10844 5044 10876
rect 5076 10844 5080 10876
rect 5040 10796 5080 10844
rect 5040 10764 5044 10796
rect 5076 10764 5080 10796
rect 5040 10716 5080 10764
rect 5040 10684 5044 10716
rect 5076 10684 5080 10716
rect 5040 10636 5080 10684
rect 5040 10604 5044 10636
rect 5076 10604 5080 10636
rect 5040 10556 5080 10604
rect 5040 10524 5044 10556
rect 5076 10524 5080 10556
rect 5040 10476 5080 10524
rect 5040 10444 5044 10476
rect 5076 10444 5080 10476
rect 5040 10396 5080 10444
rect 5040 10364 5044 10396
rect 5076 10364 5080 10396
rect 5040 10316 5080 10364
rect 5040 10284 5044 10316
rect 5076 10284 5080 10316
rect 5040 10236 5080 10284
rect 5040 10204 5044 10236
rect 5076 10204 5080 10236
rect 5040 10156 5080 10204
rect 5040 10124 5044 10156
rect 5076 10124 5080 10156
rect 5040 10076 5080 10124
rect 5040 10044 5044 10076
rect 5076 10044 5080 10076
rect 5040 9996 5080 10044
rect 5040 9964 5044 9996
rect 5076 9964 5080 9996
rect 5040 9916 5080 9964
rect 5040 9884 5044 9916
rect 5076 9884 5080 9916
rect 5040 9836 5080 9884
rect 5040 9804 5044 9836
rect 5076 9804 5080 9836
rect 5040 9756 5080 9804
rect 5040 9724 5044 9756
rect 5076 9724 5080 9756
rect 5040 9356 5080 9724
rect 5040 9324 5044 9356
rect 5076 9324 5080 9356
rect 5040 9276 5080 9324
rect 5040 9244 5044 9276
rect 5076 9244 5080 9276
rect 5040 9196 5080 9244
rect 5040 9164 5044 9196
rect 5076 9164 5080 9196
rect 5040 8876 5080 9164
rect 5040 8844 5044 8876
rect 5076 8844 5080 8876
rect 5040 8796 5080 8844
rect 5040 8764 5044 8796
rect 5076 8764 5080 8796
rect 5040 8716 5080 8764
rect 5040 8684 5044 8716
rect 5076 8684 5080 8716
rect 5040 8636 5080 8684
rect 5040 8604 5044 8636
rect 5076 8604 5080 8636
rect 5040 8556 5080 8604
rect 5040 8524 5044 8556
rect 5076 8524 5080 8556
rect 5040 8474 5080 8524
rect 5040 8446 5046 8474
rect 5074 8446 5080 8474
rect 5040 8314 5080 8446
rect 5040 8286 5046 8314
rect 5074 8286 5080 8314
rect 5040 8074 5080 8286
rect 5040 8046 5046 8074
rect 5074 8046 5080 8074
rect 5040 7754 5080 8046
rect 5040 7726 5046 7754
rect 5074 7726 5080 7754
rect 5040 7636 5080 7726
rect 5040 7604 5044 7636
rect 5076 7604 5080 7636
rect 5040 7556 5080 7604
rect 5040 7524 5044 7556
rect 5076 7524 5080 7556
rect 5040 7476 5080 7524
rect 5040 7444 5044 7476
rect 5076 7444 5080 7476
rect 5040 7396 5080 7444
rect 5040 7364 5044 7396
rect 5076 7364 5080 7396
rect 5040 7316 5080 7364
rect 5040 7284 5044 7316
rect 5076 7284 5080 7316
rect 5040 7236 5080 7284
rect 5040 7204 5044 7236
rect 5076 7204 5080 7236
rect 5040 7156 5080 7204
rect 5040 7124 5044 7156
rect 5076 7124 5080 7156
rect 5040 7076 5080 7124
rect 5040 7044 5044 7076
rect 5076 7044 5080 7076
rect 5040 6756 5080 7044
rect 5040 6724 5044 6756
rect 5076 6724 5080 6756
rect 5040 6676 5080 6724
rect 5040 6644 5044 6676
rect 5076 6644 5080 6676
rect 5040 6596 5080 6644
rect 5040 6564 5044 6596
rect 5076 6564 5080 6596
rect 5040 6516 5080 6564
rect 5040 6484 5044 6516
rect 5076 6484 5080 6516
rect 5040 6436 5080 6484
rect 5040 6404 5044 6436
rect 5076 6404 5080 6436
rect 5040 6356 5080 6404
rect 5040 6324 5044 6356
rect 5076 6324 5080 6356
rect 5040 6234 5080 6324
rect 5040 6206 5046 6234
rect 5074 6206 5080 6234
rect 5040 6074 5080 6206
rect 5040 6046 5046 6074
rect 5074 6046 5080 6074
rect 5040 5914 5080 6046
rect 5040 5886 5046 5914
rect 5074 5886 5080 5914
rect 5040 5796 5080 5886
rect 5040 5764 5044 5796
rect 5076 5764 5080 5796
rect 5040 5716 5080 5764
rect 5040 5684 5044 5716
rect 5076 5684 5080 5716
rect 5040 5636 5080 5684
rect 5040 5604 5044 5636
rect 5076 5604 5080 5636
rect 5040 5556 5080 5604
rect 5040 5524 5044 5556
rect 5076 5524 5080 5556
rect 5040 5476 5080 5524
rect 5040 5444 5044 5476
rect 5076 5444 5080 5476
rect 5040 5396 5080 5444
rect 5040 5364 5044 5396
rect 5076 5364 5080 5396
rect 5040 5316 5080 5364
rect 5040 5284 5044 5316
rect 5076 5284 5080 5316
rect 5040 5236 5080 5284
rect 5040 5204 5044 5236
rect 5076 5204 5080 5236
rect 5040 5156 5080 5204
rect 5040 5124 5044 5156
rect 5076 5124 5080 5156
rect 5040 5076 5080 5124
rect 5040 5044 5044 5076
rect 5076 5044 5080 5076
rect 5040 4996 5080 5044
rect 5040 4964 5044 4996
rect 5076 4964 5080 4996
rect 5040 4436 5080 4964
rect 5040 4404 5044 4436
rect 5076 4404 5080 4436
rect 5040 4356 5080 4404
rect 5040 4324 5044 4356
rect 5076 4324 5080 4356
rect 5040 4276 5080 4324
rect 5040 4244 5044 4276
rect 5076 4244 5080 4276
rect 5040 4196 5080 4244
rect 5040 4164 5044 4196
rect 5076 4164 5080 4196
rect 5040 4116 5080 4164
rect 5040 4084 5044 4116
rect 5076 4084 5080 4116
rect 5040 4036 5080 4084
rect 5040 4004 5044 4036
rect 5076 4004 5080 4036
rect 5040 3956 5080 4004
rect 5040 3924 5044 3956
rect 5076 3924 5080 3956
rect 5040 3156 5080 3924
rect 5040 3124 5044 3156
rect 5076 3124 5080 3156
rect 5040 3076 5080 3124
rect 5040 3044 5044 3076
rect 5076 3044 5080 3076
rect 5040 2996 5080 3044
rect 5040 2964 5044 2996
rect 5076 2964 5080 2996
rect 5040 2916 5080 2964
rect 5040 2884 5044 2916
rect 5076 2884 5080 2916
rect 5040 2836 5080 2884
rect 5040 2804 5044 2836
rect 5076 2804 5080 2836
rect 5040 2756 5080 2804
rect 5040 2724 5044 2756
rect 5076 2724 5080 2756
rect 5040 2676 5080 2724
rect 5040 2644 5044 2676
rect 5076 2644 5080 2676
rect 5040 2596 5080 2644
rect 5040 2564 5044 2596
rect 5076 2564 5080 2596
rect 5040 2516 5080 2564
rect 5040 2484 5044 2516
rect 5076 2484 5080 2516
rect 5040 2436 5080 2484
rect 5040 2404 5044 2436
rect 5076 2404 5080 2436
rect 5040 2356 5080 2404
rect 5040 2324 5044 2356
rect 5076 2324 5080 2356
rect 5040 2276 5080 2324
rect 5040 2244 5044 2276
rect 5076 2244 5080 2276
rect 5040 2196 5080 2244
rect 5040 2164 5044 2196
rect 5076 2164 5080 2196
rect 5040 2116 5080 2164
rect 5040 2084 5044 2116
rect 5076 2084 5080 2116
rect 5040 2036 5080 2084
rect 5040 2004 5044 2036
rect 5076 2004 5080 2036
rect 5040 1636 5080 2004
rect 5040 1604 5044 1636
rect 5076 1604 5080 1636
rect 5040 1556 5080 1604
rect 5040 1524 5044 1556
rect 5076 1524 5080 1556
rect 5040 1476 5080 1524
rect 5040 1444 5044 1476
rect 5076 1444 5080 1476
rect 5040 1396 5080 1444
rect 5040 1364 5044 1396
rect 5076 1364 5080 1396
rect 5040 1316 5080 1364
rect 5040 1284 5044 1316
rect 5076 1284 5080 1316
rect 5040 1236 5080 1284
rect 5040 1204 5044 1236
rect 5076 1204 5080 1236
rect 5040 1156 5080 1204
rect 5040 1124 5044 1156
rect 5076 1124 5080 1156
rect 5040 1076 5080 1124
rect 5040 1044 5044 1076
rect 5076 1044 5080 1076
rect 5040 756 5080 1044
rect 5040 724 5044 756
rect 5076 724 5080 756
rect 5040 676 5080 724
rect 5040 644 5044 676
rect 5076 644 5080 676
rect 5040 596 5080 644
rect 5040 564 5044 596
rect 5076 564 5080 596
rect 5040 196 5080 564
rect 5040 164 5044 196
rect 5076 164 5080 196
rect 5040 116 5080 164
rect 5040 84 5044 116
rect 5076 84 5080 116
rect 5040 36 5080 84
rect 5040 4 5044 36
rect 5076 4 5080 36
rect 5040 -40 5080 4
rect 5120 15396 5160 15400
rect 5120 15364 5124 15396
rect 5156 15364 5160 15396
rect 5120 14116 5160 15364
rect 5120 14084 5124 14116
rect 5156 14084 5160 14116
rect 5120 12636 5160 14084
rect 5120 12604 5124 12636
rect 5156 12604 5160 12636
rect 5120 12556 5160 12604
rect 5120 12524 5124 12556
rect 5156 12524 5160 12556
rect 5120 12476 5160 12524
rect 5120 12444 5124 12476
rect 5156 12444 5160 12476
rect 5120 12396 5160 12444
rect 5120 12364 5124 12396
rect 5156 12364 5160 12396
rect 5120 12316 5160 12364
rect 5120 12284 5124 12316
rect 5156 12284 5160 12316
rect 5120 12236 5160 12284
rect 5120 12204 5124 12236
rect 5156 12204 5160 12236
rect 5120 12156 5160 12204
rect 5120 12124 5124 12156
rect 5156 12124 5160 12156
rect 5120 11836 5160 12124
rect 5120 11804 5124 11836
rect 5156 11804 5160 11836
rect 5120 11756 5160 11804
rect 5120 11724 5124 11756
rect 5156 11724 5160 11756
rect 5120 11676 5160 11724
rect 5120 11644 5124 11676
rect 5156 11644 5160 11676
rect 5120 11596 5160 11644
rect 5120 11564 5124 11596
rect 5156 11564 5160 11596
rect 5120 11516 5160 11564
rect 5120 11484 5124 11516
rect 5156 11484 5160 11516
rect 5120 11436 5160 11484
rect 5120 11404 5124 11436
rect 5156 11404 5160 11436
rect 5120 11074 5160 11404
rect 5120 11046 5126 11074
rect 5154 11046 5160 11074
rect 5120 10876 5160 11046
rect 5120 10844 5124 10876
rect 5156 10844 5160 10876
rect 5120 10796 5160 10844
rect 5120 10764 5124 10796
rect 5156 10764 5160 10796
rect 5120 10716 5160 10764
rect 5120 10684 5124 10716
rect 5156 10684 5160 10716
rect 5120 10636 5160 10684
rect 5120 10604 5124 10636
rect 5156 10604 5160 10636
rect 5120 10556 5160 10604
rect 5120 10524 5124 10556
rect 5156 10524 5160 10556
rect 5120 10476 5160 10524
rect 5120 10444 5124 10476
rect 5156 10444 5160 10476
rect 5120 10396 5160 10444
rect 5120 10364 5124 10396
rect 5156 10364 5160 10396
rect 5120 10316 5160 10364
rect 5120 10284 5124 10316
rect 5156 10284 5160 10316
rect 5120 10236 5160 10284
rect 5120 10204 5124 10236
rect 5156 10204 5160 10236
rect 5120 10156 5160 10204
rect 5120 10124 5124 10156
rect 5156 10124 5160 10156
rect 5120 10076 5160 10124
rect 5120 10044 5124 10076
rect 5156 10044 5160 10076
rect 5120 9996 5160 10044
rect 5120 9964 5124 9996
rect 5156 9964 5160 9996
rect 5120 9916 5160 9964
rect 5120 9884 5124 9916
rect 5156 9884 5160 9916
rect 5120 9836 5160 9884
rect 5120 9804 5124 9836
rect 5156 9804 5160 9836
rect 5120 9756 5160 9804
rect 5120 9724 5124 9756
rect 5156 9724 5160 9756
rect 5120 9356 5160 9724
rect 5120 9324 5124 9356
rect 5156 9324 5160 9356
rect 5120 9276 5160 9324
rect 5120 9244 5124 9276
rect 5156 9244 5160 9276
rect 5120 9196 5160 9244
rect 5120 9164 5124 9196
rect 5156 9164 5160 9196
rect 5120 9114 5160 9164
rect 5120 9086 5126 9114
rect 5154 9086 5160 9114
rect 5120 8954 5160 9086
rect 5120 8926 5126 8954
rect 5154 8926 5160 8954
rect 5120 8876 5160 8926
rect 5120 8844 5124 8876
rect 5156 8844 5160 8876
rect 5120 8796 5160 8844
rect 5120 8764 5124 8796
rect 5156 8764 5160 8796
rect 5120 8716 5160 8764
rect 5120 8684 5124 8716
rect 5156 8684 5160 8716
rect 5120 8636 5160 8684
rect 5120 8604 5124 8636
rect 5156 8604 5160 8636
rect 5120 8556 5160 8604
rect 5120 8524 5124 8556
rect 5156 8524 5160 8556
rect 5120 7994 5160 8524
rect 5120 7966 5126 7994
rect 5154 7966 5160 7994
rect 5120 7834 5160 7966
rect 5120 7806 5126 7834
rect 5154 7806 5160 7834
rect 5120 7636 5160 7806
rect 5120 7604 5124 7636
rect 5156 7604 5160 7636
rect 5120 7556 5160 7604
rect 5120 7524 5124 7556
rect 5156 7524 5160 7556
rect 5120 7476 5160 7524
rect 5120 7444 5124 7476
rect 5156 7444 5160 7476
rect 5120 7396 5160 7444
rect 5120 7364 5124 7396
rect 5156 7364 5160 7396
rect 5120 7316 5160 7364
rect 5120 7284 5124 7316
rect 5156 7284 5160 7316
rect 5120 7236 5160 7284
rect 5120 7204 5124 7236
rect 5156 7204 5160 7236
rect 5120 7156 5160 7204
rect 5120 7124 5124 7156
rect 5156 7124 5160 7156
rect 5120 7076 5160 7124
rect 5120 7044 5124 7076
rect 5156 7044 5160 7076
rect 5120 6756 5160 7044
rect 5120 6724 5124 6756
rect 5156 6724 5160 6756
rect 5120 6676 5160 6724
rect 5120 6644 5124 6676
rect 5156 6644 5160 6676
rect 5120 6596 5160 6644
rect 5120 6564 5124 6596
rect 5156 6564 5160 6596
rect 5120 6516 5160 6564
rect 5120 6484 5124 6516
rect 5156 6484 5160 6516
rect 5120 6436 5160 6484
rect 5120 6404 5124 6436
rect 5156 6404 5160 6436
rect 5120 6356 5160 6404
rect 5120 6324 5124 6356
rect 5156 6324 5160 6356
rect 5120 5796 5160 6324
rect 5120 5764 5124 5796
rect 5156 5764 5160 5796
rect 5120 5716 5160 5764
rect 5120 5684 5124 5716
rect 5156 5684 5160 5716
rect 5120 5636 5160 5684
rect 5120 5604 5124 5636
rect 5156 5604 5160 5636
rect 5120 5556 5160 5604
rect 5120 5524 5124 5556
rect 5156 5524 5160 5556
rect 5120 5476 5160 5524
rect 5120 5444 5124 5476
rect 5156 5444 5160 5476
rect 5120 5396 5160 5444
rect 5120 5364 5124 5396
rect 5156 5364 5160 5396
rect 5120 5316 5160 5364
rect 5120 5284 5124 5316
rect 5156 5284 5160 5316
rect 5120 5236 5160 5284
rect 5120 5204 5124 5236
rect 5156 5204 5160 5236
rect 5120 5156 5160 5204
rect 5120 5124 5124 5156
rect 5156 5124 5160 5156
rect 5120 5076 5160 5124
rect 5120 5044 5124 5076
rect 5156 5044 5160 5076
rect 5120 4996 5160 5044
rect 5120 4964 5124 4996
rect 5156 4964 5160 4996
rect 5120 4436 5160 4964
rect 5120 4404 5124 4436
rect 5156 4404 5160 4436
rect 5120 4356 5160 4404
rect 5120 4324 5124 4356
rect 5156 4324 5160 4356
rect 5120 4276 5160 4324
rect 5120 4244 5124 4276
rect 5156 4244 5160 4276
rect 5120 4196 5160 4244
rect 5120 4164 5124 4196
rect 5156 4164 5160 4196
rect 5120 4116 5160 4164
rect 5120 4084 5124 4116
rect 5156 4084 5160 4116
rect 5120 4036 5160 4084
rect 5120 4004 5124 4036
rect 5156 4004 5160 4036
rect 5120 3956 5160 4004
rect 5120 3924 5124 3956
rect 5156 3924 5160 3956
rect 5120 3156 5160 3924
rect 5120 3124 5124 3156
rect 5156 3124 5160 3156
rect 5120 3076 5160 3124
rect 5120 3044 5124 3076
rect 5156 3044 5160 3076
rect 5120 2996 5160 3044
rect 5120 2964 5124 2996
rect 5156 2964 5160 2996
rect 5120 2916 5160 2964
rect 5120 2884 5124 2916
rect 5156 2884 5160 2916
rect 5120 2836 5160 2884
rect 5120 2804 5124 2836
rect 5156 2804 5160 2836
rect 5120 2756 5160 2804
rect 5120 2724 5124 2756
rect 5156 2724 5160 2756
rect 5120 2676 5160 2724
rect 5120 2644 5124 2676
rect 5156 2644 5160 2676
rect 5120 2596 5160 2644
rect 5120 2564 5124 2596
rect 5156 2564 5160 2596
rect 5120 2516 5160 2564
rect 5120 2484 5124 2516
rect 5156 2484 5160 2516
rect 5120 2436 5160 2484
rect 5120 2404 5124 2436
rect 5156 2404 5160 2436
rect 5120 2356 5160 2404
rect 5120 2324 5124 2356
rect 5156 2324 5160 2356
rect 5120 2276 5160 2324
rect 5120 2244 5124 2276
rect 5156 2244 5160 2276
rect 5120 2196 5160 2244
rect 5120 2164 5124 2196
rect 5156 2164 5160 2196
rect 5120 2116 5160 2164
rect 5120 2084 5124 2116
rect 5156 2084 5160 2116
rect 5120 2036 5160 2084
rect 5120 2004 5124 2036
rect 5156 2004 5160 2036
rect 5120 1636 5160 2004
rect 5120 1604 5124 1636
rect 5156 1604 5160 1636
rect 5120 1556 5160 1604
rect 5120 1524 5124 1556
rect 5156 1524 5160 1556
rect 5120 1476 5160 1524
rect 5120 1444 5124 1476
rect 5156 1444 5160 1476
rect 5120 1396 5160 1444
rect 5120 1364 5124 1396
rect 5156 1364 5160 1396
rect 5120 1316 5160 1364
rect 5120 1284 5124 1316
rect 5156 1284 5160 1316
rect 5120 1236 5160 1284
rect 5120 1204 5124 1236
rect 5156 1204 5160 1236
rect 5120 1156 5160 1204
rect 5120 1124 5124 1156
rect 5156 1124 5160 1156
rect 5120 1076 5160 1124
rect 5120 1044 5124 1076
rect 5156 1044 5160 1076
rect 5120 756 5160 1044
rect 5120 724 5124 756
rect 5156 724 5160 756
rect 5120 676 5160 724
rect 5120 644 5124 676
rect 5156 644 5160 676
rect 5120 596 5160 644
rect 5120 564 5124 596
rect 5156 564 5160 596
rect 5120 196 5160 564
rect 5120 164 5124 196
rect 5156 164 5160 196
rect 5120 116 5160 164
rect 5120 84 5124 116
rect 5156 84 5160 116
rect 5120 36 5160 84
rect 5120 4 5124 36
rect 5156 4 5160 36
rect 5120 -40 5160 4
rect 5200 15316 5240 15400
rect 5200 15284 5204 15316
rect 5236 15284 5240 15316
rect 5200 7914 5240 15284
rect 5200 7886 5206 7914
rect 5234 7886 5240 7914
rect 5200 -40 5240 7886
rect 5280 15396 5320 15400
rect 5280 15364 5284 15396
rect 5316 15364 5320 15396
rect 5280 14116 5320 15364
rect 5280 14084 5284 14116
rect 5316 14084 5320 14116
rect 5280 12636 5320 14084
rect 5280 12604 5284 12636
rect 5316 12604 5320 12636
rect 5280 12556 5320 12604
rect 5280 12524 5284 12556
rect 5316 12524 5320 12556
rect 5280 12476 5320 12524
rect 5280 12444 5284 12476
rect 5316 12444 5320 12476
rect 5280 12396 5320 12444
rect 5280 12364 5284 12396
rect 5316 12364 5320 12396
rect 5280 12316 5320 12364
rect 5280 12284 5284 12316
rect 5316 12284 5320 12316
rect 5280 12236 5320 12284
rect 5280 12204 5284 12236
rect 5316 12204 5320 12236
rect 5280 12156 5320 12204
rect 5280 12124 5284 12156
rect 5316 12124 5320 12156
rect 5280 11836 5320 12124
rect 5280 11804 5284 11836
rect 5316 11804 5320 11836
rect 5280 11756 5320 11804
rect 5280 11724 5284 11756
rect 5316 11724 5320 11756
rect 5280 11676 5320 11724
rect 5280 11644 5284 11676
rect 5316 11644 5320 11676
rect 5280 11596 5320 11644
rect 5280 11564 5284 11596
rect 5316 11564 5320 11596
rect 5280 11516 5320 11564
rect 5280 11484 5284 11516
rect 5316 11484 5320 11516
rect 5280 11436 5320 11484
rect 5280 11404 5284 11436
rect 5316 11404 5320 11436
rect 5280 11074 5320 11404
rect 5280 11046 5286 11074
rect 5314 11046 5320 11074
rect 5280 10876 5320 11046
rect 5280 10844 5284 10876
rect 5316 10844 5320 10876
rect 5280 10796 5320 10844
rect 5280 10764 5284 10796
rect 5316 10764 5320 10796
rect 5280 10716 5320 10764
rect 5280 10684 5284 10716
rect 5316 10684 5320 10716
rect 5280 10636 5320 10684
rect 5280 10604 5284 10636
rect 5316 10604 5320 10636
rect 5280 10556 5320 10604
rect 5280 10524 5284 10556
rect 5316 10524 5320 10556
rect 5280 10476 5320 10524
rect 5280 10444 5284 10476
rect 5316 10444 5320 10476
rect 5280 10396 5320 10444
rect 5280 10364 5284 10396
rect 5316 10364 5320 10396
rect 5280 10316 5320 10364
rect 5280 10284 5284 10316
rect 5316 10284 5320 10316
rect 5280 10236 5320 10284
rect 5280 10204 5284 10236
rect 5316 10204 5320 10236
rect 5280 10156 5320 10204
rect 5280 10124 5284 10156
rect 5316 10124 5320 10156
rect 5280 10076 5320 10124
rect 5280 10044 5284 10076
rect 5316 10044 5320 10076
rect 5280 9996 5320 10044
rect 5280 9964 5284 9996
rect 5316 9964 5320 9996
rect 5280 9916 5320 9964
rect 5280 9884 5284 9916
rect 5316 9884 5320 9916
rect 5280 9836 5320 9884
rect 5280 9804 5284 9836
rect 5316 9804 5320 9836
rect 5280 9756 5320 9804
rect 5280 9724 5284 9756
rect 5316 9724 5320 9756
rect 5280 9356 5320 9724
rect 5280 9324 5284 9356
rect 5316 9324 5320 9356
rect 5280 9276 5320 9324
rect 5280 9244 5284 9276
rect 5316 9244 5320 9276
rect 5280 9196 5320 9244
rect 5280 9164 5284 9196
rect 5316 9164 5320 9196
rect 5280 9114 5320 9164
rect 5280 9086 5286 9114
rect 5314 9086 5320 9114
rect 5280 8954 5320 9086
rect 5280 8926 5286 8954
rect 5314 8926 5320 8954
rect 5280 8876 5320 8926
rect 5280 8844 5284 8876
rect 5316 8844 5320 8876
rect 5280 8796 5320 8844
rect 5280 8764 5284 8796
rect 5316 8764 5320 8796
rect 5280 8716 5320 8764
rect 5280 8684 5284 8716
rect 5316 8684 5320 8716
rect 5280 8636 5320 8684
rect 5280 8604 5284 8636
rect 5316 8604 5320 8636
rect 5280 8556 5320 8604
rect 5280 8524 5284 8556
rect 5316 8524 5320 8556
rect 5280 7994 5320 8524
rect 5280 7966 5286 7994
rect 5314 7966 5320 7994
rect 5280 7834 5320 7966
rect 5280 7806 5286 7834
rect 5314 7806 5320 7834
rect 5280 7636 5320 7806
rect 5280 7604 5284 7636
rect 5316 7604 5320 7636
rect 5280 7556 5320 7604
rect 5280 7524 5284 7556
rect 5316 7524 5320 7556
rect 5280 7476 5320 7524
rect 5280 7444 5284 7476
rect 5316 7444 5320 7476
rect 5280 7396 5320 7444
rect 5280 7364 5284 7396
rect 5316 7364 5320 7396
rect 5280 7316 5320 7364
rect 5280 7284 5284 7316
rect 5316 7284 5320 7316
rect 5280 7236 5320 7284
rect 5280 7204 5284 7236
rect 5316 7204 5320 7236
rect 5280 7156 5320 7204
rect 5280 7124 5284 7156
rect 5316 7124 5320 7156
rect 5280 7076 5320 7124
rect 5280 7044 5284 7076
rect 5316 7044 5320 7076
rect 5280 6756 5320 7044
rect 5280 6724 5284 6756
rect 5316 6724 5320 6756
rect 5280 6676 5320 6724
rect 5280 6644 5284 6676
rect 5316 6644 5320 6676
rect 5280 6596 5320 6644
rect 5280 6564 5284 6596
rect 5316 6564 5320 6596
rect 5280 6516 5320 6564
rect 5280 6484 5284 6516
rect 5316 6484 5320 6516
rect 5280 6436 5320 6484
rect 5280 6404 5284 6436
rect 5316 6404 5320 6436
rect 5280 6356 5320 6404
rect 5280 6324 5284 6356
rect 5316 6324 5320 6356
rect 5280 5796 5320 6324
rect 5280 5764 5284 5796
rect 5316 5764 5320 5796
rect 5280 5716 5320 5764
rect 5280 5684 5284 5716
rect 5316 5684 5320 5716
rect 5280 5636 5320 5684
rect 5280 5604 5284 5636
rect 5316 5604 5320 5636
rect 5280 5556 5320 5604
rect 5280 5524 5284 5556
rect 5316 5524 5320 5556
rect 5280 5476 5320 5524
rect 5280 5444 5284 5476
rect 5316 5444 5320 5476
rect 5280 5396 5320 5444
rect 5280 5364 5284 5396
rect 5316 5364 5320 5396
rect 5280 5316 5320 5364
rect 5280 5284 5284 5316
rect 5316 5284 5320 5316
rect 5280 5236 5320 5284
rect 5280 5204 5284 5236
rect 5316 5204 5320 5236
rect 5280 5156 5320 5204
rect 5280 5124 5284 5156
rect 5316 5124 5320 5156
rect 5280 5076 5320 5124
rect 5280 5044 5284 5076
rect 5316 5044 5320 5076
rect 5280 4996 5320 5044
rect 5280 4964 5284 4996
rect 5316 4964 5320 4996
rect 5280 4436 5320 4964
rect 5280 4404 5284 4436
rect 5316 4404 5320 4436
rect 5280 4356 5320 4404
rect 5280 4324 5284 4356
rect 5316 4324 5320 4356
rect 5280 4276 5320 4324
rect 5280 4244 5284 4276
rect 5316 4244 5320 4276
rect 5280 4196 5320 4244
rect 5280 4164 5284 4196
rect 5316 4164 5320 4196
rect 5280 4116 5320 4164
rect 5280 4084 5284 4116
rect 5316 4084 5320 4116
rect 5280 4036 5320 4084
rect 5280 4004 5284 4036
rect 5316 4004 5320 4036
rect 5280 3956 5320 4004
rect 5280 3924 5284 3956
rect 5316 3924 5320 3956
rect 5280 3156 5320 3924
rect 5280 3124 5284 3156
rect 5316 3124 5320 3156
rect 5280 3076 5320 3124
rect 5280 3044 5284 3076
rect 5316 3044 5320 3076
rect 5280 2996 5320 3044
rect 5280 2964 5284 2996
rect 5316 2964 5320 2996
rect 5280 2916 5320 2964
rect 5280 2884 5284 2916
rect 5316 2884 5320 2916
rect 5280 2836 5320 2884
rect 5280 2804 5284 2836
rect 5316 2804 5320 2836
rect 5280 2756 5320 2804
rect 5280 2724 5284 2756
rect 5316 2724 5320 2756
rect 5280 2676 5320 2724
rect 5280 2644 5284 2676
rect 5316 2644 5320 2676
rect 5280 2596 5320 2644
rect 5280 2564 5284 2596
rect 5316 2564 5320 2596
rect 5280 2516 5320 2564
rect 5280 2484 5284 2516
rect 5316 2484 5320 2516
rect 5280 2436 5320 2484
rect 5280 2404 5284 2436
rect 5316 2404 5320 2436
rect 5280 2356 5320 2404
rect 5280 2324 5284 2356
rect 5316 2324 5320 2356
rect 5280 2276 5320 2324
rect 5280 2244 5284 2276
rect 5316 2244 5320 2276
rect 5280 2196 5320 2244
rect 5280 2164 5284 2196
rect 5316 2164 5320 2196
rect 5280 2116 5320 2164
rect 5280 2084 5284 2116
rect 5316 2084 5320 2116
rect 5280 2036 5320 2084
rect 5280 2004 5284 2036
rect 5316 2004 5320 2036
rect 5280 1636 5320 2004
rect 5280 1604 5284 1636
rect 5316 1604 5320 1636
rect 5280 1556 5320 1604
rect 5280 1524 5284 1556
rect 5316 1524 5320 1556
rect 5280 1476 5320 1524
rect 5280 1444 5284 1476
rect 5316 1444 5320 1476
rect 5280 1396 5320 1444
rect 5280 1364 5284 1396
rect 5316 1364 5320 1396
rect 5280 1316 5320 1364
rect 5280 1284 5284 1316
rect 5316 1284 5320 1316
rect 5280 1236 5320 1284
rect 5280 1204 5284 1236
rect 5316 1204 5320 1236
rect 5280 1156 5320 1204
rect 5280 1124 5284 1156
rect 5316 1124 5320 1156
rect 5280 1076 5320 1124
rect 5280 1044 5284 1076
rect 5316 1044 5320 1076
rect 5280 756 5320 1044
rect 5280 724 5284 756
rect 5316 724 5320 756
rect 5280 676 5320 724
rect 5280 644 5284 676
rect 5316 644 5320 676
rect 5280 596 5320 644
rect 5280 564 5284 596
rect 5316 564 5320 596
rect 5280 196 5320 564
rect 5280 164 5284 196
rect 5316 164 5320 196
rect 5280 116 5320 164
rect 5280 84 5284 116
rect 5316 84 5320 116
rect 5280 36 5320 84
rect 5280 4 5284 36
rect 5316 4 5320 36
rect 5280 -40 5320 4
rect 5360 15316 5400 15400
rect 5360 15284 5364 15316
rect 5396 15284 5400 15316
rect 5360 9034 5400 15284
rect 5360 9006 5366 9034
rect 5394 9006 5400 9034
rect 5360 -40 5400 9006
rect 5440 15396 5480 15400
rect 5440 15364 5444 15396
rect 5476 15364 5480 15396
rect 5440 14116 5480 15364
rect 5440 14084 5444 14116
rect 5476 14084 5480 14116
rect 5440 12636 5480 14084
rect 5440 12604 5444 12636
rect 5476 12604 5480 12636
rect 5440 12556 5480 12604
rect 5440 12524 5444 12556
rect 5476 12524 5480 12556
rect 5440 12476 5480 12524
rect 5440 12444 5444 12476
rect 5476 12444 5480 12476
rect 5440 12396 5480 12444
rect 5440 12364 5444 12396
rect 5476 12364 5480 12396
rect 5440 12316 5480 12364
rect 5440 12284 5444 12316
rect 5476 12284 5480 12316
rect 5440 12236 5480 12284
rect 5440 12204 5444 12236
rect 5476 12204 5480 12236
rect 5440 12156 5480 12204
rect 5440 12124 5444 12156
rect 5476 12124 5480 12156
rect 5440 11836 5480 12124
rect 5440 11804 5444 11836
rect 5476 11804 5480 11836
rect 5440 11756 5480 11804
rect 5440 11724 5444 11756
rect 5476 11724 5480 11756
rect 5440 11676 5480 11724
rect 5440 11644 5444 11676
rect 5476 11644 5480 11676
rect 5440 11596 5480 11644
rect 5440 11564 5444 11596
rect 5476 11564 5480 11596
rect 5440 11516 5480 11564
rect 5440 11484 5444 11516
rect 5476 11484 5480 11516
rect 5440 11436 5480 11484
rect 5440 11404 5444 11436
rect 5476 11404 5480 11436
rect 5440 11074 5480 11404
rect 5440 11046 5446 11074
rect 5474 11046 5480 11074
rect 5440 10876 5480 11046
rect 5440 10844 5444 10876
rect 5476 10844 5480 10876
rect 5440 10796 5480 10844
rect 5440 10764 5444 10796
rect 5476 10764 5480 10796
rect 5440 10716 5480 10764
rect 5440 10684 5444 10716
rect 5476 10684 5480 10716
rect 5440 10636 5480 10684
rect 5440 10604 5444 10636
rect 5476 10604 5480 10636
rect 5440 10556 5480 10604
rect 5440 10524 5444 10556
rect 5476 10524 5480 10556
rect 5440 10476 5480 10524
rect 5440 10444 5444 10476
rect 5476 10444 5480 10476
rect 5440 10396 5480 10444
rect 5440 10364 5444 10396
rect 5476 10364 5480 10396
rect 5440 10316 5480 10364
rect 5440 10284 5444 10316
rect 5476 10284 5480 10316
rect 5440 10236 5480 10284
rect 5440 10204 5444 10236
rect 5476 10204 5480 10236
rect 5440 10156 5480 10204
rect 5440 10124 5444 10156
rect 5476 10124 5480 10156
rect 5440 10076 5480 10124
rect 5440 10044 5444 10076
rect 5476 10044 5480 10076
rect 5440 9996 5480 10044
rect 5440 9964 5444 9996
rect 5476 9964 5480 9996
rect 5440 9916 5480 9964
rect 5440 9884 5444 9916
rect 5476 9884 5480 9916
rect 5440 9836 5480 9884
rect 5440 9804 5444 9836
rect 5476 9804 5480 9836
rect 5440 9756 5480 9804
rect 5440 9724 5444 9756
rect 5476 9724 5480 9756
rect 5440 9356 5480 9724
rect 5440 9324 5444 9356
rect 5476 9324 5480 9356
rect 5440 9276 5480 9324
rect 5440 9244 5444 9276
rect 5476 9244 5480 9276
rect 5440 9196 5480 9244
rect 5440 9164 5444 9196
rect 5476 9164 5480 9196
rect 5440 9114 5480 9164
rect 5440 9086 5446 9114
rect 5474 9086 5480 9114
rect 5440 8954 5480 9086
rect 5440 8926 5446 8954
rect 5474 8926 5480 8954
rect 5440 8876 5480 8926
rect 5440 8844 5444 8876
rect 5476 8844 5480 8876
rect 5440 8796 5480 8844
rect 5440 8764 5444 8796
rect 5476 8764 5480 8796
rect 5440 8716 5480 8764
rect 5440 8684 5444 8716
rect 5476 8684 5480 8716
rect 5440 8636 5480 8684
rect 5440 8604 5444 8636
rect 5476 8604 5480 8636
rect 5440 8556 5480 8604
rect 5440 8524 5444 8556
rect 5476 8524 5480 8556
rect 5440 7994 5480 8524
rect 5440 7966 5446 7994
rect 5474 7966 5480 7994
rect 5440 7834 5480 7966
rect 5440 7806 5446 7834
rect 5474 7806 5480 7834
rect 5440 7636 5480 7806
rect 5440 7604 5444 7636
rect 5476 7604 5480 7636
rect 5440 7556 5480 7604
rect 5440 7524 5444 7556
rect 5476 7524 5480 7556
rect 5440 7476 5480 7524
rect 5440 7444 5444 7476
rect 5476 7444 5480 7476
rect 5440 7396 5480 7444
rect 5440 7364 5444 7396
rect 5476 7364 5480 7396
rect 5440 7316 5480 7364
rect 5440 7284 5444 7316
rect 5476 7284 5480 7316
rect 5440 7236 5480 7284
rect 5440 7204 5444 7236
rect 5476 7204 5480 7236
rect 5440 7156 5480 7204
rect 5440 7124 5444 7156
rect 5476 7124 5480 7156
rect 5440 7076 5480 7124
rect 5440 7044 5444 7076
rect 5476 7044 5480 7076
rect 5440 6756 5480 7044
rect 5440 6724 5444 6756
rect 5476 6724 5480 6756
rect 5440 6676 5480 6724
rect 5440 6644 5444 6676
rect 5476 6644 5480 6676
rect 5440 6596 5480 6644
rect 5440 6564 5444 6596
rect 5476 6564 5480 6596
rect 5440 6516 5480 6564
rect 5440 6484 5444 6516
rect 5476 6484 5480 6516
rect 5440 6436 5480 6484
rect 5440 6404 5444 6436
rect 5476 6404 5480 6436
rect 5440 6356 5480 6404
rect 5440 6324 5444 6356
rect 5476 6324 5480 6356
rect 5440 5796 5480 6324
rect 5440 5764 5444 5796
rect 5476 5764 5480 5796
rect 5440 5716 5480 5764
rect 5440 5684 5444 5716
rect 5476 5684 5480 5716
rect 5440 5636 5480 5684
rect 5440 5604 5444 5636
rect 5476 5604 5480 5636
rect 5440 5556 5480 5604
rect 5440 5524 5444 5556
rect 5476 5524 5480 5556
rect 5440 5476 5480 5524
rect 5440 5444 5444 5476
rect 5476 5444 5480 5476
rect 5440 5396 5480 5444
rect 5440 5364 5444 5396
rect 5476 5364 5480 5396
rect 5440 5316 5480 5364
rect 5440 5284 5444 5316
rect 5476 5284 5480 5316
rect 5440 5236 5480 5284
rect 5440 5204 5444 5236
rect 5476 5204 5480 5236
rect 5440 5156 5480 5204
rect 5440 5124 5444 5156
rect 5476 5124 5480 5156
rect 5440 5076 5480 5124
rect 5440 5044 5444 5076
rect 5476 5044 5480 5076
rect 5440 4996 5480 5044
rect 5440 4964 5444 4996
rect 5476 4964 5480 4996
rect 5440 4436 5480 4964
rect 5440 4404 5444 4436
rect 5476 4404 5480 4436
rect 5440 4356 5480 4404
rect 5440 4324 5444 4356
rect 5476 4324 5480 4356
rect 5440 4276 5480 4324
rect 5440 4244 5444 4276
rect 5476 4244 5480 4276
rect 5440 4196 5480 4244
rect 5440 4164 5444 4196
rect 5476 4164 5480 4196
rect 5440 4116 5480 4164
rect 5440 4084 5444 4116
rect 5476 4084 5480 4116
rect 5440 4036 5480 4084
rect 5440 4004 5444 4036
rect 5476 4004 5480 4036
rect 5440 3956 5480 4004
rect 5440 3924 5444 3956
rect 5476 3924 5480 3956
rect 5440 3156 5480 3924
rect 5440 3124 5444 3156
rect 5476 3124 5480 3156
rect 5440 3076 5480 3124
rect 5440 3044 5444 3076
rect 5476 3044 5480 3076
rect 5440 2996 5480 3044
rect 5440 2964 5444 2996
rect 5476 2964 5480 2996
rect 5440 2916 5480 2964
rect 5440 2884 5444 2916
rect 5476 2884 5480 2916
rect 5440 2836 5480 2884
rect 5440 2804 5444 2836
rect 5476 2804 5480 2836
rect 5440 2756 5480 2804
rect 5440 2724 5444 2756
rect 5476 2724 5480 2756
rect 5440 2676 5480 2724
rect 5440 2644 5444 2676
rect 5476 2644 5480 2676
rect 5440 2596 5480 2644
rect 5440 2564 5444 2596
rect 5476 2564 5480 2596
rect 5440 2516 5480 2564
rect 5440 2484 5444 2516
rect 5476 2484 5480 2516
rect 5440 2436 5480 2484
rect 5440 2404 5444 2436
rect 5476 2404 5480 2436
rect 5440 2356 5480 2404
rect 5440 2324 5444 2356
rect 5476 2324 5480 2356
rect 5440 2276 5480 2324
rect 5440 2244 5444 2276
rect 5476 2244 5480 2276
rect 5440 2196 5480 2244
rect 5440 2164 5444 2196
rect 5476 2164 5480 2196
rect 5440 2116 5480 2164
rect 5440 2084 5444 2116
rect 5476 2084 5480 2116
rect 5440 2036 5480 2084
rect 5440 2004 5444 2036
rect 5476 2004 5480 2036
rect 5440 1636 5480 2004
rect 5440 1604 5444 1636
rect 5476 1604 5480 1636
rect 5440 1556 5480 1604
rect 5440 1524 5444 1556
rect 5476 1524 5480 1556
rect 5440 1476 5480 1524
rect 5440 1444 5444 1476
rect 5476 1444 5480 1476
rect 5440 1396 5480 1444
rect 5440 1364 5444 1396
rect 5476 1364 5480 1396
rect 5440 1316 5480 1364
rect 5440 1284 5444 1316
rect 5476 1284 5480 1316
rect 5440 1236 5480 1284
rect 5440 1204 5444 1236
rect 5476 1204 5480 1236
rect 5440 1156 5480 1204
rect 5440 1124 5444 1156
rect 5476 1124 5480 1156
rect 5440 1076 5480 1124
rect 5440 1044 5444 1076
rect 5476 1044 5480 1076
rect 5440 756 5480 1044
rect 5440 724 5444 756
rect 5476 724 5480 756
rect 5440 676 5480 724
rect 5440 644 5444 676
rect 5476 644 5480 676
rect 5440 596 5480 644
rect 5440 564 5444 596
rect 5476 564 5480 596
rect 5440 196 5480 564
rect 5440 164 5444 196
rect 5476 164 5480 196
rect 5440 116 5480 164
rect 5440 84 5444 116
rect 5476 84 5480 116
rect 5440 36 5480 84
rect 5440 4 5444 36
rect 5476 4 5480 36
rect 5440 -40 5480 4
rect 5520 14036 5560 15400
rect 5600 15396 5640 15400
rect 5600 15364 5604 15396
rect 5636 15364 5640 15396
rect 5600 14116 5640 15364
rect 10160 15396 10200 15400
rect 10160 15364 10164 15396
rect 10196 15364 10200 15396
rect 5680 15316 5720 15320
rect 5680 15284 5684 15316
rect 5716 15284 5720 15316
rect 5680 15240 5720 15284
rect 6720 15316 6760 15320
rect 6720 15284 6724 15316
rect 6756 15284 6760 15316
rect 6720 15240 6760 15284
rect 5680 14160 6760 15240
rect 6800 15316 6840 15320
rect 6800 15284 6804 15316
rect 6836 15284 6840 15316
rect 6800 15240 6840 15284
rect 7840 15316 7880 15320
rect 7840 15284 7844 15316
rect 7876 15284 7880 15316
rect 7840 15240 7880 15284
rect 6800 14160 7880 15240
rect 7920 15316 7960 15320
rect 7920 15284 7924 15316
rect 7956 15284 7960 15316
rect 7920 15240 7960 15284
rect 8960 15316 9000 15320
rect 8960 15284 8964 15316
rect 8996 15284 9000 15316
rect 8960 15240 9000 15284
rect 7920 14160 9000 15240
rect 9040 15316 9080 15320
rect 9040 15284 9044 15316
rect 9076 15284 9080 15316
rect 9040 15240 9080 15284
rect 10080 15316 10120 15320
rect 10080 15284 10084 15316
rect 10116 15284 10120 15316
rect 10080 15240 10120 15284
rect 9040 14160 10120 15240
rect 5600 14084 5604 14116
rect 5636 14084 5640 14116
rect 5600 14080 5640 14084
rect 10160 14116 10200 15364
rect 10160 14084 10164 14116
rect 10196 14084 10200 14116
rect 10160 14080 10200 14084
rect 5520 14004 5524 14036
rect 5556 14004 5560 14036
rect 5520 13716 5560 14004
rect 5520 13684 5524 13716
rect 5556 13684 5560 13716
rect 5520 13396 5560 13684
rect 10240 14036 10280 15444
rect 10240 14004 10244 14036
rect 10276 14004 10280 14036
rect 10240 13716 10280 14004
rect 10320 16836 10360 16920
rect 10320 16804 10324 16836
rect 10356 16804 10360 16836
rect 10320 15556 10360 16804
rect 10320 15524 10324 15556
rect 10356 15524 10360 15556
rect 10320 13956 10360 15524
rect 10320 13924 10324 13956
rect 10356 13924 10360 13956
rect 10320 13796 10360 13924
rect 10320 13764 10324 13796
rect 10356 13764 10360 13796
rect 10320 13760 10360 13764
rect 10400 16756 10440 16920
rect 10400 16724 10404 16756
rect 10436 16724 10440 16756
rect 10400 13876 10440 16724
rect 10400 13844 10404 13876
rect 10436 13844 10440 13876
rect 10400 13760 10440 13844
rect 10480 16836 10520 16920
rect 10480 16804 10484 16836
rect 10516 16804 10520 16836
rect 10480 15556 10520 16804
rect 10480 15524 10484 15556
rect 10516 15524 10520 15556
rect 10480 13956 10520 15524
rect 10480 13924 10484 13956
rect 10516 13924 10520 13956
rect 10480 13796 10520 13924
rect 10480 13764 10484 13796
rect 10516 13764 10520 13796
rect 10480 13760 10520 13764
rect 10560 16916 10600 16920
rect 10560 16884 10564 16916
rect 10596 16884 10600 16916
rect 10560 15476 10600 16884
rect 10560 15444 10564 15476
rect 10596 15444 10600 15476
rect 10560 14036 10600 15444
rect 10560 14004 10564 14036
rect 10596 14004 10600 14036
rect 10240 13684 10244 13716
rect 10276 13684 10280 13716
rect 10240 13680 10280 13684
rect 10560 13716 10600 14004
rect 10560 13684 10564 13716
rect 10596 13684 10600 13716
rect 10560 13680 10600 13684
rect 5520 13364 5524 13396
rect 5556 13364 5560 13396
rect 5520 13356 5560 13364
rect 5520 13324 5524 13356
rect 5556 13324 5560 13356
rect 5520 13316 5560 13324
rect 5520 13284 5524 13316
rect 5556 13284 5560 13316
rect 5520 13276 5560 13284
rect 5520 13244 5524 13276
rect 5556 13244 5560 13276
rect 5520 13236 5560 13244
rect 5520 13204 5524 13236
rect 5556 13204 5560 13236
rect 5520 12636 5560 13204
rect 5680 13396 5720 13400
rect 5680 13364 5684 13396
rect 5716 13364 5720 13396
rect 5680 13356 5720 13364
rect 5680 13324 5684 13356
rect 5716 13324 5720 13356
rect 5680 13316 5720 13324
rect 5680 13284 5684 13316
rect 5716 13284 5720 13316
rect 5680 13276 5720 13284
rect 5680 13244 5684 13276
rect 5716 13244 5720 13276
rect 5680 13236 5720 13244
rect 5680 13204 5684 13236
rect 5716 13204 5720 13236
rect 5520 12604 5524 12636
rect 5556 12604 5560 12636
rect 5520 12556 5560 12604
rect 5520 12524 5524 12556
rect 5556 12524 5560 12556
rect 5520 12476 5560 12524
rect 5520 12444 5524 12476
rect 5556 12444 5560 12476
rect 5520 12396 5560 12444
rect 5520 12364 5524 12396
rect 5556 12364 5560 12396
rect 5520 12316 5560 12364
rect 5520 12284 5524 12316
rect 5556 12284 5560 12316
rect 5520 12236 5560 12284
rect 5520 12204 5524 12236
rect 5556 12204 5560 12236
rect 5520 12156 5560 12204
rect 5520 12124 5524 12156
rect 5556 12124 5560 12156
rect 5520 11836 5560 12124
rect 5520 11804 5524 11836
rect 5556 11804 5560 11836
rect 5520 11756 5560 11804
rect 5520 11724 5524 11756
rect 5556 11724 5560 11756
rect 5520 11676 5560 11724
rect 5520 11644 5524 11676
rect 5556 11644 5560 11676
rect 5520 11596 5560 11644
rect 5520 11564 5524 11596
rect 5556 11564 5560 11596
rect 5520 11516 5560 11564
rect 5520 11484 5524 11516
rect 5556 11484 5560 11516
rect 5520 11436 5560 11484
rect 5520 11404 5524 11436
rect 5556 11404 5560 11436
rect 5520 11314 5560 11404
rect 5520 11286 5526 11314
rect 5554 11286 5560 11314
rect 5520 11154 5560 11286
rect 5520 11126 5526 11154
rect 5554 11126 5560 11154
rect 5520 10994 5560 11126
rect 5520 10966 5526 10994
rect 5554 10966 5560 10994
rect 5520 10876 5560 10966
rect 5520 10844 5524 10876
rect 5556 10844 5560 10876
rect 5520 10796 5560 10844
rect 5520 10764 5524 10796
rect 5556 10764 5560 10796
rect 5520 10716 5560 10764
rect 5520 10684 5524 10716
rect 5556 10684 5560 10716
rect 5520 10636 5560 10684
rect 5520 10604 5524 10636
rect 5556 10604 5560 10636
rect 5520 10556 5560 10604
rect 5520 10524 5524 10556
rect 5556 10524 5560 10556
rect 5520 10476 5560 10524
rect 5520 10444 5524 10476
rect 5556 10444 5560 10476
rect 5520 10396 5560 10444
rect 5520 10364 5524 10396
rect 5556 10364 5560 10396
rect 5520 10316 5560 10364
rect 5520 10284 5524 10316
rect 5556 10284 5560 10316
rect 5520 10236 5560 10284
rect 5520 10204 5524 10236
rect 5556 10204 5560 10236
rect 5520 10156 5560 10204
rect 5520 10124 5524 10156
rect 5556 10124 5560 10156
rect 5520 10076 5560 10124
rect 5520 10044 5524 10076
rect 5556 10044 5560 10076
rect 5520 9996 5560 10044
rect 5520 9964 5524 9996
rect 5556 9964 5560 9996
rect 5520 9916 5560 9964
rect 5520 9884 5524 9916
rect 5556 9884 5560 9916
rect 5520 9836 5560 9884
rect 5520 9804 5524 9836
rect 5556 9804 5560 9836
rect 5520 9756 5560 9804
rect 5520 9724 5524 9756
rect 5556 9724 5560 9756
rect 5520 9356 5560 9724
rect 5520 9324 5524 9356
rect 5556 9324 5560 9356
rect 5520 9276 5560 9324
rect 5520 9244 5524 9276
rect 5556 9244 5560 9276
rect 5520 9196 5560 9244
rect 5520 9164 5524 9196
rect 5556 9164 5560 9196
rect 5520 8876 5560 9164
rect 5520 8844 5524 8876
rect 5556 8844 5560 8876
rect 5520 8796 5560 8844
rect 5520 8764 5524 8796
rect 5556 8764 5560 8796
rect 5520 8716 5560 8764
rect 5520 8684 5524 8716
rect 5556 8684 5560 8716
rect 5520 8636 5560 8684
rect 5520 8604 5524 8636
rect 5556 8604 5560 8636
rect 5520 8556 5560 8604
rect 5520 8524 5524 8556
rect 5556 8524 5560 8556
rect 5520 8314 5560 8524
rect 5520 8286 5526 8314
rect 5554 8286 5560 8314
rect 5520 8154 5560 8286
rect 5520 8126 5526 8154
rect 5554 8126 5560 8154
rect 5520 8074 5560 8126
rect 5520 8046 5526 8074
rect 5554 8046 5560 8074
rect 5520 7754 5560 8046
rect 5520 7726 5526 7754
rect 5554 7726 5560 7754
rect 5520 7636 5560 7726
rect 5520 7604 5524 7636
rect 5556 7604 5560 7636
rect 5520 7556 5560 7604
rect 5520 7524 5524 7556
rect 5556 7524 5560 7556
rect 5520 7476 5560 7524
rect 5520 7444 5524 7476
rect 5556 7444 5560 7476
rect 5520 7396 5560 7444
rect 5520 7364 5524 7396
rect 5556 7364 5560 7396
rect 5520 7316 5560 7364
rect 5520 7284 5524 7316
rect 5556 7284 5560 7316
rect 5520 7236 5560 7284
rect 5520 7204 5524 7236
rect 5556 7204 5560 7236
rect 5520 7156 5560 7204
rect 5520 7124 5524 7156
rect 5556 7124 5560 7156
rect 5520 7076 5560 7124
rect 5520 7044 5524 7076
rect 5556 7044 5560 7076
rect 5520 6756 5560 7044
rect 5520 6724 5524 6756
rect 5556 6724 5560 6756
rect 5520 6676 5560 6724
rect 5520 6644 5524 6676
rect 5556 6644 5560 6676
rect 5520 6596 5560 6644
rect 5520 6564 5524 6596
rect 5556 6564 5560 6596
rect 5520 6516 5560 6564
rect 5520 6484 5524 6516
rect 5556 6484 5560 6516
rect 5520 6436 5560 6484
rect 5520 6404 5524 6436
rect 5556 6404 5560 6436
rect 5520 6356 5560 6404
rect 5520 6324 5524 6356
rect 5556 6324 5560 6356
rect 5520 5796 5560 6324
rect 5520 5764 5524 5796
rect 5556 5764 5560 5796
rect 5520 5716 5560 5764
rect 5520 5684 5524 5716
rect 5556 5684 5560 5716
rect 5520 5636 5560 5684
rect 5520 5604 5524 5636
rect 5556 5604 5560 5636
rect 5520 5556 5560 5604
rect 5520 5524 5524 5556
rect 5556 5524 5560 5556
rect 5520 5476 5560 5524
rect 5520 5444 5524 5476
rect 5556 5444 5560 5476
rect 5520 5396 5560 5444
rect 5520 5364 5524 5396
rect 5556 5364 5560 5396
rect 5520 5316 5560 5364
rect 5520 5284 5524 5316
rect 5556 5284 5560 5316
rect 5520 5236 5560 5284
rect 5520 5204 5524 5236
rect 5556 5204 5560 5236
rect 5520 5156 5560 5204
rect 5520 5124 5524 5156
rect 5556 5124 5560 5156
rect 5520 5076 5560 5124
rect 5520 5044 5524 5076
rect 5556 5044 5560 5076
rect 5520 4996 5560 5044
rect 5520 4964 5524 4996
rect 5556 4964 5560 4996
rect 5520 4436 5560 4964
rect 5520 4404 5524 4436
rect 5556 4404 5560 4436
rect 5520 4356 5560 4404
rect 5520 4324 5524 4356
rect 5556 4324 5560 4356
rect 5520 4276 5560 4324
rect 5520 4244 5524 4276
rect 5556 4244 5560 4276
rect 5520 4196 5560 4244
rect 5520 4164 5524 4196
rect 5556 4164 5560 4196
rect 5520 4116 5560 4164
rect 5520 4084 5524 4116
rect 5556 4084 5560 4116
rect 5520 4036 5560 4084
rect 5520 4004 5524 4036
rect 5556 4004 5560 4036
rect 5520 3956 5560 4004
rect 5520 3924 5524 3956
rect 5556 3924 5560 3956
rect 5520 3156 5560 3924
rect 5520 3124 5524 3156
rect 5556 3124 5560 3156
rect 5520 3076 5560 3124
rect 5520 3044 5524 3076
rect 5556 3044 5560 3076
rect 5520 2996 5560 3044
rect 5520 2964 5524 2996
rect 5556 2964 5560 2996
rect 5520 2916 5560 2964
rect 5520 2884 5524 2916
rect 5556 2884 5560 2916
rect 5520 2836 5560 2884
rect 5520 2804 5524 2836
rect 5556 2804 5560 2836
rect 5520 2756 5560 2804
rect 5520 2724 5524 2756
rect 5556 2724 5560 2756
rect 5520 2676 5560 2724
rect 5520 2644 5524 2676
rect 5556 2644 5560 2676
rect 5520 2596 5560 2644
rect 5520 2564 5524 2596
rect 5556 2564 5560 2596
rect 5520 2516 5560 2564
rect 5520 2484 5524 2516
rect 5556 2484 5560 2516
rect 5520 2436 5560 2484
rect 5520 2404 5524 2436
rect 5556 2404 5560 2436
rect 5520 2356 5560 2404
rect 5520 2324 5524 2356
rect 5556 2324 5560 2356
rect 5520 2276 5560 2324
rect 5520 2244 5524 2276
rect 5556 2244 5560 2276
rect 5520 2196 5560 2244
rect 5520 2164 5524 2196
rect 5556 2164 5560 2196
rect 5520 2116 5560 2164
rect 5520 2084 5524 2116
rect 5556 2084 5560 2116
rect 5520 2036 5560 2084
rect 5520 2004 5524 2036
rect 5556 2004 5560 2036
rect 5520 1636 5560 2004
rect 5520 1604 5524 1636
rect 5556 1604 5560 1636
rect 5520 1556 5560 1604
rect 5520 1524 5524 1556
rect 5556 1524 5560 1556
rect 5520 1476 5560 1524
rect 5520 1444 5524 1476
rect 5556 1444 5560 1476
rect 5520 1396 5560 1444
rect 5520 1364 5524 1396
rect 5556 1364 5560 1396
rect 5520 1316 5560 1364
rect 5520 1284 5524 1316
rect 5556 1284 5560 1316
rect 5520 1236 5560 1284
rect 5520 1204 5524 1236
rect 5556 1204 5560 1236
rect 5520 1156 5560 1204
rect 5520 1124 5524 1156
rect 5556 1124 5560 1156
rect 5520 1076 5560 1124
rect 5520 1044 5524 1076
rect 5556 1044 5560 1076
rect 5520 756 5560 1044
rect 5520 724 5524 756
rect 5556 724 5560 756
rect 5520 676 5560 724
rect 5520 644 5524 676
rect 5556 644 5560 676
rect 5520 596 5560 644
rect 5520 564 5524 596
rect 5556 564 5560 596
rect 5520 196 5560 564
rect 5520 164 5524 196
rect 5556 164 5560 196
rect 5520 116 5560 164
rect 5520 84 5524 116
rect 5556 84 5560 116
rect 5520 36 5560 84
rect 5520 4 5524 36
rect 5556 4 5560 36
rect 5520 -40 5560 4
rect 5600 11234 5640 12680
rect 5600 11206 5606 11234
rect 5634 11206 5640 11234
rect 5600 8234 5640 11206
rect 5600 8206 5606 8234
rect 5634 8206 5640 8234
rect 5600 -40 5640 8206
rect 5680 12636 5720 13204
rect 5840 13396 5880 13400
rect 5840 13364 5844 13396
rect 5876 13364 5880 13396
rect 5840 13356 5880 13364
rect 5840 13324 5844 13356
rect 5876 13324 5880 13356
rect 5840 13316 5880 13324
rect 5840 13284 5844 13316
rect 5876 13284 5880 13316
rect 5840 13276 5880 13284
rect 5840 13244 5844 13276
rect 5876 13244 5880 13276
rect 5840 13236 5880 13244
rect 5840 13204 5844 13236
rect 5876 13204 5880 13236
rect 5680 12604 5684 12636
rect 5716 12604 5720 12636
rect 5680 12556 5720 12604
rect 5680 12524 5684 12556
rect 5716 12524 5720 12556
rect 5680 12476 5720 12524
rect 5680 12444 5684 12476
rect 5716 12444 5720 12476
rect 5680 12396 5720 12444
rect 5680 12364 5684 12396
rect 5716 12364 5720 12396
rect 5680 12316 5720 12364
rect 5680 12284 5684 12316
rect 5716 12284 5720 12316
rect 5680 12236 5720 12284
rect 5680 12204 5684 12236
rect 5716 12204 5720 12236
rect 5680 12156 5720 12204
rect 5680 12124 5684 12156
rect 5716 12124 5720 12156
rect 5680 11836 5720 12124
rect 5680 11804 5684 11836
rect 5716 11804 5720 11836
rect 5680 11756 5720 11804
rect 5680 11724 5684 11756
rect 5716 11724 5720 11756
rect 5680 11676 5720 11724
rect 5680 11644 5684 11676
rect 5716 11644 5720 11676
rect 5680 11596 5720 11644
rect 5680 11564 5684 11596
rect 5716 11564 5720 11596
rect 5680 11516 5720 11564
rect 5680 11484 5684 11516
rect 5716 11484 5720 11516
rect 5680 11436 5720 11484
rect 5680 11404 5684 11436
rect 5716 11404 5720 11436
rect 5680 11314 5720 11404
rect 5680 11286 5686 11314
rect 5714 11286 5720 11314
rect 5680 11154 5720 11286
rect 5680 11126 5686 11154
rect 5714 11126 5720 11154
rect 5680 10876 5720 11126
rect 5680 10844 5684 10876
rect 5716 10844 5720 10876
rect 5680 10796 5720 10844
rect 5680 10764 5684 10796
rect 5716 10764 5720 10796
rect 5680 10716 5720 10764
rect 5680 10684 5684 10716
rect 5716 10684 5720 10716
rect 5680 10636 5720 10684
rect 5680 10604 5684 10636
rect 5716 10604 5720 10636
rect 5680 10556 5720 10604
rect 5680 10524 5684 10556
rect 5716 10524 5720 10556
rect 5680 10476 5720 10524
rect 5680 10444 5684 10476
rect 5716 10444 5720 10476
rect 5680 10396 5720 10444
rect 5680 10364 5684 10396
rect 5716 10364 5720 10396
rect 5680 10316 5720 10364
rect 5680 10284 5684 10316
rect 5716 10284 5720 10316
rect 5680 10236 5720 10284
rect 5680 10204 5684 10236
rect 5716 10204 5720 10236
rect 5680 10156 5720 10204
rect 5680 10124 5684 10156
rect 5716 10124 5720 10156
rect 5680 10076 5720 10124
rect 5680 10044 5684 10076
rect 5716 10044 5720 10076
rect 5680 9996 5720 10044
rect 5680 9964 5684 9996
rect 5716 9964 5720 9996
rect 5680 9916 5720 9964
rect 5680 9884 5684 9916
rect 5716 9884 5720 9916
rect 5680 9836 5720 9884
rect 5680 9804 5684 9836
rect 5716 9804 5720 9836
rect 5680 9756 5720 9804
rect 5680 9724 5684 9756
rect 5716 9724 5720 9756
rect 5680 9356 5720 9724
rect 5680 9324 5684 9356
rect 5716 9324 5720 9356
rect 5680 9276 5720 9324
rect 5680 9244 5684 9276
rect 5716 9244 5720 9276
rect 5680 9196 5720 9244
rect 5680 9164 5684 9196
rect 5716 9164 5720 9196
rect 5680 8876 5720 9164
rect 5680 8844 5684 8876
rect 5716 8844 5720 8876
rect 5680 8796 5720 8844
rect 5680 8764 5684 8796
rect 5716 8764 5720 8796
rect 5680 8716 5720 8764
rect 5680 8684 5684 8716
rect 5716 8684 5720 8716
rect 5680 8636 5720 8684
rect 5680 8604 5684 8636
rect 5716 8604 5720 8636
rect 5680 8556 5720 8604
rect 5680 8524 5684 8556
rect 5716 8524 5720 8556
rect 5680 8474 5720 8524
rect 5680 8446 5686 8474
rect 5714 8446 5720 8474
rect 5680 8314 5720 8446
rect 5680 8286 5686 8314
rect 5714 8286 5720 8314
rect 5680 8154 5720 8286
rect 5680 8126 5686 8154
rect 5714 8126 5720 8154
rect 5680 7636 5720 8126
rect 5680 7604 5684 7636
rect 5716 7604 5720 7636
rect 5680 7556 5720 7604
rect 5680 7524 5684 7556
rect 5716 7524 5720 7556
rect 5680 7476 5720 7524
rect 5680 7444 5684 7476
rect 5716 7444 5720 7476
rect 5680 7396 5720 7444
rect 5680 7364 5684 7396
rect 5716 7364 5720 7396
rect 5680 7316 5720 7364
rect 5680 7284 5684 7316
rect 5716 7284 5720 7316
rect 5680 7236 5720 7284
rect 5680 7204 5684 7236
rect 5716 7204 5720 7236
rect 5680 7156 5720 7204
rect 5680 7124 5684 7156
rect 5716 7124 5720 7156
rect 5680 7076 5720 7124
rect 5680 7044 5684 7076
rect 5716 7044 5720 7076
rect 5680 6756 5720 7044
rect 5680 6724 5684 6756
rect 5716 6724 5720 6756
rect 5680 6676 5720 6724
rect 5680 6644 5684 6676
rect 5716 6644 5720 6676
rect 5680 6596 5720 6644
rect 5680 6564 5684 6596
rect 5716 6564 5720 6596
rect 5680 6516 5720 6564
rect 5680 6484 5684 6516
rect 5716 6484 5720 6516
rect 5680 6436 5720 6484
rect 5680 6404 5684 6436
rect 5716 6404 5720 6436
rect 5680 6356 5720 6404
rect 5680 6324 5684 6356
rect 5716 6324 5720 6356
rect 5680 5796 5720 6324
rect 5680 5764 5684 5796
rect 5716 5764 5720 5796
rect 5680 5716 5720 5764
rect 5680 5684 5684 5716
rect 5716 5684 5720 5716
rect 5680 5636 5720 5684
rect 5680 5604 5684 5636
rect 5716 5604 5720 5636
rect 5680 5556 5720 5604
rect 5680 5524 5684 5556
rect 5716 5524 5720 5556
rect 5680 5476 5720 5524
rect 5680 5444 5684 5476
rect 5716 5444 5720 5476
rect 5680 5396 5720 5444
rect 5680 5364 5684 5396
rect 5716 5364 5720 5396
rect 5680 5316 5720 5364
rect 5680 5284 5684 5316
rect 5716 5284 5720 5316
rect 5680 5236 5720 5284
rect 5680 5204 5684 5236
rect 5716 5204 5720 5236
rect 5680 5156 5720 5204
rect 5680 5124 5684 5156
rect 5716 5124 5720 5156
rect 5680 5076 5720 5124
rect 5680 5044 5684 5076
rect 5716 5044 5720 5076
rect 5680 4996 5720 5044
rect 5680 4964 5684 4996
rect 5716 4964 5720 4996
rect 5680 4436 5720 4964
rect 5680 4404 5684 4436
rect 5716 4404 5720 4436
rect 5680 4356 5720 4404
rect 5680 4324 5684 4356
rect 5716 4324 5720 4356
rect 5680 4276 5720 4324
rect 5680 4244 5684 4276
rect 5716 4244 5720 4276
rect 5680 4196 5720 4244
rect 5680 4164 5684 4196
rect 5716 4164 5720 4196
rect 5680 4116 5720 4164
rect 5680 4084 5684 4116
rect 5716 4084 5720 4116
rect 5680 4036 5720 4084
rect 5680 4004 5684 4036
rect 5716 4004 5720 4036
rect 5680 3956 5720 4004
rect 5680 3924 5684 3956
rect 5716 3924 5720 3956
rect 5680 3156 5720 3924
rect 5680 3124 5684 3156
rect 5716 3124 5720 3156
rect 5680 3076 5720 3124
rect 5680 3044 5684 3076
rect 5716 3044 5720 3076
rect 5680 2996 5720 3044
rect 5680 2964 5684 2996
rect 5716 2964 5720 2996
rect 5680 2916 5720 2964
rect 5680 2884 5684 2916
rect 5716 2884 5720 2916
rect 5680 2836 5720 2884
rect 5680 2804 5684 2836
rect 5716 2804 5720 2836
rect 5680 2756 5720 2804
rect 5680 2724 5684 2756
rect 5716 2724 5720 2756
rect 5680 2676 5720 2724
rect 5680 2644 5684 2676
rect 5716 2644 5720 2676
rect 5680 2596 5720 2644
rect 5680 2564 5684 2596
rect 5716 2564 5720 2596
rect 5680 2516 5720 2564
rect 5680 2484 5684 2516
rect 5716 2484 5720 2516
rect 5680 2436 5720 2484
rect 5680 2404 5684 2436
rect 5716 2404 5720 2436
rect 5680 2356 5720 2404
rect 5680 2324 5684 2356
rect 5716 2324 5720 2356
rect 5680 2276 5720 2324
rect 5680 2244 5684 2276
rect 5716 2244 5720 2276
rect 5680 2196 5720 2244
rect 5680 2164 5684 2196
rect 5716 2164 5720 2196
rect 5680 2116 5720 2164
rect 5680 2084 5684 2116
rect 5716 2084 5720 2116
rect 5680 2036 5720 2084
rect 5680 2004 5684 2036
rect 5716 2004 5720 2036
rect 5680 1636 5720 2004
rect 5680 1604 5684 1636
rect 5716 1604 5720 1636
rect 5680 1556 5720 1604
rect 5680 1524 5684 1556
rect 5716 1524 5720 1556
rect 5680 1476 5720 1524
rect 5680 1444 5684 1476
rect 5716 1444 5720 1476
rect 5680 1396 5720 1444
rect 5680 1364 5684 1396
rect 5716 1364 5720 1396
rect 5680 1316 5720 1364
rect 5680 1284 5684 1316
rect 5716 1284 5720 1316
rect 5680 1236 5720 1284
rect 5680 1204 5684 1236
rect 5716 1204 5720 1236
rect 5680 1156 5720 1204
rect 5680 1124 5684 1156
rect 5716 1124 5720 1156
rect 5680 1076 5720 1124
rect 5680 1044 5684 1076
rect 5716 1044 5720 1076
rect 5680 756 5720 1044
rect 5680 724 5684 756
rect 5716 724 5720 756
rect 5680 676 5720 724
rect 5680 644 5684 676
rect 5716 644 5720 676
rect 5680 596 5720 644
rect 5680 564 5684 596
rect 5716 564 5720 596
rect 5680 196 5720 564
rect 5680 164 5684 196
rect 5716 164 5720 196
rect 5680 116 5720 164
rect 5680 84 5684 116
rect 5716 84 5720 116
rect 5680 36 5720 84
rect 5680 4 5684 36
rect 5716 4 5720 36
rect 5680 -40 5720 4
rect 5760 8394 5800 12680
rect 5760 8366 5766 8394
rect 5794 8366 5800 8394
rect 5760 -40 5800 8366
rect 5840 12636 5880 13204
rect 6160 13396 6200 13400
rect 6160 13364 6164 13396
rect 6196 13364 6200 13396
rect 6160 13356 6200 13364
rect 6160 13324 6164 13356
rect 6196 13324 6200 13356
rect 6160 13316 6200 13324
rect 6160 13284 6164 13316
rect 6196 13284 6200 13316
rect 6160 13276 6200 13284
rect 6160 13244 6164 13276
rect 6196 13244 6200 13276
rect 6160 13236 6200 13244
rect 6160 13204 6164 13236
rect 6196 13204 6200 13236
rect 5840 12604 5844 12636
rect 5876 12604 5880 12636
rect 5840 12556 5880 12604
rect 5840 12524 5844 12556
rect 5876 12524 5880 12556
rect 5840 12476 5880 12524
rect 5840 12444 5844 12476
rect 5876 12444 5880 12476
rect 5840 12396 5880 12444
rect 5840 12364 5844 12396
rect 5876 12364 5880 12396
rect 5840 12316 5880 12364
rect 5840 12284 5844 12316
rect 5876 12284 5880 12316
rect 5840 12236 5880 12284
rect 5840 12204 5844 12236
rect 5876 12204 5880 12236
rect 5840 12156 5880 12204
rect 5840 12124 5844 12156
rect 5876 12124 5880 12156
rect 5840 11836 5880 12124
rect 5840 11804 5844 11836
rect 5876 11804 5880 11836
rect 5840 11756 5880 11804
rect 5840 11724 5844 11756
rect 5876 11724 5880 11756
rect 5840 11676 5880 11724
rect 5840 11644 5844 11676
rect 5876 11644 5880 11676
rect 5840 11596 5880 11644
rect 5840 11564 5844 11596
rect 5876 11564 5880 11596
rect 5840 11516 5880 11564
rect 5840 11484 5844 11516
rect 5876 11484 5880 11516
rect 5840 11436 5880 11484
rect 5840 11404 5844 11436
rect 5876 11404 5880 11436
rect 5840 10876 5880 11404
rect 5840 10844 5844 10876
rect 5876 10844 5880 10876
rect 5840 10796 5880 10844
rect 5840 10764 5844 10796
rect 5876 10764 5880 10796
rect 5840 10716 5880 10764
rect 5840 10684 5844 10716
rect 5876 10684 5880 10716
rect 5840 10636 5880 10684
rect 5840 10604 5844 10636
rect 5876 10604 5880 10636
rect 5840 10556 5880 10604
rect 5840 10524 5844 10556
rect 5876 10524 5880 10556
rect 5840 10476 5880 10524
rect 5840 10444 5844 10476
rect 5876 10444 5880 10476
rect 5840 10396 5880 10444
rect 5840 10364 5844 10396
rect 5876 10364 5880 10396
rect 5840 10316 5880 10364
rect 5840 10284 5844 10316
rect 5876 10284 5880 10316
rect 5840 10236 5880 10284
rect 5840 10204 5844 10236
rect 5876 10204 5880 10236
rect 5840 10156 5880 10204
rect 5840 10124 5844 10156
rect 5876 10124 5880 10156
rect 5840 10076 5880 10124
rect 5840 10044 5844 10076
rect 5876 10044 5880 10076
rect 5840 9996 5880 10044
rect 5840 9964 5844 9996
rect 5876 9964 5880 9996
rect 5840 9916 5880 9964
rect 5840 9884 5844 9916
rect 5876 9884 5880 9916
rect 5840 9836 5880 9884
rect 5840 9804 5844 9836
rect 5876 9804 5880 9836
rect 5840 9756 5880 9804
rect 5840 9724 5844 9756
rect 5876 9724 5880 9756
rect 5840 9356 5880 9724
rect 5840 9324 5844 9356
rect 5876 9324 5880 9356
rect 5840 9276 5880 9324
rect 5840 9244 5844 9276
rect 5876 9244 5880 9276
rect 5840 9196 5880 9244
rect 5840 9164 5844 9196
rect 5876 9164 5880 9196
rect 5840 8876 5880 9164
rect 5840 8844 5844 8876
rect 5876 8844 5880 8876
rect 5840 8796 5880 8844
rect 5840 8764 5844 8796
rect 5876 8764 5880 8796
rect 5840 8716 5880 8764
rect 5840 8684 5844 8716
rect 5876 8684 5880 8716
rect 5840 8636 5880 8684
rect 5840 8604 5844 8636
rect 5876 8604 5880 8636
rect 5840 8556 5880 8604
rect 5840 8524 5844 8556
rect 5876 8524 5880 8556
rect 5840 8474 5880 8524
rect 5840 8446 5846 8474
rect 5874 8446 5880 8474
rect 5840 8314 5880 8446
rect 5840 8286 5846 8314
rect 5874 8286 5880 8314
rect 5840 7636 5880 8286
rect 5840 7604 5844 7636
rect 5876 7604 5880 7636
rect 5840 7556 5880 7604
rect 5840 7524 5844 7556
rect 5876 7524 5880 7556
rect 5840 7476 5880 7524
rect 5840 7444 5844 7476
rect 5876 7444 5880 7476
rect 5840 7396 5880 7444
rect 5840 7364 5844 7396
rect 5876 7364 5880 7396
rect 5840 7316 5880 7364
rect 5840 7284 5844 7316
rect 5876 7284 5880 7316
rect 5840 7236 5880 7284
rect 5840 7204 5844 7236
rect 5876 7204 5880 7236
rect 5840 7156 5880 7204
rect 5840 7124 5844 7156
rect 5876 7124 5880 7156
rect 5840 7076 5880 7124
rect 5840 7044 5844 7076
rect 5876 7044 5880 7076
rect 5840 6756 5880 7044
rect 5840 6724 5844 6756
rect 5876 6724 5880 6756
rect 5840 6676 5880 6724
rect 5840 6644 5844 6676
rect 5876 6644 5880 6676
rect 5840 6596 5880 6644
rect 5840 6564 5844 6596
rect 5876 6564 5880 6596
rect 5840 6516 5880 6564
rect 5840 6484 5844 6516
rect 5876 6484 5880 6516
rect 5840 6436 5880 6484
rect 5840 6404 5844 6436
rect 5876 6404 5880 6436
rect 5840 6356 5880 6404
rect 5840 6324 5844 6356
rect 5876 6324 5880 6356
rect 5840 5796 5880 6324
rect 5840 5764 5844 5796
rect 5876 5764 5880 5796
rect 5840 5716 5880 5764
rect 5840 5684 5844 5716
rect 5876 5684 5880 5716
rect 5840 5636 5880 5684
rect 5840 5604 5844 5636
rect 5876 5604 5880 5636
rect 5840 5556 5880 5604
rect 5840 5524 5844 5556
rect 5876 5524 5880 5556
rect 5840 5476 5880 5524
rect 5840 5444 5844 5476
rect 5876 5444 5880 5476
rect 5840 5396 5880 5444
rect 5840 5364 5844 5396
rect 5876 5364 5880 5396
rect 5840 5316 5880 5364
rect 5840 5284 5844 5316
rect 5876 5284 5880 5316
rect 5840 5236 5880 5284
rect 5840 5204 5844 5236
rect 5876 5204 5880 5236
rect 5840 5156 5880 5204
rect 5840 5124 5844 5156
rect 5876 5124 5880 5156
rect 5840 5076 5880 5124
rect 5840 5044 5844 5076
rect 5876 5044 5880 5076
rect 5840 4996 5880 5044
rect 5840 4964 5844 4996
rect 5876 4964 5880 4996
rect 5840 4436 5880 4964
rect 5840 4404 5844 4436
rect 5876 4404 5880 4436
rect 5840 4356 5880 4404
rect 5840 4324 5844 4356
rect 5876 4324 5880 4356
rect 5840 4276 5880 4324
rect 5840 4244 5844 4276
rect 5876 4244 5880 4276
rect 5840 4196 5880 4244
rect 5840 4164 5844 4196
rect 5876 4164 5880 4196
rect 5840 4116 5880 4164
rect 5840 4084 5844 4116
rect 5876 4084 5880 4116
rect 5840 4036 5880 4084
rect 5840 4004 5844 4036
rect 5876 4004 5880 4036
rect 5840 3956 5880 4004
rect 5840 3924 5844 3956
rect 5876 3924 5880 3956
rect 5840 3156 5880 3924
rect 5840 3124 5844 3156
rect 5876 3124 5880 3156
rect 5840 3076 5880 3124
rect 5840 3044 5844 3076
rect 5876 3044 5880 3076
rect 5840 2996 5880 3044
rect 5840 2964 5844 2996
rect 5876 2964 5880 2996
rect 5840 2916 5880 2964
rect 5840 2884 5844 2916
rect 5876 2884 5880 2916
rect 5840 2836 5880 2884
rect 5840 2804 5844 2836
rect 5876 2804 5880 2836
rect 5840 2756 5880 2804
rect 5840 2724 5844 2756
rect 5876 2724 5880 2756
rect 5840 2676 5880 2724
rect 5840 2644 5844 2676
rect 5876 2644 5880 2676
rect 5840 2596 5880 2644
rect 5840 2564 5844 2596
rect 5876 2564 5880 2596
rect 5840 2516 5880 2564
rect 5840 2484 5844 2516
rect 5876 2484 5880 2516
rect 5840 2436 5880 2484
rect 5840 2404 5844 2436
rect 5876 2404 5880 2436
rect 5840 2356 5880 2404
rect 5840 2324 5844 2356
rect 5876 2324 5880 2356
rect 5840 2276 5880 2324
rect 5840 2244 5844 2276
rect 5876 2244 5880 2276
rect 5840 2196 5880 2244
rect 5840 2164 5844 2196
rect 5876 2164 5880 2196
rect 5840 2116 5880 2164
rect 5840 2084 5844 2116
rect 5876 2084 5880 2116
rect 5840 2036 5880 2084
rect 5840 2004 5844 2036
rect 5876 2004 5880 2036
rect 5840 1636 5880 2004
rect 5840 1604 5844 1636
rect 5876 1604 5880 1636
rect 5840 1556 5880 1604
rect 5840 1524 5844 1556
rect 5876 1524 5880 1556
rect 5840 1476 5880 1524
rect 5840 1444 5844 1476
rect 5876 1444 5880 1476
rect 5840 1396 5880 1444
rect 5840 1364 5844 1396
rect 5876 1364 5880 1396
rect 5840 1316 5880 1364
rect 5840 1284 5844 1316
rect 5876 1284 5880 1316
rect 5840 1236 5880 1284
rect 5840 1204 5844 1236
rect 5876 1204 5880 1236
rect 5840 1156 5880 1204
rect 5840 1124 5844 1156
rect 5876 1124 5880 1156
rect 5840 1076 5880 1124
rect 5840 1044 5844 1076
rect 5876 1044 5880 1076
rect 5840 756 5880 1044
rect 5840 724 5844 756
rect 5876 724 5880 756
rect 5840 676 5880 724
rect 5840 644 5844 676
rect 5876 644 5880 676
rect 5840 596 5880 644
rect 5840 564 5844 596
rect 5876 564 5880 596
rect 5840 196 5880 564
rect 5840 164 5844 196
rect 5876 164 5880 196
rect 5840 116 5880 164
rect 5840 84 5844 116
rect 5876 84 5880 116
rect 5840 36 5880 84
rect 5840 4 5844 36
rect 5876 4 5880 36
rect 5840 -40 5880 4
rect 5920 12916 5960 12920
rect 5920 12884 5924 12916
rect 5956 12884 5960 12916
rect 5920 12876 5960 12884
rect 5920 12844 5924 12876
rect 5956 12844 5960 12876
rect 5920 12836 5960 12844
rect 5920 12804 5924 12836
rect 5956 12804 5960 12836
rect 5920 12796 5960 12804
rect 5920 12764 5924 12796
rect 5956 12764 5960 12796
rect 5920 12756 5960 12764
rect 5920 12724 5924 12756
rect 5956 12724 5960 12756
rect 5920 12636 5960 12724
rect 6080 12916 6120 12920
rect 6080 12884 6084 12916
rect 6116 12884 6120 12916
rect 6080 12876 6120 12884
rect 6080 12844 6084 12876
rect 6116 12844 6120 12876
rect 6080 12836 6120 12844
rect 6080 12804 6084 12836
rect 6116 12804 6120 12836
rect 6080 12796 6120 12804
rect 6080 12764 6084 12796
rect 6116 12764 6120 12796
rect 6080 12756 6120 12764
rect 6080 12724 6084 12756
rect 6116 12724 6120 12756
rect 5920 12604 5924 12636
rect 5956 12604 5960 12636
rect 5920 12556 5960 12604
rect 5920 12524 5924 12556
rect 5956 12524 5960 12556
rect 5920 12476 5960 12524
rect 5920 12444 5924 12476
rect 5956 12444 5960 12476
rect 5920 12396 5960 12444
rect 5920 12364 5924 12396
rect 5956 12364 5960 12396
rect 5920 12316 5960 12364
rect 5920 12284 5924 12316
rect 5956 12284 5960 12316
rect 5920 12236 5960 12284
rect 5920 12204 5924 12236
rect 5956 12204 5960 12236
rect 5920 12156 5960 12204
rect 5920 12124 5924 12156
rect 5956 12124 5960 12156
rect 5920 11836 5960 12124
rect 5920 11804 5924 11836
rect 5956 11804 5960 11836
rect 5920 11756 5960 11804
rect 5920 11724 5924 11756
rect 5956 11724 5960 11756
rect 5920 11676 5960 11724
rect 5920 11644 5924 11676
rect 5956 11644 5960 11676
rect 5920 11596 5960 11644
rect 5920 11564 5924 11596
rect 5956 11564 5960 11596
rect 5920 11516 5960 11564
rect 5920 11484 5924 11516
rect 5956 11484 5960 11516
rect 5920 11436 5960 11484
rect 5920 11404 5924 11436
rect 5956 11404 5960 11436
rect 5920 10876 5960 11404
rect 5920 10844 5924 10876
rect 5956 10844 5960 10876
rect 5920 10796 5960 10844
rect 5920 10764 5924 10796
rect 5956 10764 5960 10796
rect 5920 10716 5960 10764
rect 5920 10684 5924 10716
rect 5956 10684 5960 10716
rect 5920 10636 5960 10684
rect 5920 10604 5924 10636
rect 5956 10604 5960 10636
rect 5920 10556 5960 10604
rect 5920 10524 5924 10556
rect 5956 10524 5960 10556
rect 5920 10476 5960 10524
rect 5920 10444 5924 10476
rect 5956 10444 5960 10476
rect 5920 10396 5960 10444
rect 5920 10364 5924 10396
rect 5956 10364 5960 10396
rect 5920 10316 5960 10364
rect 5920 10284 5924 10316
rect 5956 10284 5960 10316
rect 5920 10236 5960 10284
rect 5920 10204 5924 10236
rect 5956 10204 5960 10236
rect 5920 10156 5960 10204
rect 5920 10124 5924 10156
rect 5956 10124 5960 10156
rect 5920 10076 5960 10124
rect 5920 10044 5924 10076
rect 5956 10044 5960 10076
rect 5920 9996 5960 10044
rect 5920 9964 5924 9996
rect 5956 9964 5960 9996
rect 5920 9916 5960 9964
rect 5920 9884 5924 9916
rect 5956 9884 5960 9916
rect 5920 9836 5960 9884
rect 5920 9804 5924 9836
rect 5956 9804 5960 9836
rect 5920 9756 5960 9804
rect 5920 9724 5924 9756
rect 5956 9724 5960 9756
rect 5920 9356 5960 9724
rect 5920 9324 5924 9356
rect 5956 9324 5960 9356
rect 5920 9276 5960 9324
rect 5920 9244 5924 9276
rect 5956 9244 5960 9276
rect 5920 9196 5960 9244
rect 5920 9164 5924 9196
rect 5956 9164 5960 9196
rect 5920 8876 5960 9164
rect 5920 8844 5924 8876
rect 5956 8844 5960 8876
rect 5920 8796 5960 8844
rect 5920 8764 5924 8796
rect 5956 8764 5960 8796
rect 5920 8716 5960 8764
rect 5920 8684 5924 8716
rect 5956 8684 5960 8716
rect 5920 8636 5960 8684
rect 5920 8604 5924 8636
rect 5956 8604 5960 8636
rect 5920 8556 5960 8604
rect 5920 8524 5924 8556
rect 5956 8524 5960 8556
rect 5920 7636 5960 8524
rect 5920 7604 5924 7636
rect 5956 7604 5960 7636
rect 5920 7556 5960 7604
rect 5920 7524 5924 7556
rect 5956 7524 5960 7556
rect 5920 7476 5960 7524
rect 5920 7444 5924 7476
rect 5956 7444 5960 7476
rect 5920 7396 5960 7444
rect 5920 7364 5924 7396
rect 5956 7364 5960 7396
rect 5920 7316 5960 7364
rect 5920 7284 5924 7316
rect 5956 7284 5960 7316
rect 5920 7236 5960 7284
rect 5920 7204 5924 7236
rect 5956 7204 5960 7236
rect 5920 7156 5960 7204
rect 5920 7124 5924 7156
rect 5956 7124 5960 7156
rect 5920 7076 5960 7124
rect 5920 7044 5924 7076
rect 5956 7044 5960 7076
rect 5920 6756 5960 7044
rect 5920 6724 5924 6756
rect 5956 6724 5960 6756
rect 5920 6676 5960 6724
rect 5920 6644 5924 6676
rect 5956 6644 5960 6676
rect 5920 6596 5960 6644
rect 5920 6564 5924 6596
rect 5956 6564 5960 6596
rect 5920 6516 5960 6564
rect 5920 6484 5924 6516
rect 5956 6484 5960 6516
rect 5920 6436 5960 6484
rect 5920 6404 5924 6436
rect 5956 6404 5960 6436
rect 5920 6356 5960 6404
rect 5920 6324 5924 6356
rect 5956 6324 5960 6356
rect 5920 5796 5960 6324
rect 5920 5764 5924 5796
rect 5956 5764 5960 5796
rect 5920 5716 5960 5764
rect 5920 5684 5924 5716
rect 5956 5684 5960 5716
rect 5920 5636 5960 5684
rect 5920 5604 5924 5636
rect 5956 5604 5960 5636
rect 5920 5556 5960 5604
rect 5920 5524 5924 5556
rect 5956 5524 5960 5556
rect 5920 5476 5960 5524
rect 5920 5444 5924 5476
rect 5956 5444 5960 5476
rect 5920 5396 5960 5444
rect 5920 5364 5924 5396
rect 5956 5364 5960 5396
rect 5920 5316 5960 5364
rect 5920 5284 5924 5316
rect 5956 5284 5960 5316
rect 5920 5236 5960 5284
rect 5920 5204 5924 5236
rect 5956 5204 5960 5236
rect 5920 5156 5960 5204
rect 5920 5124 5924 5156
rect 5956 5124 5960 5156
rect 5920 5076 5960 5124
rect 5920 5044 5924 5076
rect 5956 5044 5960 5076
rect 5920 4996 5960 5044
rect 5920 4964 5924 4996
rect 5956 4964 5960 4996
rect 5920 4914 5960 4964
rect 5920 4886 5926 4914
rect 5954 4886 5960 4914
rect 5920 4754 5960 4886
rect 5920 4726 5926 4754
rect 5954 4726 5960 4754
rect 5920 4436 5960 4726
rect 5920 4404 5924 4436
rect 5956 4404 5960 4436
rect 5920 4356 5960 4404
rect 5920 4324 5924 4356
rect 5956 4324 5960 4356
rect 5920 4276 5960 4324
rect 5920 4244 5924 4276
rect 5956 4244 5960 4276
rect 5920 4196 5960 4244
rect 5920 4164 5924 4196
rect 5956 4164 5960 4196
rect 5920 4116 5960 4164
rect 5920 4084 5924 4116
rect 5956 4084 5960 4116
rect 5920 4036 5960 4084
rect 5920 4004 5924 4036
rect 5956 4004 5960 4036
rect 5920 3956 5960 4004
rect 5920 3924 5924 3956
rect 5956 3924 5960 3956
rect 5920 3394 5960 3924
rect 5920 3366 5926 3394
rect 5954 3366 5960 3394
rect 5920 3234 5960 3366
rect 5920 3206 5926 3234
rect 5954 3206 5960 3234
rect 5920 3156 5960 3206
rect 5920 3124 5924 3156
rect 5956 3124 5960 3156
rect 5920 3076 5960 3124
rect 5920 3044 5924 3076
rect 5956 3044 5960 3076
rect 5920 2996 5960 3044
rect 5920 2964 5924 2996
rect 5956 2964 5960 2996
rect 5920 2916 5960 2964
rect 5920 2884 5924 2916
rect 5956 2884 5960 2916
rect 5920 2836 5960 2884
rect 5920 2804 5924 2836
rect 5956 2804 5960 2836
rect 5920 2756 5960 2804
rect 5920 2724 5924 2756
rect 5956 2724 5960 2756
rect 5920 2676 5960 2724
rect 5920 2644 5924 2676
rect 5956 2644 5960 2676
rect 5920 2596 5960 2644
rect 5920 2564 5924 2596
rect 5956 2564 5960 2596
rect 5920 2516 5960 2564
rect 5920 2484 5924 2516
rect 5956 2484 5960 2516
rect 5920 2436 5960 2484
rect 5920 2404 5924 2436
rect 5956 2404 5960 2436
rect 5920 2356 5960 2404
rect 5920 2324 5924 2356
rect 5956 2324 5960 2356
rect 5920 2276 5960 2324
rect 5920 2244 5924 2276
rect 5956 2244 5960 2276
rect 5920 2196 5960 2244
rect 5920 2164 5924 2196
rect 5956 2164 5960 2196
rect 5920 2116 5960 2164
rect 5920 2084 5924 2116
rect 5956 2084 5960 2116
rect 5920 2036 5960 2084
rect 5920 2004 5924 2036
rect 5956 2004 5960 2036
rect 5920 1636 5960 2004
rect 5920 1604 5924 1636
rect 5956 1604 5960 1636
rect 5920 1556 5960 1604
rect 5920 1524 5924 1556
rect 5956 1524 5960 1556
rect 5920 1476 5960 1524
rect 5920 1444 5924 1476
rect 5956 1444 5960 1476
rect 5920 1396 5960 1444
rect 5920 1364 5924 1396
rect 5956 1364 5960 1396
rect 5920 1316 5960 1364
rect 5920 1284 5924 1316
rect 5956 1284 5960 1316
rect 5920 1236 5960 1284
rect 5920 1204 5924 1236
rect 5956 1204 5960 1236
rect 5920 1156 5960 1204
rect 5920 1124 5924 1156
rect 5956 1124 5960 1156
rect 5920 1076 5960 1124
rect 5920 1044 5924 1076
rect 5956 1044 5960 1076
rect 5920 756 5960 1044
rect 5920 724 5924 756
rect 5956 724 5960 756
rect 5920 676 5960 724
rect 5920 644 5924 676
rect 5956 644 5960 676
rect 5920 596 5960 644
rect 5920 564 5924 596
rect 5956 564 5960 596
rect 5920 196 5960 564
rect 5920 164 5924 196
rect 5956 164 5960 196
rect 5920 116 5960 164
rect 5920 84 5924 116
rect 5956 84 5960 116
rect 5920 36 5960 84
rect 5920 4 5924 36
rect 5956 4 5960 36
rect 5920 -40 5960 4
rect 6000 4834 6040 12680
rect 6000 4806 6006 4834
rect 6034 4806 6040 4834
rect 6000 3314 6040 4806
rect 6000 3286 6006 3314
rect 6034 3286 6040 3314
rect 6000 -40 6040 3286
rect 6080 12636 6120 12724
rect 6080 12604 6084 12636
rect 6116 12604 6120 12636
rect 6080 12556 6120 12604
rect 6080 12524 6084 12556
rect 6116 12524 6120 12556
rect 6080 12476 6120 12524
rect 6080 12444 6084 12476
rect 6116 12444 6120 12476
rect 6080 12396 6120 12444
rect 6080 12364 6084 12396
rect 6116 12364 6120 12396
rect 6080 12316 6120 12364
rect 6080 12284 6084 12316
rect 6116 12284 6120 12316
rect 6080 12236 6120 12284
rect 6080 12204 6084 12236
rect 6116 12204 6120 12236
rect 6080 12156 6120 12204
rect 6080 12124 6084 12156
rect 6116 12124 6120 12156
rect 6080 11836 6120 12124
rect 6080 11804 6084 11836
rect 6116 11804 6120 11836
rect 6080 11756 6120 11804
rect 6080 11724 6084 11756
rect 6116 11724 6120 11756
rect 6080 11676 6120 11724
rect 6080 11644 6084 11676
rect 6116 11644 6120 11676
rect 6080 11596 6120 11644
rect 6080 11564 6084 11596
rect 6116 11564 6120 11596
rect 6080 11516 6120 11564
rect 6080 11484 6084 11516
rect 6116 11484 6120 11516
rect 6080 11436 6120 11484
rect 6080 11404 6084 11436
rect 6116 11404 6120 11436
rect 6080 10876 6120 11404
rect 6080 10844 6084 10876
rect 6116 10844 6120 10876
rect 6080 10796 6120 10844
rect 6080 10764 6084 10796
rect 6116 10764 6120 10796
rect 6080 10716 6120 10764
rect 6080 10684 6084 10716
rect 6116 10684 6120 10716
rect 6080 10636 6120 10684
rect 6080 10604 6084 10636
rect 6116 10604 6120 10636
rect 6080 10556 6120 10604
rect 6080 10524 6084 10556
rect 6116 10524 6120 10556
rect 6080 10476 6120 10524
rect 6080 10444 6084 10476
rect 6116 10444 6120 10476
rect 6080 10396 6120 10444
rect 6080 10364 6084 10396
rect 6116 10364 6120 10396
rect 6080 10316 6120 10364
rect 6080 10284 6084 10316
rect 6116 10284 6120 10316
rect 6080 10236 6120 10284
rect 6080 10204 6084 10236
rect 6116 10204 6120 10236
rect 6080 10156 6120 10204
rect 6080 10124 6084 10156
rect 6116 10124 6120 10156
rect 6080 10076 6120 10124
rect 6080 10044 6084 10076
rect 6116 10044 6120 10076
rect 6080 9996 6120 10044
rect 6080 9964 6084 9996
rect 6116 9964 6120 9996
rect 6080 9916 6120 9964
rect 6080 9884 6084 9916
rect 6116 9884 6120 9916
rect 6080 9836 6120 9884
rect 6080 9804 6084 9836
rect 6116 9804 6120 9836
rect 6080 9756 6120 9804
rect 6080 9724 6084 9756
rect 6116 9724 6120 9756
rect 6080 9356 6120 9724
rect 6080 9324 6084 9356
rect 6116 9324 6120 9356
rect 6080 9276 6120 9324
rect 6080 9244 6084 9276
rect 6116 9244 6120 9276
rect 6080 9196 6120 9244
rect 6080 9164 6084 9196
rect 6116 9164 6120 9196
rect 6080 8876 6120 9164
rect 6080 8844 6084 8876
rect 6116 8844 6120 8876
rect 6080 8796 6120 8844
rect 6080 8764 6084 8796
rect 6116 8764 6120 8796
rect 6080 8716 6120 8764
rect 6080 8684 6084 8716
rect 6116 8684 6120 8716
rect 6080 8636 6120 8684
rect 6080 8604 6084 8636
rect 6116 8604 6120 8636
rect 6080 8556 6120 8604
rect 6080 8524 6084 8556
rect 6116 8524 6120 8556
rect 6080 7636 6120 8524
rect 6080 7604 6084 7636
rect 6116 7604 6120 7636
rect 6080 7556 6120 7604
rect 6080 7524 6084 7556
rect 6116 7524 6120 7556
rect 6080 7476 6120 7524
rect 6080 7444 6084 7476
rect 6116 7444 6120 7476
rect 6080 7396 6120 7444
rect 6080 7364 6084 7396
rect 6116 7364 6120 7396
rect 6080 7316 6120 7364
rect 6080 7284 6084 7316
rect 6116 7284 6120 7316
rect 6080 7236 6120 7284
rect 6080 7204 6084 7236
rect 6116 7204 6120 7236
rect 6080 7156 6120 7204
rect 6080 7124 6084 7156
rect 6116 7124 6120 7156
rect 6080 7076 6120 7124
rect 6080 7044 6084 7076
rect 6116 7044 6120 7076
rect 6080 6756 6120 7044
rect 6080 6724 6084 6756
rect 6116 6724 6120 6756
rect 6080 6676 6120 6724
rect 6080 6644 6084 6676
rect 6116 6644 6120 6676
rect 6080 6596 6120 6644
rect 6080 6564 6084 6596
rect 6116 6564 6120 6596
rect 6080 6516 6120 6564
rect 6080 6484 6084 6516
rect 6116 6484 6120 6516
rect 6080 6436 6120 6484
rect 6080 6404 6084 6436
rect 6116 6404 6120 6436
rect 6080 6356 6120 6404
rect 6080 6324 6084 6356
rect 6116 6324 6120 6356
rect 6080 5796 6120 6324
rect 6080 5764 6084 5796
rect 6116 5764 6120 5796
rect 6080 5716 6120 5764
rect 6080 5684 6084 5716
rect 6116 5684 6120 5716
rect 6080 5636 6120 5684
rect 6080 5604 6084 5636
rect 6116 5604 6120 5636
rect 6080 5556 6120 5604
rect 6080 5524 6084 5556
rect 6116 5524 6120 5556
rect 6080 5476 6120 5524
rect 6080 5444 6084 5476
rect 6116 5444 6120 5476
rect 6080 5396 6120 5444
rect 6080 5364 6084 5396
rect 6116 5364 6120 5396
rect 6080 5316 6120 5364
rect 6080 5284 6084 5316
rect 6116 5284 6120 5316
rect 6080 5236 6120 5284
rect 6080 5204 6084 5236
rect 6116 5204 6120 5236
rect 6080 5156 6120 5204
rect 6080 5124 6084 5156
rect 6116 5124 6120 5156
rect 6080 5076 6120 5124
rect 6080 5044 6084 5076
rect 6116 5044 6120 5076
rect 6080 4996 6120 5044
rect 6080 4964 6084 4996
rect 6116 4964 6120 4996
rect 6080 4914 6120 4964
rect 6080 4886 6086 4914
rect 6114 4886 6120 4914
rect 6080 4754 6120 4886
rect 6080 4726 6086 4754
rect 6114 4726 6120 4754
rect 6080 4436 6120 4726
rect 6080 4404 6084 4436
rect 6116 4404 6120 4436
rect 6080 4356 6120 4404
rect 6080 4324 6084 4356
rect 6116 4324 6120 4356
rect 6080 4276 6120 4324
rect 6080 4244 6084 4276
rect 6116 4244 6120 4276
rect 6080 4196 6120 4244
rect 6080 4164 6084 4196
rect 6116 4164 6120 4196
rect 6080 4116 6120 4164
rect 6080 4084 6084 4116
rect 6116 4084 6120 4116
rect 6080 4036 6120 4084
rect 6080 4004 6084 4036
rect 6116 4004 6120 4036
rect 6080 3956 6120 4004
rect 6080 3924 6084 3956
rect 6116 3924 6120 3956
rect 6080 3394 6120 3924
rect 6080 3366 6086 3394
rect 6114 3366 6120 3394
rect 6080 3234 6120 3366
rect 6080 3206 6086 3234
rect 6114 3206 6120 3234
rect 6080 3156 6120 3206
rect 6080 3124 6084 3156
rect 6116 3124 6120 3156
rect 6080 3076 6120 3124
rect 6080 3044 6084 3076
rect 6116 3044 6120 3076
rect 6080 2996 6120 3044
rect 6080 2964 6084 2996
rect 6116 2964 6120 2996
rect 6080 2916 6120 2964
rect 6080 2884 6084 2916
rect 6116 2884 6120 2916
rect 6080 2836 6120 2884
rect 6080 2804 6084 2836
rect 6116 2804 6120 2836
rect 6080 2756 6120 2804
rect 6080 2724 6084 2756
rect 6116 2724 6120 2756
rect 6080 2676 6120 2724
rect 6080 2644 6084 2676
rect 6116 2644 6120 2676
rect 6080 2596 6120 2644
rect 6080 2564 6084 2596
rect 6116 2564 6120 2596
rect 6080 2516 6120 2564
rect 6080 2484 6084 2516
rect 6116 2484 6120 2516
rect 6080 2436 6120 2484
rect 6080 2404 6084 2436
rect 6116 2404 6120 2436
rect 6080 2356 6120 2404
rect 6080 2324 6084 2356
rect 6116 2324 6120 2356
rect 6080 2276 6120 2324
rect 6080 2244 6084 2276
rect 6116 2244 6120 2276
rect 6080 2196 6120 2244
rect 6080 2164 6084 2196
rect 6116 2164 6120 2196
rect 6080 2116 6120 2164
rect 6080 2084 6084 2116
rect 6116 2084 6120 2116
rect 6080 2036 6120 2084
rect 6080 2004 6084 2036
rect 6116 2004 6120 2036
rect 6080 1636 6120 2004
rect 6080 1604 6084 1636
rect 6116 1604 6120 1636
rect 6080 1556 6120 1604
rect 6080 1524 6084 1556
rect 6116 1524 6120 1556
rect 6080 1476 6120 1524
rect 6080 1444 6084 1476
rect 6116 1444 6120 1476
rect 6080 1396 6120 1444
rect 6080 1364 6084 1396
rect 6116 1364 6120 1396
rect 6080 1316 6120 1364
rect 6080 1284 6084 1316
rect 6116 1284 6120 1316
rect 6080 1236 6120 1284
rect 6080 1204 6084 1236
rect 6116 1204 6120 1236
rect 6080 1156 6120 1204
rect 6080 1124 6084 1156
rect 6116 1124 6120 1156
rect 6080 1076 6120 1124
rect 6080 1044 6084 1076
rect 6116 1044 6120 1076
rect 6080 756 6120 1044
rect 6080 724 6084 756
rect 6116 724 6120 756
rect 6080 676 6120 724
rect 6080 644 6084 676
rect 6116 644 6120 676
rect 6080 596 6120 644
rect 6080 564 6084 596
rect 6116 564 6120 596
rect 6080 196 6120 564
rect 6080 164 6084 196
rect 6116 164 6120 196
rect 6080 116 6120 164
rect 6080 84 6084 116
rect 6116 84 6120 116
rect 6080 36 6120 84
rect 6080 4 6084 36
rect 6116 4 6120 36
rect 6080 -40 6120 4
rect 6160 12636 6200 13204
rect 6320 13396 6360 13400
rect 6320 13364 6324 13396
rect 6356 13364 6360 13396
rect 6320 13356 6360 13364
rect 6320 13324 6324 13356
rect 6356 13324 6360 13356
rect 6320 13316 6360 13324
rect 6320 13284 6324 13316
rect 6356 13284 6360 13316
rect 6320 13276 6360 13284
rect 6320 13244 6324 13276
rect 6356 13244 6360 13276
rect 6320 13236 6360 13244
rect 6320 13204 6324 13236
rect 6356 13204 6360 13236
rect 6160 12604 6164 12636
rect 6196 12604 6200 12636
rect 6160 12556 6200 12604
rect 6160 12524 6164 12556
rect 6196 12524 6200 12556
rect 6160 12476 6200 12524
rect 6160 12444 6164 12476
rect 6196 12444 6200 12476
rect 6160 12396 6200 12444
rect 6160 12364 6164 12396
rect 6196 12364 6200 12396
rect 6160 12316 6200 12364
rect 6160 12284 6164 12316
rect 6196 12284 6200 12316
rect 6160 12236 6200 12284
rect 6160 12204 6164 12236
rect 6196 12204 6200 12236
rect 6160 12156 6200 12204
rect 6160 12124 6164 12156
rect 6196 12124 6200 12156
rect 6160 11836 6200 12124
rect 6160 11804 6164 11836
rect 6196 11804 6200 11836
rect 6160 11756 6200 11804
rect 6160 11724 6164 11756
rect 6196 11724 6200 11756
rect 6160 11676 6200 11724
rect 6160 11644 6164 11676
rect 6196 11644 6200 11676
rect 6160 11596 6200 11644
rect 6160 11564 6164 11596
rect 6196 11564 6200 11596
rect 6160 11516 6200 11564
rect 6160 11484 6164 11516
rect 6196 11484 6200 11516
rect 6160 11436 6200 11484
rect 6160 11404 6164 11436
rect 6196 11404 6200 11436
rect 6160 10876 6200 11404
rect 6160 10844 6164 10876
rect 6196 10844 6200 10876
rect 6160 10796 6200 10844
rect 6160 10764 6164 10796
rect 6196 10764 6200 10796
rect 6160 10716 6200 10764
rect 6160 10684 6164 10716
rect 6196 10684 6200 10716
rect 6160 10636 6200 10684
rect 6160 10604 6164 10636
rect 6196 10604 6200 10636
rect 6160 10556 6200 10604
rect 6160 10524 6164 10556
rect 6196 10524 6200 10556
rect 6160 10476 6200 10524
rect 6160 10444 6164 10476
rect 6196 10444 6200 10476
rect 6160 10396 6200 10444
rect 6160 10364 6164 10396
rect 6196 10364 6200 10396
rect 6160 10316 6200 10364
rect 6160 10284 6164 10316
rect 6196 10284 6200 10316
rect 6160 10236 6200 10284
rect 6160 10204 6164 10236
rect 6196 10204 6200 10236
rect 6160 10156 6200 10204
rect 6160 10124 6164 10156
rect 6196 10124 6200 10156
rect 6160 10076 6200 10124
rect 6160 10044 6164 10076
rect 6196 10044 6200 10076
rect 6160 9996 6200 10044
rect 6160 9964 6164 9996
rect 6196 9964 6200 9996
rect 6160 9916 6200 9964
rect 6160 9884 6164 9916
rect 6196 9884 6200 9916
rect 6160 9836 6200 9884
rect 6160 9804 6164 9836
rect 6196 9804 6200 9836
rect 6160 9756 6200 9804
rect 6160 9724 6164 9756
rect 6196 9724 6200 9756
rect 6160 9356 6200 9724
rect 6160 9324 6164 9356
rect 6196 9324 6200 9356
rect 6160 9276 6200 9324
rect 6160 9244 6164 9276
rect 6196 9244 6200 9276
rect 6160 9196 6200 9244
rect 6160 9164 6164 9196
rect 6196 9164 6200 9196
rect 6160 8876 6200 9164
rect 6160 8844 6164 8876
rect 6196 8844 6200 8876
rect 6160 8796 6200 8844
rect 6160 8764 6164 8796
rect 6196 8764 6200 8796
rect 6160 8716 6200 8764
rect 6160 8684 6164 8716
rect 6196 8684 6200 8716
rect 6160 8636 6200 8684
rect 6160 8604 6164 8636
rect 6196 8604 6200 8636
rect 6160 8556 6200 8604
rect 6160 8524 6164 8556
rect 6196 8524 6200 8556
rect 6160 7636 6200 8524
rect 6160 7604 6164 7636
rect 6196 7604 6200 7636
rect 6160 7556 6200 7604
rect 6160 7524 6164 7556
rect 6196 7524 6200 7556
rect 6160 7476 6200 7524
rect 6160 7444 6164 7476
rect 6196 7444 6200 7476
rect 6160 7396 6200 7444
rect 6160 7364 6164 7396
rect 6196 7364 6200 7396
rect 6160 7316 6200 7364
rect 6160 7284 6164 7316
rect 6196 7284 6200 7316
rect 6160 7236 6200 7284
rect 6160 7204 6164 7236
rect 6196 7204 6200 7236
rect 6160 7156 6200 7204
rect 6160 7124 6164 7156
rect 6196 7124 6200 7156
rect 6160 7076 6200 7124
rect 6160 7044 6164 7076
rect 6196 7044 6200 7076
rect 6160 6756 6200 7044
rect 6160 6724 6164 6756
rect 6196 6724 6200 6756
rect 6160 6676 6200 6724
rect 6160 6644 6164 6676
rect 6196 6644 6200 6676
rect 6160 6596 6200 6644
rect 6160 6564 6164 6596
rect 6196 6564 6200 6596
rect 6160 6516 6200 6564
rect 6160 6484 6164 6516
rect 6196 6484 6200 6516
rect 6160 6436 6200 6484
rect 6160 6404 6164 6436
rect 6196 6404 6200 6436
rect 6160 6356 6200 6404
rect 6160 6324 6164 6356
rect 6196 6324 6200 6356
rect 6160 5796 6200 6324
rect 6160 5764 6164 5796
rect 6196 5764 6200 5796
rect 6160 5716 6200 5764
rect 6160 5684 6164 5716
rect 6196 5684 6200 5716
rect 6160 5636 6200 5684
rect 6160 5604 6164 5636
rect 6196 5604 6200 5636
rect 6160 5556 6200 5604
rect 6160 5524 6164 5556
rect 6196 5524 6200 5556
rect 6160 5476 6200 5524
rect 6160 5444 6164 5476
rect 6196 5444 6200 5476
rect 6160 5396 6200 5444
rect 6160 5364 6164 5396
rect 6196 5364 6200 5396
rect 6160 5316 6200 5364
rect 6160 5284 6164 5316
rect 6196 5284 6200 5316
rect 6160 5236 6200 5284
rect 6160 5204 6164 5236
rect 6196 5204 6200 5236
rect 6160 5156 6200 5204
rect 6160 5124 6164 5156
rect 6196 5124 6200 5156
rect 6160 5076 6200 5124
rect 6160 5044 6164 5076
rect 6196 5044 6200 5076
rect 6160 4996 6200 5044
rect 6160 4964 6164 4996
rect 6196 4964 6200 4996
rect 6160 4674 6200 4964
rect 6160 4646 6166 4674
rect 6194 4646 6200 4674
rect 6160 4514 6200 4646
rect 6160 4486 6166 4514
rect 6194 4486 6200 4514
rect 6160 4436 6200 4486
rect 6160 4404 6164 4436
rect 6196 4404 6200 4436
rect 6160 4356 6200 4404
rect 6160 4324 6164 4356
rect 6196 4324 6200 4356
rect 6160 4276 6200 4324
rect 6160 4244 6164 4276
rect 6196 4244 6200 4276
rect 6160 4196 6200 4244
rect 6160 4164 6164 4196
rect 6196 4164 6200 4196
rect 6160 4116 6200 4164
rect 6160 4084 6164 4116
rect 6196 4084 6200 4116
rect 6160 4036 6200 4084
rect 6160 4004 6164 4036
rect 6196 4004 6200 4036
rect 6160 3956 6200 4004
rect 6160 3924 6164 3956
rect 6196 3924 6200 3956
rect 6160 3156 6200 3924
rect 6160 3124 6164 3156
rect 6196 3124 6200 3156
rect 6160 3076 6200 3124
rect 6160 3044 6164 3076
rect 6196 3044 6200 3076
rect 6160 2996 6200 3044
rect 6160 2964 6164 2996
rect 6196 2964 6200 2996
rect 6160 2916 6200 2964
rect 6160 2884 6164 2916
rect 6196 2884 6200 2916
rect 6160 2836 6200 2884
rect 6160 2804 6164 2836
rect 6196 2804 6200 2836
rect 6160 2756 6200 2804
rect 6160 2724 6164 2756
rect 6196 2724 6200 2756
rect 6160 2676 6200 2724
rect 6160 2644 6164 2676
rect 6196 2644 6200 2676
rect 6160 2596 6200 2644
rect 6160 2564 6164 2596
rect 6196 2564 6200 2596
rect 6160 2516 6200 2564
rect 6160 2484 6164 2516
rect 6196 2484 6200 2516
rect 6160 2436 6200 2484
rect 6160 2404 6164 2436
rect 6196 2404 6200 2436
rect 6160 2356 6200 2404
rect 6160 2324 6164 2356
rect 6196 2324 6200 2356
rect 6160 2276 6200 2324
rect 6160 2244 6164 2276
rect 6196 2244 6200 2276
rect 6160 2196 6200 2244
rect 6160 2164 6164 2196
rect 6196 2164 6200 2196
rect 6160 2116 6200 2164
rect 6160 2084 6164 2116
rect 6196 2084 6200 2116
rect 6160 2036 6200 2084
rect 6160 2004 6164 2036
rect 6196 2004 6200 2036
rect 6160 1636 6200 2004
rect 6160 1604 6164 1636
rect 6196 1604 6200 1636
rect 6160 1556 6200 1604
rect 6160 1524 6164 1556
rect 6196 1524 6200 1556
rect 6160 1476 6200 1524
rect 6160 1444 6164 1476
rect 6196 1444 6200 1476
rect 6160 1396 6200 1444
rect 6160 1364 6164 1396
rect 6196 1364 6200 1396
rect 6160 1316 6200 1364
rect 6160 1284 6164 1316
rect 6196 1284 6200 1316
rect 6160 1236 6200 1284
rect 6160 1204 6164 1236
rect 6196 1204 6200 1236
rect 6160 1156 6200 1204
rect 6160 1124 6164 1156
rect 6196 1124 6200 1156
rect 6160 1076 6200 1124
rect 6160 1044 6164 1076
rect 6196 1044 6200 1076
rect 6160 994 6200 1044
rect 6160 966 6166 994
rect 6194 966 6200 994
rect 6160 834 6200 966
rect 6160 806 6166 834
rect 6194 806 6200 834
rect 6160 756 6200 806
rect 6160 724 6164 756
rect 6196 724 6200 756
rect 6160 676 6200 724
rect 6160 644 6164 676
rect 6196 644 6200 676
rect 6160 596 6200 644
rect 6160 564 6164 596
rect 6196 564 6200 596
rect 6160 196 6200 564
rect 6160 164 6164 196
rect 6196 164 6200 196
rect 6160 116 6200 164
rect 6160 84 6164 116
rect 6196 84 6200 116
rect 6160 36 6200 84
rect 6160 4 6164 36
rect 6196 4 6200 36
rect 6160 -40 6200 4
rect 6240 4594 6280 12680
rect 6240 4566 6246 4594
rect 6274 4566 6280 4594
rect 6240 914 6280 4566
rect 6240 886 6246 914
rect 6274 886 6280 914
rect 6240 -40 6280 886
rect 6320 12636 6360 13204
rect 6320 12604 6324 12636
rect 6356 12604 6360 12636
rect 6320 12556 6360 12604
rect 6320 12524 6324 12556
rect 6356 12524 6360 12556
rect 6320 12476 6360 12524
rect 6320 12444 6324 12476
rect 6356 12444 6360 12476
rect 6320 12396 6360 12444
rect 6320 12364 6324 12396
rect 6356 12364 6360 12396
rect 6320 12316 6360 12364
rect 6320 12284 6324 12316
rect 6356 12284 6360 12316
rect 6320 12236 6360 12284
rect 6320 12204 6324 12236
rect 6356 12204 6360 12236
rect 6320 12156 6360 12204
rect 6320 12124 6324 12156
rect 6356 12124 6360 12156
rect 6320 11836 6360 12124
rect 6320 11804 6324 11836
rect 6356 11804 6360 11836
rect 6320 11756 6360 11804
rect 6320 11724 6324 11756
rect 6356 11724 6360 11756
rect 6320 11676 6360 11724
rect 6320 11644 6324 11676
rect 6356 11644 6360 11676
rect 6320 11596 6360 11644
rect 6320 11564 6324 11596
rect 6356 11564 6360 11596
rect 6320 11516 6360 11564
rect 6320 11484 6324 11516
rect 6356 11484 6360 11516
rect 6320 11436 6360 11484
rect 6320 11404 6324 11436
rect 6356 11404 6360 11436
rect 6320 10876 6360 11404
rect 6320 10844 6324 10876
rect 6356 10844 6360 10876
rect 6320 10796 6360 10844
rect 6320 10764 6324 10796
rect 6356 10764 6360 10796
rect 6320 10716 6360 10764
rect 6320 10684 6324 10716
rect 6356 10684 6360 10716
rect 6320 10636 6360 10684
rect 6320 10604 6324 10636
rect 6356 10604 6360 10636
rect 6320 10556 6360 10604
rect 6320 10524 6324 10556
rect 6356 10524 6360 10556
rect 6320 10476 6360 10524
rect 6320 10444 6324 10476
rect 6356 10444 6360 10476
rect 6320 10396 6360 10444
rect 6320 10364 6324 10396
rect 6356 10364 6360 10396
rect 6320 10316 6360 10364
rect 6320 10284 6324 10316
rect 6356 10284 6360 10316
rect 6320 10236 6360 10284
rect 6320 10204 6324 10236
rect 6356 10204 6360 10236
rect 6320 10156 6360 10204
rect 6320 10124 6324 10156
rect 6356 10124 6360 10156
rect 6320 10076 6360 10124
rect 6320 10044 6324 10076
rect 6356 10044 6360 10076
rect 6320 9996 6360 10044
rect 6320 9964 6324 9996
rect 6356 9964 6360 9996
rect 6320 9916 6360 9964
rect 6320 9884 6324 9916
rect 6356 9884 6360 9916
rect 6320 9836 6360 9884
rect 6320 9804 6324 9836
rect 6356 9804 6360 9836
rect 6320 9756 6360 9804
rect 6320 9724 6324 9756
rect 6356 9724 6360 9756
rect 6320 9356 6360 9724
rect 6320 9324 6324 9356
rect 6356 9324 6360 9356
rect 6320 9276 6360 9324
rect 6320 9244 6324 9276
rect 6356 9244 6360 9276
rect 6320 9196 6360 9244
rect 6320 9164 6324 9196
rect 6356 9164 6360 9196
rect 6320 8876 6360 9164
rect 6320 8844 6324 8876
rect 6356 8844 6360 8876
rect 6320 8796 6360 8844
rect 6320 8764 6324 8796
rect 6356 8764 6360 8796
rect 6320 8716 6360 8764
rect 6320 8684 6324 8716
rect 6356 8684 6360 8716
rect 6320 8636 6360 8684
rect 6320 8604 6324 8636
rect 6356 8604 6360 8636
rect 6320 8556 6360 8604
rect 6320 8524 6324 8556
rect 6356 8524 6360 8556
rect 6320 7636 6360 8524
rect 6320 7604 6324 7636
rect 6356 7604 6360 7636
rect 6320 7556 6360 7604
rect 6320 7524 6324 7556
rect 6356 7524 6360 7556
rect 6320 7476 6360 7524
rect 6320 7444 6324 7476
rect 6356 7444 6360 7476
rect 6320 7396 6360 7444
rect 6320 7364 6324 7396
rect 6356 7364 6360 7396
rect 6320 7316 6360 7364
rect 6320 7284 6324 7316
rect 6356 7284 6360 7316
rect 6320 7236 6360 7284
rect 6320 7204 6324 7236
rect 6356 7204 6360 7236
rect 6320 7156 6360 7204
rect 6320 7124 6324 7156
rect 6356 7124 6360 7156
rect 6320 7076 6360 7124
rect 6320 7044 6324 7076
rect 6356 7044 6360 7076
rect 6320 6756 6360 7044
rect 6320 6724 6324 6756
rect 6356 6724 6360 6756
rect 6320 6676 6360 6724
rect 6320 6644 6324 6676
rect 6356 6644 6360 6676
rect 6320 6596 6360 6644
rect 6320 6564 6324 6596
rect 6356 6564 6360 6596
rect 6320 6516 6360 6564
rect 6320 6484 6324 6516
rect 6356 6484 6360 6516
rect 6320 6436 6360 6484
rect 6320 6404 6324 6436
rect 6356 6404 6360 6436
rect 6320 6356 6360 6404
rect 6320 6324 6324 6356
rect 6356 6324 6360 6356
rect 6320 5796 6360 6324
rect 6320 5764 6324 5796
rect 6356 5764 6360 5796
rect 6320 5716 6360 5764
rect 6320 5684 6324 5716
rect 6356 5684 6360 5716
rect 6320 5636 6360 5684
rect 6320 5604 6324 5636
rect 6356 5604 6360 5636
rect 6320 5556 6360 5604
rect 6320 5524 6324 5556
rect 6356 5524 6360 5556
rect 6320 5476 6360 5524
rect 6320 5444 6324 5476
rect 6356 5444 6360 5476
rect 6320 5396 6360 5444
rect 6320 5364 6324 5396
rect 6356 5364 6360 5396
rect 6320 5316 6360 5364
rect 6320 5284 6324 5316
rect 6356 5284 6360 5316
rect 6320 5236 6360 5284
rect 6320 5204 6324 5236
rect 6356 5204 6360 5236
rect 6320 5156 6360 5204
rect 6320 5124 6324 5156
rect 6356 5124 6360 5156
rect 6320 5076 6360 5124
rect 6320 5044 6324 5076
rect 6356 5044 6360 5076
rect 6320 4996 6360 5044
rect 6320 4964 6324 4996
rect 6356 4964 6360 4996
rect 6320 4674 6360 4964
rect 6320 4646 6326 4674
rect 6354 4646 6360 4674
rect 6320 4514 6360 4646
rect 6320 4486 6326 4514
rect 6354 4486 6360 4514
rect 6320 4436 6360 4486
rect 6320 4404 6324 4436
rect 6356 4404 6360 4436
rect 6320 4356 6360 4404
rect 6320 4324 6324 4356
rect 6356 4324 6360 4356
rect 6320 4276 6360 4324
rect 6320 4244 6324 4276
rect 6356 4244 6360 4276
rect 6320 4196 6360 4244
rect 6320 4164 6324 4196
rect 6356 4164 6360 4196
rect 6320 4116 6360 4164
rect 6320 4084 6324 4116
rect 6356 4084 6360 4116
rect 6320 4036 6360 4084
rect 6320 4004 6324 4036
rect 6356 4004 6360 4036
rect 6320 3956 6360 4004
rect 6320 3924 6324 3956
rect 6356 3924 6360 3956
rect 6320 3156 6360 3924
rect 6320 3124 6324 3156
rect 6356 3124 6360 3156
rect 6320 3076 6360 3124
rect 6320 3044 6324 3076
rect 6356 3044 6360 3076
rect 6320 2996 6360 3044
rect 6320 2964 6324 2996
rect 6356 2964 6360 2996
rect 6320 2916 6360 2964
rect 6320 2884 6324 2916
rect 6356 2884 6360 2916
rect 6320 2836 6360 2884
rect 6320 2804 6324 2836
rect 6356 2804 6360 2836
rect 6320 2756 6360 2804
rect 6320 2724 6324 2756
rect 6356 2724 6360 2756
rect 6320 2676 6360 2724
rect 6320 2644 6324 2676
rect 6356 2644 6360 2676
rect 6320 2596 6360 2644
rect 6320 2564 6324 2596
rect 6356 2564 6360 2596
rect 6320 2516 6360 2564
rect 6320 2484 6324 2516
rect 6356 2484 6360 2516
rect 6320 2436 6360 2484
rect 6320 2404 6324 2436
rect 6356 2404 6360 2436
rect 6320 2356 6360 2404
rect 6320 2324 6324 2356
rect 6356 2324 6360 2356
rect 6320 2276 6360 2324
rect 6320 2244 6324 2276
rect 6356 2244 6360 2276
rect 6320 2196 6360 2244
rect 6320 2164 6324 2196
rect 6356 2164 6360 2196
rect 6320 2116 6360 2164
rect 6320 2084 6324 2116
rect 6356 2084 6360 2116
rect 6320 2036 6360 2084
rect 6320 2004 6324 2036
rect 6356 2004 6360 2036
rect 6320 1636 6360 2004
rect 6320 1604 6324 1636
rect 6356 1604 6360 1636
rect 6320 1556 6360 1604
rect 6320 1524 6324 1556
rect 6356 1524 6360 1556
rect 6320 1476 6360 1524
rect 6320 1444 6324 1476
rect 6356 1444 6360 1476
rect 6320 1396 6360 1444
rect 6320 1364 6324 1396
rect 6356 1364 6360 1396
rect 6320 1316 6360 1364
rect 6320 1284 6324 1316
rect 6356 1284 6360 1316
rect 6320 1236 6360 1284
rect 6320 1204 6324 1236
rect 6356 1204 6360 1236
rect 6320 1156 6360 1204
rect 6320 1124 6324 1156
rect 6356 1124 6360 1156
rect 6320 1076 6360 1124
rect 6320 1044 6324 1076
rect 6356 1044 6360 1076
rect 6320 994 6360 1044
rect 6320 966 6326 994
rect 6354 966 6360 994
rect 6320 834 6360 966
rect 6320 806 6326 834
rect 6354 806 6360 834
rect 6320 756 6360 806
rect 6320 724 6324 756
rect 6356 724 6360 756
rect 6320 676 6360 724
rect 6320 644 6324 676
rect 6356 644 6360 676
rect 6320 596 6360 644
rect 6320 564 6324 596
rect 6356 564 6360 596
rect 6320 196 6360 564
rect 6320 164 6324 196
rect 6356 164 6360 196
rect 6320 116 6360 164
rect 6320 84 6324 116
rect 6356 84 6360 116
rect 6320 36 6360 84
rect 6320 4 6324 36
rect 6356 4 6360 36
rect 6320 -40 6360 4
<< via3 >>
rect 4 16884 36 16916
rect 4 15444 36 15476
rect 4 14004 36 14036
rect 84 16804 116 16836
rect 84 15524 116 15556
rect 84 13924 116 13956
rect 84 13764 116 13796
rect 164 16724 196 16756
rect 164 13844 196 13876
rect 244 16804 276 16836
rect 244 15524 276 15556
rect 244 13924 276 13956
rect 244 13764 276 13796
rect 324 16884 356 16916
rect 10244 16884 10276 16916
rect 404 16804 436 16836
rect 10164 16804 10196 16836
rect 484 16724 516 16756
rect 1524 16724 1556 16756
rect 1604 16724 1636 16756
rect 2644 16724 2676 16756
rect 2724 16724 2756 16756
rect 3764 16724 3796 16756
rect 3844 16724 3876 16756
rect 4884 16724 4916 16756
rect 5684 16724 5716 16756
rect 6724 16724 6756 16756
rect 6804 16724 6836 16756
rect 7844 16724 7876 16756
rect 7924 16724 7956 16756
rect 8964 16724 8996 16756
rect 9044 16724 9076 16756
rect 10084 16724 10116 16756
rect 404 15524 436 15556
rect 10164 15524 10196 15556
rect 324 15444 356 15476
rect 10244 15444 10276 15476
rect 404 15364 436 15396
rect 4964 15364 4996 15396
rect 484 15284 516 15316
rect 1524 15284 1556 15316
rect 1604 15284 1636 15316
rect 2644 15284 2676 15316
rect 2724 15284 2756 15316
rect 3764 15284 3796 15316
rect 3844 15284 3876 15316
rect 4884 15284 4916 15316
rect 404 14084 436 14116
rect 4964 14084 4996 14116
rect 324 14004 356 14036
rect 4 13684 36 13716
rect 5044 14004 5076 14036
rect 324 13684 356 13716
rect 4484 13924 4516 13956
rect 4484 13764 4516 13796
rect 4244 13604 4276 13636
rect 4244 13564 4276 13596
rect 4244 13524 4276 13556
rect 4244 13484 4276 13516
rect 4244 13444 4276 13476
rect 4404 13604 4436 13636
rect 4404 13564 4436 13596
rect 4404 13524 4436 13556
rect 4404 13484 4436 13516
rect 4404 13444 4436 13476
rect 4244 12634 4276 12636
rect 4244 12606 4246 12634
rect 4246 12606 4274 12634
rect 4274 12606 4276 12634
rect 4244 12604 4276 12606
rect 4244 12554 4276 12556
rect 4244 12526 4246 12554
rect 4246 12526 4274 12554
rect 4274 12526 4276 12554
rect 4244 12524 4276 12526
rect 4244 12474 4276 12476
rect 4244 12446 4246 12474
rect 4246 12446 4274 12474
rect 4274 12446 4276 12474
rect 4244 12444 4276 12446
rect 4244 12394 4276 12396
rect 4244 12366 4246 12394
rect 4246 12366 4274 12394
rect 4274 12366 4276 12394
rect 4244 12364 4276 12366
rect 4244 12314 4276 12316
rect 4244 12286 4246 12314
rect 4246 12286 4274 12314
rect 4274 12286 4276 12314
rect 4244 12284 4276 12286
rect 4244 12234 4276 12236
rect 4244 12206 4246 12234
rect 4246 12206 4274 12234
rect 4274 12206 4276 12234
rect 4244 12204 4276 12206
rect 4244 12154 4276 12156
rect 4244 12126 4246 12154
rect 4246 12126 4274 12154
rect 4274 12126 4276 12154
rect 4244 12124 4276 12126
rect 4244 11834 4276 11836
rect 4244 11806 4246 11834
rect 4246 11806 4274 11834
rect 4274 11806 4276 11834
rect 4244 11804 4276 11806
rect 4244 11754 4276 11756
rect 4244 11726 4246 11754
rect 4246 11726 4274 11754
rect 4274 11726 4276 11754
rect 4244 11724 4276 11726
rect 4244 11674 4276 11676
rect 4244 11646 4246 11674
rect 4246 11646 4274 11674
rect 4274 11646 4276 11674
rect 4244 11644 4276 11646
rect 4244 11594 4276 11596
rect 4244 11566 4246 11594
rect 4246 11566 4274 11594
rect 4274 11566 4276 11594
rect 4244 11564 4276 11566
rect 4244 11514 4276 11516
rect 4244 11486 4246 11514
rect 4246 11486 4274 11514
rect 4274 11486 4276 11514
rect 4244 11484 4276 11486
rect 4244 11434 4276 11436
rect 4244 11406 4246 11434
rect 4246 11406 4274 11434
rect 4274 11406 4276 11434
rect 4244 11404 4276 11406
rect 4244 10874 4276 10876
rect 4244 10846 4246 10874
rect 4246 10846 4274 10874
rect 4274 10846 4276 10874
rect 4244 10844 4276 10846
rect 4244 10794 4276 10796
rect 4244 10766 4246 10794
rect 4246 10766 4274 10794
rect 4274 10766 4276 10794
rect 4244 10764 4276 10766
rect 4244 10714 4276 10716
rect 4244 10686 4246 10714
rect 4246 10686 4274 10714
rect 4274 10686 4276 10714
rect 4244 10684 4276 10686
rect 4244 10634 4276 10636
rect 4244 10606 4246 10634
rect 4246 10606 4274 10634
rect 4274 10606 4276 10634
rect 4244 10604 4276 10606
rect 4244 10554 4276 10556
rect 4244 10526 4246 10554
rect 4246 10526 4274 10554
rect 4274 10526 4276 10554
rect 4244 10524 4276 10526
rect 4244 10474 4276 10476
rect 4244 10446 4246 10474
rect 4246 10446 4274 10474
rect 4274 10446 4276 10474
rect 4244 10444 4276 10446
rect 4244 10394 4276 10396
rect 4244 10366 4246 10394
rect 4246 10366 4274 10394
rect 4274 10366 4276 10394
rect 4244 10364 4276 10366
rect 4244 10314 4276 10316
rect 4244 10286 4246 10314
rect 4246 10286 4274 10314
rect 4274 10286 4276 10314
rect 4244 10284 4276 10286
rect 4244 10234 4276 10236
rect 4244 10206 4246 10234
rect 4246 10206 4274 10234
rect 4274 10206 4276 10234
rect 4244 10204 4276 10206
rect 4244 10154 4276 10156
rect 4244 10126 4246 10154
rect 4246 10126 4274 10154
rect 4274 10126 4276 10154
rect 4244 10124 4276 10126
rect 4244 10074 4276 10076
rect 4244 10046 4246 10074
rect 4246 10046 4274 10074
rect 4274 10046 4276 10074
rect 4244 10044 4276 10046
rect 4244 9994 4276 9996
rect 4244 9966 4246 9994
rect 4246 9966 4274 9994
rect 4274 9966 4276 9994
rect 4244 9964 4276 9966
rect 4244 9914 4276 9916
rect 4244 9886 4246 9914
rect 4246 9886 4274 9914
rect 4274 9886 4276 9914
rect 4244 9884 4276 9886
rect 4244 9834 4276 9836
rect 4244 9806 4246 9834
rect 4246 9806 4274 9834
rect 4274 9806 4276 9834
rect 4244 9804 4276 9806
rect 4244 9754 4276 9756
rect 4244 9726 4246 9754
rect 4246 9726 4274 9754
rect 4274 9726 4276 9754
rect 4244 9724 4276 9726
rect 4244 9354 4276 9356
rect 4244 9326 4246 9354
rect 4246 9326 4274 9354
rect 4274 9326 4276 9354
rect 4244 9324 4276 9326
rect 4244 9274 4276 9276
rect 4244 9246 4246 9274
rect 4246 9246 4274 9274
rect 4274 9246 4276 9274
rect 4244 9244 4276 9246
rect 4244 9194 4276 9196
rect 4244 9166 4246 9194
rect 4246 9166 4274 9194
rect 4274 9166 4276 9194
rect 4244 9164 4276 9166
rect 4244 8874 4276 8876
rect 4244 8846 4246 8874
rect 4246 8846 4274 8874
rect 4274 8846 4276 8874
rect 4244 8844 4276 8846
rect 4244 8794 4276 8796
rect 4244 8766 4246 8794
rect 4246 8766 4274 8794
rect 4274 8766 4276 8794
rect 4244 8764 4276 8766
rect 4244 8714 4276 8716
rect 4244 8686 4246 8714
rect 4246 8686 4274 8714
rect 4274 8686 4276 8714
rect 4244 8684 4276 8686
rect 4244 8634 4276 8636
rect 4244 8606 4246 8634
rect 4246 8606 4274 8634
rect 4274 8606 4276 8634
rect 4244 8604 4276 8606
rect 4244 8554 4276 8556
rect 4244 8526 4246 8554
rect 4246 8526 4274 8554
rect 4274 8526 4276 8554
rect 4244 8524 4276 8526
rect 4244 7634 4276 7636
rect 4244 7606 4246 7634
rect 4246 7606 4274 7634
rect 4274 7606 4276 7634
rect 4244 7604 4276 7606
rect 4244 7554 4276 7556
rect 4244 7526 4246 7554
rect 4246 7526 4274 7554
rect 4274 7526 4276 7554
rect 4244 7524 4276 7526
rect 4244 7474 4276 7476
rect 4244 7446 4246 7474
rect 4246 7446 4274 7474
rect 4274 7446 4276 7474
rect 4244 7444 4276 7446
rect 4244 7394 4276 7396
rect 4244 7366 4246 7394
rect 4246 7366 4274 7394
rect 4274 7366 4276 7394
rect 4244 7364 4276 7366
rect 4244 7314 4276 7316
rect 4244 7286 4246 7314
rect 4246 7286 4274 7314
rect 4274 7286 4276 7314
rect 4244 7284 4276 7286
rect 4244 7234 4276 7236
rect 4244 7206 4246 7234
rect 4246 7206 4274 7234
rect 4274 7206 4276 7234
rect 4244 7204 4276 7206
rect 4244 7154 4276 7156
rect 4244 7126 4246 7154
rect 4246 7126 4274 7154
rect 4274 7126 4276 7154
rect 4244 7124 4276 7126
rect 4244 7074 4276 7076
rect 4244 7046 4246 7074
rect 4246 7046 4274 7074
rect 4274 7046 4276 7074
rect 4244 7044 4276 7046
rect 4244 6754 4276 6756
rect 4244 6726 4246 6754
rect 4246 6726 4274 6754
rect 4274 6726 4276 6754
rect 4244 6724 4276 6726
rect 4244 6674 4276 6676
rect 4244 6646 4246 6674
rect 4246 6646 4274 6674
rect 4274 6646 4276 6674
rect 4244 6644 4276 6646
rect 4244 6594 4276 6596
rect 4244 6566 4246 6594
rect 4246 6566 4274 6594
rect 4274 6566 4276 6594
rect 4244 6564 4276 6566
rect 4244 6514 4276 6516
rect 4244 6486 4246 6514
rect 4246 6486 4274 6514
rect 4274 6486 4276 6514
rect 4244 6484 4276 6486
rect 4244 6434 4276 6436
rect 4244 6406 4246 6434
rect 4246 6406 4274 6434
rect 4274 6406 4276 6434
rect 4244 6404 4276 6406
rect 4244 6354 4276 6356
rect 4244 6326 4246 6354
rect 4246 6326 4274 6354
rect 4274 6326 4276 6354
rect 4244 6324 4276 6326
rect 4244 5794 4276 5796
rect 4244 5766 4246 5794
rect 4246 5766 4274 5794
rect 4274 5766 4276 5794
rect 4244 5764 4276 5766
rect 4244 5714 4276 5716
rect 4244 5686 4246 5714
rect 4246 5686 4274 5714
rect 4274 5686 4276 5714
rect 4244 5684 4276 5686
rect 4244 5634 4276 5636
rect 4244 5606 4246 5634
rect 4246 5606 4274 5634
rect 4274 5606 4276 5634
rect 4244 5604 4276 5606
rect 4244 5554 4276 5556
rect 4244 5526 4246 5554
rect 4246 5526 4274 5554
rect 4274 5526 4276 5554
rect 4244 5524 4276 5526
rect 4244 5474 4276 5476
rect 4244 5446 4246 5474
rect 4246 5446 4274 5474
rect 4274 5446 4276 5474
rect 4244 5444 4276 5446
rect 4244 5394 4276 5396
rect 4244 5366 4246 5394
rect 4246 5366 4274 5394
rect 4274 5366 4276 5394
rect 4244 5364 4276 5366
rect 4244 5314 4276 5316
rect 4244 5286 4246 5314
rect 4246 5286 4274 5314
rect 4274 5286 4276 5314
rect 4244 5284 4276 5286
rect 4244 5234 4276 5236
rect 4244 5206 4246 5234
rect 4246 5206 4274 5234
rect 4274 5206 4276 5234
rect 4244 5204 4276 5206
rect 4244 5154 4276 5156
rect 4244 5126 4246 5154
rect 4246 5126 4274 5154
rect 4274 5126 4276 5154
rect 4244 5124 4276 5126
rect 4244 5074 4276 5076
rect 4244 5046 4246 5074
rect 4246 5046 4274 5074
rect 4274 5046 4276 5074
rect 4244 5044 4276 5046
rect 4244 4994 4276 4996
rect 4244 4966 4246 4994
rect 4246 4966 4274 4994
rect 4274 4966 4276 4994
rect 4244 4964 4276 4966
rect 4244 4434 4276 4436
rect 4244 4406 4246 4434
rect 4246 4406 4274 4434
rect 4274 4406 4276 4434
rect 4244 4404 4276 4406
rect 4244 4354 4276 4356
rect 4244 4326 4246 4354
rect 4246 4326 4274 4354
rect 4274 4326 4276 4354
rect 4244 4324 4276 4326
rect 4244 4274 4276 4276
rect 4244 4246 4246 4274
rect 4246 4246 4274 4274
rect 4274 4246 4276 4274
rect 4244 4244 4276 4246
rect 4244 4194 4276 4196
rect 4244 4166 4246 4194
rect 4246 4166 4274 4194
rect 4274 4166 4276 4194
rect 4244 4164 4276 4166
rect 4244 4114 4276 4116
rect 4244 4086 4246 4114
rect 4246 4086 4274 4114
rect 4274 4086 4276 4114
rect 4244 4084 4276 4086
rect 4244 4034 4276 4036
rect 4244 4006 4246 4034
rect 4246 4006 4274 4034
rect 4274 4006 4276 4034
rect 4244 4004 4276 4006
rect 4244 3954 4276 3956
rect 4244 3926 4246 3954
rect 4246 3926 4274 3954
rect 4274 3926 4276 3954
rect 4244 3924 4276 3926
rect 4244 3154 4276 3156
rect 4244 3126 4246 3154
rect 4246 3126 4274 3154
rect 4274 3126 4276 3154
rect 4244 3124 4276 3126
rect 4244 3074 4276 3076
rect 4244 3046 4246 3074
rect 4246 3046 4274 3074
rect 4274 3046 4276 3074
rect 4244 3044 4276 3046
rect 4244 2994 4276 2996
rect 4244 2966 4246 2994
rect 4246 2966 4274 2994
rect 4274 2966 4276 2994
rect 4244 2964 4276 2966
rect 4244 2914 4276 2916
rect 4244 2886 4246 2914
rect 4246 2886 4274 2914
rect 4274 2886 4276 2914
rect 4244 2884 4276 2886
rect 4244 2834 4276 2836
rect 4244 2806 4246 2834
rect 4246 2806 4274 2834
rect 4274 2806 4276 2834
rect 4244 2804 4276 2806
rect 4244 2754 4276 2756
rect 4244 2726 4246 2754
rect 4246 2726 4274 2754
rect 4274 2726 4276 2754
rect 4244 2724 4276 2726
rect 4244 2674 4276 2676
rect 4244 2646 4246 2674
rect 4246 2646 4274 2674
rect 4274 2646 4276 2674
rect 4244 2644 4276 2646
rect 4244 2594 4276 2596
rect 4244 2566 4246 2594
rect 4246 2566 4274 2594
rect 4274 2566 4276 2594
rect 4244 2564 4276 2566
rect 4244 2514 4276 2516
rect 4244 2486 4246 2514
rect 4246 2486 4274 2514
rect 4274 2486 4276 2514
rect 4244 2484 4276 2486
rect 4244 2434 4276 2436
rect 4244 2406 4246 2434
rect 4246 2406 4274 2434
rect 4274 2406 4276 2434
rect 4244 2404 4276 2406
rect 4244 2354 4276 2356
rect 4244 2326 4246 2354
rect 4246 2326 4274 2354
rect 4274 2326 4276 2354
rect 4244 2324 4276 2326
rect 4244 2274 4276 2276
rect 4244 2246 4246 2274
rect 4246 2246 4274 2274
rect 4274 2246 4276 2274
rect 4244 2244 4276 2246
rect 4244 2194 4276 2196
rect 4244 2166 4246 2194
rect 4246 2166 4274 2194
rect 4274 2166 4276 2194
rect 4244 2164 4276 2166
rect 4244 2114 4276 2116
rect 4244 2086 4246 2114
rect 4246 2086 4274 2114
rect 4274 2086 4276 2114
rect 4244 2084 4276 2086
rect 4244 2034 4276 2036
rect 4244 2006 4246 2034
rect 4246 2006 4274 2034
rect 4274 2006 4276 2034
rect 4244 2004 4276 2006
rect 4244 1634 4276 1636
rect 4244 1606 4246 1634
rect 4246 1606 4274 1634
rect 4274 1606 4276 1634
rect 4244 1604 4276 1606
rect 4244 1554 4276 1556
rect 4244 1526 4246 1554
rect 4246 1526 4274 1554
rect 4274 1526 4276 1554
rect 4244 1524 4276 1526
rect 4244 1474 4276 1476
rect 4244 1446 4246 1474
rect 4246 1446 4274 1474
rect 4274 1446 4276 1474
rect 4244 1444 4276 1446
rect 4244 1394 4276 1396
rect 4244 1366 4246 1394
rect 4246 1366 4274 1394
rect 4274 1366 4276 1394
rect 4244 1364 4276 1366
rect 4244 1314 4276 1316
rect 4244 1286 4246 1314
rect 4246 1286 4274 1314
rect 4274 1286 4276 1314
rect 4244 1284 4276 1286
rect 4244 1234 4276 1236
rect 4244 1206 4246 1234
rect 4246 1206 4274 1234
rect 4274 1206 4276 1234
rect 4244 1204 4276 1206
rect 4244 1154 4276 1156
rect 4244 1126 4246 1154
rect 4246 1126 4274 1154
rect 4274 1126 4276 1154
rect 4244 1124 4276 1126
rect 4244 1074 4276 1076
rect 4244 1046 4246 1074
rect 4246 1046 4274 1074
rect 4274 1046 4276 1074
rect 4244 1044 4276 1046
rect 4244 754 4276 756
rect 4244 726 4246 754
rect 4246 726 4274 754
rect 4274 726 4276 754
rect 4244 724 4276 726
rect 4244 674 4276 676
rect 4244 646 4246 674
rect 4246 646 4274 674
rect 4274 646 4276 674
rect 4244 644 4276 646
rect 4244 594 4276 596
rect 4244 566 4246 594
rect 4246 566 4274 594
rect 4274 566 4276 594
rect 4244 564 4276 566
rect 4244 194 4276 196
rect 4244 166 4246 194
rect 4246 166 4274 194
rect 4274 166 4276 194
rect 4244 164 4276 166
rect 4244 114 4276 116
rect 4244 86 4246 114
rect 4246 86 4274 114
rect 4274 86 4276 114
rect 4244 84 4276 86
rect 4244 34 4276 36
rect 4244 6 4246 34
rect 4246 6 4274 34
rect 4274 6 4276 34
rect 4244 4 4276 6
rect 4404 12634 4436 12636
rect 4404 12606 4406 12634
rect 4406 12606 4434 12634
rect 4434 12606 4436 12634
rect 4404 12604 4436 12606
rect 4404 12554 4436 12556
rect 4404 12526 4406 12554
rect 4406 12526 4434 12554
rect 4434 12526 4436 12554
rect 4404 12524 4436 12526
rect 4404 12474 4436 12476
rect 4404 12446 4406 12474
rect 4406 12446 4434 12474
rect 4434 12446 4436 12474
rect 4404 12444 4436 12446
rect 4404 12394 4436 12396
rect 4404 12366 4406 12394
rect 4406 12366 4434 12394
rect 4434 12366 4436 12394
rect 4404 12364 4436 12366
rect 4404 12314 4436 12316
rect 4404 12286 4406 12314
rect 4406 12286 4434 12314
rect 4434 12286 4436 12314
rect 4404 12284 4436 12286
rect 4404 12234 4436 12236
rect 4404 12206 4406 12234
rect 4406 12206 4434 12234
rect 4434 12206 4436 12234
rect 4404 12204 4436 12206
rect 4404 12154 4436 12156
rect 4404 12126 4406 12154
rect 4406 12126 4434 12154
rect 4434 12126 4436 12154
rect 4404 12124 4436 12126
rect 4404 11834 4436 11836
rect 4404 11806 4406 11834
rect 4406 11806 4434 11834
rect 4434 11806 4436 11834
rect 4404 11804 4436 11806
rect 4404 11754 4436 11756
rect 4404 11726 4406 11754
rect 4406 11726 4434 11754
rect 4434 11726 4436 11754
rect 4404 11724 4436 11726
rect 4404 11674 4436 11676
rect 4404 11646 4406 11674
rect 4406 11646 4434 11674
rect 4434 11646 4436 11674
rect 4404 11644 4436 11646
rect 4404 11594 4436 11596
rect 4404 11566 4406 11594
rect 4406 11566 4434 11594
rect 4434 11566 4436 11594
rect 4404 11564 4436 11566
rect 4404 11514 4436 11516
rect 4404 11486 4406 11514
rect 4406 11486 4434 11514
rect 4434 11486 4436 11514
rect 4404 11484 4436 11486
rect 4404 11434 4436 11436
rect 4404 11406 4406 11434
rect 4406 11406 4434 11434
rect 4434 11406 4436 11434
rect 4404 11404 4436 11406
rect 4404 10874 4436 10876
rect 4404 10846 4406 10874
rect 4406 10846 4434 10874
rect 4434 10846 4436 10874
rect 4404 10844 4436 10846
rect 4404 10794 4436 10796
rect 4404 10766 4406 10794
rect 4406 10766 4434 10794
rect 4434 10766 4436 10794
rect 4404 10764 4436 10766
rect 4404 10714 4436 10716
rect 4404 10686 4406 10714
rect 4406 10686 4434 10714
rect 4434 10686 4436 10714
rect 4404 10684 4436 10686
rect 4404 10634 4436 10636
rect 4404 10606 4406 10634
rect 4406 10606 4434 10634
rect 4434 10606 4436 10634
rect 4404 10604 4436 10606
rect 4404 10554 4436 10556
rect 4404 10526 4406 10554
rect 4406 10526 4434 10554
rect 4434 10526 4436 10554
rect 4404 10524 4436 10526
rect 4404 10474 4436 10476
rect 4404 10446 4406 10474
rect 4406 10446 4434 10474
rect 4434 10446 4436 10474
rect 4404 10444 4436 10446
rect 4404 10394 4436 10396
rect 4404 10366 4406 10394
rect 4406 10366 4434 10394
rect 4434 10366 4436 10394
rect 4404 10364 4436 10366
rect 4404 10314 4436 10316
rect 4404 10286 4406 10314
rect 4406 10286 4434 10314
rect 4434 10286 4436 10314
rect 4404 10284 4436 10286
rect 4404 10234 4436 10236
rect 4404 10206 4406 10234
rect 4406 10206 4434 10234
rect 4434 10206 4436 10234
rect 4404 10204 4436 10206
rect 4404 10154 4436 10156
rect 4404 10126 4406 10154
rect 4406 10126 4434 10154
rect 4434 10126 4436 10154
rect 4404 10124 4436 10126
rect 4404 10074 4436 10076
rect 4404 10046 4406 10074
rect 4406 10046 4434 10074
rect 4434 10046 4436 10074
rect 4404 10044 4436 10046
rect 4404 9994 4436 9996
rect 4404 9966 4406 9994
rect 4406 9966 4434 9994
rect 4434 9966 4436 9994
rect 4404 9964 4436 9966
rect 4404 9914 4436 9916
rect 4404 9886 4406 9914
rect 4406 9886 4434 9914
rect 4434 9886 4436 9914
rect 4404 9884 4436 9886
rect 4404 9834 4436 9836
rect 4404 9806 4406 9834
rect 4406 9806 4434 9834
rect 4434 9806 4436 9834
rect 4404 9804 4436 9806
rect 4404 9754 4436 9756
rect 4404 9726 4406 9754
rect 4406 9726 4434 9754
rect 4434 9726 4436 9754
rect 4404 9724 4436 9726
rect 4404 9354 4436 9356
rect 4404 9326 4406 9354
rect 4406 9326 4434 9354
rect 4434 9326 4436 9354
rect 4404 9324 4436 9326
rect 4404 9274 4436 9276
rect 4404 9246 4406 9274
rect 4406 9246 4434 9274
rect 4434 9246 4436 9274
rect 4404 9244 4436 9246
rect 4404 9194 4436 9196
rect 4404 9166 4406 9194
rect 4406 9166 4434 9194
rect 4434 9166 4436 9194
rect 4404 9164 4436 9166
rect 4404 8874 4436 8876
rect 4404 8846 4406 8874
rect 4406 8846 4434 8874
rect 4434 8846 4436 8874
rect 4404 8844 4436 8846
rect 4404 8794 4436 8796
rect 4404 8766 4406 8794
rect 4406 8766 4434 8794
rect 4434 8766 4436 8794
rect 4404 8764 4436 8766
rect 4404 8714 4436 8716
rect 4404 8686 4406 8714
rect 4406 8686 4434 8714
rect 4434 8686 4436 8714
rect 4404 8684 4436 8686
rect 4404 8634 4436 8636
rect 4404 8606 4406 8634
rect 4406 8606 4434 8634
rect 4434 8606 4436 8634
rect 4404 8604 4436 8606
rect 4404 8554 4436 8556
rect 4404 8526 4406 8554
rect 4406 8526 4434 8554
rect 4434 8526 4436 8554
rect 4404 8524 4436 8526
rect 4404 7634 4436 7636
rect 4404 7606 4406 7634
rect 4406 7606 4434 7634
rect 4434 7606 4436 7634
rect 4404 7604 4436 7606
rect 4404 7554 4436 7556
rect 4404 7526 4406 7554
rect 4406 7526 4434 7554
rect 4434 7526 4436 7554
rect 4404 7524 4436 7526
rect 4404 7474 4436 7476
rect 4404 7446 4406 7474
rect 4406 7446 4434 7474
rect 4434 7446 4436 7474
rect 4404 7444 4436 7446
rect 4404 7394 4436 7396
rect 4404 7366 4406 7394
rect 4406 7366 4434 7394
rect 4434 7366 4436 7394
rect 4404 7364 4436 7366
rect 4404 7314 4436 7316
rect 4404 7286 4406 7314
rect 4406 7286 4434 7314
rect 4434 7286 4436 7314
rect 4404 7284 4436 7286
rect 4404 7234 4436 7236
rect 4404 7206 4406 7234
rect 4406 7206 4434 7234
rect 4434 7206 4436 7234
rect 4404 7204 4436 7206
rect 4404 7154 4436 7156
rect 4404 7126 4406 7154
rect 4406 7126 4434 7154
rect 4434 7126 4436 7154
rect 4404 7124 4436 7126
rect 4404 7074 4436 7076
rect 4404 7046 4406 7074
rect 4406 7046 4434 7074
rect 4434 7046 4436 7074
rect 4404 7044 4436 7046
rect 4404 6754 4436 6756
rect 4404 6726 4406 6754
rect 4406 6726 4434 6754
rect 4434 6726 4436 6754
rect 4404 6724 4436 6726
rect 4404 6674 4436 6676
rect 4404 6646 4406 6674
rect 4406 6646 4434 6674
rect 4434 6646 4436 6674
rect 4404 6644 4436 6646
rect 4404 6594 4436 6596
rect 4404 6566 4406 6594
rect 4406 6566 4434 6594
rect 4434 6566 4436 6594
rect 4404 6564 4436 6566
rect 4404 6514 4436 6516
rect 4404 6486 4406 6514
rect 4406 6486 4434 6514
rect 4434 6486 4436 6514
rect 4404 6484 4436 6486
rect 4404 6434 4436 6436
rect 4404 6406 4406 6434
rect 4406 6406 4434 6434
rect 4434 6406 4436 6434
rect 4404 6404 4436 6406
rect 4404 6354 4436 6356
rect 4404 6326 4406 6354
rect 4406 6326 4434 6354
rect 4434 6326 4436 6354
rect 4404 6324 4436 6326
rect 4404 5794 4436 5796
rect 4404 5766 4406 5794
rect 4406 5766 4434 5794
rect 4434 5766 4436 5794
rect 4404 5764 4436 5766
rect 4404 5714 4436 5716
rect 4404 5686 4406 5714
rect 4406 5686 4434 5714
rect 4434 5686 4436 5714
rect 4404 5684 4436 5686
rect 4404 5634 4436 5636
rect 4404 5606 4406 5634
rect 4406 5606 4434 5634
rect 4434 5606 4436 5634
rect 4404 5604 4436 5606
rect 4404 5554 4436 5556
rect 4404 5526 4406 5554
rect 4406 5526 4434 5554
rect 4434 5526 4436 5554
rect 4404 5524 4436 5526
rect 4404 5474 4436 5476
rect 4404 5446 4406 5474
rect 4406 5446 4434 5474
rect 4434 5446 4436 5474
rect 4404 5444 4436 5446
rect 4404 5394 4436 5396
rect 4404 5366 4406 5394
rect 4406 5366 4434 5394
rect 4434 5366 4436 5394
rect 4404 5364 4436 5366
rect 4404 5314 4436 5316
rect 4404 5286 4406 5314
rect 4406 5286 4434 5314
rect 4434 5286 4436 5314
rect 4404 5284 4436 5286
rect 4404 5234 4436 5236
rect 4404 5206 4406 5234
rect 4406 5206 4434 5234
rect 4434 5206 4436 5234
rect 4404 5204 4436 5206
rect 4404 5154 4436 5156
rect 4404 5126 4406 5154
rect 4406 5126 4434 5154
rect 4434 5126 4436 5154
rect 4404 5124 4436 5126
rect 4404 5074 4436 5076
rect 4404 5046 4406 5074
rect 4406 5046 4434 5074
rect 4434 5046 4436 5074
rect 4404 5044 4436 5046
rect 4404 4994 4436 4996
rect 4404 4966 4406 4994
rect 4406 4966 4434 4994
rect 4434 4966 4436 4994
rect 4404 4964 4436 4966
rect 4404 4434 4436 4436
rect 4404 4406 4406 4434
rect 4406 4406 4434 4434
rect 4434 4406 4436 4434
rect 4404 4404 4436 4406
rect 4404 4354 4436 4356
rect 4404 4326 4406 4354
rect 4406 4326 4434 4354
rect 4434 4326 4436 4354
rect 4404 4324 4436 4326
rect 4404 4274 4436 4276
rect 4404 4246 4406 4274
rect 4406 4246 4434 4274
rect 4434 4246 4436 4274
rect 4404 4244 4436 4246
rect 4404 4194 4436 4196
rect 4404 4166 4406 4194
rect 4406 4166 4434 4194
rect 4434 4166 4436 4194
rect 4404 4164 4436 4166
rect 4404 4114 4436 4116
rect 4404 4086 4406 4114
rect 4406 4086 4434 4114
rect 4434 4086 4436 4114
rect 4404 4084 4436 4086
rect 4404 4034 4436 4036
rect 4404 4006 4406 4034
rect 4406 4006 4434 4034
rect 4434 4006 4436 4034
rect 4404 4004 4436 4006
rect 4404 3954 4436 3956
rect 4404 3926 4406 3954
rect 4406 3926 4434 3954
rect 4434 3926 4436 3954
rect 4404 3924 4436 3926
rect 4404 3154 4436 3156
rect 4404 3126 4406 3154
rect 4406 3126 4434 3154
rect 4434 3126 4436 3154
rect 4404 3124 4436 3126
rect 4404 3074 4436 3076
rect 4404 3046 4406 3074
rect 4406 3046 4434 3074
rect 4434 3046 4436 3074
rect 4404 3044 4436 3046
rect 4404 2994 4436 2996
rect 4404 2966 4406 2994
rect 4406 2966 4434 2994
rect 4434 2966 4436 2994
rect 4404 2964 4436 2966
rect 4404 2914 4436 2916
rect 4404 2886 4406 2914
rect 4406 2886 4434 2914
rect 4434 2886 4436 2914
rect 4404 2884 4436 2886
rect 4404 2834 4436 2836
rect 4404 2806 4406 2834
rect 4406 2806 4434 2834
rect 4434 2806 4436 2834
rect 4404 2804 4436 2806
rect 4404 2754 4436 2756
rect 4404 2726 4406 2754
rect 4406 2726 4434 2754
rect 4434 2726 4436 2754
rect 4404 2724 4436 2726
rect 4404 2674 4436 2676
rect 4404 2646 4406 2674
rect 4406 2646 4434 2674
rect 4434 2646 4436 2674
rect 4404 2644 4436 2646
rect 4404 2594 4436 2596
rect 4404 2566 4406 2594
rect 4406 2566 4434 2594
rect 4434 2566 4436 2594
rect 4404 2564 4436 2566
rect 4404 2514 4436 2516
rect 4404 2486 4406 2514
rect 4406 2486 4434 2514
rect 4434 2486 4436 2514
rect 4404 2484 4436 2486
rect 4404 2434 4436 2436
rect 4404 2406 4406 2434
rect 4406 2406 4434 2434
rect 4434 2406 4436 2434
rect 4404 2404 4436 2406
rect 4404 2354 4436 2356
rect 4404 2326 4406 2354
rect 4406 2326 4434 2354
rect 4434 2326 4436 2354
rect 4404 2324 4436 2326
rect 4404 2274 4436 2276
rect 4404 2246 4406 2274
rect 4406 2246 4434 2274
rect 4434 2246 4436 2274
rect 4404 2244 4436 2246
rect 4404 2194 4436 2196
rect 4404 2166 4406 2194
rect 4406 2166 4434 2194
rect 4434 2166 4436 2194
rect 4404 2164 4436 2166
rect 4404 2114 4436 2116
rect 4404 2086 4406 2114
rect 4406 2086 4434 2114
rect 4434 2086 4436 2114
rect 4404 2084 4436 2086
rect 4404 2034 4436 2036
rect 4404 2006 4406 2034
rect 4406 2006 4434 2034
rect 4434 2006 4436 2034
rect 4404 2004 4436 2006
rect 4404 1634 4436 1636
rect 4404 1606 4406 1634
rect 4406 1606 4434 1634
rect 4434 1606 4436 1634
rect 4404 1604 4436 1606
rect 4404 1554 4436 1556
rect 4404 1526 4406 1554
rect 4406 1526 4434 1554
rect 4434 1526 4436 1554
rect 4404 1524 4436 1526
rect 4404 1474 4436 1476
rect 4404 1446 4406 1474
rect 4406 1446 4434 1474
rect 4434 1446 4436 1474
rect 4404 1444 4436 1446
rect 4404 1394 4436 1396
rect 4404 1366 4406 1394
rect 4406 1366 4434 1394
rect 4434 1366 4436 1394
rect 4404 1364 4436 1366
rect 4404 1314 4436 1316
rect 4404 1286 4406 1314
rect 4406 1286 4434 1314
rect 4434 1286 4436 1314
rect 4404 1284 4436 1286
rect 4404 1234 4436 1236
rect 4404 1206 4406 1234
rect 4406 1206 4434 1234
rect 4434 1206 4436 1234
rect 4404 1204 4436 1206
rect 4404 1154 4436 1156
rect 4404 1126 4406 1154
rect 4406 1126 4434 1154
rect 4434 1126 4436 1154
rect 4404 1124 4436 1126
rect 4404 1074 4436 1076
rect 4404 1046 4406 1074
rect 4406 1046 4434 1074
rect 4434 1046 4436 1074
rect 4404 1044 4436 1046
rect 4404 754 4436 756
rect 4404 726 4406 754
rect 4406 726 4434 754
rect 4434 726 4436 754
rect 4404 724 4436 726
rect 4404 674 4436 676
rect 4404 646 4406 674
rect 4406 646 4434 674
rect 4434 646 4436 674
rect 4404 644 4436 646
rect 4404 594 4436 596
rect 4404 566 4406 594
rect 4406 566 4434 594
rect 4434 566 4436 594
rect 4404 564 4436 566
rect 4404 194 4436 196
rect 4404 166 4406 194
rect 4406 166 4434 194
rect 4434 166 4436 194
rect 4404 164 4436 166
rect 4404 114 4436 116
rect 4404 86 4406 114
rect 4406 86 4434 114
rect 4434 86 4436 114
rect 4404 84 4436 86
rect 4404 34 4436 36
rect 4404 6 4406 34
rect 4406 6 4434 34
rect 4434 6 4436 34
rect 4404 4 4436 6
rect 4484 13124 4516 13156
rect 4484 13084 4516 13116
rect 4484 13044 4516 13076
rect 4484 13004 4516 13036
rect 4484 12964 4516 12996
rect 4484 12634 4516 12636
rect 4484 12606 4486 12634
rect 4486 12606 4514 12634
rect 4514 12606 4516 12634
rect 4484 12604 4516 12606
rect 4484 12554 4516 12556
rect 4484 12526 4486 12554
rect 4486 12526 4514 12554
rect 4514 12526 4516 12554
rect 4484 12524 4516 12526
rect 4484 12474 4516 12476
rect 4484 12446 4486 12474
rect 4486 12446 4514 12474
rect 4514 12446 4516 12474
rect 4484 12444 4516 12446
rect 4484 12394 4516 12396
rect 4484 12366 4486 12394
rect 4486 12366 4514 12394
rect 4514 12366 4516 12394
rect 4484 12364 4516 12366
rect 4484 12314 4516 12316
rect 4484 12286 4486 12314
rect 4486 12286 4514 12314
rect 4514 12286 4516 12314
rect 4484 12284 4516 12286
rect 4484 12234 4516 12236
rect 4484 12206 4486 12234
rect 4486 12206 4514 12234
rect 4514 12206 4516 12234
rect 4484 12204 4516 12206
rect 4484 12154 4516 12156
rect 4484 12126 4486 12154
rect 4486 12126 4514 12154
rect 4514 12126 4516 12154
rect 4484 12124 4516 12126
rect 4484 11834 4516 11836
rect 4484 11806 4486 11834
rect 4486 11806 4514 11834
rect 4514 11806 4516 11834
rect 4484 11804 4516 11806
rect 4484 11754 4516 11756
rect 4484 11726 4486 11754
rect 4486 11726 4514 11754
rect 4514 11726 4516 11754
rect 4484 11724 4516 11726
rect 4484 11674 4516 11676
rect 4484 11646 4486 11674
rect 4486 11646 4514 11674
rect 4514 11646 4516 11674
rect 4484 11644 4516 11646
rect 4484 11594 4516 11596
rect 4484 11566 4486 11594
rect 4486 11566 4514 11594
rect 4514 11566 4516 11594
rect 4484 11564 4516 11566
rect 4484 11514 4516 11516
rect 4484 11486 4486 11514
rect 4486 11486 4514 11514
rect 4514 11486 4516 11514
rect 4484 11484 4516 11486
rect 4484 11434 4516 11436
rect 4484 11406 4486 11434
rect 4486 11406 4514 11434
rect 4514 11406 4516 11434
rect 4484 11404 4516 11406
rect 4484 10874 4516 10876
rect 4484 10846 4486 10874
rect 4486 10846 4514 10874
rect 4514 10846 4516 10874
rect 4484 10844 4516 10846
rect 4484 10794 4516 10796
rect 4484 10766 4486 10794
rect 4486 10766 4514 10794
rect 4514 10766 4516 10794
rect 4484 10764 4516 10766
rect 4484 10714 4516 10716
rect 4484 10686 4486 10714
rect 4486 10686 4514 10714
rect 4514 10686 4516 10714
rect 4484 10684 4516 10686
rect 4484 10634 4516 10636
rect 4484 10606 4486 10634
rect 4486 10606 4514 10634
rect 4514 10606 4516 10634
rect 4484 10604 4516 10606
rect 4484 10554 4516 10556
rect 4484 10526 4486 10554
rect 4486 10526 4514 10554
rect 4514 10526 4516 10554
rect 4484 10524 4516 10526
rect 4484 10474 4516 10476
rect 4484 10446 4486 10474
rect 4486 10446 4514 10474
rect 4514 10446 4516 10474
rect 4484 10444 4516 10446
rect 4484 10394 4516 10396
rect 4484 10366 4486 10394
rect 4486 10366 4514 10394
rect 4514 10366 4516 10394
rect 4484 10364 4516 10366
rect 4484 10314 4516 10316
rect 4484 10286 4486 10314
rect 4486 10286 4514 10314
rect 4514 10286 4516 10314
rect 4484 10284 4516 10286
rect 4484 10234 4516 10236
rect 4484 10206 4486 10234
rect 4486 10206 4514 10234
rect 4514 10206 4516 10234
rect 4484 10204 4516 10206
rect 4484 10154 4516 10156
rect 4484 10126 4486 10154
rect 4486 10126 4514 10154
rect 4514 10126 4516 10154
rect 4484 10124 4516 10126
rect 4484 10074 4516 10076
rect 4484 10046 4486 10074
rect 4486 10046 4514 10074
rect 4514 10046 4516 10074
rect 4484 10044 4516 10046
rect 4484 9994 4516 9996
rect 4484 9966 4486 9994
rect 4486 9966 4514 9994
rect 4514 9966 4516 9994
rect 4484 9964 4516 9966
rect 4484 9914 4516 9916
rect 4484 9886 4486 9914
rect 4486 9886 4514 9914
rect 4514 9886 4516 9914
rect 4484 9884 4516 9886
rect 4484 9834 4516 9836
rect 4484 9806 4486 9834
rect 4486 9806 4514 9834
rect 4514 9806 4516 9834
rect 4484 9804 4516 9806
rect 4484 9754 4516 9756
rect 4484 9726 4486 9754
rect 4486 9726 4514 9754
rect 4514 9726 4516 9754
rect 4484 9724 4516 9726
rect 4484 9354 4516 9356
rect 4484 9326 4486 9354
rect 4486 9326 4514 9354
rect 4514 9326 4516 9354
rect 4484 9324 4516 9326
rect 4484 9274 4516 9276
rect 4484 9246 4486 9274
rect 4486 9246 4514 9274
rect 4514 9246 4516 9274
rect 4484 9244 4516 9246
rect 4484 9194 4516 9196
rect 4484 9166 4486 9194
rect 4486 9166 4514 9194
rect 4514 9166 4516 9194
rect 4484 9164 4516 9166
rect 4484 8874 4516 8876
rect 4484 8846 4486 8874
rect 4486 8846 4514 8874
rect 4514 8846 4516 8874
rect 4484 8844 4516 8846
rect 4484 8794 4516 8796
rect 4484 8766 4486 8794
rect 4486 8766 4514 8794
rect 4514 8766 4516 8794
rect 4484 8764 4516 8766
rect 4484 8714 4516 8716
rect 4484 8686 4486 8714
rect 4486 8686 4514 8714
rect 4514 8686 4516 8714
rect 4484 8684 4516 8686
rect 4484 8634 4516 8636
rect 4484 8606 4486 8634
rect 4486 8606 4514 8634
rect 4514 8606 4516 8634
rect 4484 8604 4516 8606
rect 4484 8554 4516 8556
rect 4484 8526 4486 8554
rect 4486 8526 4514 8554
rect 4514 8526 4516 8554
rect 4484 8524 4516 8526
rect 4484 7634 4516 7636
rect 4484 7606 4486 7634
rect 4486 7606 4514 7634
rect 4514 7606 4516 7634
rect 4484 7604 4516 7606
rect 4484 7554 4516 7556
rect 4484 7526 4486 7554
rect 4486 7526 4514 7554
rect 4514 7526 4516 7554
rect 4484 7524 4516 7526
rect 4484 7474 4516 7476
rect 4484 7446 4486 7474
rect 4486 7446 4514 7474
rect 4514 7446 4516 7474
rect 4484 7444 4516 7446
rect 4484 7394 4516 7396
rect 4484 7366 4486 7394
rect 4486 7366 4514 7394
rect 4514 7366 4516 7394
rect 4484 7364 4516 7366
rect 4484 7314 4516 7316
rect 4484 7286 4486 7314
rect 4486 7286 4514 7314
rect 4514 7286 4516 7314
rect 4484 7284 4516 7286
rect 4484 7234 4516 7236
rect 4484 7206 4486 7234
rect 4486 7206 4514 7234
rect 4514 7206 4516 7234
rect 4484 7204 4516 7206
rect 4484 7154 4516 7156
rect 4484 7126 4486 7154
rect 4486 7126 4514 7154
rect 4514 7126 4516 7154
rect 4484 7124 4516 7126
rect 4484 7074 4516 7076
rect 4484 7046 4486 7074
rect 4486 7046 4514 7074
rect 4514 7046 4516 7074
rect 4484 7044 4516 7046
rect 4484 6754 4516 6756
rect 4484 6726 4486 6754
rect 4486 6726 4514 6754
rect 4514 6726 4516 6754
rect 4484 6724 4516 6726
rect 4484 6674 4516 6676
rect 4484 6646 4486 6674
rect 4486 6646 4514 6674
rect 4514 6646 4516 6674
rect 4484 6644 4516 6646
rect 4484 6594 4516 6596
rect 4484 6566 4486 6594
rect 4486 6566 4514 6594
rect 4514 6566 4516 6594
rect 4484 6564 4516 6566
rect 4484 6514 4516 6516
rect 4484 6486 4486 6514
rect 4486 6486 4514 6514
rect 4514 6486 4516 6514
rect 4484 6484 4516 6486
rect 4484 6434 4516 6436
rect 4484 6406 4486 6434
rect 4486 6406 4514 6434
rect 4514 6406 4516 6434
rect 4484 6404 4516 6406
rect 4484 6354 4516 6356
rect 4484 6326 4486 6354
rect 4486 6326 4514 6354
rect 4514 6326 4516 6354
rect 4484 6324 4516 6326
rect 4484 5794 4516 5796
rect 4484 5766 4486 5794
rect 4486 5766 4514 5794
rect 4514 5766 4516 5794
rect 4484 5764 4516 5766
rect 4484 5714 4516 5716
rect 4484 5686 4486 5714
rect 4486 5686 4514 5714
rect 4514 5686 4516 5714
rect 4484 5684 4516 5686
rect 4484 5634 4516 5636
rect 4484 5606 4486 5634
rect 4486 5606 4514 5634
rect 4514 5606 4516 5634
rect 4484 5604 4516 5606
rect 4484 5554 4516 5556
rect 4484 5526 4486 5554
rect 4486 5526 4514 5554
rect 4514 5526 4516 5554
rect 4484 5524 4516 5526
rect 4484 5474 4516 5476
rect 4484 5446 4486 5474
rect 4486 5446 4514 5474
rect 4514 5446 4516 5474
rect 4484 5444 4516 5446
rect 4484 5394 4516 5396
rect 4484 5366 4486 5394
rect 4486 5366 4514 5394
rect 4514 5366 4516 5394
rect 4484 5364 4516 5366
rect 4484 5314 4516 5316
rect 4484 5286 4486 5314
rect 4486 5286 4514 5314
rect 4514 5286 4516 5314
rect 4484 5284 4516 5286
rect 4484 5234 4516 5236
rect 4484 5206 4486 5234
rect 4486 5206 4514 5234
rect 4514 5206 4516 5234
rect 4484 5204 4516 5206
rect 4484 5154 4516 5156
rect 4484 5126 4486 5154
rect 4486 5126 4514 5154
rect 4514 5126 4516 5154
rect 4484 5124 4516 5126
rect 4484 5074 4516 5076
rect 4484 5046 4486 5074
rect 4486 5046 4514 5074
rect 4514 5046 4516 5074
rect 4484 5044 4516 5046
rect 4484 4994 4516 4996
rect 4484 4966 4486 4994
rect 4486 4966 4514 4994
rect 4514 4966 4516 4994
rect 4484 4964 4516 4966
rect 4484 4434 4516 4436
rect 4484 4406 4486 4434
rect 4486 4406 4514 4434
rect 4514 4406 4516 4434
rect 4484 4404 4516 4406
rect 4484 4354 4516 4356
rect 4484 4326 4486 4354
rect 4486 4326 4514 4354
rect 4514 4326 4516 4354
rect 4484 4324 4516 4326
rect 4484 4274 4516 4276
rect 4484 4246 4486 4274
rect 4486 4246 4514 4274
rect 4514 4246 4516 4274
rect 4484 4244 4516 4246
rect 4484 4194 4516 4196
rect 4484 4166 4486 4194
rect 4486 4166 4514 4194
rect 4514 4166 4516 4194
rect 4484 4164 4516 4166
rect 4484 4114 4516 4116
rect 4484 4086 4486 4114
rect 4486 4086 4514 4114
rect 4514 4086 4516 4114
rect 4484 4084 4516 4086
rect 4484 4034 4516 4036
rect 4484 4006 4486 4034
rect 4486 4006 4514 4034
rect 4514 4006 4516 4034
rect 4484 4004 4516 4006
rect 4484 3954 4516 3956
rect 4484 3926 4486 3954
rect 4486 3926 4514 3954
rect 4514 3926 4516 3954
rect 4484 3924 4516 3926
rect 4484 3154 4516 3156
rect 4484 3126 4486 3154
rect 4486 3126 4514 3154
rect 4514 3126 4516 3154
rect 4484 3124 4516 3126
rect 4484 3074 4516 3076
rect 4484 3046 4486 3074
rect 4486 3046 4514 3074
rect 4514 3046 4516 3074
rect 4484 3044 4516 3046
rect 4484 2994 4516 2996
rect 4484 2966 4486 2994
rect 4486 2966 4514 2994
rect 4514 2966 4516 2994
rect 4484 2964 4516 2966
rect 4484 2914 4516 2916
rect 4484 2886 4486 2914
rect 4486 2886 4514 2914
rect 4514 2886 4516 2914
rect 4484 2884 4516 2886
rect 4484 2834 4516 2836
rect 4484 2806 4486 2834
rect 4486 2806 4514 2834
rect 4514 2806 4516 2834
rect 4484 2804 4516 2806
rect 4484 2754 4516 2756
rect 4484 2726 4486 2754
rect 4486 2726 4514 2754
rect 4514 2726 4516 2754
rect 4484 2724 4516 2726
rect 4484 2674 4516 2676
rect 4484 2646 4486 2674
rect 4486 2646 4514 2674
rect 4514 2646 4516 2674
rect 4484 2644 4516 2646
rect 4484 2594 4516 2596
rect 4484 2566 4486 2594
rect 4486 2566 4514 2594
rect 4514 2566 4516 2594
rect 4484 2564 4516 2566
rect 4484 2514 4516 2516
rect 4484 2486 4486 2514
rect 4486 2486 4514 2514
rect 4514 2486 4516 2514
rect 4484 2484 4516 2486
rect 4484 2434 4516 2436
rect 4484 2406 4486 2434
rect 4486 2406 4514 2434
rect 4514 2406 4516 2434
rect 4484 2404 4516 2406
rect 4484 2354 4516 2356
rect 4484 2326 4486 2354
rect 4486 2326 4514 2354
rect 4514 2326 4516 2354
rect 4484 2324 4516 2326
rect 4484 2274 4516 2276
rect 4484 2246 4486 2274
rect 4486 2246 4514 2274
rect 4514 2246 4516 2274
rect 4484 2244 4516 2246
rect 4484 2194 4516 2196
rect 4484 2166 4486 2194
rect 4486 2166 4514 2194
rect 4514 2166 4516 2194
rect 4484 2164 4516 2166
rect 4484 2114 4516 2116
rect 4484 2086 4486 2114
rect 4486 2086 4514 2114
rect 4514 2086 4516 2114
rect 4484 2084 4516 2086
rect 4484 2034 4516 2036
rect 4484 2006 4486 2034
rect 4486 2006 4514 2034
rect 4514 2006 4516 2034
rect 4484 2004 4516 2006
rect 4484 1634 4516 1636
rect 4484 1606 4486 1634
rect 4486 1606 4514 1634
rect 4514 1606 4516 1634
rect 4484 1604 4516 1606
rect 4484 1554 4516 1556
rect 4484 1526 4486 1554
rect 4486 1526 4514 1554
rect 4514 1526 4516 1554
rect 4484 1524 4516 1526
rect 4484 1474 4516 1476
rect 4484 1446 4486 1474
rect 4486 1446 4514 1474
rect 4514 1446 4516 1474
rect 4484 1444 4516 1446
rect 4484 1394 4516 1396
rect 4484 1366 4486 1394
rect 4486 1366 4514 1394
rect 4514 1366 4516 1394
rect 4484 1364 4516 1366
rect 4484 1314 4516 1316
rect 4484 1286 4486 1314
rect 4486 1286 4514 1314
rect 4514 1286 4516 1314
rect 4484 1284 4516 1286
rect 4484 1234 4516 1236
rect 4484 1206 4486 1234
rect 4486 1206 4514 1234
rect 4514 1206 4516 1234
rect 4484 1204 4516 1206
rect 4484 1154 4516 1156
rect 4484 1126 4486 1154
rect 4486 1126 4514 1154
rect 4514 1126 4516 1154
rect 4484 1124 4516 1126
rect 4484 1074 4516 1076
rect 4484 1046 4486 1074
rect 4486 1046 4514 1074
rect 4514 1046 4516 1074
rect 4484 1044 4516 1046
rect 4484 754 4516 756
rect 4484 726 4486 754
rect 4486 726 4514 754
rect 4514 726 4516 754
rect 4484 724 4516 726
rect 4484 674 4516 676
rect 4484 646 4486 674
rect 4486 646 4514 674
rect 4514 646 4516 674
rect 4484 644 4516 646
rect 4484 594 4516 596
rect 4484 566 4486 594
rect 4486 566 4514 594
rect 4514 566 4516 594
rect 4484 564 4516 566
rect 4484 194 4516 196
rect 4484 166 4486 194
rect 4486 166 4514 194
rect 4514 166 4516 194
rect 4484 164 4516 166
rect 4484 114 4516 116
rect 4484 86 4486 114
rect 4486 86 4514 114
rect 4514 86 4516 114
rect 4484 84 4516 86
rect 4484 34 4516 36
rect 4484 6 4486 34
rect 4486 6 4514 34
rect 4514 6 4516 34
rect 4484 4 4516 6
rect 4564 13844 4596 13876
rect 4644 13924 4676 13956
rect 4644 13764 4676 13796
rect 5044 13684 5076 13716
rect 4644 13124 4676 13156
rect 4644 13084 4676 13116
rect 4644 13044 4676 13076
rect 4644 13004 4676 13036
rect 4644 12964 4676 12996
rect 4644 12634 4676 12636
rect 4644 12606 4646 12634
rect 4646 12606 4674 12634
rect 4674 12606 4676 12634
rect 4644 12604 4676 12606
rect 4644 12554 4676 12556
rect 4644 12526 4646 12554
rect 4646 12526 4674 12554
rect 4674 12526 4676 12554
rect 4644 12524 4676 12526
rect 4644 12474 4676 12476
rect 4644 12446 4646 12474
rect 4646 12446 4674 12474
rect 4674 12446 4676 12474
rect 4644 12444 4676 12446
rect 4644 12394 4676 12396
rect 4644 12366 4646 12394
rect 4646 12366 4674 12394
rect 4674 12366 4676 12394
rect 4644 12364 4676 12366
rect 4644 12314 4676 12316
rect 4644 12286 4646 12314
rect 4646 12286 4674 12314
rect 4674 12286 4676 12314
rect 4644 12284 4676 12286
rect 4644 12234 4676 12236
rect 4644 12206 4646 12234
rect 4646 12206 4674 12234
rect 4674 12206 4676 12234
rect 4644 12204 4676 12206
rect 4644 12154 4676 12156
rect 4644 12126 4646 12154
rect 4646 12126 4674 12154
rect 4674 12126 4676 12154
rect 4644 12124 4676 12126
rect 4644 11834 4676 11836
rect 4644 11806 4646 11834
rect 4646 11806 4674 11834
rect 4674 11806 4676 11834
rect 4644 11804 4676 11806
rect 4644 11754 4676 11756
rect 4644 11726 4646 11754
rect 4646 11726 4674 11754
rect 4674 11726 4676 11754
rect 4644 11724 4676 11726
rect 4644 11674 4676 11676
rect 4644 11646 4646 11674
rect 4646 11646 4674 11674
rect 4674 11646 4676 11674
rect 4644 11644 4676 11646
rect 4644 11594 4676 11596
rect 4644 11566 4646 11594
rect 4646 11566 4674 11594
rect 4674 11566 4676 11594
rect 4644 11564 4676 11566
rect 4644 11514 4676 11516
rect 4644 11486 4646 11514
rect 4646 11486 4674 11514
rect 4674 11486 4676 11514
rect 4644 11484 4676 11486
rect 4644 11434 4676 11436
rect 4644 11406 4646 11434
rect 4646 11406 4674 11434
rect 4674 11406 4676 11434
rect 4644 11404 4676 11406
rect 4644 10874 4676 10876
rect 4644 10846 4646 10874
rect 4646 10846 4674 10874
rect 4674 10846 4676 10874
rect 4644 10844 4676 10846
rect 4644 10794 4676 10796
rect 4644 10766 4646 10794
rect 4646 10766 4674 10794
rect 4674 10766 4676 10794
rect 4644 10764 4676 10766
rect 4644 10714 4676 10716
rect 4644 10686 4646 10714
rect 4646 10686 4674 10714
rect 4674 10686 4676 10714
rect 4644 10684 4676 10686
rect 4644 10634 4676 10636
rect 4644 10606 4646 10634
rect 4646 10606 4674 10634
rect 4674 10606 4676 10634
rect 4644 10604 4676 10606
rect 4644 10554 4676 10556
rect 4644 10526 4646 10554
rect 4646 10526 4674 10554
rect 4674 10526 4676 10554
rect 4644 10524 4676 10526
rect 4644 10474 4676 10476
rect 4644 10446 4646 10474
rect 4646 10446 4674 10474
rect 4674 10446 4676 10474
rect 4644 10444 4676 10446
rect 4644 10394 4676 10396
rect 4644 10366 4646 10394
rect 4646 10366 4674 10394
rect 4674 10366 4676 10394
rect 4644 10364 4676 10366
rect 4644 10314 4676 10316
rect 4644 10286 4646 10314
rect 4646 10286 4674 10314
rect 4674 10286 4676 10314
rect 4644 10284 4676 10286
rect 4644 10234 4676 10236
rect 4644 10206 4646 10234
rect 4646 10206 4674 10234
rect 4674 10206 4676 10234
rect 4644 10204 4676 10206
rect 4644 10154 4676 10156
rect 4644 10126 4646 10154
rect 4646 10126 4674 10154
rect 4674 10126 4676 10154
rect 4644 10124 4676 10126
rect 4644 10074 4676 10076
rect 4644 10046 4646 10074
rect 4646 10046 4674 10074
rect 4674 10046 4676 10074
rect 4644 10044 4676 10046
rect 4644 9994 4676 9996
rect 4644 9966 4646 9994
rect 4646 9966 4674 9994
rect 4674 9966 4676 9994
rect 4644 9964 4676 9966
rect 4644 9914 4676 9916
rect 4644 9886 4646 9914
rect 4646 9886 4674 9914
rect 4674 9886 4676 9914
rect 4644 9884 4676 9886
rect 4644 9834 4676 9836
rect 4644 9806 4646 9834
rect 4646 9806 4674 9834
rect 4674 9806 4676 9834
rect 4644 9804 4676 9806
rect 4644 9754 4676 9756
rect 4644 9726 4646 9754
rect 4646 9726 4674 9754
rect 4674 9726 4676 9754
rect 4644 9724 4676 9726
rect 4644 9354 4676 9356
rect 4644 9326 4646 9354
rect 4646 9326 4674 9354
rect 4674 9326 4676 9354
rect 4644 9324 4676 9326
rect 4644 9274 4676 9276
rect 4644 9246 4646 9274
rect 4646 9246 4674 9274
rect 4674 9246 4676 9274
rect 4644 9244 4676 9246
rect 4644 9194 4676 9196
rect 4644 9166 4646 9194
rect 4646 9166 4674 9194
rect 4674 9166 4676 9194
rect 4644 9164 4676 9166
rect 4644 8874 4676 8876
rect 4644 8846 4646 8874
rect 4646 8846 4674 8874
rect 4674 8846 4676 8874
rect 4644 8844 4676 8846
rect 4644 8794 4676 8796
rect 4644 8766 4646 8794
rect 4646 8766 4674 8794
rect 4674 8766 4676 8794
rect 4644 8764 4676 8766
rect 4644 8714 4676 8716
rect 4644 8686 4646 8714
rect 4646 8686 4674 8714
rect 4674 8686 4676 8714
rect 4644 8684 4676 8686
rect 4644 8634 4676 8636
rect 4644 8606 4646 8634
rect 4646 8606 4674 8634
rect 4674 8606 4676 8634
rect 4644 8604 4676 8606
rect 4644 8554 4676 8556
rect 4644 8526 4646 8554
rect 4646 8526 4674 8554
rect 4674 8526 4676 8554
rect 4644 8524 4676 8526
rect 4644 7634 4676 7636
rect 4644 7606 4646 7634
rect 4646 7606 4674 7634
rect 4674 7606 4676 7634
rect 4644 7604 4676 7606
rect 4644 7554 4676 7556
rect 4644 7526 4646 7554
rect 4646 7526 4674 7554
rect 4674 7526 4676 7554
rect 4644 7524 4676 7526
rect 4644 7474 4676 7476
rect 4644 7446 4646 7474
rect 4646 7446 4674 7474
rect 4674 7446 4676 7474
rect 4644 7444 4676 7446
rect 4644 7394 4676 7396
rect 4644 7366 4646 7394
rect 4646 7366 4674 7394
rect 4674 7366 4676 7394
rect 4644 7364 4676 7366
rect 4644 7314 4676 7316
rect 4644 7286 4646 7314
rect 4646 7286 4674 7314
rect 4674 7286 4676 7314
rect 4644 7284 4676 7286
rect 4644 7234 4676 7236
rect 4644 7206 4646 7234
rect 4646 7206 4674 7234
rect 4674 7206 4676 7234
rect 4644 7204 4676 7206
rect 4644 7154 4676 7156
rect 4644 7126 4646 7154
rect 4646 7126 4674 7154
rect 4674 7126 4676 7154
rect 4644 7124 4676 7126
rect 4644 7074 4676 7076
rect 4644 7046 4646 7074
rect 4646 7046 4674 7074
rect 4674 7046 4676 7074
rect 4644 7044 4676 7046
rect 4644 6754 4676 6756
rect 4644 6726 4646 6754
rect 4646 6726 4674 6754
rect 4674 6726 4676 6754
rect 4644 6724 4676 6726
rect 4644 6674 4676 6676
rect 4644 6646 4646 6674
rect 4646 6646 4674 6674
rect 4674 6646 4676 6674
rect 4644 6644 4676 6646
rect 4644 6594 4676 6596
rect 4644 6566 4646 6594
rect 4646 6566 4674 6594
rect 4674 6566 4676 6594
rect 4644 6564 4676 6566
rect 4644 6514 4676 6516
rect 4644 6486 4646 6514
rect 4646 6486 4674 6514
rect 4674 6486 4676 6514
rect 4644 6484 4676 6486
rect 4644 6434 4676 6436
rect 4644 6406 4646 6434
rect 4646 6406 4674 6434
rect 4674 6406 4676 6434
rect 4644 6404 4676 6406
rect 4644 6354 4676 6356
rect 4644 6326 4646 6354
rect 4646 6326 4674 6354
rect 4674 6326 4676 6354
rect 4644 6324 4676 6326
rect 4644 5794 4676 5796
rect 4644 5766 4646 5794
rect 4646 5766 4674 5794
rect 4674 5766 4676 5794
rect 4644 5764 4676 5766
rect 4644 5714 4676 5716
rect 4644 5686 4646 5714
rect 4646 5686 4674 5714
rect 4674 5686 4676 5714
rect 4644 5684 4676 5686
rect 4644 5634 4676 5636
rect 4644 5606 4646 5634
rect 4646 5606 4674 5634
rect 4674 5606 4676 5634
rect 4644 5604 4676 5606
rect 4644 5554 4676 5556
rect 4644 5526 4646 5554
rect 4646 5526 4674 5554
rect 4674 5526 4676 5554
rect 4644 5524 4676 5526
rect 4644 5474 4676 5476
rect 4644 5446 4646 5474
rect 4646 5446 4674 5474
rect 4674 5446 4676 5474
rect 4644 5444 4676 5446
rect 4644 5394 4676 5396
rect 4644 5366 4646 5394
rect 4646 5366 4674 5394
rect 4674 5366 4676 5394
rect 4644 5364 4676 5366
rect 4644 5314 4676 5316
rect 4644 5286 4646 5314
rect 4646 5286 4674 5314
rect 4674 5286 4676 5314
rect 4644 5284 4676 5286
rect 4644 5234 4676 5236
rect 4644 5206 4646 5234
rect 4646 5206 4674 5234
rect 4674 5206 4676 5234
rect 4644 5204 4676 5206
rect 4644 5154 4676 5156
rect 4644 5126 4646 5154
rect 4646 5126 4674 5154
rect 4674 5126 4676 5154
rect 4644 5124 4676 5126
rect 4644 5074 4676 5076
rect 4644 5046 4646 5074
rect 4646 5046 4674 5074
rect 4674 5046 4676 5074
rect 4644 5044 4676 5046
rect 4644 4994 4676 4996
rect 4644 4966 4646 4994
rect 4646 4966 4674 4994
rect 4674 4966 4676 4994
rect 4644 4964 4676 4966
rect 4644 4434 4676 4436
rect 4644 4406 4646 4434
rect 4646 4406 4674 4434
rect 4674 4406 4676 4434
rect 4644 4404 4676 4406
rect 4644 4354 4676 4356
rect 4644 4326 4646 4354
rect 4646 4326 4674 4354
rect 4674 4326 4676 4354
rect 4644 4324 4676 4326
rect 4644 4274 4676 4276
rect 4644 4246 4646 4274
rect 4646 4246 4674 4274
rect 4674 4246 4676 4274
rect 4644 4244 4676 4246
rect 4644 4194 4676 4196
rect 4644 4166 4646 4194
rect 4646 4166 4674 4194
rect 4674 4166 4676 4194
rect 4644 4164 4676 4166
rect 4644 4114 4676 4116
rect 4644 4086 4646 4114
rect 4646 4086 4674 4114
rect 4674 4086 4676 4114
rect 4644 4084 4676 4086
rect 4644 4034 4676 4036
rect 4644 4006 4646 4034
rect 4646 4006 4674 4034
rect 4674 4006 4676 4034
rect 4644 4004 4676 4006
rect 4644 3954 4676 3956
rect 4644 3926 4646 3954
rect 4646 3926 4674 3954
rect 4674 3926 4676 3954
rect 4644 3924 4676 3926
rect 4644 3154 4676 3156
rect 4644 3126 4646 3154
rect 4646 3126 4674 3154
rect 4674 3126 4676 3154
rect 4644 3124 4676 3126
rect 4644 3074 4676 3076
rect 4644 3046 4646 3074
rect 4646 3046 4674 3074
rect 4674 3046 4676 3074
rect 4644 3044 4676 3046
rect 4644 2994 4676 2996
rect 4644 2966 4646 2994
rect 4646 2966 4674 2994
rect 4674 2966 4676 2994
rect 4644 2964 4676 2966
rect 4644 2914 4676 2916
rect 4644 2886 4646 2914
rect 4646 2886 4674 2914
rect 4674 2886 4676 2914
rect 4644 2884 4676 2886
rect 4644 2834 4676 2836
rect 4644 2806 4646 2834
rect 4646 2806 4674 2834
rect 4674 2806 4676 2834
rect 4644 2804 4676 2806
rect 4644 2754 4676 2756
rect 4644 2726 4646 2754
rect 4646 2726 4674 2754
rect 4674 2726 4676 2754
rect 4644 2724 4676 2726
rect 4644 2674 4676 2676
rect 4644 2646 4646 2674
rect 4646 2646 4674 2674
rect 4674 2646 4676 2674
rect 4644 2644 4676 2646
rect 4644 2594 4676 2596
rect 4644 2566 4646 2594
rect 4646 2566 4674 2594
rect 4674 2566 4676 2594
rect 4644 2564 4676 2566
rect 4644 2514 4676 2516
rect 4644 2486 4646 2514
rect 4646 2486 4674 2514
rect 4674 2486 4676 2514
rect 4644 2484 4676 2486
rect 4644 2434 4676 2436
rect 4644 2406 4646 2434
rect 4646 2406 4674 2434
rect 4674 2406 4676 2434
rect 4644 2404 4676 2406
rect 4644 2354 4676 2356
rect 4644 2326 4646 2354
rect 4646 2326 4674 2354
rect 4674 2326 4676 2354
rect 4644 2324 4676 2326
rect 4644 2274 4676 2276
rect 4644 2246 4646 2274
rect 4646 2246 4674 2274
rect 4674 2246 4676 2274
rect 4644 2244 4676 2246
rect 4644 2194 4676 2196
rect 4644 2166 4646 2194
rect 4646 2166 4674 2194
rect 4674 2166 4676 2194
rect 4644 2164 4676 2166
rect 4644 2114 4676 2116
rect 4644 2086 4646 2114
rect 4646 2086 4674 2114
rect 4674 2086 4676 2114
rect 4644 2084 4676 2086
rect 4644 2034 4676 2036
rect 4644 2006 4646 2034
rect 4646 2006 4674 2034
rect 4674 2006 4676 2034
rect 4644 2004 4676 2006
rect 4644 1634 4676 1636
rect 4644 1606 4646 1634
rect 4646 1606 4674 1634
rect 4674 1606 4676 1634
rect 4644 1604 4676 1606
rect 4644 1554 4676 1556
rect 4644 1526 4646 1554
rect 4646 1526 4674 1554
rect 4674 1526 4676 1554
rect 4644 1524 4676 1526
rect 4644 1474 4676 1476
rect 4644 1446 4646 1474
rect 4646 1446 4674 1474
rect 4674 1446 4676 1474
rect 4644 1444 4676 1446
rect 4644 1394 4676 1396
rect 4644 1366 4646 1394
rect 4646 1366 4674 1394
rect 4674 1366 4676 1394
rect 4644 1364 4676 1366
rect 4644 1314 4676 1316
rect 4644 1286 4646 1314
rect 4646 1286 4674 1314
rect 4674 1286 4676 1314
rect 4644 1284 4676 1286
rect 4644 1234 4676 1236
rect 4644 1206 4646 1234
rect 4646 1206 4674 1234
rect 4674 1206 4676 1234
rect 4644 1204 4676 1206
rect 4644 1154 4676 1156
rect 4644 1126 4646 1154
rect 4646 1126 4674 1154
rect 4674 1126 4676 1154
rect 4644 1124 4676 1126
rect 4644 1074 4676 1076
rect 4644 1046 4646 1074
rect 4646 1046 4674 1074
rect 4674 1046 4676 1074
rect 4644 1044 4676 1046
rect 4644 754 4676 756
rect 4644 726 4646 754
rect 4646 726 4674 754
rect 4674 726 4676 754
rect 4644 724 4676 726
rect 4644 674 4676 676
rect 4644 646 4646 674
rect 4646 646 4674 674
rect 4674 646 4676 674
rect 4644 644 4676 646
rect 4644 594 4676 596
rect 4644 566 4646 594
rect 4646 566 4674 594
rect 4674 566 4676 594
rect 4644 564 4676 566
rect 4644 194 4676 196
rect 4644 166 4646 194
rect 4646 166 4674 194
rect 4674 166 4676 194
rect 4644 164 4676 166
rect 4644 114 4676 116
rect 4644 86 4646 114
rect 4646 86 4674 114
rect 4674 86 4676 114
rect 4644 84 4676 86
rect 4644 34 4676 36
rect 4644 6 4646 34
rect 4646 6 4674 34
rect 4674 6 4676 34
rect 4644 4 4676 6
rect 4724 13364 4756 13396
rect 4724 13324 4756 13356
rect 4724 13284 4756 13316
rect 4724 13244 4756 13276
rect 4724 13204 4756 13236
rect 4884 13364 4916 13396
rect 4884 13324 4916 13356
rect 4884 13284 4916 13316
rect 4884 13244 4916 13276
rect 4884 13204 4916 13236
rect 4724 12634 4756 12636
rect 4724 12606 4726 12634
rect 4726 12606 4754 12634
rect 4754 12606 4756 12634
rect 4724 12604 4756 12606
rect 4724 12554 4756 12556
rect 4724 12526 4726 12554
rect 4726 12526 4754 12554
rect 4754 12526 4756 12554
rect 4724 12524 4756 12526
rect 4724 12474 4756 12476
rect 4724 12446 4726 12474
rect 4726 12446 4754 12474
rect 4754 12446 4756 12474
rect 4724 12444 4756 12446
rect 4724 12394 4756 12396
rect 4724 12366 4726 12394
rect 4726 12366 4754 12394
rect 4754 12366 4756 12394
rect 4724 12364 4756 12366
rect 4724 12314 4756 12316
rect 4724 12286 4726 12314
rect 4726 12286 4754 12314
rect 4754 12286 4756 12314
rect 4724 12284 4756 12286
rect 4724 12234 4756 12236
rect 4724 12206 4726 12234
rect 4726 12206 4754 12234
rect 4754 12206 4756 12234
rect 4724 12204 4756 12206
rect 4724 12154 4756 12156
rect 4724 12126 4726 12154
rect 4726 12126 4754 12154
rect 4754 12126 4756 12154
rect 4724 12124 4756 12126
rect 4724 11834 4756 11836
rect 4724 11806 4726 11834
rect 4726 11806 4754 11834
rect 4754 11806 4756 11834
rect 4724 11804 4756 11806
rect 4724 11754 4756 11756
rect 4724 11726 4726 11754
rect 4726 11726 4754 11754
rect 4754 11726 4756 11754
rect 4724 11724 4756 11726
rect 4724 11674 4756 11676
rect 4724 11646 4726 11674
rect 4726 11646 4754 11674
rect 4754 11646 4756 11674
rect 4724 11644 4756 11646
rect 4724 11594 4756 11596
rect 4724 11566 4726 11594
rect 4726 11566 4754 11594
rect 4754 11566 4756 11594
rect 4724 11564 4756 11566
rect 4724 11514 4756 11516
rect 4724 11486 4726 11514
rect 4726 11486 4754 11514
rect 4754 11486 4756 11514
rect 4724 11484 4756 11486
rect 4724 11434 4756 11436
rect 4724 11406 4726 11434
rect 4726 11406 4754 11434
rect 4754 11406 4756 11434
rect 4724 11404 4756 11406
rect 4724 10874 4756 10876
rect 4724 10846 4726 10874
rect 4726 10846 4754 10874
rect 4754 10846 4756 10874
rect 4724 10844 4756 10846
rect 4724 10794 4756 10796
rect 4724 10766 4726 10794
rect 4726 10766 4754 10794
rect 4754 10766 4756 10794
rect 4724 10764 4756 10766
rect 4724 10714 4756 10716
rect 4724 10686 4726 10714
rect 4726 10686 4754 10714
rect 4754 10686 4756 10714
rect 4724 10684 4756 10686
rect 4724 10634 4756 10636
rect 4724 10606 4726 10634
rect 4726 10606 4754 10634
rect 4754 10606 4756 10634
rect 4724 10604 4756 10606
rect 4724 10554 4756 10556
rect 4724 10526 4726 10554
rect 4726 10526 4754 10554
rect 4754 10526 4756 10554
rect 4724 10524 4756 10526
rect 4724 10474 4756 10476
rect 4724 10446 4726 10474
rect 4726 10446 4754 10474
rect 4754 10446 4756 10474
rect 4724 10444 4756 10446
rect 4724 10394 4756 10396
rect 4724 10366 4726 10394
rect 4726 10366 4754 10394
rect 4754 10366 4756 10394
rect 4724 10364 4756 10366
rect 4724 10314 4756 10316
rect 4724 10286 4726 10314
rect 4726 10286 4754 10314
rect 4754 10286 4756 10314
rect 4724 10284 4756 10286
rect 4724 10234 4756 10236
rect 4724 10206 4726 10234
rect 4726 10206 4754 10234
rect 4754 10206 4756 10234
rect 4724 10204 4756 10206
rect 4724 10154 4756 10156
rect 4724 10126 4726 10154
rect 4726 10126 4754 10154
rect 4754 10126 4756 10154
rect 4724 10124 4756 10126
rect 4724 10074 4756 10076
rect 4724 10046 4726 10074
rect 4726 10046 4754 10074
rect 4754 10046 4756 10074
rect 4724 10044 4756 10046
rect 4724 9994 4756 9996
rect 4724 9966 4726 9994
rect 4726 9966 4754 9994
rect 4754 9966 4756 9994
rect 4724 9964 4756 9966
rect 4724 9914 4756 9916
rect 4724 9886 4726 9914
rect 4726 9886 4754 9914
rect 4754 9886 4756 9914
rect 4724 9884 4756 9886
rect 4724 9834 4756 9836
rect 4724 9806 4726 9834
rect 4726 9806 4754 9834
rect 4754 9806 4756 9834
rect 4724 9804 4756 9806
rect 4724 9754 4756 9756
rect 4724 9726 4726 9754
rect 4726 9726 4754 9754
rect 4754 9726 4756 9754
rect 4724 9724 4756 9726
rect 4724 9354 4756 9356
rect 4724 9326 4726 9354
rect 4726 9326 4754 9354
rect 4754 9326 4756 9354
rect 4724 9324 4756 9326
rect 4724 9274 4756 9276
rect 4724 9246 4726 9274
rect 4726 9246 4754 9274
rect 4754 9246 4756 9274
rect 4724 9244 4756 9246
rect 4724 9194 4756 9196
rect 4724 9166 4726 9194
rect 4726 9166 4754 9194
rect 4754 9166 4756 9194
rect 4724 9164 4756 9166
rect 4724 8874 4756 8876
rect 4724 8846 4726 8874
rect 4726 8846 4754 8874
rect 4754 8846 4756 8874
rect 4724 8844 4756 8846
rect 4724 8794 4756 8796
rect 4724 8766 4726 8794
rect 4726 8766 4754 8794
rect 4754 8766 4756 8794
rect 4724 8764 4756 8766
rect 4724 8714 4756 8716
rect 4724 8686 4726 8714
rect 4726 8686 4754 8714
rect 4754 8686 4756 8714
rect 4724 8684 4756 8686
rect 4724 8634 4756 8636
rect 4724 8606 4726 8634
rect 4726 8606 4754 8634
rect 4754 8606 4756 8634
rect 4724 8604 4756 8606
rect 4724 8554 4756 8556
rect 4724 8526 4726 8554
rect 4726 8526 4754 8554
rect 4754 8526 4756 8554
rect 4724 8524 4756 8526
rect 4724 7634 4756 7636
rect 4724 7606 4726 7634
rect 4726 7606 4754 7634
rect 4754 7606 4756 7634
rect 4724 7604 4756 7606
rect 4724 7554 4756 7556
rect 4724 7526 4726 7554
rect 4726 7526 4754 7554
rect 4754 7526 4756 7554
rect 4724 7524 4756 7526
rect 4724 7474 4756 7476
rect 4724 7446 4726 7474
rect 4726 7446 4754 7474
rect 4754 7446 4756 7474
rect 4724 7444 4756 7446
rect 4724 7394 4756 7396
rect 4724 7366 4726 7394
rect 4726 7366 4754 7394
rect 4754 7366 4756 7394
rect 4724 7364 4756 7366
rect 4724 7314 4756 7316
rect 4724 7286 4726 7314
rect 4726 7286 4754 7314
rect 4754 7286 4756 7314
rect 4724 7284 4756 7286
rect 4724 7234 4756 7236
rect 4724 7206 4726 7234
rect 4726 7206 4754 7234
rect 4754 7206 4756 7234
rect 4724 7204 4756 7206
rect 4724 7154 4756 7156
rect 4724 7126 4726 7154
rect 4726 7126 4754 7154
rect 4754 7126 4756 7154
rect 4724 7124 4756 7126
rect 4724 7074 4756 7076
rect 4724 7046 4726 7074
rect 4726 7046 4754 7074
rect 4754 7046 4756 7074
rect 4724 7044 4756 7046
rect 4724 6754 4756 6756
rect 4724 6726 4726 6754
rect 4726 6726 4754 6754
rect 4754 6726 4756 6754
rect 4724 6724 4756 6726
rect 4724 6674 4756 6676
rect 4724 6646 4726 6674
rect 4726 6646 4754 6674
rect 4754 6646 4756 6674
rect 4724 6644 4756 6646
rect 4724 6594 4756 6596
rect 4724 6566 4726 6594
rect 4726 6566 4754 6594
rect 4754 6566 4756 6594
rect 4724 6564 4756 6566
rect 4724 6514 4756 6516
rect 4724 6486 4726 6514
rect 4726 6486 4754 6514
rect 4754 6486 4756 6514
rect 4724 6484 4756 6486
rect 4724 6434 4756 6436
rect 4724 6406 4726 6434
rect 4726 6406 4754 6434
rect 4754 6406 4756 6434
rect 4724 6404 4756 6406
rect 4724 6354 4756 6356
rect 4724 6326 4726 6354
rect 4726 6326 4754 6354
rect 4754 6326 4756 6354
rect 4724 6324 4756 6326
rect 4724 5794 4756 5796
rect 4724 5766 4726 5794
rect 4726 5766 4754 5794
rect 4754 5766 4756 5794
rect 4724 5764 4756 5766
rect 4724 5714 4756 5716
rect 4724 5686 4726 5714
rect 4726 5686 4754 5714
rect 4754 5686 4756 5714
rect 4724 5684 4756 5686
rect 4724 5634 4756 5636
rect 4724 5606 4726 5634
rect 4726 5606 4754 5634
rect 4754 5606 4756 5634
rect 4724 5604 4756 5606
rect 4724 5554 4756 5556
rect 4724 5526 4726 5554
rect 4726 5526 4754 5554
rect 4754 5526 4756 5554
rect 4724 5524 4756 5526
rect 4724 5474 4756 5476
rect 4724 5446 4726 5474
rect 4726 5446 4754 5474
rect 4754 5446 4756 5474
rect 4724 5444 4756 5446
rect 4724 5394 4756 5396
rect 4724 5366 4726 5394
rect 4726 5366 4754 5394
rect 4754 5366 4756 5394
rect 4724 5364 4756 5366
rect 4724 5314 4756 5316
rect 4724 5286 4726 5314
rect 4726 5286 4754 5314
rect 4754 5286 4756 5314
rect 4724 5284 4756 5286
rect 4724 5234 4756 5236
rect 4724 5206 4726 5234
rect 4726 5206 4754 5234
rect 4754 5206 4756 5234
rect 4724 5204 4756 5206
rect 4724 5154 4756 5156
rect 4724 5126 4726 5154
rect 4726 5126 4754 5154
rect 4754 5126 4756 5154
rect 4724 5124 4756 5126
rect 4724 5074 4756 5076
rect 4724 5046 4726 5074
rect 4726 5046 4754 5074
rect 4754 5046 4756 5074
rect 4724 5044 4756 5046
rect 4724 4994 4756 4996
rect 4724 4966 4726 4994
rect 4726 4966 4754 4994
rect 4754 4966 4756 4994
rect 4724 4964 4756 4966
rect 4724 4434 4756 4436
rect 4724 4406 4726 4434
rect 4726 4406 4754 4434
rect 4754 4406 4756 4434
rect 4724 4404 4756 4406
rect 4724 4354 4756 4356
rect 4724 4326 4726 4354
rect 4726 4326 4754 4354
rect 4754 4326 4756 4354
rect 4724 4324 4756 4326
rect 4724 4274 4756 4276
rect 4724 4246 4726 4274
rect 4726 4246 4754 4274
rect 4754 4246 4756 4274
rect 4724 4244 4756 4246
rect 4724 4194 4756 4196
rect 4724 4166 4726 4194
rect 4726 4166 4754 4194
rect 4754 4166 4756 4194
rect 4724 4164 4756 4166
rect 4724 4114 4756 4116
rect 4724 4086 4726 4114
rect 4726 4086 4754 4114
rect 4754 4086 4756 4114
rect 4724 4084 4756 4086
rect 4724 4034 4756 4036
rect 4724 4006 4726 4034
rect 4726 4006 4754 4034
rect 4754 4006 4756 4034
rect 4724 4004 4756 4006
rect 4724 3954 4756 3956
rect 4724 3926 4726 3954
rect 4726 3926 4754 3954
rect 4754 3926 4756 3954
rect 4724 3924 4756 3926
rect 4724 3154 4756 3156
rect 4724 3126 4726 3154
rect 4726 3126 4754 3154
rect 4754 3126 4756 3154
rect 4724 3124 4756 3126
rect 4724 3074 4756 3076
rect 4724 3046 4726 3074
rect 4726 3046 4754 3074
rect 4754 3046 4756 3074
rect 4724 3044 4756 3046
rect 4724 2994 4756 2996
rect 4724 2966 4726 2994
rect 4726 2966 4754 2994
rect 4754 2966 4756 2994
rect 4724 2964 4756 2966
rect 4724 2914 4756 2916
rect 4724 2886 4726 2914
rect 4726 2886 4754 2914
rect 4754 2886 4756 2914
rect 4724 2884 4756 2886
rect 4724 2834 4756 2836
rect 4724 2806 4726 2834
rect 4726 2806 4754 2834
rect 4754 2806 4756 2834
rect 4724 2804 4756 2806
rect 4724 2754 4756 2756
rect 4724 2726 4726 2754
rect 4726 2726 4754 2754
rect 4754 2726 4756 2754
rect 4724 2724 4756 2726
rect 4724 2674 4756 2676
rect 4724 2646 4726 2674
rect 4726 2646 4754 2674
rect 4754 2646 4756 2674
rect 4724 2644 4756 2646
rect 4724 2594 4756 2596
rect 4724 2566 4726 2594
rect 4726 2566 4754 2594
rect 4754 2566 4756 2594
rect 4724 2564 4756 2566
rect 4724 2514 4756 2516
rect 4724 2486 4726 2514
rect 4726 2486 4754 2514
rect 4754 2486 4756 2514
rect 4724 2484 4756 2486
rect 4724 2434 4756 2436
rect 4724 2406 4726 2434
rect 4726 2406 4754 2434
rect 4754 2406 4756 2434
rect 4724 2404 4756 2406
rect 4724 2354 4756 2356
rect 4724 2326 4726 2354
rect 4726 2326 4754 2354
rect 4754 2326 4756 2354
rect 4724 2324 4756 2326
rect 4724 2274 4756 2276
rect 4724 2246 4726 2274
rect 4726 2246 4754 2274
rect 4754 2246 4756 2274
rect 4724 2244 4756 2246
rect 4724 2194 4756 2196
rect 4724 2166 4726 2194
rect 4726 2166 4754 2194
rect 4754 2166 4756 2194
rect 4724 2164 4756 2166
rect 4724 2114 4756 2116
rect 4724 2086 4726 2114
rect 4726 2086 4754 2114
rect 4754 2086 4756 2114
rect 4724 2084 4756 2086
rect 4724 2034 4756 2036
rect 4724 2006 4726 2034
rect 4726 2006 4754 2034
rect 4754 2006 4756 2034
rect 4724 2004 4756 2006
rect 4724 1634 4756 1636
rect 4724 1606 4726 1634
rect 4726 1606 4754 1634
rect 4754 1606 4756 1634
rect 4724 1604 4756 1606
rect 4724 1554 4756 1556
rect 4724 1526 4726 1554
rect 4726 1526 4754 1554
rect 4754 1526 4756 1554
rect 4724 1524 4756 1526
rect 4724 1474 4756 1476
rect 4724 1446 4726 1474
rect 4726 1446 4754 1474
rect 4754 1446 4756 1474
rect 4724 1444 4756 1446
rect 4724 1394 4756 1396
rect 4724 1366 4726 1394
rect 4726 1366 4754 1394
rect 4754 1366 4756 1394
rect 4724 1364 4756 1366
rect 4724 1314 4756 1316
rect 4724 1286 4726 1314
rect 4726 1286 4754 1314
rect 4754 1286 4756 1314
rect 4724 1284 4756 1286
rect 4724 1234 4756 1236
rect 4724 1206 4726 1234
rect 4726 1206 4754 1234
rect 4754 1206 4756 1234
rect 4724 1204 4756 1206
rect 4724 1154 4756 1156
rect 4724 1126 4726 1154
rect 4726 1126 4754 1154
rect 4754 1126 4756 1154
rect 4724 1124 4756 1126
rect 4724 1074 4756 1076
rect 4724 1046 4726 1074
rect 4726 1046 4754 1074
rect 4754 1046 4756 1074
rect 4724 1044 4756 1046
rect 4724 754 4756 756
rect 4724 726 4726 754
rect 4726 726 4754 754
rect 4754 726 4756 754
rect 4724 724 4756 726
rect 4724 674 4756 676
rect 4724 646 4726 674
rect 4726 646 4754 674
rect 4754 646 4756 674
rect 4724 644 4756 646
rect 4724 594 4756 596
rect 4724 566 4726 594
rect 4726 566 4754 594
rect 4754 566 4756 594
rect 4724 564 4756 566
rect 4724 194 4756 196
rect 4724 166 4726 194
rect 4726 166 4754 194
rect 4754 166 4756 194
rect 4724 164 4756 166
rect 4724 114 4756 116
rect 4724 86 4726 114
rect 4726 86 4754 114
rect 4754 86 4756 114
rect 4724 84 4756 86
rect 4724 34 4756 36
rect 4724 6 4726 34
rect 4726 6 4754 34
rect 4754 6 4756 34
rect 4724 4 4756 6
rect 5044 13364 5076 13396
rect 5044 13324 5076 13356
rect 5044 13284 5076 13316
rect 5044 13244 5076 13276
rect 5044 13204 5076 13236
rect 4884 12634 4916 12636
rect 4884 12606 4886 12634
rect 4886 12606 4914 12634
rect 4914 12606 4916 12634
rect 4884 12604 4916 12606
rect 4884 12554 4916 12556
rect 4884 12526 4886 12554
rect 4886 12526 4914 12554
rect 4914 12526 4916 12554
rect 4884 12524 4916 12526
rect 4884 12474 4916 12476
rect 4884 12446 4886 12474
rect 4886 12446 4914 12474
rect 4914 12446 4916 12474
rect 4884 12444 4916 12446
rect 4884 12394 4916 12396
rect 4884 12366 4886 12394
rect 4886 12366 4914 12394
rect 4914 12366 4916 12394
rect 4884 12364 4916 12366
rect 4884 12314 4916 12316
rect 4884 12286 4886 12314
rect 4886 12286 4914 12314
rect 4914 12286 4916 12314
rect 4884 12284 4916 12286
rect 4884 12234 4916 12236
rect 4884 12206 4886 12234
rect 4886 12206 4914 12234
rect 4914 12206 4916 12234
rect 4884 12204 4916 12206
rect 4884 12154 4916 12156
rect 4884 12126 4886 12154
rect 4886 12126 4914 12154
rect 4914 12126 4916 12154
rect 4884 12124 4916 12126
rect 4884 11834 4916 11836
rect 4884 11806 4886 11834
rect 4886 11806 4914 11834
rect 4914 11806 4916 11834
rect 4884 11804 4916 11806
rect 4884 11754 4916 11756
rect 4884 11726 4886 11754
rect 4886 11726 4914 11754
rect 4914 11726 4916 11754
rect 4884 11724 4916 11726
rect 4884 11674 4916 11676
rect 4884 11646 4886 11674
rect 4886 11646 4914 11674
rect 4914 11646 4916 11674
rect 4884 11644 4916 11646
rect 4884 11594 4916 11596
rect 4884 11566 4886 11594
rect 4886 11566 4914 11594
rect 4914 11566 4916 11594
rect 4884 11564 4916 11566
rect 4884 11514 4916 11516
rect 4884 11486 4886 11514
rect 4886 11486 4914 11514
rect 4914 11486 4916 11514
rect 4884 11484 4916 11486
rect 4884 11434 4916 11436
rect 4884 11406 4886 11434
rect 4886 11406 4914 11434
rect 4914 11406 4916 11434
rect 4884 11404 4916 11406
rect 4884 10874 4916 10876
rect 4884 10846 4886 10874
rect 4886 10846 4914 10874
rect 4914 10846 4916 10874
rect 4884 10844 4916 10846
rect 4884 10794 4916 10796
rect 4884 10766 4886 10794
rect 4886 10766 4914 10794
rect 4914 10766 4916 10794
rect 4884 10764 4916 10766
rect 4884 10714 4916 10716
rect 4884 10686 4886 10714
rect 4886 10686 4914 10714
rect 4914 10686 4916 10714
rect 4884 10684 4916 10686
rect 4884 10634 4916 10636
rect 4884 10606 4886 10634
rect 4886 10606 4914 10634
rect 4914 10606 4916 10634
rect 4884 10604 4916 10606
rect 4884 10554 4916 10556
rect 4884 10526 4886 10554
rect 4886 10526 4914 10554
rect 4914 10526 4916 10554
rect 4884 10524 4916 10526
rect 4884 10474 4916 10476
rect 4884 10446 4886 10474
rect 4886 10446 4914 10474
rect 4914 10446 4916 10474
rect 4884 10444 4916 10446
rect 4884 10394 4916 10396
rect 4884 10366 4886 10394
rect 4886 10366 4914 10394
rect 4914 10366 4916 10394
rect 4884 10364 4916 10366
rect 4884 10314 4916 10316
rect 4884 10286 4886 10314
rect 4886 10286 4914 10314
rect 4914 10286 4916 10314
rect 4884 10284 4916 10286
rect 4884 10234 4916 10236
rect 4884 10206 4886 10234
rect 4886 10206 4914 10234
rect 4914 10206 4916 10234
rect 4884 10204 4916 10206
rect 4884 10154 4916 10156
rect 4884 10126 4886 10154
rect 4886 10126 4914 10154
rect 4914 10126 4916 10154
rect 4884 10124 4916 10126
rect 4884 10074 4916 10076
rect 4884 10046 4886 10074
rect 4886 10046 4914 10074
rect 4914 10046 4916 10074
rect 4884 10044 4916 10046
rect 4884 9994 4916 9996
rect 4884 9966 4886 9994
rect 4886 9966 4914 9994
rect 4914 9966 4916 9994
rect 4884 9964 4916 9966
rect 4884 9914 4916 9916
rect 4884 9886 4886 9914
rect 4886 9886 4914 9914
rect 4914 9886 4916 9914
rect 4884 9884 4916 9886
rect 4884 9834 4916 9836
rect 4884 9806 4886 9834
rect 4886 9806 4914 9834
rect 4914 9806 4916 9834
rect 4884 9804 4916 9806
rect 4884 9754 4916 9756
rect 4884 9726 4886 9754
rect 4886 9726 4914 9754
rect 4914 9726 4916 9754
rect 4884 9724 4916 9726
rect 4884 9354 4916 9356
rect 4884 9326 4886 9354
rect 4886 9326 4914 9354
rect 4914 9326 4916 9354
rect 4884 9324 4916 9326
rect 4884 9274 4916 9276
rect 4884 9246 4886 9274
rect 4886 9246 4914 9274
rect 4914 9246 4916 9274
rect 4884 9244 4916 9246
rect 4884 9194 4916 9196
rect 4884 9166 4886 9194
rect 4886 9166 4914 9194
rect 4914 9166 4916 9194
rect 4884 9164 4916 9166
rect 4884 8874 4916 8876
rect 4884 8846 4886 8874
rect 4886 8846 4914 8874
rect 4914 8846 4916 8874
rect 4884 8844 4916 8846
rect 4884 8794 4916 8796
rect 4884 8766 4886 8794
rect 4886 8766 4914 8794
rect 4914 8766 4916 8794
rect 4884 8764 4916 8766
rect 4884 8714 4916 8716
rect 4884 8686 4886 8714
rect 4886 8686 4914 8714
rect 4914 8686 4916 8714
rect 4884 8684 4916 8686
rect 4884 8634 4916 8636
rect 4884 8606 4886 8634
rect 4886 8606 4914 8634
rect 4914 8606 4916 8634
rect 4884 8604 4916 8606
rect 4884 8554 4916 8556
rect 4884 8526 4886 8554
rect 4886 8526 4914 8554
rect 4914 8526 4916 8554
rect 4884 8524 4916 8526
rect 4884 7634 4916 7636
rect 4884 7606 4886 7634
rect 4886 7606 4914 7634
rect 4914 7606 4916 7634
rect 4884 7604 4916 7606
rect 4884 7554 4916 7556
rect 4884 7526 4886 7554
rect 4886 7526 4914 7554
rect 4914 7526 4916 7554
rect 4884 7524 4916 7526
rect 4884 7474 4916 7476
rect 4884 7446 4886 7474
rect 4886 7446 4914 7474
rect 4914 7446 4916 7474
rect 4884 7444 4916 7446
rect 4884 7394 4916 7396
rect 4884 7366 4886 7394
rect 4886 7366 4914 7394
rect 4914 7366 4916 7394
rect 4884 7364 4916 7366
rect 4884 7314 4916 7316
rect 4884 7286 4886 7314
rect 4886 7286 4914 7314
rect 4914 7286 4916 7314
rect 4884 7284 4916 7286
rect 4884 7234 4916 7236
rect 4884 7206 4886 7234
rect 4886 7206 4914 7234
rect 4914 7206 4916 7234
rect 4884 7204 4916 7206
rect 4884 7154 4916 7156
rect 4884 7126 4886 7154
rect 4886 7126 4914 7154
rect 4914 7126 4916 7154
rect 4884 7124 4916 7126
rect 4884 7074 4916 7076
rect 4884 7046 4886 7074
rect 4886 7046 4914 7074
rect 4914 7046 4916 7074
rect 4884 7044 4916 7046
rect 4884 6754 4916 6756
rect 4884 6726 4886 6754
rect 4886 6726 4914 6754
rect 4914 6726 4916 6754
rect 4884 6724 4916 6726
rect 4884 6674 4916 6676
rect 4884 6646 4886 6674
rect 4886 6646 4914 6674
rect 4914 6646 4916 6674
rect 4884 6644 4916 6646
rect 4884 6594 4916 6596
rect 4884 6566 4886 6594
rect 4886 6566 4914 6594
rect 4914 6566 4916 6594
rect 4884 6564 4916 6566
rect 4884 6514 4916 6516
rect 4884 6486 4886 6514
rect 4886 6486 4914 6514
rect 4914 6486 4916 6514
rect 4884 6484 4916 6486
rect 4884 6434 4916 6436
rect 4884 6406 4886 6434
rect 4886 6406 4914 6434
rect 4914 6406 4916 6434
rect 4884 6404 4916 6406
rect 4884 6354 4916 6356
rect 4884 6326 4886 6354
rect 4886 6326 4914 6354
rect 4914 6326 4916 6354
rect 4884 6324 4916 6326
rect 4884 5794 4916 5796
rect 4884 5766 4886 5794
rect 4886 5766 4914 5794
rect 4914 5766 4916 5794
rect 4884 5764 4916 5766
rect 4884 5714 4916 5716
rect 4884 5686 4886 5714
rect 4886 5686 4914 5714
rect 4914 5686 4916 5714
rect 4884 5684 4916 5686
rect 4884 5634 4916 5636
rect 4884 5606 4886 5634
rect 4886 5606 4914 5634
rect 4914 5606 4916 5634
rect 4884 5604 4916 5606
rect 4884 5554 4916 5556
rect 4884 5526 4886 5554
rect 4886 5526 4914 5554
rect 4914 5526 4916 5554
rect 4884 5524 4916 5526
rect 4884 5474 4916 5476
rect 4884 5446 4886 5474
rect 4886 5446 4914 5474
rect 4914 5446 4916 5474
rect 4884 5444 4916 5446
rect 4884 5394 4916 5396
rect 4884 5366 4886 5394
rect 4886 5366 4914 5394
rect 4914 5366 4916 5394
rect 4884 5364 4916 5366
rect 4884 5314 4916 5316
rect 4884 5286 4886 5314
rect 4886 5286 4914 5314
rect 4914 5286 4916 5314
rect 4884 5284 4916 5286
rect 4884 5234 4916 5236
rect 4884 5206 4886 5234
rect 4886 5206 4914 5234
rect 4914 5206 4916 5234
rect 4884 5204 4916 5206
rect 4884 5154 4916 5156
rect 4884 5126 4886 5154
rect 4886 5126 4914 5154
rect 4914 5126 4916 5154
rect 4884 5124 4916 5126
rect 4884 5074 4916 5076
rect 4884 5046 4886 5074
rect 4886 5046 4914 5074
rect 4914 5046 4916 5074
rect 4884 5044 4916 5046
rect 4884 4994 4916 4996
rect 4884 4966 4886 4994
rect 4886 4966 4914 4994
rect 4914 4966 4916 4994
rect 4884 4964 4916 4966
rect 4884 4434 4916 4436
rect 4884 4406 4886 4434
rect 4886 4406 4914 4434
rect 4914 4406 4916 4434
rect 4884 4404 4916 4406
rect 4884 4354 4916 4356
rect 4884 4326 4886 4354
rect 4886 4326 4914 4354
rect 4914 4326 4916 4354
rect 4884 4324 4916 4326
rect 4884 4274 4916 4276
rect 4884 4246 4886 4274
rect 4886 4246 4914 4274
rect 4914 4246 4916 4274
rect 4884 4244 4916 4246
rect 4884 4194 4916 4196
rect 4884 4166 4886 4194
rect 4886 4166 4914 4194
rect 4914 4166 4916 4194
rect 4884 4164 4916 4166
rect 4884 4114 4916 4116
rect 4884 4086 4886 4114
rect 4886 4086 4914 4114
rect 4914 4086 4916 4114
rect 4884 4084 4916 4086
rect 4884 4034 4916 4036
rect 4884 4006 4886 4034
rect 4886 4006 4914 4034
rect 4914 4006 4916 4034
rect 4884 4004 4916 4006
rect 4884 3954 4916 3956
rect 4884 3926 4886 3954
rect 4886 3926 4914 3954
rect 4914 3926 4916 3954
rect 4884 3924 4916 3926
rect 4884 3154 4916 3156
rect 4884 3126 4886 3154
rect 4886 3126 4914 3154
rect 4914 3126 4916 3154
rect 4884 3124 4916 3126
rect 4884 3074 4916 3076
rect 4884 3046 4886 3074
rect 4886 3046 4914 3074
rect 4914 3046 4916 3074
rect 4884 3044 4916 3046
rect 4884 2994 4916 2996
rect 4884 2966 4886 2994
rect 4886 2966 4914 2994
rect 4914 2966 4916 2994
rect 4884 2964 4916 2966
rect 4884 2914 4916 2916
rect 4884 2886 4886 2914
rect 4886 2886 4914 2914
rect 4914 2886 4916 2914
rect 4884 2884 4916 2886
rect 4884 2834 4916 2836
rect 4884 2806 4886 2834
rect 4886 2806 4914 2834
rect 4914 2806 4916 2834
rect 4884 2804 4916 2806
rect 4884 2754 4916 2756
rect 4884 2726 4886 2754
rect 4886 2726 4914 2754
rect 4914 2726 4916 2754
rect 4884 2724 4916 2726
rect 4884 2674 4916 2676
rect 4884 2646 4886 2674
rect 4886 2646 4914 2674
rect 4914 2646 4916 2674
rect 4884 2644 4916 2646
rect 4884 2594 4916 2596
rect 4884 2566 4886 2594
rect 4886 2566 4914 2594
rect 4914 2566 4916 2594
rect 4884 2564 4916 2566
rect 4884 2514 4916 2516
rect 4884 2486 4886 2514
rect 4886 2486 4914 2514
rect 4914 2486 4916 2514
rect 4884 2484 4916 2486
rect 4884 2434 4916 2436
rect 4884 2406 4886 2434
rect 4886 2406 4914 2434
rect 4914 2406 4916 2434
rect 4884 2404 4916 2406
rect 4884 2354 4916 2356
rect 4884 2326 4886 2354
rect 4886 2326 4914 2354
rect 4914 2326 4916 2354
rect 4884 2324 4916 2326
rect 4884 2274 4916 2276
rect 4884 2246 4886 2274
rect 4886 2246 4914 2274
rect 4914 2246 4916 2274
rect 4884 2244 4916 2246
rect 4884 2194 4916 2196
rect 4884 2166 4886 2194
rect 4886 2166 4914 2194
rect 4914 2166 4916 2194
rect 4884 2164 4916 2166
rect 4884 2114 4916 2116
rect 4884 2086 4886 2114
rect 4886 2086 4914 2114
rect 4914 2086 4916 2114
rect 4884 2084 4916 2086
rect 4884 2034 4916 2036
rect 4884 2006 4886 2034
rect 4886 2006 4914 2034
rect 4914 2006 4916 2034
rect 4884 2004 4916 2006
rect 4884 1634 4916 1636
rect 4884 1606 4886 1634
rect 4886 1606 4914 1634
rect 4914 1606 4916 1634
rect 4884 1604 4916 1606
rect 4884 1554 4916 1556
rect 4884 1526 4886 1554
rect 4886 1526 4914 1554
rect 4914 1526 4916 1554
rect 4884 1524 4916 1526
rect 4884 1474 4916 1476
rect 4884 1446 4886 1474
rect 4886 1446 4914 1474
rect 4914 1446 4916 1474
rect 4884 1444 4916 1446
rect 4884 1394 4916 1396
rect 4884 1366 4886 1394
rect 4886 1366 4914 1394
rect 4914 1366 4916 1394
rect 4884 1364 4916 1366
rect 4884 1314 4916 1316
rect 4884 1286 4886 1314
rect 4886 1286 4914 1314
rect 4914 1286 4916 1314
rect 4884 1284 4916 1286
rect 4884 1234 4916 1236
rect 4884 1206 4886 1234
rect 4886 1206 4914 1234
rect 4914 1206 4916 1234
rect 4884 1204 4916 1206
rect 4884 1154 4916 1156
rect 4884 1126 4886 1154
rect 4886 1126 4914 1154
rect 4914 1126 4916 1154
rect 4884 1124 4916 1126
rect 4884 1074 4916 1076
rect 4884 1046 4886 1074
rect 4886 1046 4914 1074
rect 4914 1046 4916 1074
rect 4884 1044 4916 1046
rect 4884 754 4916 756
rect 4884 726 4886 754
rect 4886 726 4914 754
rect 4914 726 4916 754
rect 4884 724 4916 726
rect 4884 674 4916 676
rect 4884 646 4886 674
rect 4886 646 4914 674
rect 4914 646 4916 674
rect 4884 644 4916 646
rect 4884 594 4916 596
rect 4884 566 4886 594
rect 4886 566 4914 594
rect 4914 566 4916 594
rect 4884 564 4916 566
rect 4884 194 4916 196
rect 4884 166 4886 194
rect 4886 166 4914 194
rect 4914 166 4916 194
rect 4884 164 4916 166
rect 4884 114 4916 116
rect 4884 86 4886 114
rect 4886 86 4914 114
rect 4914 86 4916 114
rect 4884 84 4916 86
rect 4884 34 4916 36
rect 4884 6 4886 34
rect 4886 6 4914 34
rect 4914 6 4916 34
rect 4884 4 4916 6
rect 5044 12634 5076 12636
rect 5044 12606 5046 12634
rect 5046 12606 5074 12634
rect 5074 12606 5076 12634
rect 5044 12604 5076 12606
rect 5044 12554 5076 12556
rect 5044 12526 5046 12554
rect 5046 12526 5074 12554
rect 5074 12526 5076 12554
rect 5044 12524 5076 12526
rect 5044 12474 5076 12476
rect 5044 12446 5046 12474
rect 5046 12446 5074 12474
rect 5074 12446 5076 12474
rect 5044 12444 5076 12446
rect 5044 12394 5076 12396
rect 5044 12366 5046 12394
rect 5046 12366 5074 12394
rect 5074 12366 5076 12394
rect 5044 12364 5076 12366
rect 5044 12314 5076 12316
rect 5044 12286 5046 12314
rect 5046 12286 5074 12314
rect 5074 12286 5076 12314
rect 5044 12284 5076 12286
rect 5044 12234 5076 12236
rect 5044 12206 5046 12234
rect 5046 12206 5074 12234
rect 5074 12206 5076 12234
rect 5044 12204 5076 12206
rect 5044 12154 5076 12156
rect 5044 12126 5046 12154
rect 5046 12126 5074 12154
rect 5074 12126 5076 12154
rect 5044 12124 5076 12126
rect 5044 11834 5076 11836
rect 5044 11806 5046 11834
rect 5046 11806 5074 11834
rect 5074 11806 5076 11834
rect 5044 11804 5076 11806
rect 5044 11754 5076 11756
rect 5044 11726 5046 11754
rect 5046 11726 5074 11754
rect 5074 11726 5076 11754
rect 5044 11724 5076 11726
rect 5044 11674 5076 11676
rect 5044 11646 5046 11674
rect 5046 11646 5074 11674
rect 5074 11646 5076 11674
rect 5044 11644 5076 11646
rect 5044 11594 5076 11596
rect 5044 11566 5046 11594
rect 5046 11566 5074 11594
rect 5074 11566 5076 11594
rect 5044 11564 5076 11566
rect 5044 11514 5076 11516
rect 5044 11486 5046 11514
rect 5046 11486 5074 11514
rect 5074 11486 5076 11514
rect 5044 11484 5076 11486
rect 5044 11434 5076 11436
rect 5044 11406 5046 11434
rect 5046 11406 5074 11434
rect 5074 11406 5076 11434
rect 5044 11404 5076 11406
rect 5044 10874 5076 10876
rect 5044 10846 5046 10874
rect 5046 10846 5074 10874
rect 5074 10846 5076 10874
rect 5044 10844 5076 10846
rect 5044 10794 5076 10796
rect 5044 10766 5046 10794
rect 5046 10766 5074 10794
rect 5074 10766 5076 10794
rect 5044 10764 5076 10766
rect 5044 10714 5076 10716
rect 5044 10686 5046 10714
rect 5046 10686 5074 10714
rect 5074 10686 5076 10714
rect 5044 10684 5076 10686
rect 5044 10634 5076 10636
rect 5044 10606 5046 10634
rect 5046 10606 5074 10634
rect 5074 10606 5076 10634
rect 5044 10604 5076 10606
rect 5044 10554 5076 10556
rect 5044 10526 5046 10554
rect 5046 10526 5074 10554
rect 5074 10526 5076 10554
rect 5044 10524 5076 10526
rect 5044 10474 5076 10476
rect 5044 10446 5046 10474
rect 5046 10446 5074 10474
rect 5074 10446 5076 10474
rect 5044 10444 5076 10446
rect 5044 10394 5076 10396
rect 5044 10366 5046 10394
rect 5046 10366 5074 10394
rect 5074 10366 5076 10394
rect 5044 10364 5076 10366
rect 5044 10314 5076 10316
rect 5044 10286 5046 10314
rect 5046 10286 5074 10314
rect 5074 10286 5076 10314
rect 5044 10284 5076 10286
rect 5044 10234 5076 10236
rect 5044 10206 5046 10234
rect 5046 10206 5074 10234
rect 5074 10206 5076 10234
rect 5044 10204 5076 10206
rect 5044 10154 5076 10156
rect 5044 10126 5046 10154
rect 5046 10126 5074 10154
rect 5074 10126 5076 10154
rect 5044 10124 5076 10126
rect 5044 10074 5076 10076
rect 5044 10046 5046 10074
rect 5046 10046 5074 10074
rect 5074 10046 5076 10074
rect 5044 10044 5076 10046
rect 5044 9994 5076 9996
rect 5044 9966 5046 9994
rect 5046 9966 5074 9994
rect 5074 9966 5076 9994
rect 5044 9964 5076 9966
rect 5044 9914 5076 9916
rect 5044 9886 5046 9914
rect 5046 9886 5074 9914
rect 5074 9886 5076 9914
rect 5044 9884 5076 9886
rect 5044 9834 5076 9836
rect 5044 9806 5046 9834
rect 5046 9806 5074 9834
rect 5074 9806 5076 9834
rect 5044 9804 5076 9806
rect 5044 9754 5076 9756
rect 5044 9726 5046 9754
rect 5046 9726 5074 9754
rect 5074 9726 5076 9754
rect 5044 9724 5076 9726
rect 5044 9354 5076 9356
rect 5044 9326 5046 9354
rect 5046 9326 5074 9354
rect 5074 9326 5076 9354
rect 5044 9324 5076 9326
rect 5044 9274 5076 9276
rect 5044 9246 5046 9274
rect 5046 9246 5074 9274
rect 5074 9246 5076 9274
rect 5044 9244 5076 9246
rect 5044 9194 5076 9196
rect 5044 9166 5046 9194
rect 5046 9166 5074 9194
rect 5074 9166 5076 9194
rect 5044 9164 5076 9166
rect 5044 8874 5076 8876
rect 5044 8846 5046 8874
rect 5046 8846 5074 8874
rect 5074 8846 5076 8874
rect 5044 8844 5076 8846
rect 5044 8794 5076 8796
rect 5044 8766 5046 8794
rect 5046 8766 5074 8794
rect 5074 8766 5076 8794
rect 5044 8764 5076 8766
rect 5044 8714 5076 8716
rect 5044 8686 5046 8714
rect 5046 8686 5074 8714
rect 5074 8686 5076 8714
rect 5044 8684 5076 8686
rect 5044 8634 5076 8636
rect 5044 8606 5046 8634
rect 5046 8606 5074 8634
rect 5074 8606 5076 8634
rect 5044 8604 5076 8606
rect 5044 8554 5076 8556
rect 5044 8526 5046 8554
rect 5046 8526 5074 8554
rect 5074 8526 5076 8554
rect 5044 8524 5076 8526
rect 5044 7634 5076 7636
rect 5044 7606 5046 7634
rect 5046 7606 5074 7634
rect 5074 7606 5076 7634
rect 5044 7604 5076 7606
rect 5044 7554 5076 7556
rect 5044 7526 5046 7554
rect 5046 7526 5074 7554
rect 5074 7526 5076 7554
rect 5044 7524 5076 7526
rect 5044 7474 5076 7476
rect 5044 7446 5046 7474
rect 5046 7446 5074 7474
rect 5074 7446 5076 7474
rect 5044 7444 5076 7446
rect 5044 7394 5076 7396
rect 5044 7366 5046 7394
rect 5046 7366 5074 7394
rect 5074 7366 5076 7394
rect 5044 7364 5076 7366
rect 5044 7314 5076 7316
rect 5044 7286 5046 7314
rect 5046 7286 5074 7314
rect 5074 7286 5076 7314
rect 5044 7284 5076 7286
rect 5044 7234 5076 7236
rect 5044 7206 5046 7234
rect 5046 7206 5074 7234
rect 5074 7206 5076 7234
rect 5044 7204 5076 7206
rect 5044 7154 5076 7156
rect 5044 7126 5046 7154
rect 5046 7126 5074 7154
rect 5074 7126 5076 7154
rect 5044 7124 5076 7126
rect 5044 7074 5076 7076
rect 5044 7046 5046 7074
rect 5046 7046 5074 7074
rect 5074 7046 5076 7074
rect 5044 7044 5076 7046
rect 5044 6754 5076 6756
rect 5044 6726 5046 6754
rect 5046 6726 5074 6754
rect 5074 6726 5076 6754
rect 5044 6724 5076 6726
rect 5044 6674 5076 6676
rect 5044 6646 5046 6674
rect 5046 6646 5074 6674
rect 5074 6646 5076 6674
rect 5044 6644 5076 6646
rect 5044 6594 5076 6596
rect 5044 6566 5046 6594
rect 5046 6566 5074 6594
rect 5074 6566 5076 6594
rect 5044 6564 5076 6566
rect 5044 6514 5076 6516
rect 5044 6486 5046 6514
rect 5046 6486 5074 6514
rect 5074 6486 5076 6514
rect 5044 6484 5076 6486
rect 5044 6434 5076 6436
rect 5044 6406 5046 6434
rect 5046 6406 5074 6434
rect 5074 6406 5076 6434
rect 5044 6404 5076 6406
rect 5044 6354 5076 6356
rect 5044 6326 5046 6354
rect 5046 6326 5074 6354
rect 5074 6326 5076 6354
rect 5044 6324 5076 6326
rect 5044 5794 5076 5796
rect 5044 5766 5046 5794
rect 5046 5766 5074 5794
rect 5074 5766 5076 5794
rect 5044 5764 5076 5766
rect 5044 5714 5076 5716
rect 5044 5686 5046 5714
rect 5046 5686 5074 5714
rect 5074 5686 5076 5714
rect 5044 5684 5076 5686
rect 5044 5634 5076 5636
rect 5044 5606 5046 5634
rect 5046 5606 5074 5634
rect 5074 5606 5076 5634
rect 5044 5604 5076 5606
rect 5044 5554 5076 5556
rect 5044 5526 5046 5554
rect 5046 5526 5074 5554
rect 5074 5526 5076 5554
rect 5044 5524 5076 5526
rect 5044 5474 5076 5476
rect 5044 5446 5046 5474
rect 5046 5446 5074 5474
rect 5074 5446 5076 5474
rect 5044 5444 5076 5446
rect 5044 5394 5076 5396
rect 5044 5366 5046 5394
rect 5046 5366 5074 5394
rect 5074 5366 5076 5394
rect 5044 5364 5076 5366
rect 5044 5314 5076 5316
rect 5044 5286 5046 5314
rect 5046 5286 5074 5314
rect 5074 5286 5076 5314
rect 5044 5284 5076 5286
rect 5044 5234 5076 5236
rect 5044 5206 5046 5234
rect 5046 5206 5074 5234
rect 5074 5206 5076 5234
rect 5044 5204 5076 5206
rect 5044 5154 5076 5156
rect 5044 5126 5046 5154
rect 5046 5126 5074 5154
rect 5074 5126 5076 5154
rect 5044 5124 5076 5126
rect 5044 5074 5076 5076
rect 5044 5046 5046 5074
rect 5046 5046 5074 5074
rect 5074 5046 5076 5074
rect 5044 5044 5076 5046
rect 5044 4994 5076 4996
rect 5044 4966 5046 4994
rect 5046 4966 5074 4994
rect 5074 4966 5076 4994
rect 5044 4964 5076 4966
rect 5044 4434 5076 4436
rect 5044 4406 5046 4434
rect 5046 4406 5074 4434
rect 5074 4406 5076 4434
rect 5044 4404 5076 4406
rect 5044 4354 5076 4356
rect 5044 4326 5046 4354
rect 5046 4326 5074 4354
rect 5074 4326 5076 4354
rect 5044 4324 5076 4326
rect 5044 4274 5076 4276
rect 5044 4246 5046 4274
rect 5046 4246 5074 4274
rect 5074 4246 5076 4274
rect 5044 4244 5076 4246
rect 5044 4194 5076 4196
rect 5044 4166 5046 4194
rect 5046 4166 5074 4194
rect 5074 4166 5076 4194
rect 5044 4164 5076 4166
rect 5044 4114 5076 4116
rect 5044 4086 5046 4114
rect 5046 4086 5074 4114
rect 5074 4086 5076 4114
rect 5044 4084 5076 4086
rect 5044 4034 5076 4036
rect 5044 4006 5046 4034
rect 5046 4006 5074 4034
rect 5074 4006 5076 4034
rect 5044 4004 5076 4006
rect 5044 3954 5076 3956
rect 5044 3926 5046 3954
rect 5046 3926 5074 3954
rect 5074 3926 5076 3954
rect 5044 3924 5076 3926
rect 5044 3154 5076 3156
rect 5044 3126 5046 3154
rect 5046 3126 5074 3154
rect 5074 3126 5076 3154
rect 5044 3124 5076 3126
rect 5044 3074 5076 3076
rect 5044 3046 5046 3074
rect 5046 3046 5074 3074
rect 5074 3046 5076 3074
rect 5044 3044 5076 3046
rect 5044 2994 5076 2996
rect 5044 2966 5046 2994
rect 5046 2966 5074 2994
rect 5074 2966 5076 2994
rect 5044 2964 5076 2966
rect 5044 2914 5076 2916
rect 5044 2886 5046 2914
rect 5046 2886 5074 2914
rect 5074 2886 5076 2914
rect 5044 2884 5076 2886
rect 5044 2834 5076 2836
rect 5044 2806 5046 2834
rect 5046 2806 5074 2834
rect 5074 2806 5076 2834
rect 5044 2804 5076 2806
rect 5044 2754 5076 2756
rect 5044 2726 5046 2754
rect 5046 2726 5074 2754
rect 5074 2726 5076 2754
rect 5044 2724 5076 2726
rect 5044 2674 5076 2676
rect 5044 2646 5046 2674
rect 5046 2646 5074 2674
rect 5074 2646 5076 2674
rect 5044 2644 5076 2646
rect 5044 2594 5076 2596
rect 5044 2566 5046 2594
rect 5046 2566 5074 2594
rect 5074 2566 5076 2594
rect 5044 2564 5076 2566
rect 5044 2514 5076 2516
rect 5044 2486 5046 2514
rect 5046 2486 5074 2514
rect 5074 2486 5076 2514
rect 5044 2484 5076 2486
rect 5044 2434 5076 2436
rect 5044 2406 5046 2434
rect 5046 2406 5074 2434
rect 5074 2406 5076 2434
rect 5044 2404 5076 2406
rect 5044 2354 5076 2356
rect 5044 2326 5046 2354
rect 5046 2326 5074 2354
rect 5074 2326 5076 2354
rect 5044 2324 5076 2326
rect 5044 2274 5076 2276
rect 5044 2246 5046 2274
rect 5046 2246 5074 2274
rect 5074 2246 5076 2274
rect 5044 2244 5076 2246
rect 5044 2194 5076 2196
rect 5044 2166 5046 2194
rect 5046 2166 5074 2194
rect 5074 2166 5076 2194
rect 5044 2164 5076 2166
rect 5044 2114 5076 2116
rect 5044 2086 5046 2114
rect 5046 2086 5074 2114
rect 5074 2086 5076 2114
rect 5044 2084 5076 2086
rect 5044 2034 5076 2036
rect 5044 2006 5046 2034
rect 5046 2006 5074 2034
rect 5074 2006 5076 2034
rect 5044 2004 5076 2006
rect 5044 1634 5076 1636
rect 5044 1606 5046 1634
rect 5046 1606 5074 1634
rect 5074 1606 5076 1634
rect 5044 1604 5076 1606
rect 5044 1554 5076 1556
rect 5044 1526 5046 1554
rect 5046 1526 5074 1554
rect 5074 1526 5076 1554
rect 5044 1524 5076 1526
rect 5044 1474 5076 1476
rect 5044 1446 5046 1474
rect 5046 1446 5074 1474
rect 5074 1446 5076 1474
rect 5044 1444 5076 1446
rect 5044 1394 5076 1396
rect 5044 1366 5046 1394
rect 5046 1366 5074 1394
rect 5074 1366 5076 1394
rect 5044 1364 5076 1366
rect 5044 1314 5076 1316
rect 5044 1286 5046 1314
rect 5046 1286 5074 1314
rect 5074 1286 5076 1314
rect 5044 1284 5076 1286
rect 5044 1234 5076 1236
rect 5044 1206 5046 1234
rect 5046 1206 5074 1234
rect 5074 1206 5076 1234
rect 5044 1204 5076 1206
rect 5044 1154 5076 1156
rect 5044 1126 5046 1154
rect 5046 1126 5074 1154
rect 5074 1126 5076 1154
rect 5044 1124 5076 1126
rect 5044 1074 5076 1076
rect 5044 1046 5046 1074
rect 5046 1046 5074 1074
rect 5074 1046 5076 1074
rect 5044 1044 5076 1046
rect 5044 754 5076 756
rect 5044 726 5046 754
rect 5046 726 5074 754
rect 5074 726 5076 754
rect 5044 724 5076 726
rect 5044 674 5076 676
rect 5044 646 5046 674
rect 5046 646 5074 674
rect 5074 646 5076 674
rect 5044 644 5076 646
rect 5044 594 5076 596
rect 5044 566 5046 594
rect 5046 566 5074 594
rect 5074 566 5076 594
rect 5044 564 5076 566
rect 5044 194 5076 196
rect 5044 166 5046 194
rect 5046 166 5074 194
rect 5074 166 5076 194
rect 5044 164 5076 166
rect 5044 114 5076 116
rect 5044 86 5046 114
rect 5046 86 5074 114
rect 5074 86 5076 114
rect 5044 84 5076 86
rect 5044 34 5076 36
rect 5044 6 5046 34
rect 5046 6 5074 34
rect 5074 6 5076 34
rect 5044 4 5076 6
rect 5124 15364 5156 15396
rect 5124 14084 5156 14116
rect 5124 12634 5156 12636
rect 5124 12606 5126 12634
rect 5126 12606 5154 12634
rect 5154 12606 5156 12634
rect 5124 12604 5156 12606
rect 5124 12554 5156 12556
rect 5124 12526 5126 12554
rect 5126 12526 5154 12554
rect 5154 12526 5156 12554
rect 5124 12524 5156 12526
rect 5124 12474 5156 12476
rect 5124 12446 5126 12474
rect 5126 12446 5154 12474
rect 5154 12446 5156 12474
rect 5124 12444 5156 12446
rect 5124 12394 5156 12396
rect 5124 12366 5126 12394
rect 5126 12366 5154 12394
rect 5154 12366 5156 12394
rect 5124 12364 5156 12366
rect 5124 12314 5156 12316
rect 5124 12286 5126 12314
rect 5126 12286 5154 12314
rect 5154 12286 5156 12314
rect 5124 12284 5156 12286
rect 5124 12234 5156 12236
rect 5124 12206 5126 12234
rect 5126 12206 5154 12234
rect 5154 12206 5156 12234
rect 5124 12204 5156 12206
rect 5124 12154 5156 12156
rect 5124 12126 5126 12154
rect 5126 12126 5154 12154
rect 5154 12126 5156 12154
rect 5124 12124 5156 12126
rect 5124 11834 5156 11836
rect 5124 11806 5126 11834
rect 5126 11806 5154 11834
rect 5154 11806 5156 11834
rect 5124 11804 5156 11806
rect 5124 11754 5156 11756
rect 5124 11726 5126 11754
rect 5126 11726 5154 11754
rect 5154 11726 5156 11754
rect 5124 11724 5156 11726
rect 5124 11674 5156 11676
rect 5124 11646 5126 11674
rect 5126 11646 5154 11674
rect 5154 11646 5156 11674
rect 5124 11644 5156 11646
rect 5124 11594 5156 11596
rect 5124 11566 5126 11594
rect 5126 11566 5154 11594
rect 5154 11566 5156 11594
rect 5124 11564 5156 11566
rect 5124 11514 5156 11516
rect 5124 11486 5126 11514
rect 5126 11486 5154 11514
rect 5154 11486 5156 11514
rect 5124 11484 5156 11486
rect 5124 11434 5156 11436
rect 5124 11406 5126 11434
rect 5126 11406 5154 11434
rect 5154 11406 5156 11434
rect 5124 11404 5156 11406
rect 5124 10874 5156 10876
rect 5124 10846 5126 10874
rect 5126 10846 5154 10874
rect 5154 10846 5156 10874
rect 5124 10844 5156 10846
rect 5124 10794 5156 10796
rect 5124 10766 5126 10794
rect 5126 10766 5154 10794
rect 5154 10766 5156 10794
rect 5124 10764 5156 10766
rect 5124 10714 5156 10716
rect 5124 10686 5126 10714
rect 5126 10686 5154 10714
rect 5154 10686 5156 10714
rect 5124 10684 5156 10686
rect 5124 10634 5156 10636
rect 5124 10606 5126 10634
rect 5126 10606 5154 10634
rect 5154 10606 5156 10634
rect 5124 10604 5156 10606
rect 5124 10554 5156 10556
rect 5124 10526 5126 10554
rect 5126 10526 5154 10554
rect 5154 10526 5156 10554
rect 5124 10524 5156 10526
rect 5124 10474 5156 10476
rect 5124 10446 5126 10474
rect 5126 10446 5154 10474
rect 5154 10446 5156 10474
rect 5124 10444 5156 10446
rect 5124 10394 5156 10396
rect 5124 10366 5126 10394
rect 5126 10366 5154 10394
rect 5154 10366 5156 10394
rect 5124 10364 5156 10366
rect 5124 10314 5156 10316
rect 5124 10286 5126 10314
rect 5126 10286 5154 10314
rect 5154 10286 5156 10314
rect 5124 10284 5156 10286
rect 5124 10234 5156 10236
rect 5124 10206 5126 10234
rect 5126 10206 5154 10234
rect 5154 10206 5156 10234
rect 5124 10204 5156 10206
rect 5124 10154 5156 10156
rect 5124 10126 5126 10154
rect 5126 10126 5154 10154
rect 5154 10126 5156 10154
rect 5124 10124 5156 10126
rect 5124 10074 5156 10076
rect 5124 10046 5126 10074
rect 5126 10046 5154 10074
rect 5154 10046 5156 10074
rect 5124 10044 5156 10046
rect 5124 9994 5156 9996
rect 5124 9966 5126 9994
rect 5126 9966 5154 9994
rect 5154 9966 5156 9994
rect 5124 9964 5156 9966
rect 5124 9914 5156 9916
rect 5124 9886 5126 9914
rect 5126 9886 5154 9914
rect 5154 9886 5156 9914
rect 5124 9884 5156 9886
rect 5124 9834 5156 9836
rect 5124 9806 5126 9834
rect 5126 9806 5154 9834
rect 5154 9806 5156 9834
rect 5124 9804 5156 9806
rect 5124 9754 5156 9756
rect 5124 9726 5126 9754
rect 5126 9726 5154 9754
rect 5154 9726 5156 9754
rect 5124 9724 5156 9726
rect 5124 9354 5156 9356
rect 5124 9326 5126 9354
rect 5126 9326 5154 9354
rect 5154 9326 5156 9354
rect 5124 9324 5156 9326
rect 5124 9274 5156 9276
rect 5124 9246 5126 9274
rect 5126 9246 5154 9274
rect 5154 9246 5156 9274
rect 5124 9244 5156 9246
rect 5124 9194 5156 9196
rect 5124 9166 5126 9194
rect 5126 9166 5154 9194
rect 5154 9166 5156 9194
rect 5124 9164 5156 9166
rect 5124 8874 5156 8876
rect 5124 8846 5126 8874
rect 5126 8846 5154 8874
rect 5154 8846 5156 8874
rect 5124 8844 5156 8846
rect 5124 8794 5156 8796
rect 5124 8766 5126 8794
rect 5126 8766 5154 8794
rect 5154 8766 5156 8794
rect 5124 8764 5156 8766
rect 5124 8714 5156 8716
rect 5124 8686 5126 8714
rect 5126 8686 5154 8714
rect 5154 8686 5156 8714
rect 5124 8684 5156 8686
rect 5124 8634 5156 8636
rect 5124 8606 5126 8634
rect 5126 8606 5154 8634
rect 5154 8606 5156 8634
rect 5124 8604 5156 8606
rect 5124 8554 5156 8556
rect 5124 8526 5126 8554
rect 5126 8526 5154 8554
rect 5154 8526 5156 8554
rect 5124 8524 5156 8526
rect 5124 7634 5156 7636
rect 5124 7606 5126 7634
rect 5126 7606 5154 7634
rect 5154 7606 5156 7634
rect 5124 7604 5156 7606
rect 5124 7554 5156 7556
rect 5124 7526 5126 7554
rect 5126 7526 5154 7554
rect 5154 7526 5156 7554
rect 5124 7524 5156 7526
rect 5124 7474 5156 7476
rect 5124 7446 5126 7474
rect 5126 7446 5154 7474
rect 5154 7446 5156 7474
rect 5124 7444 5156 7446
rect 5124 7394 5156 7396
rect 5124 7366 5126 7394
rect 5126 7366 5154 7394
rect 5154 7366 5156 7394
rect 5124 7364 5156 7366
rect 5124 7314 5156 7316
rect 5124 7286 5126 7314
rect 5126 7286 5154 7314
rect 5154 7286 5156 7314
rect 5124 7284 5156 7286
rect 5124 7234 5156 7236
rect 5124 7206 5126 7234
rect 5126 7206 5154 7234
rect 5154 7206 5156 7234
rect 5124 7204 5156 7206
rect 5124 7154 5156 7156
rect 5124 7126 5126 7154
rect 5126 7126 5154 7154
rect 5154 7126 5156 7154
rect 5124 7124 5156 7126
rect 5124 7074 5156 7076
rect 5124 7046 5126 7074
rect 5126 7046 5154 7074
rect 5154 7046 5156 7074
rect 5124 7044 5156 7046
rect 5124 6754 5156 6756
rect 5124 6726 5126 6754
rect 5126 6726 5154 6754
rect 5154 6726 5156 6754
rect 5124 6724 5156 6726
rect 5124 6674 5156 6676
rect 5124 6646 5126 6674
rect 5126 6646 5154 6674
rect 5154 6646 5156 6674
rect 5124 6644 5156 6646
rect 5124 6594 5156 6596
rect 5124 6566 5126 6594
rect 5126 6566 5154 6594
rect 5154 6566 5156 6594
rect 5124 6564 5156 6566
rect 5124 6514 5156 6516
rect 5124 6486 5126 6514
rect 5126 6486 5154 6514
rect 5154 6486 5156 6514
rect 5124 6484 5156 6486
rect 5124 6434 5156 6436
rect 5124 6406 5126 6434
rect 5126 6406 5154 6434
rect 5154 6406 5156 6434
rect 5124 6404 5156 6406
rect 5124 6354 5156 6356
rect 5124 6326 5126 6354
rect 5126 6326 5154 6354
rect 5154 6326 5156 6354
rect 5124 6324 5156 6326
rect 5124 5794 5156 5796
rect 5124 5766 5126 5794
rect 5126 5766 5154 5794
rect 5154 5766 5156 5794
rect 5124 5764 5156 5766
rect 5124 5714 5156 5716
rect 5124 5686 5126 5714
rect 5126 5686 5154 5714
rect 5154 5686 5156 5714
rect 5124 5684 5156 5686
rect 5124 5634 5156 5636
rect 5124 5606 5126 5634
rect 5126 5606 5154 5634
rect 5154 5606 5156 5634
rect 5124 5604 5156 5606
rect 5124 5554 5156 5556
rect 5124 5526 5126 5554
rect 5126 5526 5154 5554
rect 5154 5526 5156 5554
rect 5124 5524 5156 5526
rect 5124 5474 5156 5476
rect 5124 5446 5126 5474
rect 5126 5446 5154 5474
rect 5154 5446 5156 5474
rect 5124 5444 5156 5446
rect 5124 5394 5156 5396
rect 5124 5366 5126 5394
rect 5126 5366 5154 5394
rect 5154 5366 5156 5394
rect 5124 5364 5156 5366
rect 5124 5314 5156 5316
rect 5124 5286 5126 5314
rect 5126 5286 5154 5314
rect 5154 5286 5156 5314
rect 5124 5284 5156 5286
rect 5124 5234 5156 5236
rect 5124 5206 5126 5234
rect 5126 5206 5154 5234
rect 5154 5206 5156 5234
rect 5124 5204 5156 5206
rect 5124 5154 5156 5156
rect 5124 5126 5126 5154
rect 5126 5126 5154 5154
rect 5154 5126 5156 5154
rect 5124 5124 5156 5126
rect 5124 5074 5156 5076
rect 5124 5046 5126 5074
rect 5126 5046 5154 5074
rect 5154 5046 5156 5074
rect 5124 5044 5156 5046
rect 5124 4994 5156 4996
rect 5124 4966 5126 4994
rect 5126 4966 5154 4994
rect 5154 4966 5156 4994
rect 5124 4964 5156 4966
rect 5124 4434 5156 4436
rect 5124 4406 5126 4434
rect 5126 4406 5154 4434
rect 5154 4406 5156 4434
rect 5124 4404 5156 4406
rect 5124 4354 5156 4356
rect 5124 4326 5126 4354
rect 5126 4326 5154 4354
rect 5154 4326 5156 4354
rect 5124 4324 5156 4326
rect 5124 4274 5156 4276
rect 5124 4246 5126 4274
rect 5126 4246 5154 4274
rect 5154 4246 5156 4274
rect 5124 4244 5156 4246
rect 5124 4194 5156 4196
rect 5124 4166 5126 4194
rect 5126 4166 5154 4194
rect 5154 4166 5156 4194
rect 5124 4164 5156 4166
rect 5124 4114 5156 4116
rect 5124 4086 5126 4114
rect 5126 4086 5154 4114
rect 5154 4086 5156 4114
rect 5124 4084 5156 4086
rect 5124 4034 5156 4036
rect 5124 4006 5126 4034
rect 5126 4006 5154 4034
rect 5154 4006 5156 4034
rect 5124 4004 5156 4006
rect 5124 3954 5156 3956
rect 5124 3926 5126 3954
rect 5126 3926 5154 3954
rect 5154 3926 5156 3954
rect 5124 3924 5156 3926
rect 5124 3154 5156 3156
rect 5124 3126 5126 3154
rect 5126 3126 5154 3154
rect 5154 3126 5156 3154
rect 5124 3124 5156 3126
rect 5124 3074 5156 3076
rect 5124 3046 5126 3074
rect 5126 3046 5154 3074
rect 5154 3046 5156 3074
rect 5124 3044 5156 3046
rect 5124 2994 5156 2996
rect 5124 2966 5126 2994
rect 5126 2966 5154 2994
rect 5154 2966 5156 2994
rect 5124 2964 5156 2966
rect 5124 2914 5156 2916
rect 5124 2886 5126 2914
rect 5126 2886 5154 2914
rect 5154 2886 5156 2914
rect 5124 2884 5156 2886
rect 5124 2834 5156 2836
rect 5124 2806 5126 2834
rect 5126 2806 5154 2834
rect 5154 2806 5156 2834
rect 5124 2804 5156 2806
rect 5124 2754 5156 2756
rect 5124 2726 5126 2754
rect 5126 2726 5154 2754
rect 5154 2726 5156 2754
rect 5124 2724 5156 2726
rect 5124 2674 5156 2676
rect 5124 2646 5126 2674
rect 5126 2646 5154 2674
rect 5154 2646 5156 2674
rect 5124 2644 5156 2646
rect 5124 2594 5156 2596
rect 5124 2566 5126 2594
rect 5126 2566 5154 2594
rect 5154 2566 5156 2594
rect 5124 2564 5156 2566
rect 5124 2514 5156 2516
rect 5124 2486 5126 2514
rect 5126 2486 5154 2514
rect 5154 2486 5156 2514
rect 5124 2484 5156 2486
rect 5124 2434 5156 2436
rect 5124 2406 5126 2434
rect 5126 2406 5154 2434
rect 5154 2406 5156 2434
rect 5124 2404 5156 2406
rect 5124 2354 5156 2356
rect 5124 2326 5126 2354
rect 5126 2326 5154 2354
rect 5154 2326 5156 2354
rect 5124 2324 5156 2326
rect 5124 2274 5156 2276
rect 5124 2246 5126 2274
rect 5126 2246 5154 2274
rect 5154 2246 5156 2274
rect 5124 2244 5156 2246
rect 5124 2194 5156 2196
rect 5124 2166 5126 2194
rect 5126 2166 5154 2194
rect 5154 2166 5156 2194
rect 5124 2164 5156 2166
rect 5124 2114 5156 2116
rect 5124 2086 5126 2114
rect 5126 2086 5154 2114
rect 5154 2086 5156 2114
rect 5124 2084 5156 2086
rect 5124 2034 5156 2036
rect 5124 2006 5126 2034
rect 5126 2006 5154 2034
rect 5154 2006 5156 2034
rect 5124 2004 5156 2006
rect 5124 1634 5156 1636
rect 5124 1606 5126 1634
rect 5126 1606 5154 1634
rect 5154 1606 5156 1634
rect 5124 1604 5156 1606
rect 5124 1554 5156 1556
rect 5124 1526 5126 1554
rect 5126 1526 5154 1554
rect 5154 1526 5156 1554
rect 5124 1524 5156 1526
rect 5124 1474 5156 1476
rect 5124 1446 5126 1474
rect 5126 1446 5154 1474
rect 5154 1446 5156 1474
rect 5124 1444 5156 1446
rect 5124 1394 5156 1396
rect 5124 1366 5126 1394
rect 5126 1366 5154 1394
rect 5154 1366 5156 1394
rect 5124 1364 5156 1366
rect 5124 1314 5156 1316
rect 5124 1286 5126 1314
rect 5126 1286 5154 1314
rect 5154 1286 5156 1314
rect 5124 1284 5156 1286
rect 5124 1234 5156 1236
rect 5124 1206 5126 1234
rect 5126 1206 5154 1234
rect 5154 1206 5156 1234
rect 5124 1204 5156 1206
rect 5124 1154 5156 1156
rect 5124 1126 5126 1154
rect 5126 1126 5154 1154
rect 5154 1126 5156 1154
rect 5124 1124 5156 1126
rect 5124 1074 5156 1076
rect 5124 1046 5126 1074
rect 5126 1046 5154 1074
rect 5154 1046 5156 1074
rect 5124 1044 5156 1046
rect 5124 754 5156 756
rect 5124 726 5126 754
rect 5126 726 5154 754
rect 5154 726 5156 754
rect 5124 724 5156 726
rect 5124 674 5156 676
rect 5124 646 5126 674
rect 5126 646 5154 674
rect 5154 646 5156 674
rect 5124 644 5156 646
rect 5124 594 5156 596
rect 5124 566 5126 594
rect 5126 566 5154 594
rect 5154 566 5156 594
rect 5124 564 5156 566
rect 5124 194 5156 196
rect 5124 166 5126 194
rect 5126 166 5154 194
rect 5154 166 5156 194
rect 5124 164 5156 166
rect 5124 114 5156 116
rect 5124 86 5126 114
rect 5126 86 5154 114
rect 5154 86 5156 114
rect 5124 84 5156 86
rect 5124 34 5156 36
rect 5124 6 5126 34
rect 5126 6 5154 34
rect 5154 6 5156 34
rect 5124 4 5156 6
rect 5204 15284 5236 15316
rect 5284 15364 5316 15396
rect 5284 14084 5316 14116
rect 5284 12634 5316 12636
rect 5284 12606 5286 12634
rect 5286 12606 5314 12634
rect 5314 12606 5316 12634
rect 5284 12604 5316 12606
rect 5284 12554 5316 12556
rect 5284 12526 5286 12554
rect 5286 12526 5314 12554
rect 5314 12526 5316 12554
rect 5284 12524 5316 12526
rect 5284 12474 5316 12476
rect 5284 12446 5286 12474
rect 5286 12446 5314 12474
rect 5314 12446 5316 12474
rect 5284 12444 5316 12446
rect 5284 12394 5316 12396
rect 5284 12366 5286 12394
rect 5286 12366 5314 12394
rect 5314 12366 5316 12394
rect 5284 12364 5316 12366
rect 5284 12314 5316 12316
rect 5284 12286 5286 12314
rect 5286 12286 5314 12314
rect 5314 12286 5316 12314
rect 5284 12284 5316 12286
rect 5284 12234 5316 12236
rect 5284 12206 5286 12234
rect 5286 12206 5314 12234
rect 5314 12206 5316 12234
rect 5284 12204 5316 12206
rect 5284 12154 5316 12156
rect 5284 12126 5286 12154
rect 5286 12126 5314 12154
rect 5314 12126 5316 12154
rect 5284 12124 5316 12126
rect 5284 11834 5316 11836
rect 5284 11806 5286 11834
rect 5286 11806 5314 11834
rect 5314 11806 5316 11834
rect 5284 11804 5316 11806
rect 5284 11754 5316 11756
rect 5284 11726 5286 11754
rect 5286 11726 5314 11754
rect 5314 11726 5316 11754
rect 5284 11724 5316 11726
rect 5284 11674 5316 11676
rect 5284 11646 5286 11674
rect 5286 11646 5314 11674
rect 5314 11646 5316 11674
rect 5284 11644 5316 11646
rect 5284 11594 5316 11596
rect 5284 11566 5286 11594
rect 5286 11566 5314 11594
rect 5314 11566 5316 11594
rect 5284 11564 5316 11566
rect 5284 11514 5316 11516
rect 5284 11486 5286 11514
rect 5286 11486 5314 11514
rect 5314 11486 5316 11514
rect 5284 11484 5316 11486
rect 5284 11434 5316 11436
rect 5284 11406 5286 11434
rect 5286 11406 5314 11434
rect 5314 11406 5316 11434
rect 5284 11404 5316 11406
rect 5284 10874 5316 10876
rect 5284 10846 5286 10874
rect 5286 10846 5314 10874
rect 5314 10846 5316 10874
rect 5284 10844 5316 10846
rect 5284 10794 5316 10796
rect 5284 10766 5286 10794
rect 5286 10766 5314 10794
rect 5314 10766 5316 10794
rect 5284 10764 5316 10766
rect 5284 10714 5316 10716
rect 5284 10686 5286 10714
rect 5286 10686 5314 10714
rect 5314 10686 5316 10714
rect 5284 10684 5316 10686
rect 5284 10634 5316 10636
rect 5284 10606 5286 10634
rect 5286 10606 5314 10634
rect 5314 10606 5316 10634
rect 5284 10604 5316 10606
rect 5284 10554 5316 10556
rect 5284 10526 5286 10554
rect 5286 10526 5314 10554
rect 5314 10526 5316 10554
rect 5284 10524 5316 10526
rect 5284 10474 5316 10476
rect 5284 10446 5286 10474
rect 5286 10446 5314 10474
rect 5314 10446 5316 10474
rect 5284 10444 5316 10446
rect 5284 10394 5316 10396
rect 5284 10366 5286 10394
rect 5286 10366 5314 10394
rect 5314 10366 5316 10394
rect 5284 10364 5316 10366
rect 5284 10314 5316 10316
rect 5284 10286 5286 10314
rect 5286 10286 5314 10314
rect 5314 10286 5316 10314
rect 5284 10284 5316 10286
rect 5284 10234 5316 10236
rect 5284 10206 5286 10234
rect 5286 10206 5314 10234
rect 5314 10206 5316 10234
rect 5284 10204 5316 10206
rect 5284 10154 5316 10156
rect 5284 10126 5286 10154
rect 5286 10126 5314 10154
rect 5314 10126 5316 10154
rect 5284 10124 5316 10126
rect 5284 10074 5316 10076
rect 5284 10046 5286 10074
rect 5286 10046 5314 10074
rect 5314 10046 5316 10074
rect 5284 10044 5316 10046
rect 5284 9994 5316 9996
rect 5284 9966 5286 9994
rect 5286 9966 5314 9994
rect 5314 9966 5316 9994
rect 5284 9964 5316 9966
rect 5284 9914 5316 9916
rect 5284 9886 5286 9914
rect 5286 9886 5314 9914
rect 5314 9886 5316 9914
rect 5284 9884 5316 9886
rect 5284 9834 5316 9836
rect 5284 9806 5286 9834
rect 5286 9806 5314 9834
rect 5314 9806 5316 9834
rect 5284 9804 5316 9806
rect 5284 9754 5316 9756
rect 5284 9726 5286 9754
rect 5286 9726 5314 9754
rect 5314 9726 5316 9754
rect 5284 9724 5316 9726
rect 5284 9354 5316 9356
rect 5284 9326 5286 9354
rect 5286 9326 5314 9354
rect 5314 9326 5316 9354
rect 5284 9324 5316 9326
rect 5284 9274 5316 9276
rect 5284 9246 5286 9274
rect 5286 9246 5314 9274
rect 5314 9246 5316 9274
rect 5284 9244 5316 9246
rect 5284 9194 5316 9196
rect 5284 9166 5286 9194
rect 5286 9166 5314 9194
rect 5314 9166 5316 9194
rect 5284 9164 5316 9166
rect 5284 8874 5316 8876
rect 5284 8846 5286 8874
rect 5286 8846 5314 8874
rect 5314 8846 5316 8874
rect 5284 8844 5316 8846
rect 5284 8794 5316 8796
rect 5284 8766 5286 8794
rect 5286 8766 5314 8794
rect 5314 8766 5316 8794
rect 5284 8764 5316 8766
rect 5284 8714 5316 8716
rect 5284 8686 5286 8714
rect 5286 8686 5314 8714
rect 5314 8686 5316 8714
rect 5284 8684 5316 8686
rect 5284 8634 5316 8636
rect 5284 8606 5286 8634
rect 5286 8606 5314 8634
rect 5314 8606 5316 8634
rect 5284 8604 5316 8606
rect 5284 8554 5316 8556
rect 5284 8526 5286 8554
rect 5286 8526 5314 8554
rect 5314 8526 5316 8554
rect 5284 8524 5316 8526
rect 5284 7634 5316 7636
rect 5284 7606 5286 7634
rect 5286 7606 5314 7634
rect 5314 7606 5316 7634
rect 5284 7604 5316 7606
rect 5284 7554 5316 7556
rect 5284 7526 5286 7554
rect 5286 7526 5314 7554
rect 5314 7526 5316 7554
rect 5284 7524 5316 7526
rect 5284 7474 5316 7476
rect 5284 7446 5286 7474
rect 5286 7446 5314 7474
rect 5314 7446 5316 7474
rect 5284 7444 5316 7446
rect 5284 7394 5316 7396
rect 5284 7366 5286 7394
rect 5286 7366 5314 7394
rect 5314 7366 5316 7394
rect 5284 7364 5316 7366
rect 5284 7314 5316 7316
rect 5284 7286 5286 7314
rect 5286 7286 5314 7314
rect 5314 7286 5316 7314
rect 5284 7284 5316 7286
rect 5284 7234 5316 7236
rect 5284 7206 5286 7234
rect 5286 7206 5314 7234
rect 5314 7206 5316 7234
rect 5284 7204 5316 7206
rect 5284 7154 5316 7156
rect 5284 7126 5286 7154
rect 5286 7126 5314 7154
rect 5314 7126 5316 7154
rect 5284 7124 5316 7126
rect 5284 7074 5316 7076
rect 5284 7046 5286 7074
rect 5286 7046 5314 7074
rect 5314 7046 5316 7074
rect 5284 7044 5316 7046
rect 5284 6754 5316 6756
rect 5284 6726 5286 6754
rect 5286 6726 5314 6754
rect 5314 6726 5316 6754
rect 5284 6724 5316 6726
rect 5284 6674 5316 6676
rect 5284 6646 5286 6674
rect 5286 6646 5314 6674
rect 5314 6646 5316 6674
rect 5284 6644 5316 6646
rect 5284 6594 5316 6596
rect 5284 6566 5286 6594
rect 5286 6566 5314 6594
rect 5314 6566 5316 6594
rect 5284 6564 5316 6566
rect 5284 6514 5316 6516
rect 5284 6486 5286 6514
rect 5286 6486 5314 6514
rect 5314 6486 5316 6514
rect 5284 6484 5316 6486
rect 5284 6434 5316 6436
rect 5284 6406 5286 6434
rect 5286 6406 5314 6434
rect 5314 6406 5316 6434
rect 5284 6404 5316 6406
rect 5284 6354 5316 6356
rect 5284 6326 5286 6354
rect 5286 6326 5314 6354
rect 5314 6326 5316 6354
rect 5284 6324 5316 6326
rect 5284 5794 5316 5796
rect 5284 5766 5286 5794
rect 5286 5766 5314 5794
rect 5314 5766 5316 5794
rect 5284 5764 5316 5766
rect 5284 5714 5316 5716
rect 5284 5686 5286 5714
rect 5286 5686 5314 5714
rect 5314 5686 5316 5714
rect 5284 5684 5316 5686
rect 5284 5634 5316 5636
rect 5284 5606 5286 5634
rect 5286 5606 5314 5634
rect 5314 5606 5316 5634
rect 5284 5604 5316 5606
rect 5284 5554 5316 5556
rect 5284 5526 5286 5554
rect 5286 5526 5314 5554
rect 5314 5526 5316 5554
rect 5284 5524 5316 5526
rect 5284 5474 5316 5476
rect 5284 5446 5286 5474
rect 5286 5446 5314 5474
rect 5314 5446 5316 5474
rect 5284 5444 5316 5446
rect 5284 5394 5316 5396
rect 5284 5366 5286 5394
rect 5286 5366 5314 5394
rect 5314 5366 5316 5394
rect 5284 5364 5316 5366
rect 5284 5314 5316 5316
rect 5284 5286 5286 5314
rect 5286 5286 5314 5314
rect 5314 5286 5316 5314
rect 5284 5284 5316 5286
rect 5284 5234 5316 5236
rect 5284 5206 5286 5234
rect 5286 5206 5314 5234
rect 5314 5206 5316 5234
rect 5284 5204 5316 5206
rect 5284 5154 5316 5156
rect 5284 5126 5286 5154
rect 5286 5126 5314 5154
rect 5314 5126 5316 5154
rect 5284 5124 5316 5126
rect 5284 5074 5316 5076
rect 5284 5046 5286 5074
rect 5286 5046 5314 5074
rect 5314 5046 5316 5074
rect 5284 5044 5316 5046
rect 5284 4994 5316 4996
rect 5284 4966 5286 4994
rect 5286 4966 5314 4994
rect 5314 4966 5316 4994
rect 5284 4964 5316 4966
rect 5284 4434 5316 4436
rect 5284 4406 5286 4434
rect 5286 4406 5314 4434
rect 5314 4406 5316 4434
rect 5284 4404 5316 4406
rect 5284 4354 5316 4356
rect 5284 4326 5286 4354
rect 5286 4326 5314 4354
rect 5314 4326 5316 4354
rect 5284 4324 5316 4326
rect 5284 4274 5316 4276
rect 5284 4246 5286 4274
rect 5286 4246 5314 4274
rect 5314 4246 5316 4274
rect 5284 4244 5316 4246
rect 5284 4194 5316 4196
rect 5284 4166 5286 4194
rect 5286 4166 5314 4194
rect 5314 4166 5316 4194
rect 5284 4164 5316 4166
rect 5284 4114 5316 4116
rect 5284 4086 5286 4114
rect 5286 4086 5314 4114
rect 5314 4086 5316 4114
rect 5284 4084 5316 4086
rect 5284 4034 5316 4036
rect 5284 4006 5286 4034
rect 5286 4006 5314 4034
rect 5314 4006 5316 4034
rect 5284 4004 5316 4006
rect 5284 3954 5316 3956
rect 5284 3926 5286 3954
rect 5286 3926 5314 3954
rect 5314 3926 5316 3954
rect 5284 3924 5316 3926
rect 5284 3154 5316 3156
rect 5284 3126 5286 3154
rect 5286 3126 5314 3154
rect 5314 3126 5316 3154
rect 5284 3124 5316 3126
rect 5284 3074 5316 3076
rect 5284 3046 5286 3074
rect 5286 3046 5314 3074
rect 5314 3046 5316 3074
rect 5284 3044 5316 3046
rect 5284 2994 5316 2996
rect 5284 2966 5286 2994
rect 5286 2966 5314 2994
rect 5314 2966 5316 2994
rect 5284 2964 5316 2966
rect 5284 2914 5316 2916
rect 5284 2886 5286 2914
rect 5286 2886 5314 2914
rect 5314 2886 5316 2914
rect 5284 2884 5316 2886
rect 5284 2834 5316 2836
rect 5284 2806 5286 2834
rect 5286 2806 5314 2834
rect 5314 2806 5316 2834
rect 5284 2804 5316 2806
rect 5284 2754 5316 2756
rect 5284 2726 5286 2754
rect 5286 2726 5314 2754
rect 5314 2726 5316 2754
rect 5284 2724 5316 2726
rect 5284 2674 5316 2676
rect 5284 2646 5286 2674
rect 5286 2646 5314 2674
rect 5314 2646 5316 2674
rect 5284 2644 5316 2646
rect 5284 2594 5316 2596
rect 5284 2566 5286 2594
rect 5286 2566 5314 2594
rect 5314 2566 5316 2594
rect 5284 2564 5316 2566
rect 5284 2514 5316 2516
rect 5284 2486 5286 2514
rect 5286 2486 5314 2514
rect 5314 2486 5316 2514
rect 5284 2484 5316 2486
rect 5284 2434 5316 2436
rect 5284 2406 5286 2434
rect 5286 2406 5314 2434
rect 5314 2406 5316 2434
rect 5284 2404 5316 2406
rect 5284 2354 5316 2356
rect 5284 2326 5286 2354
rect 5286 2326 5314 2354
rect 5314 2326 5316 2354
rect 5284 2324 5316 2326
rect 5284 2274 5316 2276
rect 5284 2246 5286 2274
rect 5286 2246 5314 2274
rect 5314 2246 5316 2274
rect 5284 2244 5316 2246
rect 5284 2194 5316 2196
rect 5284 2166 5286 2194
rect 5286 2166 5314 2194
rect 5314 2166 5316 2194
rect 5284 2164 5316 2166
rect 5284 2114 5316 2116
rect 5284 2086 5286 2114
rect 5286 2086 5314 2114
rect 5314 2086 5316 2114
rect 5284 2084 5316 2086
rect 5284 2034 5316 2036
rect 5284 2006 5286 2034
rect 5286 2006 5314 2034
rect 5314 2006 5316 2034
rect 5284 2004 5316 2006
rect 5284 1634 5316 1636
rect 5284 1606 5286 1634
rect 5286 1606 5314 1634
rect 5314 1606 5316 1634
rect 5284 1604 5316 1606
rect 5284 1554 5316 1556
rect 5284 1526 5286 1554
rect 5286 1526 5314 1554
rect 5314 1526 5316 1554
rect 5284 1524 5316 1526
rect 5284 1474 5316 1476
rect 5284 1446 5286 1474
rect 5286 1446 5314 1474
rect 5314 1446 5316 1474
rect 5284 1444 5316 1446
rect 5284 1394 5316 1396
rect 5284 1366 5286 1394
rect 5286 1366 5314 1394
rect 5314 1366 5316 1394
rect 5284 1364 5316 1366
rect 5284 1314 5316 1316
rect 5284 1286 5286 1314
rect 5286 1286 5314 1314
rect 5314 1286 5316 1314
rect 5284 1284 5316 1286
rect 5284 1234 5316 1236
rect 5284 1206 5286 1234
rect 5286 1206 5314 1234
rect 5314 1206 5316 1234
rect 5284 1204 5316 1206
rect 5284 1154 5316 1156
rect 5284 1126 5286 1154
rect 5286 1126 5314 1154
rect 5314 1126 5316 1154
rect 5284 1124 5316 1126
rect 5284 1074 5316 1076
rect 5284 1046 5286 1074
rect 5286 1046 5314 1074
rect 5314 1046 5316 1074
rect 5284 1044 5316 1046
rect 5284 754 5316 756
rect 5284 726 5286 754
rect 5286 726 5314 754
rect 5314 726 5316 754
rect 5284 724 5316 726
rect 5284 674 5316 676
rect 5284 646 5286 674
rect 5286 646 5314 674
rect 5314 646 5316 674
rect 5284 644 5316 646
rect 5284 594 5316 596
rect 5284 566 5286 594
rect 5286 566 5314 594
rect 5314 566 5316 594
rect 5284 564 5316 566
rect 5284 194 5316 196
rect 5284 166 5286 194
rect 5286 166 5314 194
rect 5314 166 5316 194
rect 5284 164 5316 166
rect 5284 114 5316 116
rect 5284 86 5286 114
rect 5286 86 5314 114
rect 5314 86 5316 114
rect 5284 84 5316 86
rect 5284 34 5316 36
rect 5284 6 5286 34
rect 5286 6 5314 34
rect 5314 6 5316 34
rect 5284 4 5316 6
rect 5364 15284 5396 15316
rect 5444 15364 5476 15396
rect 5444 14084 5476 14116
rect 5444 12634 5476 12636
rect 5444 12606 5446 12634
rect 5446 12606 5474 12634
rect 5474 12606 5476 12634
rect 5444 12604 5476 12606
rect 5444 12554 5476 12556
rect 5444 12526 5446 12554
rect 5446 12526 5474 12554
rect 5474 12526 5476 12554
rect 5444 12524 5476 12526
rect 5444 12474 5476 12476
rect 5444 12446 5446 12474
rect 5446 12446 5474 12474
rect 5474 12446 5476 12474
rect 5444 12444 5476 12446
rect 5444 12394 5476 12396
rect 5444 12366 5446 12394
rect 5446 12366 5474 12394
rect 5474 12366 5476 12394
rect 5444 12364 5476 12366
rect 5444 12314 5476 12316
rect 5444 12286 5446 12314
rect 5446 12286 5474 12314
rect 5474 12286 5476 12314
rect 5444 12284 5476 12286
rect 5444 12234 5476 12236
rect 5444 12206 5446 12234
rect 5446 12206 5474 12234
rect 5474 12206 5476 12234
rect 5444 12204 5476 12206
rect 5444 12154 5476 12156
rect 5444 12126 5446 12154
rect 5446 12126 5474 12154
rect 5474 12126 5476 12154
rect 5444 12124 5476 12126
rect 5444 11834 5476 11836
rect 5444 11806 5446 11834
rect 5446 11806 5474 11834
rect 5474 11806 5476 11834
rect 5444 11804 5476 11806
rect 5444 11754 5476 11756
rect 5444 11726 5446 11754
rect 5446 11726 5474 11754
rect 5474 11726 5476 11754
rect 5444 11724 5476 11726
rect 5444 11674 5476 11676
rect 5444 11646 5446 11674
rect 5446 11646 5474 11674
rect 5474 11646 5476 11674
rect 5444 11644 5476 11646
rect 5444 11594 5476 11596
rect 5444 11566 5446 11594
rect 5446 11566 5474 11594
rect 5474 11566 5476 11594
rect 5444 11564 5476 11566
rect 5444 11514 5476 11516
rect 5444 11486 5446 11514
rect 5446 11486 5474 11514
rect 5474 11486 5476 11514
rect 5444 11484 5476 11486
rect 5444 11434 5476 11436
rect 5444 11406 5446 11434
rect 5446 11406 5474 11434
rect 5474 11406 5476 11434
rect 5444 11404 5476 11406
rect 5444 10874 5476 10876
rect 5444 10846 5446 10874
rect 5446 10846 5474 10874
rect 5474 10846 5476 10874
rect 5444 10844 5476 10846
rect 5444 10794 5476 10796
rect 5444 10766 5446 10794
rect 5446 10766 5474 10794
rect 5474 10766 5476 10794
rect 5444 10764 5476 10766
rect 5444 10714 5476 10716
rect 5444 10686 5446 10714
rect 5446 10686 5474 10714
rect 5474 10686 5476 10714
rect 5444 10684 5476 10686
rect 5444 10634 5476 10636
rect 5444 10606 5446 10634
rect 5446 10606 5474 10634
rect 5474 10606 5476 10634
rect 5444 10604 5476 10606
rect 5444 10554 5476 10556
rect 5444 10526 5446 10554
rect 5446 10526 5474 10554
rect 5474 10526 5476 10554
rect 5444 10524 5476 10526
rect 5444 10474 5476 10476
rect 5444 10446 5446 10474
rect 5446 10446 5474 10474
rect 5474 10446 5476 10474
rect 5444 10444 5476 10446
rect 5444 10394 5476 10396
rect 5444 10366 5446 10394
rect 5446 10366 5474 10394
rect 5474 10366 5476 10394
rect 5444 10364 5476 10366
rect 5444 10314 5476 10316
rect 5444 10286 5446 10314
rect 5446 10286 5474 10314
rect 5474 10286 5476 10314
rect 5444 10284 5476 10286
rect 5444 10234 5476 10236
rect 5444 10206 5446 10234
rect 5446 10206 5474 10234
rect 5474 10206 5476 10234
rect 5444 10204 5476 10206
rect 5444 10154 5476 10156
rect 5444 10126 5446 10154
rect 5446 10126 5474 10154
rect 5474 10126 5476 10154
rect 5444 10124 5476 10126
rect 5444 10074 5476 10076
rect 5444 10046 5446 10074
rect 5446 10046 5474 10074
rect 5474 10046 5476 10074
rect 5444 10044 5476 10046
rect 5444 9994 5476 9996
rect 5444 9966 5446 9994
rect 5446 9966 5474 9994
rect 5474 9966 5476 9994
rect 5444 9964 5476 9966
rect 5444 9914 5476 9916
rect 5444 9886 5446 9914
rect 5446 9886 5474 9914
rect 5474 9886 5476 9914
rect 5444 9884 5476 9886
rect 5444 9834 5476 9836
rect 5444 9806 5446 9834
rect 5446 9806 5474 9834
rect 5474 9806 5476 9834
rect 5444 9804 5476 9806
rect 5444 9754 5476 9756
rect 5444 9726 5446 9754
rect 5446 9726 5474 9754
rect 5474 9726 5476 9754
rect 5444 9724 5476 9726
rect 5444 9354 5476 9356
rect 5444 9326 5446 9354
rect 5446 9326 5474 9354
rect 5474 9326 5476 9354
rect 5444 9324 5476 9326
rect 5444 9274 5476 9276
rect 5444 9246 5446 9274
rect 5446 9246 5474 9274
rect 5474 9246 5476 9274
rect 5444 9244 5476 9246
rect 5444 9194 5476 9196
rect 5444 9166 5446 9194
rect 5446 9166 5474 9194
rect 5474 9166 5476 9194
rect 5444 9164 5476 9166
rect 5444 8874 5476 8876
rect 5444 8846 5446 8874
rect 5446 8846 5474 8874
rect 5474 8846 5476 8874
rect 5444 8844 5476 8846
rect 5444 8794 5476 8796
rect 5444 8766 5446 8794
rect 5446 8766 5474 8794
rect 5474 8766 5476 8794
rect 5444 8764 5476 8766
rect 5444 8714 5476 8716
rect 5444 8686 5446 8714
rect 5446 8686 5474 8714
rect 5474 8686 5476 8714
rect 5444 8684 5476 8686
rect 5444 8634 5476 8636
rect 5444 8606 5446 8634
rect 5446 8606 5474 8634
rect 5474 8606 5476 8634
rect 5444 8604 5476 8606
rect 5444 8554 5476 8556
rect 5444 8526 5446 8554
rect 5446 8526 5474 8554
rect 5474 8526 5476 8554
rect 5444 8524 5476 8526
rect 5444 7634 5476 7636
rect 5444 7606 5446 7634
rect 5446 7606 5474 7634
rect 5474 7606 5476 7634
rect 5444 7604 5476 7606
rect 5444 7554 5476 7556
rect 5444 7526 5446 7554
rect 5446 7526 5474 7554
rect 5474 7526 5476 7554
rect 5444 7524 5476 7526
rect 5444 7474 5476 7476
rect 5444 7446 5446 7474
rect 5446 7446 5474 7474
rect 5474 7446 5476 7474
rect 5444 7444 5476 7446
rect 5444 7394 5476 7396
rect 5444 7366 5446 7394
rect 5446 7366 5474 7394
rect 5474 7366 5476 7394
rect 5444 7364 5476 7366
rect 5444 7314 5476 7316
rect 5444 7286 5446 7314
rect 5446 7286 5474 7314
rect 5474 7286 5476 7314
rect 5444 7284 5476 7286
rect 5444 7234 5476 7236
rect 5444 7206 5446 7234
rect 5446 7206 5474 7234
rect 5474 7206 5476 7234
rect 5444 7204 5476 7206
rect 5444 7154 5476 7156
rect 5444 7126 5446 7154
rect 5446 7126 5474 7154
rect 5474 7126 5476 7154
rect 5444 7124 5476 7126
rect 5444 7074 5476 7076
rect 5444 7046 5446 7074
rect 5446 7046 5474 7074
rect 5474 7046 5476 7074
rect 5444 7044 5476 7046
rect 5444 6754 5476 6756
rect 5444 6726 5446 6754
rect 5446 6726 5474 6754
rect 5474 6726 5476 6754
rect 5444 6724 5476 6726
rect 5444 6674 5476 6676
rect 5444 6646 5446 6674
rect 5446 6646 5474 6674
rect 5474 6646 5476 6674
rect 5444 6644 5476 6646
rect 5444 6594 5476 6596
rect 5444 6566 5446 6594
rect 5446 6566 5474 6594
rect 5474 6566 5476 6594
rect 5444 6564 5476 6566
rect 5444 6514 5476 6516
rect 5444 6486 5446 6514
rect 5446 6486 5474 6514
rect 5474 6486 5476 6514
rect 5444 6484 5476 6486
rect 5444 6434 5476 6436
rect 5444 6406 5446 6434
rect 5446 6406 5474 6434
rect 5474 6406 5476 6434
rect 5444 6404 5476 6406
rect 5444 6354 5476 6356
rect 5444 6326 5446 6354
rect 5446 6326 5474 6354
rect 5474 6326 5476 6354
rect 5444 6324 5476 6326
rect 5444 5794 5476 5796
rect 5444 5766 5446 5794
rect 5446 5766 5474 5794
rect 5474 5766 5476 5794
rect 5444 5764 5476 5766
rect 5444 5714 5476 5716
rect 5444 5686 5446 5714
rect 5446 5686 5474 5714
rect 5474 5686 5476 5714
rect 5444 5684 5476 5686
rect 5444 5634 5476 5636
rect 5444 5606 5446 5634
rect 5446 5606 5474 5634
rect 5474 5606 5476 5634
rect 5444 5604 5476 5606
rect 5444 5554 5476 5556
rect 5444 5526 5446 5554
rect 5446 5526 5474 5554
rect 5474 5526 5476 5554
rect 5444 5524 5476 5526
rect 5444 5474 5476 5476
rect 5444 5446 5446 5474
rect 5446 5446 5474 5474
rect 5474 5446 5476 5474
rect 5444 5444 5476 5446
rect 5444 5394 5476 5396
rect 5444 5366 5446 5394
rect 5446 5366 5474 5394
rect 5474 5366 5476 5394
rect 5444 5364 5476 5366
rect 5444 5314 5476 5316
rect 5444 5286 5446 5314
rect 5446 5286 5474 5314
rect 5474 5286 5476 5314
rect 5444 5284 5476 5286
rect 5444 5234 5476 5236
rect 5444 5206 5446 5234
rect 5446 5206 5474 5234
rect 5474 5206 5476 5234
rect 5444 5204 5476 5206
rect 5444 5154 5476 5156
rect 5444 5126 5446 5154
rect 5446 5126 5474 5154
rect 5474 5126 5476 5154
rect 5444 5124 5476 5126
rect 5444 5074 5476 5076
rect 5444 5046 5446 5074
rect 5446 5046 5474 5074
rect 5474 5046 5476 5074
rect 5444 5044 5476 5046
rect 5444 4994 5476 4996
rect 5444 4966 5446 4994
rect 5446 4966 5474 4994
rect 5474 4966 5476 4994
rect 5444 4964 5476 4966
rect 5444 4434 5476 4436
rect 5444 4406 5446 4434
rect 5446 4406 5474 4434
rect 5474 4406 5476 4434
rect 5444 4404 5476 4406
rect 5444 4354 5476 4356
rect 5444 4326 5446 4354
rect 5446 4326 5474 4354
rect 5474 4326 5476 4354
rect 5444 4324 5476 4326
rect 5444 4274 5476 4276
rect 5444 4246 5446 4274
rect 5446 4246 5474 4274
rect 5474 4246 5476 4274
rect 5444 4244 5476 4246
rect 5444 4194 5476 4196
rect 5444 4166 5446 4194
rect 5446 4166 5474 4194
rect 5474 4166 5476 4194
rect 5444 4164 5476 4166
rect 5444 4114 5476 4116
rect 5444 4086 5446 4114
rect 5446 4086 5474 4114
rect 5474 4086 5476 4114
rect 5444 4084 5476 4086
rect 5444 4034 5476 4036
rect 5444 4006 5446 4034
rect 5446 4006 5474 4034
rect 5474 4006 5476 4034
rect 5444 4004 5476 4006
rect 5444 3954 5476 3956
rect 5444 3926 5446 3954
rect 5446 3926 5474 3954
rect 5474 3926 5476 3954
rect 5444 3924 5476 3926
rect 5444 3154 5476 3156
rect 5444 3126 5446 3154
rect 5446 3126 5474 3154
rect 5474 3126 5476 3154
rect 5444 3124 5476 3126
rect 5444 3074 5476 3076
rect 5444 3046 5446 3074
rect 5446 3046 5474 3074
rect 5474 3046 5476 3074
rect 5444 3044 5476 3046
rect 5444 2994 5476 2996
rect 5444 2966 5446 2994
rect 5446 2966 5474 2994
rect 5474 2966 5476 2994
rect 5444 2964 5476 2966
rect 5444 2914 5476 2916
rect 5444 2886 5446 2914
rect 5446 2886 5474 2914
rect 5474 2886 5476 2914
rect 5444 2884 5476 2886
rect 5444 2834 5476 2836
rect 5444 2806 5446 2834
rect 5446 2806 5474 2834
rect 5474 2806 5476 2834
rect 5444 2804 5476 2806
rect 5444 2754 5476 2756
rect 5444 2726 5446 2754
rect 5446 2726 5474 2754
rect 5474 2726 5476 2754
rect 5444 2724 5476 2726
rect 5444 2674 5476 2676
rect 5444 2646 5446 2674
rect 5446 2646 5474 2674
rect 5474 2646 5476 2674
rect 5444 2644 5476 2646
rect 5444 2594 5476 2596
rect 5444 2566 5446 2594
rect 5446 2566 5474 2594
rect 5474 2566 5476 2594
rect 5444 2564 5476 2566
rect 5444 2514 5476 2516
rect 5444 2486 5446 2514
rect 5446 2486 5474 2514
rect 5474 2486 5476 2514
rect 5444 2484 5476 2486
rect 5444 2434 5476 2436
rect 5444 2406 5446 2434
rect 5446 2406 5474 2434
rect 5474 2406 5476 2434
rect 5444 2404 5476 2406
rect 5444 2354 5476 2356
rect 5444 2326 5446 2354
rect 5446 2326 5474 2354
rect 5474 2326 5476 2354
rect 5444 2324 5476 2326
rect 5444 2274 5476 2276
rect 5444 2246 5446 2274
rect 5446 2246 5474 2274
rect 5474 2246 5476 2274
rect 5444 2244 5476 2246
rect 5444 2194 5476 2196
rect 5444 2166 5446 2194
rect 5446 2166 5474 2194
rect 5474 2166 5476 2194
rect 5444 2164 5476 2166
rect 5444 2114 5476 2116
rect 5444 2086 5446 2114
rect 5446 2086 5474 2114
rect 5474 2086 5476 2114
rect 5444 2084 5476 2086
rect 5444 2034 5476 2036
rect 5444 2006 5446 2034
rect 5446 2006 5474 2034
rect 5474 2006 5476 2034
rect 5444 2004 5476 2006
rect 5444 1634 5476 1636
rect 5444 1606 5446 1634
rect 5446 1606 5474 1634
rect 5474 1606 5476 1634
rect 5444 1604 5476 1606
rect 5444 1554 5476 1556
rect 5444 1526 5446 1554
rect 5446 1526 5474 1554
rect 5474 1526 5476 1554
rect 5444 1524 5476 1526
rect 5444 1474 5476 1476
rect 5444 1446 5446 1474
rect 5446 1446 5474 1474
rect 5474 1446 5476 1474
rect 5444 1444 5476 1446
rect 5444 1394 5476 1396
rect 5444 1366 5446 1394
rect 5446 1366 5474 1394
rect 5474 1366 5476 1394
rect 5444 1364 5476 1366
rect 5444 1314 5476 1316
rect 5444 1286 5446 1314
rect 5446 1286 5474 1314
rect 5474 1286 5476 1314
rect 5444 1284 5476 1286
rect 5444 1234 5476 1236
rect 5444 1206 5446 1234
rect 5446 1206 5474 1234
rect 5474 1206 5476 1234
rect 5444 1204 5476 1206
rect 5444 1154 5476 1156
rect 5444 1126 5446 1154
rect 5446 1126 5474 1154
rect 5474 1126 5476 1154
rect 5444 1124 5476 1126
rect 5444 1074 5476 1076
rect 5444 1046 5446 1074
rect 5446 1046 5474 1074
rect 5474 1046 5476 1074
rect 5444 1044 5476 1046
rect 5444 754 5476 756
rect 5444 726 5446 754
rect 5446 726 5474 754
rect 5474 726 5476 754
rect 5444 724 5476 726
rect 5444 674 5476 676
rect 5444 646 5446 674
rect 5446 646 5474 674
rect 5474 646 5476 674
rect 5444 644 5476 646
rect 5444 594 5476 596
rect 5444 566 5446 594
rect 5446 566 5474 594
rect 5474 566 5476 594
rect 5444 564 5476 566
rect 5444 194 5476 196
rect 5444 166 5446 194
rect 5446 166 5474 194
rect 5474 166 5476 194
rect 5444 164 5476 166
rect 5444 114 5476 116
rect 5444 86 5446 114
rect 5446 86 5474 114
rect 5474 86 5476 114
rect 5444 84 5476 86
rect 5444 34 5476 36
rect 5444 6 5446 34
rect 5446 6 5474 34
rect 5474 6 5476 34
rect 5444 4 5476 6
rect 5604 15364 5636 15396
rect 10164 15364 10196 15396
rect 5684 15284 5716 15316
rect 6724 15284 6756 15316
rect 6804 15284 6836 15316
rect 7844 15284 7876 15316
rect 7924 15284 7956 15316
rect 8964 15284 8996 15316
rect 9044 15284 9076 15316
rect 10084 15284 10116 15316
rect 5604 14084 5636 14116
rect 10164 14084 10196 14116
rect 5524 14004 5556 14036
rect 5524 13684 5556 13716
rect 10244 14004 10276 14036
rect 10324 16804 10356 16836
rect 10324 15524 10356 15556
rect 10324 13924 10356 13956
rect 10324 13764 10356 13796
rect 10404 16724 10436 16756
rect 10404 13844 10436 13876
rect 10484 16804 10516 16836
rect 10484 15524 10516 15556
rect 10484 13924 10516 13956
rect 10484 13764 10516 13796
rect 10564 16884 10596 16916
rect 10564 15444 10596 15476
rect 10564 14004 10596 14036
rect 10244 13684 10276 13716
rect 10564 13684 10596 13716
rect 5524 13364 5556 13396
rect 5524 13324 5556 13356
rect 5524 13284 5556 13316
rect 5524 13244 5556 13276
rect 5524 13204 5556 13236
rect 5684 13364 5716 13396
rect 5684 13324 5716 13356
rect 5684 13284 5716 13316
rect 5684 13244 5716 13276
rect 5684 13204 5716 13236
rect 5524 12634 5556 12636
rect 5524 12606 5526 12634
rect 5526 12606 5554 12634
rect 5554 12606 5556 12634
rect 5524 12604 5556 12606
rect 5524 12554 5556 12556
rect 5524 12526 5526 12554
rect 5526 12526 5554 12554
rect 5554 12526 5556 12554
rect 5524 12524 5556 12526
rect 5524 12474 5556 12476
rect 5524 12446 5526 12474
rect 5526 12446 5554 12474
rect 5554 12446 5556 12474
rect 5524 12444 5556 12446
rect 5524 12394 5556 12396
rect 5524 12366 5526 12394
rect 5526 12366 5554 12394
rect 5554 12366 5556 12394
rect 5524 12364 5556 12366
rect 5524 12314 5556 12316
rect 5524 12286 5526 12314
rect 5526 12286 5554 12314
rect 5554 12286 5556 12314
rect 5524 12284 5556 12286
rect 5524 12234 5556 12236
rect 5524 12206 5526 12234
rect 5526 12206 5554 12234
rect 5554 12206 5556 12234
rect 5524 12204 5556 12206
rect 5524 12154 5556 12156
rect 5524 12126 5526 12154
rect 5526 12126 5554 12154
rect 5554 12126 5556 12154
rect 5524 12124 5556 12126
rect 5524 11834 5556 11836
rect 5524 11806 5526 11834
rect 5526 11806 5554 11834
rect 5554 11806 5556 11834
rect 5524 11804 5556 11806
rect 5524 11754 5556 11756
rect 5524 11726 5526 11754
rect 5526 11726 5554 11754
rect 5554 11726 5556 11754
rect 5524 11724 5556 11726
rect 5524 11674 5556 11676
rect 5524 11646 5526 11674
rect 5526 11646 5554 11674
rect 5554 11646 5556 11674
rect 5524 11644 5556 11646
rect 5524 11594 5556 11596
rect 5524 11566 5526 11594
rect 5526 11566 5554 11594
rect 5554 11566 5556 11594
rect 5524 11564 5556 11566
rect 5524 11514 5556 11516
rect 5524 11486 5526 11514
rect 5526 11486 5554 11514
rect 5554 11486 5556 11514
rect 5524 11484 5556 11486
rect 5524 11434 5556 11436
rect 5524 11406 5526 11434
rect 5526 11406 5554 11434
rect 5554 11406 5556 11434
rect 5524 11404 5556 11406
rect 5524 10874 5556 10876
rect 5524 10846 5526 10874
rect 5526 10846 5554 10874
rect 5554 10846 5556 10874
rect 5524 10844 5556 10846
rect 5524 10794 5556 10796
rect 5524 10766 5526 10794
rect 5526 10766 5554 10794
rect 5554 10766 5556 10794
rect 5524 10764 5556 10766
rect 5524 10714 5556 10716
rect 5524 10686 5526 10714
rect 5526 10686 5554 10714
rect 5554 10686 5556 10714
rect 5524 10684 5556 10686
rect 5524 10634 5556 10636
rect 5524 10606 5526 10634
rect 5526 10606 5554 10634
rect 5554 10606 5556 10634
rect 5524 10604 5556 10606
rect 5524 10554 5556 10556
rect 5524 10526 5526 10554
rect 5526 10526 5554 10554
rect 5554 10526 5556 10554
rect 5524 10524 5556 10526
rect 5524 10474 5556 10476
rect 5524 10446 5526 10474
rect 5526 10446 5554 10474
rect 5554 10446 5556 10474
rect 5524 10444 5556 10446
rect 5524 10394 5556 10396
rect 5524 10366 5526 10394
rect 5526 10366 5554 10394
rect 5554 10366 5556 10394
rect 5524 10364 5556 10366
rect 5524 10314 5556 10316
rect 5524 10286 5526 10314
rect 5526 10286 5554 10314
rect 5554 10286 5556 10314
rect 5524 10284 5556 10286
rect 5524 10234 5556 10236
rect 5524 10206 5526 10234
rect 5526 10206 5554 10234
rect 5554 10206 5556 10234
rect 5524 10204 5556 10206
rect 5524 10154 5556 10156
rect 5524 10126 5526 10154
rect 5526 10126 5554 10154
rect 5554 10126 5556 10154
rect 5524 10124 5556 10126
rect 5524 10074 5556 10076
rect 5524 10046 5526 10074
rect 5526 10046 5554 10074
rect 5554 10046 5556 10074
rect 5524 10044 5556 10046
rect 5524 9994 5556 9996
rect 5524 9966 5526 9994
rect 5526 9966 5554 9994
rect 5554 9966 5556 9994
rect 5524 9964 5556 9966
rect 5524 9914 5556 9916
rect 5524 9886 5526 9914
rect 5526 9886 5554 9914
rect 5554 9886 5556 9914
rect 5524 9884 5556 9886
rect 5524 9834 5556 9836
rect 5524 9806 5526 9834
rect 5526 9806 5554 9834
rect 5554 9806 5556 9834
rect 5524 9804 5556 9806
rect 5524 9754 5556 9756
rect 5524 9726 5526 9754
rect 5526 9726 5554 9754
rect 5554 9726 5556 9754
rect 5524 9724 5556 9726
rect 5524 9354 5556 9356
rect 5524 9326 5526 9354
rect 5526 9326 5554 9354
rect 5554 9326 5556 9354
rect 5524 9324 5556 9326
rect 5524 9274 5556 9276
rect 5524 9246 5526 9274
rect 5526 9246 5554 9274
rect 5554 9246 5556 9274
rect 5524 9244 5556 9246
rect 5524 9194 5556 9196
rect 5524 9166 5526 9194
rect 5526 9166 5554 9194
rect 5554 9166 5556 9194
rect 5524 9164 5556 9166
rect 5524 8874 5556 8876
rect 5524 8846 5526 8874
rect 5526 8846 5554 8874
rect 5554 8846 5556 8874
rect 5524 8844 5556 8846
rect 5524 8794 5556 8796
rect 5524 8766 5526 8794
rect 5526 8766 5554 8794
rect 5554 8766 5556 8794
rect 5524 8764 5556 8766
rect 5524 8714 5556 8716
rect 5524 8686 5526 8714
rect 5526 8686 5554 8714
rect 5554 8686 5556 8714
rect 5524 8684 5556 8686
rect 5524 8634 5556 8636
rect 5524 8606 5526 8634
rect 5526 8606 5554 8634
rect 5554 8606 5556 8634
rect 5524 8604 5556 8606
rect 5524 8554 5556 8556
rect 5524 8526 5526 8554
rect 5526 8526 5554 8554
rect 5554 8526 5556 8554
rect 5524 8524 5556 8526
rect 5524 7634 5556 7636
rect 5524 7606 5526 7634
rect 5526 7606 5554 7634
rect 5554 7606 5556 7634
rect 5524 7604 5556 7606
rect 5524 7554 5556 7556
rect 5524 7526 5526 7554
rect 5526 7526 5554 7554
rect 5554 7526 5556 7554
rect 5524 7524 5556 7526
rect 5524 7474 5556 7476
rect 5524 7446 5526 7474
rect 5526 7446 5554 7474
rect 5554 7446 5556 7474
rect 5524 7444 5556 7446
rect 5524 7394 5556 7396
rect 5524 7366 5526 7394
rect 5526 7366 5554 7394
rect 5554 7366 5556 7394
rect 5524 7364 5556 7366
rect 5524 7314 5556 7316
rect 5524 7286 5526 7314
rect 5526 7286 5554 7314
rect 5554 7286 5556 7314
rect 5524 7284 5556 7286
rect 5524 7234 5556 7236
rect 5524 7206 5526 7234
rect 5526 7206 5554 7234
rect 5554 7206 5556 7234
rect 5524 7204 5556 7206
rect 5524 7154 5556 7156
rect 5524 7126 5526 7154
rect 5526 7126 5554 7154
rect 5554 7126 5556 7154
rect 5524 7124 5556 7126
rect 5524 7074 5556 7076
rect 5524 7046 5526 7074
rect 5526 7046 5554 7074
rect 5554 7046 5556 7074
rect 5524 7044 5556 7046
rect 5524 6754 5556 6756
rect 5524 6726 5526 6754
rect 5526 6726 5554 6754
rect 5554 6726 5556 6754
rect 5524 6724 5556 6726
rect 5524 6674 5556 6676
rect 5524 6646 5526 6674
rect 5526 6646 5554 6674
rect 5554 6646 5556 6674
rect 5524 6644 5556 6646
rect 5524 6594 5556 6596
rect 5524 6566 5526 6594
rect 5526 6566 5554 6594
rect 5554 6566 5556 6594
rect 5524 6564 5556 6566
rect 5524 6514 5556 6516
rect 5524 6486 5526 6514
rect 5526 6486 5554 6514
rect 5554 6486 5556 6514
rect 5524 6484 5556 6486
rect 5524 6434 5556 6436
rect 5524 6406 5526 6434
rect 5526 6406 5554 6434
rect 5554 6406 5556 6434
rect 5524 6404 5556 6406
rect 5524 6354 5556 6356
rect 5524 6326 5526 6354
rect 5526 6326 5554 6354
rect 5554 6326 5556 6354
rect 5524 6324 5556 6326
rect 5524 5794 5556 5796
rect 5524 5766 5526 5794
rect 5526 5766 5554 5794
rect 5554 5766 5556 5794
rect 5524 5764 5556 5766
rect 5524 5714 5556 5716
rect 5524 5686 5526 5714
rect 5526 5686 5554 5714
rect 5554 5686 5556 5714
rect 5524 5684 5556 5686
rect 5524 5634 5556 5636
rect 5524 5606 5526 5634
rect 5526 5606 5554 5634
rect 5554 5606 5556 5634
rect 5524 5604 5556 5606
rect 5524 5554 5556 5556
rect 5524 5526 5526 5554
rect 5526 5526 5554 5554
rect 5554 5526 5556 5554
rect 5524 5524 5556 5526
rect 5524 5474 5556 5476
rect 5524 5446 5526 5474
rect 5526 5446 5554 5474
rect 5554 5446 5556 5474
rect 5524 5444 5556 5446
rect 5524 5394 5556 5396
rect 5524 5366 5526 5394
rect 5526 5366 5554 5394
rect 5554 5366 5556 5394
rect 5524 5364 5556 5366
rect 5524 5314 5556 5316
rect 5524 5286 5526 5314
rect 5526 5286 5554 5314
rect 5554 5286 5556 5314
rect 5524 5284 5556 5286
rect 5524 5234 5556 5236
rect 5524 5206 5526 5234
rect 5526 5206 5554 5234
rect 5554 5206 5556 5234
rect 5524 5204 5556 5206
rect 5524 5154 5556 5156
rect 5524 5126 5526 5154
rect 5526 5126 5554 5154
rect 5554 5126 5556 5154
rect 5524 5124 5556 5126
rect 5524 5074 5556 5076
rect 5524 5046 5526 5074
rect 5526 5046 5554 5074
rect 5554 5046 5556 5074
rect 5524 5044 5556 5046
rect 5524 4994 5556 4996
rect 5524 4966 5526 4994
rect 5526 4966 5554 4994
rect 5554 4966 5556 4994
rect 5524 4964 5556 4966
rect 5524 4434 5556 4436
rect 5524 4406 5526 4434
rect 5526 4406 5554 4434
rect 5554 4406 5556 4434
rect 5524 4404 5556 4406
rect 5524 4354 5556 4356
rect 5524 4326 5526 4354
rect 5526 4326 5554 4354
rect 5554 4326 5556 4354
rect 5524 4324 5556 4326
rect 5524 4274 5556 4276
rect 5524 4246 5526 4274
rect 5526 4246 5554 4274
rect 5554 4246 5556 4274
rect 5524 4244 5556 4246
rect 5524 4194 5556 4196
rect 5524 4166 5526 4194
rect 5526 4166 5554 4194
rect 5554 4166 5556 4194
rect 5524 4164 5556 4166
rect 5524 4114 5556 4116
rect 5524 4086 5526 4114
rect 5526 4086 5554 4114
rect 5554 4086 5556 4114
rect 5524 4084 5556 4086
rect 5524 4034 5556 4036
rect 5524 4006 5526 4034
rect 5526 4006 5554 4034
rect 5554 4006 5556 4034
rect 5524 4004 5556 4006
rect 5524 3954 5556 3956
rect 5524 3926 5526 3954
rect 5526 3926 5554 3954
rect 5554 3926 5556 3954
rect 5524 3924 5556 3926
rect 5524 3154 5556 3156
rect 5524 3126 5526 3154
rect 5526 3126 5554 3154
rect 5554 3126 5556 3154
rect 5524 3124 5556 3126
rect 5524 3074 5556 3076
rect 5524 3046 5526 3074
rect 5526 3046 5554 3074
rect 5554 3046 5556 3074
rect 5524 3044 5556 3046
rect 5524 2994 5556 2996
rect 5524 2966 5526 2994
rect 5526 2966 5554 2994
rect 5554 2966 5556 2994
rect 5524 2964 5556 2966
rect 5524 2914 5556 2916
rect 5524 2886 5526 2914
rect 5526 2886 5554 2914
rect 5554 2886 5556 2914
rect 5524 2884 5556 2886
rect 5524 2834 5556 2836
rect 5524 2806 5526 2834
rect 5526 2806 5554 2834
rect 5554 2806 5556 2834
rect 5524 2804 5556 2806
rect 5524 2754 5556 2756
rect 5524 2726 5526 2754
rect 5526 2726 5554 2754
rect 5554 2726 5556 2754
rect 5524 2724 5556 2726
rect 5524 2674 5556 2676
rect 5524 2646 5526 2674
rect 5526 2646 5554 2674
rect 5554 2646 5556 2674
rect 5524 2644 5556 2646
rect 5524 2594 5556 2596
rect 5524 2566 5526 2594
rect 5526 2566 5554 2594
rect 5554 2566 5556 2594
rect 5524 2564 5556 2566
rect 5524 2514 5556 2516
rect 5524 2486 5526 2514
rect 5526 2486 5554 2514
rect 5554 2486 5556 2514
rect 5524 2484 5556 2486
rect 5524 2434 5556 2436
rect 5524 2406 5526 2434
rect 5526 2406 5554 2434
rect 5554 2406 5556 2434
rect 5524 2404 5556 2406
rect 5524 2354 5556 2356
rect 5524 2326 5526 2354
rect 5526 2326 5554 2354
rect 5554 2326 5556 2354
rect 5524 2324 5556 2326
rect 5524 2274 5556 2276
rect 5524 2246 5526 2274
rect 5526 2246 5554 2274
rect 5554 2246 5556 2274
rect 5524 2244 5556 2246
rect 5524 2194 5556 2196
rect 5524 2166 5526 2194
rect 5526 2166 5554 2194
rect 5554 2166 5556 2194
rect 5524 2164 5556 2166
rect 5524 2114 5556 2116
rect 5524 2086 5526 2114
rect 5526 2086 5554 2114
rect 5554 2086 5556 2114
rect 5524 2084 5556 2086
rect 5524 2034 5556 2036
rect 5524 2006 5526 2034
rect 5526 2006 5554 2034
rect 5554 2006 5556 2034
rect 5524 2004 5556 2006
rect 5524 1634 5556 1636
rect 5524 1606 5526 1634
rect 5526 1606 5554 1634
rect 5554 1606 5556 1634
rect 5524 1604 5556 1606
rect 5524 1554 5556 1556
rect 5524 1526 5526 1554
rect 5526 1526 5554 1554
rect 5554 1526 5556 1554
rect 5524 1524 5556 1526
rect 5524 1474 5556 1476
rect 5524 1446 5526 1474
rect 5526 1446 5554 1474
rect 5554 1446 5556 1474
rect 5524 1444 5556 1446
rect 5524 1394 5556 1396
rect 5524 1366 5526 1394
rect 5526 1366 5554 1394
rect 5554 1366 5556 1394
rect 5524 1364 5556 1366
rect 5524 1314 5556 1316
rect 5524 1286 5526 1314
rect 5526 1286 5554 1314
rect 5554 1286 5556 1314
rect 5524 1284 5556 1286
rect 5524 1234 5556 1236
rect 5524 1206 5526 1234
rect 5526 1206 5554 1234
rect 5554 1206 5556 1234
rect 5524 1204 5556 1206
rect 5524 1154 5556 1156
rect 5524 1126 5526 1154
rect 5526 1126 5554 1154
rect 5554 1126 5556 1154
rect 5524 1124 5556 1126
rect 5524 1074 5556 1076
rect 5524 1046 5526 1074
rect 5526 1046 5554 1074
rect 5554 1046 5556 1074
rect 5524 1044 5556 1046
rect 5524 754 5556 756
rect 5524 726 5526 754
rect 5526 726 5554 754
rect 5554 726 5556 754
rect 5524 724 5556 726
rect 5524 674 5556 676
rect 5524 646 5526 674
rect 5526 646 5554 674
rect 5554 646 5556 674
rect 5524 644 5556 646
rect 5524 594 5556 596
rect 5524 566 5526 594
rect 5526 566 5554 594
rect 5554 566 5556 594
rect 5524 564 5556 566
rect 5524 194 5556 196
rect 5524 166 5526 194
rect 5526 166 5554 194
rect 5554 166 5556 194
rect 5524 164 5556 166
rect 5524 114 5556 116
rect 5524 86 5526 114
rect 5526 86 5554 114
rect 5554 86 5556 114
rect 5524 84 5556 86
rect 5524 34 5556 36
rect 5524 6 5526 34
rect 5526 6 5554 34
rect 5554 6 5556 34
rect 5524 4 5556 6
rect 5844 13364 5876 13396
rect 5844 13324 5876 13356
rect 5844 13284 5876 13316
rect 5844 13244 5876 13276
rect 5844 13204 5876 13236
rect 5684 12634 5716 12636
rect 5684 12606 5686 12634
rect 5686 12606 5714 12634
rect 5714 12606 5716 12634
rect 5684 12604 5716 12606
rect 5684 12554 5716 12556
rect 5684 12526 5686 12554
rect 5686 12526 5714 12554
rect 5714 12526 5716 12554
rect 5684 12524 5716 12526
rect 5684 12474 5716 12476
rect 5684 12446 5686 12474
rect 5686 12446 5714 12474
rect 5714 12446 5716 12474
rect 5684 12444 5716 12446
rect 5684 12394 5716 12396
rect 5684 12366 5686 12394
rect 5686 12366 5714 12394
rect 5714 12366 5716 12394
rect 5684 12364 5716 12366
rect 5684 12314 5716 12316
rect 5684 12286 5686 12314
rect 5686 12286 5714 12314
rect 5714 12286 5716 12314
rect 5684 12284 5716 12286
rect 5684 12234 5716 12236
rect 5684 12206 5686 12234
rect 5686 12206 5714 12234
rect 5714 12206 5716 12234
rect 5684 12204 5716 12206
rect 5684 12154 5716 12156
rect 5684 12126 5686 12154
rect 5686 12126 5714 12154
rect 5714 12126 5716 12154
rect 5684 12124 5716 12126
rect 5684 11834 5716 11836
rect 5684 11806 5686 11834
rect 5686 11806 5714 11834
rect 5714 11806 5716 11834
rect 5684 11804 5716 11806
rect 5684 11754 5716 11756
rect 5684 11726 5686 11754
rect 5686 11726 5714 11754
rect 5714 11726 5716 11754
rect 5684 11724 5716 11726
rect 5684 11674 5716 11676
rect 5684 11646 5686 11674
rect 5686 11646 5714 11674
rect 5714 11646 5716 11674
rect 5684 11644 5716 11646
rect 5684 11594 5716 11596
rect 5684 11566 5686 11594
rect 5686 11566 5714 11594
rect 5714 11566 5716 11594
rect 5684 11564 5716 11566
rect 5684 11514 5716 11516
rect 5684 11486 5686 11514
rect 5686 11486 5714 11514
rect 5714 11486 5716 11514
rect 5684 11484 5716 11486
rect 5684 11434 5716 11436
rect 5684 11406 5686 11434
rect 5686 11406 5714 11434
rect 5714 11406 5716 11434
rect 5684 11404 5716 11406
rect 5684 10874 5716 10876
rect 5684 10846 5686 10874
rect 5686 10846 5714 10874
rect 5714 10846 5716 10874
rect 5684 10844 5716 10846
rect 5684 10794 5716 10796
rect 5684 10766 5686 10794
rect 5686 10766 5714 10794
rect 5714 10766 5716 10794
rect 5684 10764 5716 10766
rect 5684 10714 5716 10716
rect 5684 10686 5686 10714
rect 5686 10686 5714 10714
rect 5714 10686 5716 10714
rect 5684 10684 5716 10686
rect 5684 10634 5716 10636
rect 5684 10606 5686 10634
rect 5686 10606 5714 10634
rect 5714 10606 5716 10634
rect 5684 10604 5716 10606
rect 5684 10554 5716 10556
rect 5684 10526 5686 10554
rect 5686 10526 5714 10554
rect 5714 10526 5716 10554
rect 5684 10524 5716 10526
rect 5684 10474 5716 10476
rect 5684 10446 5686 10474
rect 5686 10446 5714 10474
rect 5714 10446 5716 10474
rect 5684 10444 5716 10446
rect 5684 10394 5716 10396
rect 5684 10366 5686 10394
rect 5686 10366 5714 10394
rect 5714 10366 5716 10394
rect 5684 10364 5716 10366
rect 5684 10314 5716 10316
rect 5684 10286 5686 10314
rect 5686 10286 5714 10314
rect 5714 10286 5716 10314
rect 5684 10284 5716 10286
rect 5684 10234 5716 10236
rect 5684 10206 5686 10234
rect 5686 10206 5714 10234
rect 5714 10206 5716 10234
rect 5684 10204 5716 10206
rect 5684 10154 5716 10156
rect 5684 10126 5686 10154
rect 5686 10126 5714 10154
rect 5714 10126 5716 10154
rect 5684 10124 5716 10126
rect 5684 10074 5716 10076
rect 5684 10046 5686 10074
rect 5686 10046 5714 10074
rect 5714 10046 5716 10074
rect 5684 10044 5716 10046
rect 5684 9994 5716 9996
rect 5684 9966 5686 9994
rect 5686 9966 5714 9994
rect 5714 9966 5716 9994
rect 5684 9964 5716 9966
rect 5684 9914 5716 9916
rect 5684 9886 5686 9914
rect 5686 9886 5714 9914
rect 5714 9886 5716 9914
rect 5684 9884 5716 9886
rect 5684 9834 5716 9836
rect 5684 9806 5686 9834
rect 5686 9806 5714 9834
rect 5714 9806 5716 9834
rect 5684 9804 5716 9806
rect 5684 9754 5716 9756
rect 5684 9726 5686 9754
rect 5686 9726 5714 9754
rect 5714 9726 5716 9754
rect 5684 9724 5716 9726
rect 5684 9354 5716 9356
rect 5684 9326 5686 9354
rect 5686 9326 5714 9354
rect 5714 9326 5716 9354
rect 5684 9324 5716 9326
rect 5684 9274 5716 9276
rect 5684 9246 5686 9274
rect 5686 9246 5714 9274
rect 5714 9246 5716 9274
rect 5684 9244 5716 9246
rect 5684 9194 5716 9196
rect 5684 9166 5686 9194
rect 5686 9166 5714 9194
rect 5714 9166 5716 9194
rect 5684 9164 5716 9166
rect 5684 8874 5716 8876
rect 5684 8846 5686 8874
rect 5686 8846 5714 8874
rect 5714 8846 5716 8874
rect 5684 8844 5716 8846
rect 5684 8794 5716 8796
rect 5684 8766 5686 8794
rect 5686 8766 5714 8794
rect 5714 8766 5716 8794
rect 5684 8764 5716 8766
rect 5684 8714 5716 8716
rect 5684 8686 5686 8714
rect 5686 8686 5714 8714
rect 5714 8686 5716 8714
rect 5684 8684 5716 8686
rect 5684 8634 5716 8636
rect 5684 8606 5686 8634
rect 5686 8606 5714 8634
rect 5714 8606 5716 8634
rect 5684 8604 5716 8606
rect 5684 8554 5716 8556
rect 5684 8526 5686 8554
rect 5686 8526 5714 8554
rect 5714 8526 5716 8554
rect 5684 8524 5716 8526
rect 5684 7634 5716 7636
rect 5684 7606 5686 7634
rect 5686 7606 5714 7634
rect 5714 7606 5716 7634
rect 5684 7604 5716 7606
rect 5684 7554 5716 7556
rect 5684 7526 5686 7554
rect 5686 7526 5714 7554
rect 5714 7526 5716 7554
rect 5684 7524 5716 7526
rect 5684 7474 5716 7476
rect 5684 7446 5686 7474
rect 5686 7446 5714 7474
rect 5714 7446 5716 7474
rect 5684 7444 5716 7446
rect 5684 7394 5716 7396
rect 5684 7366 5686 7394
rect 5686 7366 5714 7394
rect 5714 7366 5716 7394
rect 5684 7364 5716 7366
rect 5684 7314 5716 7316
rect 5684 7286 5686 7314
rect 5686 7286 5714 7314
rect 5714 7286 5716 7314
rect 5684 7284 5716 7286
rect 5684 7234 5716 7236
rect 5684 7206 5686 7234
rect 5686 7206 5714 7234
rect 5714 7206 5716 7234
rect 5684 7204 5716 7206
rect 5684 7154 5716 7156
rect 5684 7126 5686 7154
rect 5686 7126 5714 7154
rect 5714 7126 5716 7154
rect 5684 7124 5716 7126
rect 5684 7074 5716 7076
rect 5684 7046 5686 7074
rect 5686 7046 5714 7074
rect 5714 7046 5716 7074
rect 5684 7044 5716 7046
rect 5684 6754 5716 6756
rect 5684 6726 5686 6754
rect 5686 6726 5714 6754
rect 5714 6726 5716 6754
rect 5684 6724 5716 6726
rect 5684 6674 5716 6676
rect 5684 6646 5686 6674
rect 5686 6646 5714 6674
rect 5714 6646 5716 6674
rect 5684 6644 5716 6646
rect 5684 6594 5716 6596
rect 5684 6566 5686 6594
rect 5686 6566 5714 6594
rect 5714 6566 5716 6594
rect 5684 6564 5716 6566
rect 5684 6514 5716 6516
rect 5684 6486 5686 6514
rect 5686 6486 5714 6514
rect 5714 6486 5716 6514
rect 5684 6484 5716 6486
rect 5684 6434 5716 6436
rect 5684 6406 5686 6434
rect 5686 6406 5714 6434
rect 5714 6406 5716 6434
rect 5684 6404 5716 6406
rect 5684 6354 5716 6356
rect 5684 6326 5686 6354
rect 5686 6326 5714 6354
rect 5714 6326 5716 6354
rect 5684 6324 5716 6326
rect 5684 5794 5716 5796
rect 5684 5766 5686 5794
rect 5686 5766 5714 5794
rect 5714 5766 5716 5794
rect 5684 5764 5716 5766
rect 5684 5714 5716 5716
rect 5684 5686 5686 5714
rect 5686 5686 5714 5714
rect 5714 5686 5716 5714
rect 5684 5684 5716 5686
rect 5684 5634 5716 5636
rect 5684 5606 5686 5634
rect 5686 5606 5714 5634
rect 5714 5606 5716 5634
rect 5684 5604 5716 5606
rect 5684 5554 5716 5556
rect 5684 5526 5686 5554
rect 5686 5526 5714 5554
rect 5714 5526 5716 5554
rect 5684 5524 5716 5526
rect 5684 5474 5716 5476
rect 5684 5446 5686 5474
rect 5686 5446 5714 5474
rect 5714 5446 5716 5474
rect 5684 5444 5716 5446
rect 5684 5394 5716 5396
rect 5684 5366 5686 5394
rect 5686 5366 5714 5394
rect 5714 5366 5716 5394
rect 5684 5364 5716 5366
rect 5684 5314 5716 5316
rect 5684 5286 5686 5314
rect 5686 5286 5714 5314
rect 5714 5286 5716 5314
rect 5684 5284 5716 5286
rect 5684 5234 5716 5236
rect 5684 5206 5686 5234
rect 5686 5206 5714 5234
rect 5714 5206 5716 5234
rect 5684 5204 5716 5206
rect 5684 5154 5716 5156
rect 5684 5126 5686 5154
rect 5686 5126 5714 5154
rect 5714 5126 5716 5154
rect 5684 5124 5716 5126
rect 5684 5074 5716 5076
rect 5684 5046 5686 5074
rect 5686 5046 5714 5074
rect 5714 5046 5716 5074
rect 5684 5044 5716 5046
rect 5684 4994 5716 4996
rect 5684 4966 5686 4994
rect 5686 4966 5714 4994
rect 5714 4966 5716 4994
rect 5684 4964 5716 4966
rect 5684 4434 5716 4436
rect 5684 4406 5686 4434
rect 5686 4406 5714 4434
rect 5714 4406 5716 4434
rect 5684 4404 5716 4406
rect 5684 4354 5716 4356
rect 5684 4326 5686 4354
rect 5686 4326 5714 4354
rect 5714 4326 5716 4354
rect 5684 4324 5716 4326
rect 5684 4274 5716 4276
rect 5684 4246 5686 4274
rect 5686 4246 5714 4274
rect 5714 4246 5716 4274
rect 5684 4244 5716 4246
rect 5684 4194 5716 4196
rect 5684 4166 5686 4194
rect 5686 4166 5714 4194
rect 5714 4166 5716 4194
rect 5684 4164 5716 4166
rect 5684 4114 5716 4116
rect 5684 4086 5686 4114
rect 5686 4086 5714 4114
rect 5714 4086 5716 4114
rect 5684 4084 5716 4086
rect 5684 4034 5716 4036
rect 5684 4006 5686 4034
rect 5686 4006 5714 4034
rect 5714 4006 5716 4034
rect 5684 4004 5716 4006
rect 5684 3954 5716 3956
rect 5684 3926 5686 3954
rect 5686 3926 5714 3954
rect 5714 3926 5716 3954
rect 5684 3924 5716 3926
rect 5684 3154 5716 3156
rect 5684 3126 5686 3154
rect 5686 3126 5714 3154
rect 5714 3126 5716 3154
rect 5684 3124 5716 3126
rect 5684 3074 5716 3076
rect 5684 3046 5686 3074
rect 5686 3046 5714 3074
rect 5714 3046 5716 3074
rect 5684 3044 5716 3046
rect 5684 2994 5716 2996
rect 5684 2966 5686 2994
rect 5686 2966 5714 2994
rect 5714 2966 5716 2994
rect 5684 2964 5716 2966
rect 5684 2914 5716 2916
rect 5684 2886 5686 2914
rect 5686 2886 5714 2914
rect 5714 2886 5716 2914
rect 5684 2884 5716 2886
rect 5684 2834 5716 2836
rect 5684 2806 5686 2834
rect 5686 2806 5714 2834
rect 5714 2806 5716 2834
rect 5684 2804 5716 2806
rect 5684 2754 5716 2756
rect 5684 2726 5686 2754
rect 5686 2726 5714 2754
rect 5714 2726 5716 2754
rect 5684 2724 5716 2726
rect 5684 2674 5716 2676
rect 5684 2646 5686 2674
rect 5686 2646 5714 2674
rect 5714 2646 5716 2674
rect 5684 2644 5716 2646
rect 5684 2594 5716 2596
rect 5684 2566 5686 2594
rect 5686 2566 5714 2594
rect 5714 2566 5716 2594
rect 5684 2564 5716 2566
rect 5684 2514 5716 2516
rect 5684 2486 5686 2514
rect 5686 2486 5714 2514
rect 5714 2486 5716 2514
rect 5684 2484 5716 2486
rect 5684 2434 5716 2436
rect 5684 2406 5686 2434
rect 5686 2406 5714 2434
rect 5714 2406 5716 2434
rect 5684 2404 5716 2406
rect 5684 2354 5716 2356
rect 5684 2326 5686 2354
rect 5686 2326 5714 2354
rect 5714 2326 5716 2354
rect 5684 2324 5716 2326
rect 5684 2274 5716 2276
rect 5684 2246 5686 2274
rect 5686 2246 5714 2274
rect 5714 2246 5716 2274
rect 5684 2244 5716 2246
rect 5684 2194 5716 2196
rect 5684 2166 5686 2194
rect 5686 2166 5714 2194
rect 5714 2166 5716 2194
rect 5684 2164 5716 2166
rect 5684 2114 5716 2116
rect 5684 2086 5686 2114
rect 5686 2086 5714 2114
rect 5714 2086 5716 2114
rect 5684 2084 5716 2086
rect 5684 2034 5716 2036
rect 5684 2006 5686 2034
rect 5686 2006 5714 2034
rect 5714 2006 5716 2034
rect 5684 2004 5716 2006
rect 5684 1634 5716 1636
rect 5684 1606 5686 1634
rect 5686 1606 5714 1634
rect 5714 1606 5716 1634
rect 5684 1604 5716 1606
rect 5684 1554 5716 1556
rect 5684 1526 5686 1554
rect 5686 1526 5714 1554
rect 5714 1526 5716 1554
rect 5684 1524 5716 1526
rect 5684 1474 5716 1476
rect 5684 1446 5686 1474
rect 5686 1446 5714 1474
rect 5714 1446 5716 1474
rect 5684 1444 5716 1446
rect 5684 1394 5716 1396
rect 5684 1366 5686 1394
rect 5686 1366 5714 1394
rect 5714 1366 5716 1394
rect 5684 1364 5716 1366
rect 5684 1314 5716 1316
rect 5684 1286 5686 1314
rect 5686 1286 5714 1314
rect 5714 1286 5716 1314
rect 5684 1284 5716 1286
rect 5684 1234 5716 1236
rect 5684 1206 5686 1234
rect 5686 1206 5714 1234
rect 5714 1206 5716 1234
rect 5684 1204 5716 1206
rect 5684 1154 5716 1156
rect 5684 1126 5686 1154
rect 5686 1126 5714 1154
rect 5714 1126 5716 1154
rect 5684 1124 5716 1126
rect 5684 1074 5716 1076
rect 5684 1046 5686 1074
rect 5686 1046 5714 1074
rect 5714 1046 5716 1074
rect 5684 1044 5716 1046
rect 5684 754 5716 756
rect 5684 726 5686 754
rect 5686 726 5714 754
rect 5714 726 5716 754
rect 5684 724 5716 726
rect 5684 674 5716 676
rect 5684 646 5686 674
rect 5686 646 5714 674
rect 5714 646 5716 674
rect 5684 644 5716 646
rect 5684 594 5716 596
rect 5684 566 5686 594
rect 5686 566 5714 594
rect 5714 566 5716 594
rect 5684 564 5716 566
rect 5684 194 5716 196
rect 5684 166 5686 194
rect 5686 166 5714 194
rect 5714 166 5716 194
rect 5684 164 5716 166
rect 5684 114 5716 116
rect 5684 86 5686 114
rect 5686 86 5714 114
rect 5714 86 5716 114
rect 5684 84 5716 86
rect 5684 34 5716 36
rect 5684 6 5686 34
rect 5686 6 5714 34
rect 5714 6 5716 34
rect 5684 4 5716 6
rect 6164 13364 6196 13396
rect 6164 13324 6196 13356
rect 6164 13284 6196 13316
rect 6164 13244 6196 13276
rect 6164 13204 6196 13236
rect 5844 12634 5876 12636
rect 5844 12606 5846 12634
rect 5846 12606 5874 12634
rect 5874 12606 5876 12634
rect 5844 12604 5876 12606
rect 5844 12554 5876 12556
rect 5844 12526 5846 12554
rect 5846 12526 5874 12554
rect 5874 12526 5876 12554
rect 5844 12524 5876 12526
rect 5844 12474 5876 12476
rect 5844 12446 5846 12474
rect 5846 12446 5874 12474
rect 5874 12446 5876 12474
rect 5844 12444 5876 12446
rect 5844 12394 5876 12396
rect 5844 12366 5846 12394
rect 5846 12366 5874 12394
rect 5874 12366 5876 12394
rect 5844 12364 5876 12366
rect 5844 12314 5876 12316
rect 5844 12286 5846 12314
rect 5846 12286 5874 12314
rect 5874 12286 5876 12314
rect 5844 12284 5876 12286
rect 5844 12234 5876 12236
rect 5844 12206 5846 12234
rect 5846 12206 5874 12234
rect 5874 12206 5876 12234
rect 5844 12204 5876 12206
rect 5844 12154 5876 12156
rect 5844 12126 5846 12154
rect 5846 12126 5874 12154
rect 5874 12126 5876 12154
rect 5844 12124 5876 12126
rect 5844 11834 5876 11836
rect 5844 11806 5846 11834
rect 5846 11806 5874 11834
rect 5874 11806 5876 11834
rect 5844 11804 5876 11806
rect 5844 11754 5876 11756
rect 5844 11726 5846 11754
rect 5846 11726 5874 11754
rect 5874 11726 5876 11754
rect 5844 11724 5876 11726
rect 5844 11674 5876 11676
rect 5844 11646 5846 11674
rect 5846 11646 5874 11674
rect 5874 11646 5876 11674
rect 5844 11644 5876 11646
rect 5844 11594 5876 11596
rect 5844 11566 5846 11594
rect 5846 11566 5874 11594
rect 5874 11566 5876 11594
rect 5844 11564 5876 11566
rect 5844 11514 5876 11516
rect 5844 11486 5846 11514
rect 5846 11486 5874 11514
rect 5874 11486 5876 11514
rect 5844 11484 5876 11486
rect 5844 11434 5876 11436
rect 5844 11406 5846 11434
rect 5846 11406 5874 11434
rect 5874 11406 5876 11434
rect 5844 11404 5876 11406
rect 5844 10874 5876 10876
rect 5844 10846 5846 10874
rect 5846 10846 5874 10874
rect 5874 10846 5876 10874
rect 5844 10844 5876 10846
rect 5844 10794 5876 10796
rect 5844 10766 5846 10794
rect 5846 10766 5874 10794
rect 5874 10766 5876 10794
rect 5844 10764 5876 10766
rect 5844 10714 5876 10716
rect 5844 10686 5846 10714
rect 5846 10686 5874 10714
rect 5874 10686 5876 10714
rect 5844 10684 5876 10686
rect 5844 10634 5876 10636
rect 5844 10606 5846 10634
rect 5846 10606 5874 10634
rect 5874 10606 5876 10634
rect 5844 10604 5876 10606
rect 5844 10554 5876 10556
rect 5844 10526 5846 10554
rect 5846 10526 5874 10554
rect 5874 10526 5876 10554
rect 5844 10524 5876 10526
rect 5844 10474 5876 10476
rect 5844 10446 5846 10474
rect 5846 10446 5874 10474
rect 5874 10446 5876 10474
rect 5844 10444 5876 10446
rect 5844 10394 5876 10396
rect 5844 10366 5846 10394
rect 5846 10366 5874 10394
rect 5874 10366 5876 10394
rect 5844 10364 5876 10366
rect 5844 10314 5876 10316
rect 5844 10286 5846 10314
rect 5846 10286 5874 10314
rect 5874 10286 5876 10314
rect 5844 10284 5876 10286
rect 5844 10234 5876 10236
rect 5844 10206 5846 10234
rect 5846 10206 5874 10234
rect 5874 10206 5876 10234
rect 5844 10204 5876 10206
rect 5844 10154 5876 10156
rect 5844 10126 5846 10154
rect 5846 10126 5874 10154
rect 5874 10126 5876 10154
rect 5844 10124 5876 10126
rect 5844 10074 5876 10076
rect 5844 10046 5846 10074
rect 5846 10046 5874 10074
rect 5874 10046 5876 10074
rect 5844 10044 5876 10046
rect 5844 9994 5876 9996
rect 5844 9966 5846 9994
rect 5846 9966 5874 9994
rect 5874 9966 5876 9994
rect 5844 9964 5876 9966
rect 5844 9914 5876 9916
rect 5844 9886 5846 9914
rect 5846 9886 5874 9914
rect 5874 9886 5876 9914
rect 5844 9884 5876 9886
rect 5844 9834 5876 9836
rect 5844 9806 5846 9834
rect 5846 9806 5874 9834
rect 5874 9806 5876 9834
rect 5844 9804 5876 9806
rect 5844 9754 5876 9756
rect 5844 9726 5846 9754
rect 5846 9726 5874 9754
rect 5874 9726 5876 9754
rect 5844 9724 5876 9726
rect 5844 9354 5876 9356
rect 5844 9326 5846 9354
rect 5846 9326 5874 9354
rect 5874 9326 5876 9354
rect 5844 9324 5876 9326
rect 5844 9274 5876 9276
rect 5844 9246 5846 9274
rect 5846 9246 5874 9274
rect 5874 9246 5876 9274
rect 5844 9244 5876 9246
rect 5844 9194 5876 9196
rect 5844 9166 5846 9194
rect 5846 9166 5874 9194
rect 5874 9166 5876 9194
rect 5844 9164 5876 9166
rect 5844 8874 5876 8876
rect 5844 8846 5846 8874
rect 5846 8846 5874 8874
rect 5874 8846 5876 8874
rect 5844 8844 5876 8846
rect 5844 8794 5876 8796
rect 5844 8766 5846 8794
rect 5846 8766 5874 8794
rect 5874 8766 5876 8794
rect 5844 8764 5876 8766
rect 5844 8714 5876 8716
rect 5844 8686 5846 8714
rect 5846 8686 5874 8714
rect 5874 8686 5876 8714
rect 5844 8684 5876 8686
rect 5844 8634 5876 8636
rect 5844 8606 5846 8634
rect 5846 8606 5874 8634
rect 5874 8606 5876 8634
rect 5844 8604 5876 8606
rect 5844 8554 5876 8556
rect 5844 8526 5846 8554
rect 5846 8526 5874 8554
rect 5874 8526 5876 8554
rect 5844 8524 5876 8526
rect 5844 7634 5876 7636
rect 5844 7606 5846 7634
rect 5846 7606 5874 7634
rect 5874 7606 5876 7634
rect 5844 7604 5876 7606
rect 5844 7554 5876 7556
rect 5844 7526 5846 7554
rect 5846 7526 5874 7554
rect 5874 7526 5876 7554
rect 5844 7524 5876 7526
rect 5844 7474 5876 7476
rect 5844 7446 5846 7474
rect 5846 7446 5874 7474
rect 5874 7446 5876 7474
rect 5844 7444 5876 7446
rect 5844 7394 5876 7396
rect 5844 7366 5846 7394
rect 5846 7366 5874 7394
rect 5874 7366 5876 7394
rect 5844 7364 5876 7366
rect 5844 7314 5876 7316
rect 5844 7286 5846 7314
rect 5846 7286 5874 7314
rect 5874 7286 5876 7314
rect 5844 7284 5876 7286
rect 5844 7234 5876 7236
rect 5844 7206 5846 7234
rect 5846 7206 5874 7234
rect 5874 7206 5876 7234
rect 5844 7204 5876 7206
rect 5844 7154 5876 7156
rect 5844 7126 5846 7154
rect 5846 7126 5874 7154
rect 5874 7126 5876 7154
rect 5844 7124 5876 7126
rect 5844 7074 5876 7076
rect 5844 7046 5846 7074
rect 5846 7046 5874 7074
rect 5874 7046 5876 7074
rect 5844 7044 5876 7046
rect 5844 6754 5876 6756
rect 5844 6726 5846 6754
rect 5846 6726 5874 6754
rect 5874 6726 5876 6754
rect 5844 6724 5876 6726
rect 5844 6674 5876 6676
rect 5844 6646 5846 6674
rect 5846 6646 5874 6674
rect 5874 6646 5876 6674
rect 5844 6644 5876 6646
rect 5844 6594 5876 6596
rect 5844 6566 5846 6594
rect 5846 6566 5874 6594
rect 5874 6566 5876 6594
rect 5844 6564 5876 6566
rect 5844 6514 5876 6516
rect 5844 6486 5846 6514
rect 5846 6486 5874 6514
rect 5874 6486 5876 6514
rect 5844 6484 5876 6486
rect 5844 6434 5876 6436
rect 5844 6406 5846 6434
rect 5846 6406 5874 6434
rect 5874 6406 5876 6434
rect 5844 6404 5876 6406
rect 5844 6354 5876 6356
rect 5844 6326 5846 6354
rect 5846 6326 5874 6354
rect 5874 6326 5876 6354
rect 5844 6324 5876 6326
rect 5844 5794 5876 5796
rect 5844 5766 5846 5794
rect 5846 5766 5874 5794
rect 5874 5766 5876 5794
rect 5844 5764 5876 5766
rect 5844 5714 5876 5716
rect 5844 5686 5846 5714
rect 5846 5686 5874 5714
rect 5874 5686 5876 5714
rect 5844 5684 5876 5686
rect 5844 5634 5876 5636
rect 5844 5606 5846 5634
rect 5846 5606 5874 5634
rect 5874 5606 5876 5634
rect 5844 5604 5876 5606
rect 5844 5554 5876 5556
rect 5844 5526 5846 5554
rect 5846 5526 5874 5554
rect 5874 5526 5876 5554
rect 5844 5524 5876 5526
rect 5844 5474 5876 5476
rect 5844 5446 5846 5474
rect 5846 5446 5874 5474
rect 5874 5446 5876 5474
rect 5844 5444 5876 5446
rect 5844 5394 5876 5396
rect 5844 5366 5846 5394
rect 5846 5366 5874 5394
rect 5874 5366 5876 5394
rect 5844 5364 5876 5366
rect 5844 5314 5876 5316
rect 5844 5286 5846 5314
rect 5846 5286 5874 5314
rect 5874 5286 5876 5314
rect 5844 5284 5876 5286
rect 5844 5234 5876 5236
rect 5844 5206 5846 5234
rect 5846 5206 5874 5234
rect 5874 5206 5876 5234
rect 5844 5204 5876 5206
rect 5844 5154 5876 5156
rect 5844 5126 5846 5154
rect 5846 5126 5874 5154
rect 5874 5126 5876 5154
rect 5844 5124 5876 5126
rect 5844 5074 5876 5076
rect 5844 5046 5846 5074
rect 5846 5046 5874 5074
rect 5874 5046 5876 5074
rect 5844 5044 5876 5046
rect 5844 4994 5876 4996
rect 5844 4966 5846 4994
rect 5846 4966 5874 4994
rect 5874 4966 5876 4994
rect 5844 4964 5876 4966
rect 5844 4434 5876 4436
rect 5844 4406 5846 4434
rect 5846 4406 5874 4434
rect 5874 4406 5876 4434
rect 5844 4404 5876 4406
rect 5844 4354 5876 4356
rect 5844 4326 5846 4354
rect 5846 4326 5874 4354
rect 5874 4326 5876 4354
rect 5844 4324 5876 4326
rect 5844 4274 5876 4276
rect 5844 4246 5846 4274
rect 5846 4246 5874 4274
rect 5874 4246 5876 4274
rect 5844 4244 5876 4246
rect 5844 4194 5876 4196
rect 5844 4166 5846 4194
rect 5846 4166 5874 4194
rect 5874 4166 5876 4194
rect 5844 4164 5876 4166
rect 5844 4114 5876 4116
rect 5844 4086 5846 4114
rect 5846 4086 5874 4114
rect 5874 4086 5876 4114
rect 5844 4084 5876 4086
rect 5844 4034 5876 4036
rect 5844 4006 5846 4034
rect 5846 4006 5874 4034
rect 5874 4006 5876 4034
rect 5844 4004 5876 4006
rect 5844 3954 5876 3956
rect 5844 3926 5846 3954
rect 5846 3926 5874 3954
rect 5874 3926 5876 3954
rect 5844 3924 5876 3926
rect 5844 3154 5876 3156
rect 5844 3126 5846 3154
rect 5846 3126 5874 3154
rect 5874 3126 5876 3154
rect 5844 3124 5876 3126
rect 5844 3074 5876 3076
rect 5844 3046 5846 3074
rect 5846 3046 5874 3074
rect 5874 3046 5876 3074
rect 5844 3044 5876 3046
rect 5844 2994 5876 2996
rect 5844 2966 5846 2994
rect 5846 2966 5874 2994
rect 5874 2966 5876 2994
rect 5844 2964 5876 2966
rect 5844 2914 5876 2916
rect 5844 2886 5846 2914
rect 5846 2886 5874 2914
rect 5874 2886 5876 2914
rect 5844 2884 5876 2886
rect 5844 2834 5876 2836
rect 5844 2806 5846 2834
rect 5846 2806 5874 2834
rect 5874 2806 5876 2834
rect 5844 2804 5876 2806
rect 5844 2754 5876 2756
rect 5844 2726 5846 2754
rect 5846 2726 5874 2754
rect 5874 2726 5876 2754
rect 5844 2724 5876 2726
rect 5844 2674 5876 2676
rect 5844 2646 5846 2674
rect 5846 2646 5874 2674
rect 5874 2646 5876 2674
rect 5844 2644 5876 2646
rect 5844 2594 5876 2596
rect 5844 2566 5846 2594
rect 5846 2566 5874 2594
rect 5874 2566 5876 2594
rect 5844 2564 5876 2566
rect 5844 2514 5876 2516
rect 5844 2486 5846 2514
rect 5846 2486 5874 2514
rect 5874 2486 5876 2514
rect 5844 2484 5876 2486
rect 5844 2434 5876 2436
rect 5844 2406 5846 2434
rect 5846 2406 5874 2434
rect 5874 2406 5876 2434
rect 5844 2404 5876 2406
rect 5844 2354 5876 2356
rect 5844 2326 5846 2354
rect 5846 2326 5874 2354
rect 5874 2326 5876 2354
rect 5844 2324 5876 2326
rect 5844 2274 5876 2276
rect 5844 2246 5846 2274
rect 5846 2246 5874 2274
rect 5874 2246 5876 2274
rect 5844 2244 5876 2246
rect 5844 2194 5876 2196
rect 5844 2166 5846 2194
rect 5846 2166 5874 2194
rect 5874 2166 5876 2194
rect 5844 2164 5876 2166
rect 5844 2114 5876 2116
rect 5844 2086 5846 2114
rect 5846 2086 5874 2114
rect 5874 2086 5876 2114
rect 5844 2084 5876 2086
rect 5844 2034 5876 2036
rect 5844 2006 5846 2034
rect 5846 2006 5874 2034
rect 5874 2006 5876 2034
rect 5844 2004 5876 2006
rect 5844 1634 5876 1636
rect 5844 1606 5846 1634
rect 5846 1606 5874 1634
rect 5874 1606 5876 1634
rect 5844 1604 5876 1606
rect 5844 1554 5876 1556
rect 5844 1526 5846 1554
rect 5846 1526 5874 1554
rect 5874 1526 5876 1554
rect 5844 1524 5876 1526
rect 5844 1474 5876 1476
rect 5844 1446 5846 1474
rect 5846 1446 5874 1474
rect 5874 1446 5876 1474
rect 5844 1444 5876 1446
rect 5844 1394 5876 1396
rect 5844 1366 5846 1394
rect 5846 1366 5874 1394
rect 5874 1366 5876 1394
rect 5844 1364 5876 1366
rect 5844 1314 5876 1316
rect 5844 1286 5846 1314
rect 5846 1286 5874 1314
rect 5874 1286 5876 1314
rect 5844 1284 5876 1286
rect 5844 1234 5876 1236
rect 5844 1206 5846 1234
rect 5846 1206 5874 1234
rect 5874 1206 5876 1234
rect 5844 1204 5876 1206
rect 5844 1154 5876 1156
rect 5844 1126 5846 1154
rect 5846 1126 5874 1154
rect 5874 1126 5876 1154
rect 5844 1124 5876 1126
rect 5844 1074 5876 1076
rect 5844 1046 5846 1074
rect 5846 1046 5874 1074
rect 5874 1046 5876 1074
rect 5844 1044 5876 1046
rect 5844 754 5876 756
rect 5844 726 5846 754
rect 5846 726 5874 754
rect 5874 726 5876 754
rect 5844 724 5876 726
rect 5844 674 5876 676
rect 5844 646 5846 674
rect 5846 646 5874 674
rect 5874 646 5876 674
rect 5844 644 5876 646
rect 5844 594 5876 596
rect 5844 566 5846 594
rect 5846 566 5874 594
rect 5874 566 5876 594
rect 5844 564 5876 566
rect 5844 194 5876 196
rect 5844 166 5846 194
rect 5846 166 5874 194
rect 5874 166 5876 194
rect 5844 164 5876 166
rect 5844 114 5876 116
rect 5844 86 5846 114
rect 5846 86 5874 114
rect 5874 86 5876 114
rect 5844 84 5876 86
rect 5844 34 5876 36
rect 5844 6 5846 34
rect 5846 6 5874 34
rect 5874 6 5876 34
rect 5844 4 5876 6
rect 5924 12884 5956 12916
rect 5924 12844 5956 12876
rect 5924 12804 5956 12836
rect 5924 12764 5956 12796
rect 5924 12724 5956 12756
rect 6084 12884 6116 12916
rect 6084 12844 6116 12876
rect 6084 12804 6116 12836
rect 6084 12764 6116 12796
rect 6084 12724 6116 12756
rect 5924 12634 5956 12636
rect 5924 12606 5926 12634
rect 5926 12606 5954 12634
rect 5954 12606 5956 12634
rect 5924 12604 5956 12606
rect 5924 12554 5956 12556
rect 5924 12526 5926 12554
rect 5926 12526 5954 12554
rect 5954 12526 5956 12554
rect 5924 12524 5956 12526
rect 5924 12474 5956 12476
rect 5924 12446 5926 12474
rect 5926 12446 5954 12474
rect 5954 12446 5956 12474
rect 5924 12444 5956 12446
rect 5924 12394 5956 12396
rect 5924 12366 5926 12394
rect 5926 12366 5954 12394
rect 5954 12366 5956 12394
rect 5924 12364 5956 12366
rect 5924 12314 5956 12316
rect 5924 12286 5926 12314
rect 5926 12286 5954 12314
rect 5954 12286 5956 12314
rect 5924 12284 5956 12286
rect 5924 12234 5956 12236
rect 5924 12206 5926 12234
rect 5926 12206 5954 12234
rect 5954 12206 5956 12234
rect 5924 12204 5956 12206
rect 5924 12154 5956 12156
rect 5924 12126 5926 12154
rect 5926 12126 5954 12154
rect 5954 12126 5956 12154
rect 5924 12124 5956 12126
rect 5924 11834 5956 11836
rect 5924 11806 5926 11834
rect 5926 11806 5954 11834
rect 5954 11806 5956 11834
rect 5924 11804 5956 11806
rect 5924 11754 5956 11756
rect 5924 11726 5926 11754
rect 5926 11726 5954 11754
rect 5954 11726 5956 11754
rect 5924 11724 5956 11726
rect 5924 11674 5956 11676
rect 5924 11646 5926 11674
rect 5926 11646 5954 11674
rect 5954 11646 5956 11674
rect 5924 11644 5956 11646
rect 5924 11594 5956 11596
rect 5924 11566 5926 11594
rect 5926 11566 5954 11594
rect 5954 11566 5956 11594
rect 5924 11564 5956 11566
rect 5924 11514 5956 11516
rect 5924 11486 5926 11514
rect 5926 11486 5954 11514
rect 5954 11486 5956 11514
rect 5924 11484 5956 11486
rect 5924 11434 5956 11436
rect 5924 11406 5926 11434
rect 5926 11406 5954 11434
rect 5954 11406 5956 11434
rect 5924 11404 5956 11406
rect 5924 10874 5956 10876
rect 5924 10846 5926 10874
rect 5926 10846 5954 10874
rect 5954 10846 5956 10874
rect 5924 10844 5956 10846
rect 5924 10794 5956 10796
rect 5924 10766 5926 10794
rect 5926 10766 5954 10794
rect 5954 10766 5956 10794
rect 5924 10764 5956 10766
rect 5924 10714 5956 10716
rect 5924 10686 5926 10714
rect 5926 10686 5954 10714
rect 5954 10686 5956 10714
rect 5924 10684 5956 10686
rect 5924 10634 5956 10636
rect 5924 10606 5926 10634
rect 5926 10606 5954 10634
rect 5954 10606 5956 10634
rect 5924 10604 5956 10606
rect 5924 10554 5956 10556
rect 5924 10526 5926 10554
rect 5926 10526 5954 10554
rect 5954 10526 5956 10554
rect 5924 10524 5956 10526
rect 5924 10474 5956 10476
rect 5924 10446 5926 10474
rect 5926 10446 5954 10474
rect 5954 10446 5956 10474
rect 5924 10444 5956 10446
rect 5924 10394 5956 10396
rect 5924 10366 5926 10394
rect 5926 10366 5954 10394
rect 5954 10366 5956 10394
rect 5924 10364 5956 10366
rect 5924 10314 5956 10316
rect 5924 10286 5926 10314
rect 5926 10286 5954 10314
rect 5954 10286 5956 10314
rect 5924 10284 5956 10286
rect 5924 10234 5956 10236
rect 5924 10206 5926 10234
rect 5926 10206 5954 10234
rect 5954 10206 5956 10234
rect 5924 10204 5956 10206
rect 5924 10154 5956 10156
rect 5924 10126 5926 10154
rect 5926 10126 5954 10154
rect 5954 10126 5956 10154
rect 5924 10124 5956 10126
rect 5924 10074 5956 10076
rect 5924 10046 5926 10074
rect 5926 10046 5954 10074
rect 5954 10046 5956 10074
rect 5924 10044 5956 10046
rect 5924 9994 5956 9996
rect 5924 9966 5926 9994
rect 5926 9966 5954 9994
rect 5954 9966 5956 9994
rect 5924 9964 5956 9966
rect 5924 9914 5956 9916
rect 5924 9886 5926 9914
rect 5926 9886 5954 9914
rect 5954 9886 5956 9914
rect 5924 9884 5956 9886
rect 5924 9834 5956 9836
rect 5924 9806 5926 9834
rect 5926 9806 5954 9834
rect 5954 9806 5956 9834
rect 5924 9804 5956 9806
rect 5924 9754 5956 9756
rect 5924 9726 5926 9754
rect 5926 9726 5954 9754
rect 5954 9726 5956 9754
rect 5924 9724 5956 9726
rect 5924 9354 5956 9356
rect 5924 9326 5926 9354
rect 5926 9326 5954 9354
rect 5954 9326 5956 9354
rect 5924 9324 5956 9326
rect 5924 9274 5956 9276
rect 5924 9246 5926 9274
rect 5926 9246 5954 9274
rect 5954 9246 5956 9274
rect 5924 9244 5956 9246
rect 5924 9194 5956 9196
rect 5924 9166 5926 9194
rect 5926 9166 5954 9194
rect 5954 9166 5956 9194
rect 5924 9164 5956 9166
rect 5924 8874 5956 8876
rect 5924 8846 5926 8874
rect 5926 8846 5954 8874
rect 5954 8846 5956 8874
rect 5924 8844 5956 8846
rect 5924 8794 5956 8796
rect 5924 8766 5926 8794
rect 5926 8766 5954 8794
rect 5954 8766 5956 8794
rect 5924 8764 5956 8766
rect 5924 8714 5956 8716
rect 5924 8686 5926 8714
rect 5926 8686 5954 8714
rect 5954 8686 5956 8714
rect 5924 8684 5956 8686
rect 5924 8634 5956 8636
rect 5924 8606 5926 8634
rect 5926 8606 5954 8634
rect 5954 8606 5956 8634
rect 5924 8604 5956 8606
rect 5924 8554 5956 8556
rect 5924 8526 5926 8554
rect 5926 8526 5954 8554
rect 5954 8526 5956 8554
rect 5924 8524 5956 8526
rect 5924 7634 5956 7636
rect 5924 7606 5926 7634
rect 5926 7606 5954 7634
rect 5954 7606 5956 7634
rect 5924 7604 5956 7606
rect 5924 7554 5956 7556
rect 5924 7526 5926 7554
rect 5926 7526 5954 7554
rect 5954 7526 5956 7554
rect 5924 7524 5956 7526
rect 5924 7474 5956 7476
rect 5924 7446 5926 7474
rect 5926 7446 5954 7474
rect 5954 7446 5956 7474
rect 5924 7444 5956 7446
rect 5924 7394 5956 7396
rect 5924 7366 5926 7394
rect 5926 7366 5954 7394
rect 5954 7366 5956 7394
rect 5924 7364 5956 7366
rect 5924 7314 5956 7316
rect 5924 7286 5926 7314
rect 5926 7286 5954 7314
rect 5954 7286 5956 7314
rect 5924 7284 5956 7286
rect 5924 7234 5956 7236
rect 5924 7206 5926 7234
rect 5926 7206 5954 7234
rect 5954 7206 5956 7234
rect 5924 7204 5956 7206
rect 5924 7154 5956 7156
rect 5924 7126 5926 7154
rect 5926 7126 5954 7154
rect 5954 7126 5956 7154
rect 5924 7124 5956 7126
rect 5924 7074 5956 7076
rect 5924 7046 5926 7074
rect 5926 7046 5954 7074
rect 5954 7046 5956 7074
rect 5924 7044 5956 7046
rect 5924 6754 5956 6756
rect 5924 6726 5926 6754
rect 5926 6726 5954 6754
rect 5954 6726 5956 6754
rect 5924 6724 5956 6726
rect 5924 6674 5956 6676
rect 5924 6646 5926 6674
rect 5926 6646 5954 6674
rect 5954 6646 5956 6674
rect 5924 6644 5956 6646
rect 5924 6594 5956 6596
rect 5924 6566 5926 6594
rect 5926 6566 5954 6594
rect 5954 6566 5956 6594
rect 5924 6564 5956 6566
rect 5924 6514 5956 6516
rect 5924 6486 5926 6514
rect 5926 6486 5954 6514
rect 5954 6486 5956 6514
rect 5924 6484 5956 6486
rect 5924 6434 5956 6436
rect 5924 6406 5926 6434
rect 5926 6406 5954 6434
rect 5954 6406 5956 6434
rect 5924 6404 5956 6406
rect 5924 6354 5956 6356
rect 5924 6326 5926 6354
rect 5926 6326 5954 6354
rect 5954 6326 5956 6354
rect 5924 6324 5956 6326
rect 5924 5794 5956 5796
rect 5924 5766 5926 5794
rect 5926 5766 5954 5794
rect 5954 5766 5956 5794
rect 5924 5764 5956 5766
rect 5924 5714 5956 5716
rect 5924 5686 5926 5714
rect 5926 5686 5954 5714
rect 5954 5686 5956 5714
rect 5924 5684 5956 5686
rect 5924 5634 5956 5636
rect 5924 5606 5926 5634
rect 5926 5606 5954 5634
rect 5954 5606 5956 5634
rect 5924 5604 5956 5606
rect 5924 5554 5956 5556
rect 5924 5526 5926 5554
rect 5926 5526 5954 5554
rect 5954 5526 5956 5554
rect 5924 5524 5956 5526
rect 5924 5474 5956 5476
rect 5924 5446 5926 5474
rect 5926 5446 5954 5474
rect 5954 5446 5956 5474
rect 5924 5444 5956 5446
rect 5924 5394 5956 5396
rect 5924 5366 5926 5394
rect 5926 5366 5954 5394
rect 5954 5366 5956 5394
rect 5924 5364 5956 5366
rect 5924 5314 5956 5316
rect 5924 5286 5926 5314
rect 5926 5286 5954 5314
rect 5954 5286 5956 5314
rect 5924 5284 5956 5286
rect 5924 5234 5956 5236
rect 5924 5206 5926 5234
rect 5926 5206 5954 5234
rect 5954 5206 5956 5234
rect 5924 5204 5956 5206
rect 5924 5154 5956 5156
rect 5924 5126 5926 5154
rect 5926 5126 5954 5154
rect 5954 5126 5956 5154
rect 5924 5124 5956 5126
rect 5924 5074 5956 5076
rect 5924 5046 5926 5074
rect 5926 5046 5954 5074
rect 5954 5046 5956 5074
rect 5924 5044 5956 5046
rect 5924 4994 5956 4996
rect 5924 4966 5926 4994
rect 5926 4966 5954 4994
rect 5954 4966 5956 4994
rect 5924 4964 5956 4966
rect 5924 4434 5956 4436
rect 5924 4406 5926 4434
rect 5926 4406 5954 4434
rect 5954 4406 5956 4434
rect 5924 4404 5956 4406
rect 5924 4354 5956 4356
rect 5924 4326 5926 4354
rect 5926 4326 5954 4354
rect 5954 4326 5956 4354
rect 5924 4324 5956 4326
rect 5924 4274 5956 4276
rect 5924 4246 5926 4274
rect 5926 4246 5954 4274
rect 5954 4246 5956 4274
rect 5924 4244 5956 4246
rect 5924 4194 5956 4196
rect 5924 4166 5926 4194
rect 5926 4166 5954 4194
rect 5954 4166 5956 4194
rect 5924 4164 5956 4166
rect 5924 4114 5956 4116
rect 5924 4086 5926 4114
rect 5926 4086 5954 4114
rect 5954 4086 5956 4114
rect 5924 4084 5956 4086
rect 5924 4034 5956 4036
rect 5924 4006 5926 4034
rect 5926 4006 5954 4034
rect 5954 4006 5956 4034
rect 5924 4004 5956 4006
rect 5924 3954 5956 3956
rect 5924 3926 5926 3954
rect 5926 3926 5954 3954
rect 5954 3926 5956 3954
rect 5924 3924 5956 3926
rect 5924 3154 5956 3156
rect 5924 3126 5926 3154
rect 5926 3126 5954 3154
rect 5954 3126 5956 3154
rect 5924 3124 5956 3126
rect 5924 3074 5956 3076
rect 5924 3046 5926 3074
rect 5926 3046 5954 3074
rect 5954 3046 5956 3074
rect 5924 3044 5956 3046
rect 5924 2994 5956 2996
rect 5924 2966 5926 2994
rect 5926 2966 5954 2994
rect 5954 2966 5956 2994
rect 5924 2964 5956 2966
rect 5924 2914 5956 2916
rect 5924 2886 5926 2914
rect 5926 2886 5954 2914
rect 5954 2886 5956 2914
rect 5924 2884 5956 2886
rect 5924 2834 5956 2836
rect 5924 2806 5926 2834
rect 5926 2806 5954 2834
rect 5954 2806 5956 2834
rect 5924 2804 5956 2806
rect 5924 2754 5956 2756
rect 5924 2726 5926 2754
rect 5926 2726 5954 2754
rect 5954 2726 5956 2754
rect 5924 2724 5956 2726
rect 5924 2674 5956 2676
rect 5924 2646 5926 2674
rect 5926 2646 5954 2674
rect 5954 2646 5956 2674
rect 5924 2644 5956 2646
rect 5924 2594 5956 2596
rect 5924 2566 5926 2594
rect 5926 2566 5954 2594
rect 5954 2566 5956 2594
rect 5924 2564 5956 2566
rect 5924 2514 5956 2516
rect 5924 2486 5926 2514
rect 5926 2486 5954 2514
rect 5954 2486 5956 2514
rect 5924 2484 5956 2486
rect 5924 2434 5956 2436
rect 5924 2406 5926 2434
rect 5926 2406 5954 2434
rect 5954 2406 5956 2434
rect 5924 2404 5956 2406
rect 5924 2354 5956 2356
rect 5924 2326 5926 2354
rect 5926 2326 5954 2354
rect 5954 2326 5956 2354
rect 5924 2324 5956 2326
rect 5924 2274 5956 2276
rect 5924 2246 5926 2274
rect 5926 2246 5954 2274
rect 5954 2246 5956 2274
rect 5924 2244 5956 2246
rect 5924 2194 5956 2196
rect 5924 2166 5926 2194
rect 5926 2166 5954 2194
rect 5954 2166 5956 2194
rect 5924 2164 5956 2166
rect 5924 2114 5956 2116
rect 5924 2086 5926 2114
rect 5926 2086 5954 2114
rect 5954 2086 5956 2114
rect 5924 2084 5956 2086
rect 5924 2034 5956 2036
rect 5924 2006 5926 2034
rect 5926 2006 5954 2034
rect 5954 2006 5956 2034
rect 5924 2004 5956 2006
rect 5924 1634 5956 1636
rect 5924 1606 5926 1634
rect 5926 1606 5954 1634
rect 5954 1606 5956 1634
rect 5924 1604 5956 1606
rect 5924 1554 5956 1556
rect 5924 1526 5926 1554
rect 5926 1526 5954 1554
rect 5954 1526 5956 1554
rect 5924 1524 5956 1526
rect 5924 1474 5956 1476
rect 5924 1446 5926 1474
rect 5926 1446 5954 1474
rect 5954 1446 5956 1474
rect 5924 1444 5956 1446
rect 5924 1394 5956 1396
rect 5924 1366 5926 1394
rect 5926 1366 5954 1394
rect 5954 1366 5956 1394
rect 5924 1364 5956 1366
rect 5924 1314 5956 1316
rect 5924 1286 5926 1314
rect 5926 1286 5954 1314
rect 5954 1286 5956 1314
rect 5924 1284 5956 1286
rect 5924 1234 5956 1236
rect 5924 1206 5926 1234
rect 5926 1206 5954 1234
rect 5954 1206 5956 1234
rect 5924 1204 5956 1206
rect 5924 1154 5956 1156
rect 5924 1126 5926 1154
rect 5926 1126 5954 1154
rect 5954 1126 5956 1154
rect 5924 1124 5956 1126
rect 5924 1074 5956 1076
rect 5924 1046 5926 1074
rect 5926 1046 5954 1074
rect 5954 1046 5956 1074
rect 5924 1044 5956 1046
rect 5924 754 5956 756
rect 5924 726 5926 754
rect 5926 726 5954 754
rect 5954 726 5956 754
rect 5924 724 5956 726
rect 5924 674 5956 676
rect 5924 646 5926 674
rect 5926 646 5954 674
rect 5954 646 5956 674
rect 5924 644 5956 646
rect 5924 594 5956 596
rect 5924 566 5926 594
rect 5926 566 5954 594
rect 5954 566 5956 594
rect 5924 564 5956 566
rect 5924 194 5956 196
rect 5924 166 5926 194
rect 5926 166 5954 194
rect 5954 166 5956 194
rect 5924 164 5956 166
rect 5924 114 5956 116
rect 5924 86 5926 114
rect 5926 86 5954 114
rect 5954 86 5956 114
rect 5924 84 5956 86
rect 5924 34 5956 36
rect 5924 6 5926 34
rect 5926 6 5954 34
rect 5954 6 5956 34
rect 5924 4 5956 6
rect 6084 12634 6116 12636
rect 6084 12606 6086 12634
rect 6086 12606 6114 12634
rect 6114 12606 6116 12634
rect 6084 12604 6116 12606
rect 6084 12554 6116 12556
rect 6084 12526 6086 12554
rect 6086 12526 6114 12554
rect 6114 12526 6116 12554
rect 6084 12524 6116 12526
rect 6084 12474 6116 12476
rect 6084 12446 6086 12474
rect 6086 12446 6114 12474
rect 6114 12446 6116 12474
rect 6084 12444 6116 12446
rect 6084 12394 6116 12396
rect 6084 12366 6086 12394
rect 6086 12366 6114 12394
rect 6114 12366 6116 12394
rect 6084 12364 6116 12366
rect 6084 12314 6116 12316
rect 6084 12286 6086 12314
rect 6086 12286 6114 12314
rect 6114 12286 6116 12314
rect 6084 12284 6116 12286
rect 6084 12234 6116 12236
rect 6084 12206 6086 12234
rect 6086 12206 6114 12234
rect 6114 12206 6116 12234
rect 6084 12204 6116 12206
rect 6084 12154 6116 12156
rect 6084 12126 6086 12154
rect 6086 12126 6114 12154
rect 6114 12126 6116 12154
rect 6084 12124 6116 12126
rect 6084 11834 6116 11836
rect 6084 11806 6086 11834
rect 6086 11806 6114 11834
rect 6114 11806 6116 11834
rect 6084 11804 6116 11806
rect 6084 11754 6116 11756
rect 6084 11726 6086 11754
rect 6086 11726 6114 11754
rect 6114 11726 6116 11754
rect 6084 11724 6116 11726
rect 6084 11674 6116 11676
rect 6084 11646 6086 11674
rect 6086 11646 6114 11674
rect 6114 11646 6116 11674
rect 6084 11644 6116 11646
rect 6084 11594 6116 11596
rect 6084 11566 6086 11594
rect 6086 11566 6114 11594
rect 6114 11566 6116 11594
rect 6084 11564 6116 11566
rect 6084 11514 6116 11516
rect 6084 11486 6086 11514
rect 6086 11486 6114 11514
rect 6114 11486 6116 11514
rect 6084 11484 6116 11486
rect 6084 11434 6116 11436
rect 6084 11406 6086 11434
rect 6086 11406 6114 11434
rect 6114 11406 6116 11434
rect 6084 11404 6116 11406
rect 6084 10874 6116 10876
rect 6084 10846 6086 10874
rect 6086 10846 6114 10874
rect 6114 10846 6116 10874
rect 6084 10844 6116 10846
rect 6084 10794 6116 10796
rect 6084 10766 6086 10794
rect 6086 10766 6114 10794
rect 6114 10766 6116 10794
rect 6084 10764 6116 10766
rect 6084 10714 6116 10716
rect 6084 10686 6086 10714
rect 6086 10686 6114 10714
rect 6114 10686 6116 10714
rect 6084 10684 6116 10686
rect 6084 10634 6116 10636
rect 6084 10606 6086 10634
rect 6086 10606 6114 10634
rect 6114 10606 6116 10634
rect 6084 10604 6116 10606
rect 6084 10554 6116 10556
rect 6084 10526 6086 10554
rect 6086 10526 6114 10554
rect 6114 10526 6116 10554
rect 6084 10524 6116 10526
rect 6084 10474 6116 10476
rect 6084 10446 6086 10474
rect 6086 10446 6114 10474
rect 6114 10446 6116 10474
rect 6084 10444 6116 10446
rect 6084 10394 6116 10396
rect 6084 10366 6086 10394
rect 6086 10366 6114 10394
rect 6114 10366 6116 10394
rect 6084 10364 6116 10366
rect 6084 10314 6116 10316
rect 6084 10286 6086 10314
rect 6086 10286 6114 10314
rect 6114 10286 6116 10314
rect 6084 10284 6116 10286
rect 6084 10234 6116 10236
rect 6084 10206 6086 10234
rect 6086 10206 6114 10234
rect 6114 10206 6116 10234
rect 6084 10204 6116 10206
rect 6084 10154 6116 10156
rect 6084 10126 6086 10154
rect 6086 10126 6114 10154
rect 6114 10126 6116 10154
rect 6084 10124 6116 10126
rect 6084 10074 6116 10076
rect 6084 10046 6086 10074
rect 6086 10046 6114 10074
rect 6114 10046 6116 10074
rect 6084 10044 6116 10046
rect 6084 9994 6116 9996
rect 6084 9966 6086 9994
rect 6086 9966 6114 9994
rect 6114 9966 6116 9994
rect 6084 9964 6116 9966
rect 6084 9914 6116 9916
rect 6084 9886 6086 9914
rect 6086 9886 6114 9914
rect 6114 9886 6116 9914
rect 6084 9884 6116 9886
rect 6084 9834 6116 9836
rect 6084 9806 6086 9834
rect 6086 9806 6114 9834
rect 6114 9806 6116 9834
rect 6084 9804 6116 9806
rect 6084 9754 6116 9756
rect 6084 9726 6086 9754
rect 6086 9726 6114 9754
rect 6114 9726 6116 9754
rect 6084 9724 6116 9726
rect 6084 9354 6116 9356
rect 6084 9326 6086 9354
rect 6086 9326 6114 9354
rect 6114 9326 6116 9354
rect 6084 9324 6116 9326
rect 6084 9274 6116 9276
rect 6084 9246 6086 9274
rect 6086 9246 6114 9274
rect 6114 9246 6116 9274
rect 6084 9244 6116 9246
rect 6084 9194 6116 9196
rect 6084 9166 6086 9194
rect 6086 9166 6114 9194
rect 6114 9166 6116 9194
rect 6084 9164 6116 9166
rect 6084 8874 6116 8876
rect 6084 8846 6086 8874
rect 6086 8846 6114 8874
rect 6114 8846 6116 8874
rect 6084 8844 6116 8846
rect 6084 8794 6116 8796
rect 6084 8766 6086 8794
rect 6086 8766 6114 8794
rect 6114 8766 6116 8794
rect 6084 8764 6116 8766
rect 6084 8714 6116 8716
rect 6084 8686 6086 8714
rect 6086 8686 6114 8714
rect 6114 8686 6116 8714
rect 6084 8684 6116 8686
rect 6084 8634 6116 8636
rect 6084 8606 6086 8634
rect 6086 8606 6114 8634
rect 6114 8606 6116 8634
rect 6084 8604 6116 8606
rect 6084 8554 6116 8556
rect 6084 8526 6086 8554
rect 6086 8526 6114 8554
rect 6114 8526 6116 8554
rect 6084 8524 6116 8526
rect 6084 7634 6116 7636
rect 6084 7606 6086 7634
rect 6086 7606 6114 7634
rect 6114 7606 6116 7634
rect 6084 7604 6116 7606
rect 6084 7554 6116 7556
rect 6084 7526 6086 7554
rect 6086 7526 6114 7554
rect 6114 7526 6116 7554
rect 6084 7524 6116 7526
rect 6084 7474 6116 7476
rect 6084 7446 6086 7474
rect 6086 7446 6114 7474
rect 6114 7446 6116 7474
rect 6084 7444 6116 7446
rect 6084 7394 6116 7396
rect 6084 7366 6086 7394
rect 6086 7366 6114 7394
rect 6114 7366 6116 7394
rect 6084 7364 6116 7366
rect 6084 7314 6116 7316
rect 6084 7286 6086 7314
rect 6086 7286 6114 7314
rect 6114 7286 6116 7314
rect 6084 7284 6116 7286
rect 6084 7234 6116 7236
rect 6084 7206 6086 7234
rect 6086 7206 6114 7234
rect 6114 7206 6116 7234
rect 6084 7204 6116 7206
rect 6084 7154 6116 7156
rect 6084 7126 6086 7154
rect 6086 7126 6114 7154
rect 6114 7126 6116 7154
rect 6084 7124 6116 7126
rect 6084 7074 6116 7076
rect 6084 7046 6086 7074
rect 6086 7046 6114 7074
rect 6114 7046 6116 7074
rect 6084 7044 6116 7046
rect 6084 6754 6116 6756
rect 6084 6726 6086 6754
rect 6086 6726 6114 6754
rect 6114 6726 6116 6754
rect 6084 6724 6116 6726
rect 6084 6674 6116 6676
rect 6084 6646 6086 6674
rect 6086 6646 6114 6674
rect 6114 6646 6116 6674
rect 6084 6644 6116 6646
rect 6084 6594 6116 6596
rect 6084 6566 6086 6594
rect 6086 6566 6114 6594
rect 6114 6566 6116 6594
rect 6084 6564 6116 6566
rect 6084 6514 6116 6516
rect 6084 6486 6086 6514
rect 6086 6486 6114 6514
rect 6114 6486 6116 6514
rect 6084 6484 6116 6486
rect 6084 6434 6116 6436
rect 6084 6406 6086 6434
rect 6086 6406 6114 6434
rect 6114 6406 6116 6434
rect 6084 6404 6116 6406
rect 6084 6354 6116 6356
rect 6084 6326 6086 6354
rect 6086 6326 6114 6354
rect 6114 6326 6116 6354
rect 6084 6324 6116 6326
rect 6084 5794 6116 5796
rect 6084 5766 6086 5794
rect 6086 5766 6114 5794
rect 6114 5766 6116 5794
rect 6084 5764 6116 5766
rect 6084 5714 6116 5716
rect 6084 5686 6086 5714
rect 6086 5686 6114 5714
rect 6114 5686 6116 5714
rect 6084 5684 6116 5686
rect 6084 5634 6116 5636
rect 6084 5606 6086 5634
rect 6086 5606 6114 5634
rect 6114 5606 6116 5634
rect 6084 5604 6116 5606
rect 6084 5554 6116 5556
rect 6084 5526 6086 5554
rect 6086 5526 6114 5554
rect 6114 5526 6116 5554
rect 6084 5524 6116 5526
rect 6084 5474 6116 5476
rect 6084 5446 6086 5474
rect 6086 5446 6114 5474
rect 6114 5446 6116 5474
rect 6084 5444 6116 5446
rect 6084 5394 6116 5396
rect 6084 5366 6086 5394
rect 6086 5366 6114 5394
rect 6114 5366 6116 5394
rect 6084 5364 6116 5366
rect 6084 5314 6116 5316
rect 6084 5286 6086 5314
rect 6086 5286 6114 5314
rect 6114 5286 6116 5314
rect 6084 5284 6116 5286
rect 6084 5234 6116 5236
rect 6084 5206 6086 5234
rect 6086 5206 6114 5234
rect 6114 5206 6116 5234
rect 6084 5204 6116 5206
rect 6084 5154 6116 5156
rect 6084 5126 6086 5154
rect 6086 5126 6114 5154
rect 6114 5126 6116 5154
rect 6084 5124 6116 5126
rect 6084 5074 6116 5076
rect 6084 5046 6086 5074
rect 6086 5046 6114 5074
rect 6114 5046 6116 5074
rect 6084 5044 6116 5046
rect 6084 4994 6116 4996
rect 6084 4966 6086 4994
rect 6086 4966 6114 4994
rect 6114 4966 6116 4994
rect 6084 4964 6116 4966
rect 6084 4434 6116 4436
rect 6084 4406 6086 4434
rect 6086 4406 6114 4434
rect 6114 4406 6116 4434
rect 6084 4404 6116 4406
rect 6084 4354 6116 4356
rect 6084 4326 6086 4354
rect 6086 4326 6114 4354
rect 6114 4326 6116 4354
rect 6084 4324 6116 4326
rect 6084 4274 6116 4276
rect 6084 4246 6086 4274
rect 6086 4246 6114 4274
rect 6114 4246 6116 4274
rect 6084 4244 6116 4246
rect 6084 4194 6116 4196
rect 6084 4166 6086 4194
rect 6086 4166 6114 4194
rect 6114 4166 6116 4194
rect 6084 4164 6116 4166
rect 6084 4114 6116 4116
rect 6084 4086 6086 4114
rect 6086 4086 6114 4114
rect 6114 4086 6116 4114
rect 6084 4084 6116 4086
rect 6084 4034 6116 4036
rect 6084 4006 6086 4034
rect 6086 4006 6114 4034
rect 6114 4006 6116 4034
rect 6084 4004 6116 4006
rect 6084 3954 6116 3956
rect 6084 3926 6086 3954
rect 6086 3926 6114 3954
rect 6114 3926 6116 3954
rect 6084 3924 6116 3926
rect 6084 3154 6116 3156
rect 6084 3126 6086 3154
rect 6086 3126 6114 3154
rect 6114 3126 6116 3154
rect 6084 3124 6116 3126
rect 6084 3074 6116 3076
rect 6084 3046 6086 3074
rect 6086 3046 6114 3074
rect 6114 3046 6116 3074
rect 6084 3044 6116 3046
rect 6084 2994 6116 2996
rect 6084 2966 6086 2994
rect 6086 2966 6114 2994
rect 6114 2966 6116 2994
rect 6084 2964 6116 2966
rect 6084 2914 6116 2916
rect 6084 2886 6086 2914
rect 6086 2886 6114 2914
rect 6114 2886 6116 2914
rect 6084 2884 6116 2886
rect 6084 2834 6116 2836
rect 6084 2806 6086 2834
rect 6086 2806 6114 2834
rect 6114 2806 6116 2834
rect 6084 2804 6116 2806
rect 6084 2754 6116 2756
rect 6084 2726 6086 2754
rect 6086 2726 6114 2754
rect 6114 2726 6116 2754
rect 6084 2724 6116 2726
rect 6084 2674 6116 2676
rect 6084 2646 6086 2674
rect 6086 2646 6114 2674
rect 6114 2646 6116 2674
rect 6084 2644 6116 2646
rect 6084 2594 6116 2596
rect 6084 2566 6086 2594
rect 6086 2566 6114 2594
rect 6114 2566 6116 2594
rect 6084 2564 6116 2566
rect 6084 2514 6116 2516
rect 6084 2486 6086 2514
rect 6086 2486 6114 2514
rect 6114 2486 6116 2514
rect 6084 2484 6116 2486
rect 6084 2434 6116 2436
rect 6084 2406 6086 2434
rect 6086 2406 6114 2434
rect 6114 2406 6116 2434
rect 6084 2404 6116 2406
rect 6084 2354 6116 2356
rect 6084 2326 6086 2354
rect 6086 2326 6114 2354
rect 6114 2326 6116 2354
rect 6084 2324 6116 2326
rect 6084 2274 6116 2276
rect 6084 2246 6086 2274
rect 6086 2246 6114 2274
rect 6114 2246 6116 2274
rect 6084 2244 6116 2246
rect 6084 2194 6116 2196
rect 6084 2166 6086 2194
rect 6086 2166 6114 2194
rect 6114 2166 6116 2194
rect 6084 2164 6116 2166
rect 6084 2114 6116 2116
rect 6084 2086 6086 2114
rect 6086 2086 6114 2114
rect 6114 2086 6116 2114
rect 6084 2084 6116 2086
rect 6084 2034 6116 2036
rect 6084 2006 6086 2034
rect 6086 2006 6114 2034
rect 6114 2006 6116 2034
rect 6084 2004 6116 2006
rect 6084 1634 6116 1636
rect 6084 1606 6086 1634
rect 6086 1606 6114 1634
rect 6114 1606 6116 1634
rect 6084 1604 6116 1606
rect 6084 1554 6116 1556
rect 6084 1526 6086 1554
rect 6086 1526 6114 1554
rect 6114 1526 6116 1554
rect 6084 1524 6116 1526
rect 6084 1474 6116 1476
rect 6084 1446 6086 1474
rect 6086 1446 6114 1474
rect 6114 1446 6116 1474
rect 6084 1444 6116 1446
rect 6084 1394 6116 1396
rect 6084 1366 6086 1394
rect 6086 1366 6114 1394
rect 6114 1366 6116 1394
rect 6084 1364 6116 1366
rect 6084 1314 6116 1316
rect 6084 1286 6086 1314
rect 6086 1286 6114 1314
rect 6114 1286 6116 1314
rect 6084 1284 6116 1286
rect 6084 1234 6116 1236
rect 6084 1206 6086 1234
rect 6086 1206 6114 1234
rect 6114 1206 6116 1234
rect 6084 1204 6116 1206
rect 6084 1154 6116 1156
rect 6084 1126 6086 1154
rect 6086 1126 6114 1154
rect 6114 1126 6116 1154
rect 6084 1124 6116 1126
rect 6084 1074 6116 1076
rect 6084 1046 6086 1074
rect 6086 1046 6114 1074
rect 6114 1046 6116 1074
rect 6084 1044 6116 1046
rect 6084 754 6116 756
rect 6084 726 6086 754
rect 6086 726 6114 754
rect 6114 726 6116 754
rect 6084 724 6116 726
rect 6084 674 6116 676
rect 6084 646 6086 674
rect 6086 646 6114 674
rect 6114 646 6116 674
rect 6084 644 6116 646
rect 6084 594 6116 596
rect 6084 566 6086 594
rect 6086 566 6114 594
rect 6114 566 6116 594
rect 6084 564 6116 566
rect 6084 194 6116 196
rect 6084 166 6086 194
rect 6086 166 6114 194
rect 6114 166 6116 194
rect 6084 164 6116 166
rect 6084 114 6116 116
rect 6084 86 6086 114
rect 6086 86 6114 114
rect 6114 86 6116 114
rect 6084 84 6116 86
rect 6084 34 6116 36
rect 6084 6 6086 34
rect 6086 6 6114 34
rect 6114 6 6116 34
rect 6084 4 6116 6
rect 6324 13364 6356 13396
rect 6324 13324 6356 13356
rect 6324 13284 6356 13316
rect 6324 13244 6356 13276
rect 6324 13204 6356 13236
rect 6164 12634 6196 12636
rect 6164 12606 6166 12634
rect 6166 12606 6194 12634
rect 6194 12606 6196 12634
rect 6164 12604 6196 12606
rect 6164 12554 6196 12556
rect 6164 12526 6166 12554
rect 6166 12526 6194 12554
rect 6194 12526 6196 12554
rect 6164 12524 6196 12526
rect 6164 12474 6196 12476
rect 6164 12446 6166 12474
rect 6166 12446 6194 12474
rect 6194 12446 6196 12474
rect 6164 12444 6196 12446
rect 6164 12394 6196 12396
rect 6164 12366 6166 12394
rect 6166 12366 6194 12394
rect 6194 12366 6196 12394
rect 6164 12364 6196 12366
rect 6164 12314 6196 12316
rect 6164 12286 6166 12314
rect 6166 12286 6194 12314
rect 6194 12286 6196 12314
rect 6164 12284 6196 12286
rect 6164 12234 6196 12236
rect 6164 12206 6166 12234
rect 6166 12206 6194 12234
rect 6194 12206 6196 12234
rect 6164 12204 6196 12206
rect 6164 12154 6196 12156
rect 6164 12126 6166 12154
rect 6166 12126 6194 12154
rect 6194 12126 6196 12154
rect 6164 12124 6196 12126
rect 6164 11834 6196 11836
rect 6164 11806 6166 11834
rect 6166 11806 6194 11834
rect 6194 11806 6196 11834
rect 6164 11804 6196 11806
rect 6164 11754 6196 11756
rect 6164 11726 6166 11754
rect 6166 11726 6194 11754
rect 6194 11726 6196 11754
rect 6164 11724 6196 11726
rect 6164 11674 6196 11676
rect 6164 11646 6166 11674
rect 6166 11646 6194 11674
rect 6194 11646 6196 11674
rect 6164 11644 6196 11646
rect 6164 11594 6196 11596
rect 6164 11566 6166 11594
rect 6166 11566 6194 11594
rect 6194 11566 6196 11594
rect 6164 11564 6196 11566
rect 6164 11514 6196 11516
rect 6164 11486 6166 11514
rect 6166 11486 6194 11514
rect 6194 11486 6196 11514
rect 6164 11484 6196 11486
rect 6164 11434 6196 11436
rect 6164 11406 6166 11434
rect 6166 11406 6194 11434
rect 6194 11406 6196 11434
rect 6164 11404 6196 11406
rect 6164 10874 6196 10876
rect 6164 10846 6166 10874
rect 6166 10846 6194 10874
rect 6194 10846 6196 10874
rect 6164 10844 6196 10846
rect 6164 10794 6196 10796
rect 6164 10766 6166 10794
rect 6166 10766 6194 10794
rect 6194 10766 6196 10794
rect 6164 10764 6196 10766
rect 6164 10714 6196 10716
rect 6164 10686 6166 10714
rect 6166 10686 6194 10714
rect 6194 10686 6196 10714
rect 6164 10684 6196 10686
rect 6164 10634 6196 10636
rect 6164 10606 6166 10634
rect 6166 10606 6194 10634
rect 6194 10606 6196 10634
rect 6164 10604 6196 10606
rect 6164 10554 6196 10556
rect 6164 10526 6166 10554
rect 6166 10526 6194 10554
rect 6194 10526 6196 10554
rect 6164 10524 6196 10526
rect 6164 10474 6196 10476
rect 6164 10446 6166 10474
rect 6166 10446 6194 10474
rect 6194 10446 6196 10474
rect 6164 10444 6196 10446
rect 6164 10394 6196 10396
rect 6164 10366 6166 10394
rect 6166 10366 6194 10394
rect 6194 10366 6196 10394
rect 6164 10364 6196 10366
rect 6164 10314 6196 10316
rect 6164 10286 6166 10314
rect 6166 10286 6194 10314
rect 6194 10286 6196 10314
rect 6164 10284 6196 10286
rect 6164 10234 6196 10236
rect 6164 10206 6166 10234
rect 6166 10206 6194 10234
rect 6194 10206 6196 10234
rect 6164 10204 6196 10206
rect 6164 10154 6196 10156
rect 6164 10126 6166 10154
rect 6166 10126 6194 10154
rect 6194 10126 6196 10154
rect 6164 10124 6196 10126
rect 6164 10074 6196 10076
rect 6164 10046 6166 10074
rect 6166 10046 6194 10074
rect 6194 10046 6196 10074
rect 6164 10044 6196 10046
rect 6164 9994 6196 9996
rect 6164 9966 6166 9994
rect 6166 9966 6194 9994
rect 6194 9966 6196 9994
rect 6164 9964 6196 9966
rect 6164 9914 6196 9916
rect 6164 9886 6166 9914
rect 6166 9886 6194 9914
rect 6194 9886 6196 9914
rect 6164 9884 6196 9886
rect 6164 9834 6196 9836
rect 6164 9806 6166 9834
rect 6166 9806 6194 9834
rect 6194 9806 6196 9834
rect 6164 9804 6196 9806
rect 6164 9754 6196 9756
rect 6164 9726 6166 9754
rect 6166 9726 6194 9754
rect 6194 9726 6196 9754
rect 6164 9724 6196 9726
rect 6164 9354 6196 9356
rect 6164 9326 6166 9354
rect 6166 9326 6194 9354
rect 6194 9326 6196 9354
rect 6164 9324 6196 9326
rect 6164 9274 6196 9276
rect 6164 9246 6166 9274
rect 6166 9246 6194 9274
rect 6194 9246 6196 9274
rect 6164 9244 6196 9246
rect 6164 9194 6196 9196
rect 6164 9166 6166 9194
rect 6166 9166 6194 9194
rect 6194 9166 6196 9194
rect 6164 9164 6196 9166
rect 6164 8874 6196 8876
rect 6164 8846 6166 8874
rect 6166 8846 6194 8874
rect 6194 8846 6196 8874
rect 6164 8844 6196 8846
rect 6164 8794 6196 8796
rect 6164 8766 6166 8794
rect 6166 8766 6194 8794
rect 6194 8766 6196 8794
rect 6164 8764 6196 8766
rect 6164 8714 6196 8716
rect 6164 8686 6166 8714
rect 6166 8686 6194 8714
rect 6194 8686 6196 8714
rect 6164 8684 6196 8686
rect 6164 8634 6196 8636
rect 6164 8606 6166 8634
rect 6166 8606 6194 8634
rect 6194 8606 6196 8634
rect 6164 8604 6196 8606
rect 6164 8554 6196 8556
rect 6164 8526 6166 8554
rect 6166 8526 6194 8554
rect 6194 8526 6196 8554
rect 6164 8524 6196 8526
rect 6164 7634 6196 7636
rect 6164 7606 6166 7634
rect 6166 7606 6194 7634
rect 6194 7606 6196 7634
rect 6164 7604 6196 7606
rect 6164 7554 6196 7556
rect 6164 7526 6166 7554
rect 6166 7526 6194 7554
rect 6194 7526 6196 7554
rect 6164 7524 6196 7526
rect 6164 7474 6196 7476
rect 6164 7446 6166 7474
rect 6166 7446 6194 7474
rect 6194 7446 6196 7474
rect 6164 7444 6196 7446
rect 6164 7394 6196 7396
rect 6164 7366 6166 7394
rect 6166 7366 6194 7394
rect 6194 7366 6196 7394
rect 6164 7364 6196 7366
rect 6164 7314 6196 7316
rect 6164 7286 6166 7314
rect 6166 7286 6194 7314
rect 6194 7286 6196 7314
rect 6164 7284 6196 7286
rect 6164 7234 6196 7236
rect 6164 7206 6166 7234
rect 6166 7206 6194 7234
rect 6194 7206 6196 7234
rect 6164 7204 6196 7206
rect 6164 7154 6196 7156
rect 6164 7126 6166 7154
rect 6166 7126 6194 7154
rect 6194 7126 6196 7154
rect 6164 7124 6196 7126
rect 6164 7074 6196 7076
rect 6164 7046 6166 7074
rect 6166 7046 6194 7074
rect 6194 7046 6196 7074
rect 6164 7044 6196 7046
rect 6164 6754 6196 6756
rect 6164 6726 6166 6754
rect 6166 6726 6194 6754
rect 6194 6726 6196 6754
rect 6164 6724 6196 6726
rect 6164 6674 6196 6676
rect 6164 6646 6166 6674
rect 6166 6646 6194 6674
rect 6194 6646 6196 6674
rect 6164 6644 6196 6646
rect 6164 6594 6196 6596
rect 6164 6566 6166 6594
rect 6166 6566 6194 6594
rect 6194 6566 6196 6594
rect 6164 6564 6196 6566
rect 6164 6514 6196 6516
rect 6164 6486 6166 6514
rect 6166 6486 6194 6514
rect 6194 6486 6196 6514
rect 6164 6484 6196 6486
rect 6164 6434 6196 6436
rect 6164 6406 6166 6434
rect 6166 6406 6194 6434
rect 6194 6406 6196 6434
rect 6164 6404 6196 6406
rect 6164 6354 6196 6356
rect 6164 6326 6166 6354
rect 6166 6326 6194 6354
rect 6194 6326 6196 6354
rect 6164 6324 6196 6326
rect 6164 5794 6196 5796
rect 6164 5766 6166 5794
rect 6166 5766 6194 5794
rect 6194 5766 6196 5794
rect 6164 5764 6196 5766
rect 6164 5714 6196 5716
rect 6164 5686 6166 5714
rect 6166 5686 6194 5714
rect 6194 5686 6196 5714
rect 6164 5684 6196 5686
rect 6164 5634 6196 5636
rect 6164 5606 6166 5634
rect 6166 5606 6194 5634
rect 6194 5606 6196 5634
rect 6164 5604 6196 5606
rect 6164 5554 6196 5556
rect 6164 5526 6166 5554
rect 6166 5526 6194 5554
rect 6194 5526 6196 5554
rect 6164 5524 6196 5526
rect 6164 5474 6196 5476
rect 6164 5446 6166 5474
rect 6166 5446 6194 5474
rect 6194 5446 6196 5474
rect 6164 5444 6196 5446
rect 6164 5394 6196 5396
rect 6164 5366 6166 5394
rect 6166 5366 6194 5394
rect 6194 5366 6196 5394
rect 6164 5364 6196 5366
rect 6164 5314 6196 5316
rect 6164 5286 6166 5314
rect 6166 5286 6194 5314
rect 6194 5286 6196 5314
rect 6164 5284 6196 5286
rect 6164 5234 6196 5236
rect 6164 5206 6166 5234
rect 6166 5206 6194 5234
rect 6194 5206 6196 5234
rect 6164 5204 6196 5206
rect 6164 5154 6196 5156
rect 6164 5126 6166 5154
rect 6166 5126 6194 5154
rect 6194 5126 6196 5154
rect 6164 5124 6196 5126
rect 6164 5074 6196 5076
rect 6164 5046 6166 5074
rect 6166 5046 6194 5074
rect 6194 5046 6196 5074
rect 6164 5044 6196 5046
rect 6164 4994 6196 4996
rect 6164 4966 6166 4994
rect 6166 4966 6194 4994
rect 6194 4966 6196 4994
rect 6164 4964 6196 4966
rect 6164 4434 6196 4436
rect 6164 4406 6166 4434
rect 6166 4406 6194 4434
rect 6194 4406 6196 4434
rect 6164 4404 6196 4406
rect 6164 4354 6196 4356
rect 6164 4326 6166 4354
rect 6166 4326 6194 4354
rect 6194 4326 6196 4354
rect 6164 4324 6196 4326
rect 6164 4274 6196 4276
rect 6164 4246 6166 4274
rect 6166 4246 6194 4274
rect 6194 4246 6196 4274
rect 6164 4244 6196 4246
rect 6164 4194 6196 4196
rect 6164 4166 6166 4194
rect 6166 4166 6194 4194
rect 6194 4166 6196 4194
rect 6164 4164 6196 4166
rect 6164 4114 6196 4116
rect 6164 4086 6166 4114
rect 6166 4086 6194 4114
rect 6194 4086 6196 4114
rect 6164 4084 6196 4086
rect 6164 4034 6196 4036
rect 6164 4006 6166 4034
rect 6166 4006 6194 4034
rect 6194 4006 6196 4034
rect 6164 4004 6196 4006
rect 6164 3954 6196 3956
rect 6164 3926 6166 3954
rect 6166 3926 6194 3954
rect 6194 3926 6196 3954
rect 6164 3924 6196 3926
rect 6164 3154 6196 3156
rect 6164 3126 6166 3154
rect 6166 3126 6194 3154
rect 6194 3126 6196 3154
rect 6164 3124 6196 3126
rect 6164 3074 6196 3076
rect 6164 3046 6166 3074
rect 6166 3046 6194 3074
rect 6194 3046 6196 3074
rect 6164 3044 6196 3046
rect 6164 2994 6196 2996
rect 6164 2966 6166 2994
rect 6166 2966 6194 2994
rect 6194 2966 6196 2994
rect 6164 2964 6196 2966
rect 6164 2914 6196 2916
rect 6164 2886 6166 2914
rect 6166 2886 6194 2914
rect 6194 2886 6196 2914
rect 6164 2884 6196 2886
rect 6164 2834 6196 2836
rect 6164 2806 6166 2834
rect 6166 2806 6194 2834
rect 6194 2806 6196 2834
rect 6164 2804 6196 2806
rect 6164 2754 6196 2756
rect 6164 2726 6166 2754
rect 6166 2726 6194 2754
rect 6194 2726 6196 2754
rect 6164 2724 6196 2726
rect 6164 2674 6196 2676
rect 6164 2646 6166 2674
rect 6166 2646 6194 2674
rect 6194 2646 6196 2674
rect 6164 2644 6196 2646
rect 6164 2594 6196 2596
rect 6164 2566 6166 2594
rect 6166 2566 6194 2594
rect 6194 2566 6196 2594
rect 6164 2564 6196 2566
rect 6164 2514 6196 2516
rect 6164 2486 6166 2514
rect 6166 2486 6194 2514
rect 6194 2486 6196 2514
rect 6164 2484 6196 2486
rect 6164 2434 6196 2436
rect 6164 2406 6166 2434
rect 6166 2406 6194 2434
rect 6194 2406 6196 2434
rect 6164 2404 6196 2406
rect 6164 2354 6196 2356
rect 6164 2326 6166 2354
rect 6166 2326 6194 2354
rect 6194 2326 6196 2354
rect 6164 2324 6196 2326
rect 6164 2274 6196 2276
rect 6164 2246 6166 2274
rect 6166 2246 6194 2274
rect 6194 2246 6196 2274
rect 6164 2244 6196 2246
rect 6164 2194 6196 2196
rect 6164 2166 6166 2194
rect 6166 2166 6194 2194
rect 6194 2166 6196 2194
rect 6164 2164 6196 2166
rect 6164 2114 6196 2116
rect 6164 2086 6166 2114
rect 6166 2086 6194 2114
rect 6194 2086 6196 2114
rect 6164 2084 6196 2086
rect 6164 2034 6196 2036
rect 6164 2006 6166 2034
rect 6166 2006 6194 2034
rect 6194 2006 6196 2034
rect 6164 2004 6196 2006
rect 6164 1634 6196 1636
rect 6164 1606 6166 1634
rect 6166 1606 6194 1634
rect 6194 1606 6196 1634
rect 6164 1604 6196 1606
rect 6164 1554 6196 1556
rect 6164 1526 6166 1554
rect 6166 1526 6194 1554
rect 6194 1526 6196 1554
rect 6164 1524 6196 1526
rect 6164 1474 6196 1476
rect 6164 1446 6166 1474
rect 6166 1446 6194 1474
rect 6194 1446 6196 1474
rect 6164 1444 6196 1446
rect 6164 1394 6196 1396
rect 6164 1366 6166 1394
rect 6166 1366 6194 1394
rect 6194 1366 6196 1394
rect 6164 1364 6196 1366
rect 6164 1314 6196 1316
rect 6164 1286 6166 1314
rect 6166 1286 6194 1314
rect 6194 1286 6196 1314
rect 6164 1284 6196 1286
rect 6164 1234 6196 1236
rect 6164 1206 6166 1234
rect 6166 1206 6194 1234
rect 6194 1206 6196 1234
rect 6164 1204 6196 1206
rect 6164 1154 6196 1156
rect 6164 1126 6166 1154
rect 6166 1126 6194 1154
rect 6194 1126 6196 1154
rect 6164 1124 6196 1126
rect 6164 1074 6196 1076
rect 6164 1046 6166 1074
rect 6166 1046 6194 1074
rect 6194 1046 6196 1074
rect 6164 1044 6196 1046
rect 6164 754 6196 756
rect 6164 726 6166 754
rect 6166 726 6194 754
rect 6194 726 6196 754
rect 6164 724 6196 726
rect 6164 674 6196 676
rect 6164 646 6166 674
rect 6166 646 6194 674
rect 6194 646 6196 674
rect 6164 644 6196 646
rect 6164 594 6196 596
rect 6164 566 6166 594
rect 6166 566 6194 594
rect 6194 566 6196 594
rect 6164 564 6196 566
rect 6164 194 6196 196
rect 6164 166 6166 194
rect 6166 166 6194 194
rect 6194 166 6196 194
rect 6164 164 6196 166
rect 6164 114 6196 116
rect 6164 86 6166 114
rect 6166 86 6194 114
rect 6194 86 6196 114
rect 6164 84 6196 86
rect 6164 34 6196 36
rect 6164 6 6166 34
rect 6166 6 6194 34
rect 6194 6 6196 34
rect 6164 4 6196 6
rect 6324 12634 6356 12636
rect 6324 12606 6326 12634
rect 6326 12606 6354 12634
rect 6354 12606 6356 12634
rect 6324 12604 6356 12606
rect 6324 12554 6356 12556
rect 6324 12526 6326 12554
rect 6326 12526 6354 12554
rect 6354 12526 6356 12554
rect 6324 12524 6356 12526
rect 6324 12474 6356 12476
rect 6324 12446 6326 12474
rect 6326 12446 6354 12474
rect 6354 12446 6356 12474
rect 6324 12444 6356 12446
rect 6324 12394 6356 12396
rect 6324 12366 6326 12394
rect 6326 12366 6354 12394
rect 6354 12366 6356 12394
rect 6324 12364 6356 12366
rect 6324 12314 6356 12316
rect 6324 12286 6326 12314
rect 6326 12286 6354 12314
rect 6354 12286 6356 12314
rect 6324 12284 6356 12286
rect 6324 12234 6356 12236
rect 6324 12206 6326 12234
rect 6326 12206 6354 12234
rect 6354 12206 6356 12234
rect 6324 12204 6356 12206
rect 6324 12154 6356 12156
rect 6324 12126 6326 12154
rect 6326 12126 6354 12154
rect 6354 12126 6356 12154
rect 6324 12124 6356 12126
rect 6324 11834 6356 11836
rect 6324 11806 6326 11834
rect 6326 11806 6354 11834
rect 6354 11806 6356 11834
rect 6324 11804 6356 11806
rect 6324 11754 6356 11756
rect 6324 11726 6326 11754
rect 6326 11726 6354 11754
rect 6354 11726 6356 11754
rect 6324 11724 6356 11726
rect 6324 11674 6356 11676
rect 6324 11646 6326 11674
rect 6326 11646 6354 11674
rect 6354 11646 6356 11674
rect 6324 11644 6356 11646
rect 6324 11594 6356 11596
rect 6324 11566 6326 11594
rect 6326 11566 6354 11594
rect 6354 11566 6356 11594
rect 6324 11564 6356 11566
rect 6324 11514 6356 11516
rect 6324 11486 6326 11514
rect 6326 11486 6354 11514
rect 6354 11486 6356 11514
rect 6324 11484 6356 11486
rect 6324 11434 6356 11436
rect 6324 11406 6326 11434
rect 6326 11406 6354 11434
rect 6354 11406 6356 11434
rect 6324 11404 6356 11406
rect 6324 10874 6356 10876
rect 6324 10846 6326 10874
rect 6326 10846 6354 10874
rect 6354 10846 6356 10874
rect 6324 10844 6356 10846
rect 6324 10794 6356 10796
rect 6324 10766 6326 10794
rect 6326 10766 6354 10794
rect 6354 10766 6356 10794
rect 6324 10764 6356 10766
rect 6324 10714 6356 10716
rect 6324 10686 6326 10714
rect 6326 10686 6354 10714
rect 6354 10686 6356 10714
rect 6324 10684 6356 10686
rect 6324 10634 6356 10636
rect 6324 10606 6326 10634
rect 6326 10606 6354 10634
rect 6354 10606 6356 10634
rect 6324 10604 6356 10606
rect 6324 10554 6356 10556
rect 6324 10526 6326 10554
rect 6326 10526 6354 10554
rect 6354 10526 6356 10554
rect 6324 10524 6356 10526
rect 6324 10474 6356 10476
rect 6324 10446 6326 10474
rect 6326 10446 6354 10474
rect 6354 10446 6356 10474
rect 6324 10444 6356 10446
rect 6324 10394 6356 10396
rect 6324 10366 6326 10394
rect 6326 10366 6354 10394
rect 6354 10366 6356 10394
rect 6324 10364 6356 10366
rect 6324 10314 6356 10316
rect 6324 10286 6326 10314
rect 6326 10286 6354 10314
rect 6354 10286 6356 10314
rect 6324 10284 6356 10286
rect 6324 10234 6356 10236
rect 6324 10206 6326 10234
rect 6326 10206 6354 10234
rect 6354 10206 6356 10234
rect 6324 10204 6356 10206
rect 6324 10154 6356 10156
rect 6324 10126 6326 10154
rect 6326 10126 6354 10154
rect 6354 10126 6356 10154
rect 6324 10124 6356 10126
rect 6324 10074 6356 10076
rect 6324 10046 6326 10074
rect 6326 10046 6354 10074
rect 6354 10046 6356 10074
rect 6324 10044 6356 10046
rect 6324 9994 6356 9996
rect 6324 9966 6326 9994
rect 6326 9966 6354 9994
rect 6354 9966 6356 9994
rect 6324 9964 6356 9966
rect 6324 9914 6356 9916
rect 6324 9886 6326 9914
rect 6326 9886 6354 9914
rect 6354 9886 6356 9914
rect 6324 9884 6356 9886
rect 6324 9834 6356 9836
rect 6324 9806 6326 9834
rect 6326 9806 6354 9834
rect 6354 9806 6356 9834
rect 6324 9804 6356 9806
rect 6324 9754 6356 9756
rect 6324 9726 6326 9754
rect 6326 9726 6354 9754
rect 6354 9726 6356 9754
rect 6324 9724 6356 9726
rect 6324 9354 6356 9356
rect 6324 9326 6326 9354
rect 6326 9326 6354 9354
rect 6354 9326 6356 9354
rect 6324 9324 6356 9326
rect 6324 9274 6356 9276
rect 6324 9246 6326 9274
rect 6326 9246 6354 9274
rect 6354 9246 6356 9274
rect 6324 9244 6356 9246
rect 6324 9194 6356 9196
rect 6324 9166 6326 9194
rect 6326 9166 6354 9194
rect 6354 9166 6356 9194
rect 6324 9164 6356 9166
rect 6324 8874 6356 8876
rect 6324 8846 6326 8874
rect 6326 8846 6354 8874
rect 6354 8846 6356 8874
rect 6324 8844 6356 8846
rect 6324 8794 6356 8796
rect 6324 8766 6326 8794
rect 6326 8766 6354 8794
rect 6354 8766 6356 8794
rect 6324 8764 6356 8766
rect 6324 8714 6356 8716
rect 6324 8686 6326 8714
rect 6326 8686 6354 8714
rect 6354 8686 6356 8714
rect 6324 8684 6356 8686
rect 6324 8634 6356 8636
rect 6324 8606 6326 8634
rect 6326 8606 6354 8634
rect 6354 8606 6356 8634
rect 6324 8604 6356 8606
rect 6324 8554 6356 8556
rect 6324 8526 6326 8554
rect 6326 8526 6354 8554
rect 6354 8526 6356 8554
rect 6324 8524 6356 8526
rect 6324 7634 6356 7636
rect 6324 7606 6326 7634
rect 6326 7606 6354 7634
rect 6354 7606 6356 7634
rect 6324 7604 6356 7606
rect 6324 7554 6356 7556
rect 6324 7526 6326 7554
rect 6326 7526 6354 7554
rect 6354 7526 6356 7554
rect 6324 7524 6356 7526
rect 6324 7474 6356 7476
rect 6324 7446 6326 7474
rect 6326 7446 6354 7474
rect 6354 7446 6356 7474
rect 6324 7444 6356 7446
rect 6324 7394 6356 7396
rect 6324 7366 6326 7394
rect 6326 7366 6354 7394
rect 6354 7366 6356 7394
rect 6324 7364 6356 7366
rect 6324 7314 6356 7316
rect 6324 7286 6326 7314
rect 6326 7286 6354 7314
rect 6354 7286 6356 7314
rect 6324 7284 6356 7286
rect 6324 7234 6356 7236
rect 6324 7206 6326 7234
rect 6326 7206 6354 7234
rect 6354 7206 6356 7234
rect 6324 7204 6356 7206
rect 6324 7154 6356 7156
rect 6324 7126 6326 7154
rect 6326 7126 6354 7154
rect 6354 7126 6356 7154
rect 6324 7124 6356 7126
rect 6324 7074 6356 7076
rect 6324 7046 6326 7074
rect 6326 7046 6354 7074
rect 6354 7046 6356 7074
rect 6324 7044 6356 7046
rect 6324 6754 6356 6756
rect 6324 6726 6326 6754
rect 6326 6726 6354 6754
rect 6354 6726 6356 6754
rect 6324 6724 6356 6726
rect 6324 6674 6356 6676
rect 6324 6646 6326 6674
rect 6326 6646 6354 6674
rect 6354 6646 6356 6674
rect 6324 6644 6356 6646
rect 6324 6594 6356 6596
rect 6324 6566 6326 6594
rect 6326 6566 6354 6594
rect 6354 6566 6356 6594
rect 6324 6564 6356 6566
rect 6324 6514 6356 6516
rect 6324 6486 6326 6514
rect 6326 6486 6354 6514
rect 6354 6486 6356 6514
rect 6324 6484 6356 6486
rect 6324 6434 6356 6436
rect 6324 6406 6326 6434
rect 6326 6406 6354 6434
rect 6354 6406 6356 6434
rect 6324 6404 6356 6406
rect 6324 6354 6356 6356
rect 6324 6326 6326 6354
rect 6326 6326 6354 6354
rect 6354 6326 6356 6354
rect 6324 6324 6356 6326
rect 6324 5794 6356 5796
rect 6324 5766 6326 5794
rect 6326 5766 6354 5794
rect 6354 5766 6356 5794
rect 6324 5764 6356 5766
rect 6324 5714 6356 5716
rect 6324 5686 6326 5714
rect 6326 5686 6354 5714
rect 6354 5686 6356 5714
rect 6324 5684 6356 5686
rect 6324 5634 6356 5636
rect 6324 5606 6326 5634
rect 6326 5606 6354 5634
rect 6354 5606 6356 5634
rect 6324 5604 6356 5606
rect 6324 5554 6356 5556
rect 6324 5526 6326 5554
rect 6326 5526 6354 5554
rect 6354 5526 6356 5554
rect 6324 5524 6356 5526
rect 6324 5474 6356 5476
rect 6324 5446 6326 5474
rect 6326 5446 6354 5474
rect 6354 5446 6356 5474
rect 6324 5444 6356 5446
rect 6324 5394 6356 5396
rect 6324 5366 6326 5394
rect 6326 5366 6354 5394
rect 6354 5366 6356 5394
rect 6324 5364 6356 5366
rect 6324 5314 6356 5316
rect 6324 5286 6326 5314
rect 6326 5286 6354 5314
rect 6354 5286 6356 5314
rect 6324 5284 6356 5286
rect 6324 5234 6356 5236
rect 6324 5206 6326 5234
rect 6326 5206 6354 5234
rect 6354 5206 6356 5234
rect 6324 5204 6356 5206
rect 6324 5154 6356 5156
rect 6324 5126 6326 5154
rect 6326 5126 6354 5154
rect 6354 5126 6356 5154
rect 6324 5124 6356 5126
rect 6324 5074 6356 5076
rect 6324 5046 6326 5074
rect 6326 5046 6354 5074
rect 6354 5046 6356 5074
rect 6324 5044 6356 5046
rect 6324 4994 6356 4996
rect 6324 4966 6326 4994
rect 6326 4966 6354 4994
rect 6354 4966 6356 4994
rect 6324 4964 6356 4966
rect 6324 4434 6356 4436
rect 6324 4406 6326 4434
rect 6326 4406 6354 4434
rect 6354 4406 6356 4434
rect 6324 4404 6356 4406
rect 6324 4354 6356 4356
rect 6324 4326 6326 4354
rect 6326 4326 6354 4354
rect 6354 4326 6356 4354
rect 6324 4324 6356 4326
rect 6324 4274 6356 4276
rect 6324 4246 6326 4274
rect 6326 4246 6354 4274
rect 6354 4246 6356 4274
rect 6324 4244 6356 4246
rect 6324 4194 6356 4196
rect 6324 4166 6326 4194
rect 6326 4166 6354 4194
rect 6354 4166 6356 4194
rect 6324 4164 6356 4166
rect 6324 4114 6356 4116
rect 6324 4086 6326 4114
rect 6326 4086 6354 4114
rect 6354 4086 6356 4114
rect 6324 4084 6356 4086
rect 6324 4034 6356 4036
rect 6324 4006 6326 4034
rect 6326 4006 6354 4034
rect 6354 4006 6356 4034
rect 6324 4004 6356 4006
rect 6324 3954 6356 3956
rect 6324 3926 6326 3954
rect 6326 3926 6354 3954
rect 6354 3926 6356 3954
rect 6324 3924 6356 3926
rect 6324 3154 6356 3156
rect 6324 3126 6326 3154
rect 6326 3126 6354 3154
rect 6354 3126 6356 3154
rect 6324 3124 6356 3126
rect 6324 3074 6356 3076
rect 6324 3046 6326 3074
rect 6326 3046 6354 3074
rect 6354 3046 6356 3074
rect 6324 3044 6356 3046
rect 6324 2994 6356 2996
rect 6324 2966 6326 2994
rect 6326 2966 6354 2994
rect 6354 2966 6356 2994
rect 6324 2964 6356 2966
rect 6324 2914 6356 2916
rect 6324 2886 6326 2914
rect 6326 2886 6354 2914
rect 6354 2886 6356 2914
rect 6324 2884 6356 2886
rect 6324 2834 6356 2836
rect 6324 2806 6326 2834
rect 6326 2806 6354 2834
rect 6354 2806 6356 2834
rect 6324 2804 6356 2806
rect 6324 2754 6356 2756
rect 6324 2726 6326 2754
rect 6326 2726 6354 2754
rect 6354 2726 6356 2754
rect 6324 2724 6356 2726
rect 6324 2674 6356 2676
rect 6324 2646 6326 2674
rect 6326 2646 6354 2674
rect 6354 2646 6356 2674
rect 6324 2644 6356 2646
rect 6324 2594 6356 2596
rect 6324 2566 6326 2594
rect 6326 2566 6354 2594
rect 6354 2566 6356 2594
rect 6324 2564 6356 2566
rect 6324 2514 6356 2516
rect 6324 2486 6326 2514
rect 6326 2486 6354 2514
rect 6354 2486 6356 2514
rect 6324 2484 6356 2486
rect 6324 2434 6356 2436
rect 6324 2406 6326 2434
rect 6326 2406 6354 2434
rect 6354 2406 6356 2434
rect 6324 2404 6356 2406
rect 6324 2354 6356 2356
rect 6324 2326 6326 2354
rect 6326 2326 6354 2354
rect 6354 2326 6356 2354
rect 6324 2324 6356 2326
rect 6324 2274 6356 2276
rect 6324 2246 6326 2274
rect 6326 2246 6354 2274
rect 6354 2246 6356 2274
rect 6324 2244 6356 2246
rect 6324 2194 6356 2196
rect 6324 2166 6326 2194
rect 6326 2166 6354 2194
rect 6354 2166 6356 2194
rect 6324 2164 6356 2166
rect 6324 2114 6356 2116
rect 6324 2086 6326 2114
rect 6326 2086 6354 2114
rect 6354 2086 6356 2114
rect 6324 2084 6356 2086
rect 6324 2034 6356 2036
rect 6324 2006 6326 2034
rect 6326 2006 6354 2034
rect 6354 2006 6356 2034
rect 6324 2004 6356 2006
rect 6324 1634 6356 1636
rect 6324 1606 6326 1634
rect 6326 1606 6354 1634
rect 6354 1606 6356 1634
rect 6324 1604 6356 1606
rect 6324 1554 6356 1556
rect 6324 1526 6326 1554
rect 6326 1526 6354 1554
rect 6354 1526 6356 1554
rect 6324 1524 6356 1526
rect 6324 1474 6356 1476
rect 6324 1446 6326 1474
rect 6326 1446 6354 1474
rect 6354 1446 6356 1474
rect 6324 1444 6356 1446
rect 6324 1394 6356 1396
rect 6324 1366 6326 1394
rect 6326 1366 6354 1394
rect 6354 1366 6356 1394
rect 6324 1364 6356 1366
rect 6324 1314 6356 1316
rect 6324 1286 6326 1314
rect 6326 1286 6354 1314
rect 6354 1286 6356 1314
rect 6324 1284 6356 1286
rect 6324 1234 6356 1236
rect 6324 1206 6326 1234
rect 6326 1206 6354 1234
rect 6354 1206 6356 1234
rect 6324 1204 6356 1206
rect 6324 1154 6356 1156
rect 6324 1126 6326 1154
rect 6326 1126 6354 1154
rect 6354 1126 6356 1154
rect 6324 1124 6356 1126
rect 6324 1074 6356 1076
rect 6324 1046 6326 1074
rect 6326 1046 6354 1074
rect 6354 1046 6356 1074
rect 6324 1044 6356 1046
rect 6324 754 6356 756
rect 6324 726 6326 754
rect 6326 726 6354 754
rect 6354 726 6356 754
rect 6324 724 6356 726
rect 6324 674 6356 676
rect 6324 646 6326 674
rect 6326 646 6354 674
rect 6354 646 6356 674
rect 6324 644 6356 646
rect 6324 594 6356 596
rect 6324 566 6326 594
rect 6326 566 6354 594
rect 6354 566 6356 594
rect 6324 564 6356 566
rect 6324 194 6356 196
rect 6324 166 6326 194
rect 6326 166 6354 194
rect 6354 166 6356 194
rect 6324 164 6356 166
rect 6324 114 6356 116
rect 6324 86 6326 114
rect 6326 86 6354 114
rect 6354 86 6356 114
rect 6324 84 6356 86
rect 6324 34 6356 36
rect 6324 6 6326 34
rect 6326 6 6354 34
rect 6354 6 6356 34
rect 6324 4 6356 6
<< mimcap >>
rect 520 16596 1520 16640
rect 520 15684 564 16596
rect 1476 15684 1520 16596
rect 520 15640 1520 15684
rect 1640 16596 2640 16640
rect 1640 15684 1684 16596
rect 2596 15684 2640 16596
rect 1640 15640 2640 15684
rect 2760 16596 3760 16640
rect 2760 15684 2804 16596
rect 3716 15684 3760 16596
rect 2760 15640 3760 15684
rect 3880 16596 4880 16640
rect 3880 15684 3924 16596
rect 4836 15684 4880 16596
rect 3880 15640 4880 15684
rect 5720 16596 6720 16640
rect 5720 15684 5764 16596
rect 6676 15684 6720 16596
rect 5720 15640 6720 15684
rect 6840 16596 7840 16640
rect 6840 15684 6884 16596
rect 7796 15684 7840 16596
rect 6840 15640 7840 15684
rect 7960 16596 8960 16640
rect 7960 15684 8004 16596
rect 8916 15684 8960 16596
rect 7960 15640 8960 15684
rect 9080 16596 10080 16640
rect 9080 15684 9124 16596
rect 10036 15684 10080 16596
rect 9080 15640 10080 15684
rect 520 15156 1520 15200
rect 520 14244 564 15156
rect 1476 14244 1520 15156
rect 520 14200 1520 14244
rect 1640 15156 2640 15200
rect 1640 14244 1684 15156
rect 2596 14244 2640 15156
rect 1640 14200 2640 14244
rect 2760 15156 3760 15200
rect 2760 14244 2804 15156
rect 3716 14244 3760 15156
rect 2760 14200 3760 14244
rect 3880 15156 4880 15200
rect 3880 14244 3924 15156
rect 4836 14244 4880 15156
rect 3880 14200 4880 14244
rect 5720 15156 6720 15200
rect 5720 14244 5764 15156
rect 6676 14244 6720 15156
rect 5720 14200 6720 14244
rect 6840 15156 7840 15200
rect 6840 14244 6884 15156
rect 7796 14244 7840 15156
rect 6840 14200 7840 14244
rect 7960 15156 8960 15200
rect 7960 14244 8004 15156
rect 8916 14244 8960 15156
rect 7960 14200 8960 14244
rect 9080 15156 10080 15200
rect 9080 14244 9124 15156
rect 10036 14244 10080 15156
rect 9080 14200 10080 14244
<< mimcapcontact >>
rect 564 15684 1476 16596
rect 1684 15684 2596 16596
rect 2804 15684 3716 16596
rect 3924 15684 4836 16596
rect 5764 15684 6676 16596
rect 6884 15684 7796 16596
rect 8004 15684 8916 16596
rect 9124 15684 10036 16596
rect 564 14244 1476 15156
rect 1684 14244 2596 15156
rect 2804 14244 3716 15156
rect 3924 14244 4836 15156
rect 5764 14244 6676 15156
rect 6884 14244 7796 15156
rect 8004 14244 8916 15156
rect 9124 14244 10036 15156
<< metal4 >>
rect 0 16916 10600 16920
rect 0 16884 4 16916
rect 36 16884 324 16916
rect 356 16884 10244 16916
rect 10276 16884 10564 16916
rect 10596 16884 10600 16916
rect 0 16880 10600 16884
rect 0 16836 10600 16840
rect 0 16804 84 16836
rect 116 16804 244 16836
rect 276 16804 404 16836
rect 436 16804 10164 16836
rect 10196 16804 10324 16836
rect 10356 16804 10484 16836
rect 10516 16804 10600 16836
rect 0 16800 10600 16804
rect 80 16756 10520 16760
rect 80 16724 164 16756
rect 196 16724 484 16756
rect 516 16724 1524 16756
rect 1556 16724 1604 16756
rect 1636 16724 2644 16756
rect 2676 16724 2724 16756
rect 2756 16724 3764 16756
rect 3796 16724 3844 16756
rect 3876 16724 4884 16756
rect 4916 16724 5684 16756
rect 5716 16724 6724 16756
rect 6756 16724 6804 16756
rect 6836 16724 7844 16756
rect 7876 16724 7924 16756
rect 7956 16724 8964 16756
rect 8996 16724 9044 16756
rect 9076 16724 10084 16756
rect 10116 16724 10404 16756
rect 10436 16724 10520 16756
rect 80 16720 10520 16724
rect 480 16596 1560 16680
rect 480 15684 564 16596
rect 1476 15684 1560 16596
rect 480 15600 1560 15684
rect 480 15560 520 15600
rect 1520 15560 1560 15600
rect 1600 16596 2680 16680
rect 1600 15684 1684 16596
rect 2596 15684 2680 16596
rect 1600 15600 2680 15684
rect 1600 15560 1640 15600
rect 2640 15560 2680 15600
rect 2720 16596 3800 16680
rect 2720 15684 2804 16596
rect 3716 15684 3800 16596
rect 2720 15600 3800 15684
rect 2720 15560 2760 15600
rect 3760 15560 3800 15600
rect 3840 16596 4920 16680
rect 3840 15684 3924 16596
rect 4836 15684 4920 16596
rect 3840 15600 4920 15684
rect 3840 15560 3880 15600
rect 4880 15560 4920 15600
rect 5680 16596 6760 16680
rect 5680 15684 5764 16596
rect 6676 15684 6760 16596
rect 5680 15600 6760 15684
rect 5680 15560 5720 15600
rect 6720 15560 6760 15600
rect 6800 16596 7880 16680
rect 6800 15684 6884 16596
rect 7796 15684 7880 16596
rect 6800 15600 7880 15684
rect 6800 15560 6840 15600
rect 7840 15560 7880 15600
rect 7920 16596 9000 16680
rect 7920 15684 8004 16596
rect 8916 15684 9000 16596
rect 7920 15600 9000 15684
rect 7920 15560 7960 15600
rect 8960 15560 9000 15600
rect 9040 16596 10120 16680
rect 9040 15684 9124 16596
rect 10036 15684 10120 16596
rect 9040 15600 10120 15684
rect 9040 15560 9080 15600
rect 10080 15560 10120 15600
rect 0 15556 10600 15560
rect 0 15524 84 15556
rect 116 15524 244 15556
rect 276 15524 404 15556
rect 436 15524 10164 15556
rect 10196 15524 10324 15556
rect 10356 15524 10484 15556
rect 10516 15524 10600 15556
rect 0 15520 10600 15524
rect 0 15476 10600 15480
rect 0 15444 4 15476
rect 36 15444 324 15476
rect 356 15444 10244 15476
rect 10276 15444 10564 15476
rect 10596 15444 10600 15476
rect 0 15440 10600 15444
rect 400 15396 10200 15400
rect 400 15364 404 15396
rect 436 15364 4964 15396
rect 4996 15364 5124 15396
rect 5156 15364 5284 15396
rect 5316 15364 5444 15396
rect 5476 15364 5604 15396
rect 5636 15364 10164 15396
rect 10196 15364 10200 15396
rect 400 15360 10200 15364
rect 480 15316 5240 15320
rect 480 15284 484 15316
rect 516 15284 1524 15316
rect 1556 15284 1604 15316
rect 1636 15284 2644 15316
rect 2676 15284 2724 15316
rect 2756 15284 3764 15316
rect 3796 15284 3844 15316
rect 3876 15284 4884 15316
rect 4916 15284 5204 15316
rect 5236 15284 5240 15316
rect 480 15280 5240 15284
rect 5360 15316 10160 15320
rect 5360 15284 5364 15316
rect 5396 15284 5684 15316
rect 5716 15284 6724 15316
rect 6756 15284 6804 15316
rect 6836 15284 7844 15316
rect 7876 15284 7924 15316
rect 7956 15284 8964 15316
rect 8996 15284 9044 15316
rect 9076 15284 10084 15316
rect 10116 15284 10160 15316
rect 5360 15280 10160 15284
rect 480 15156 1560 15240
rect 480 14244 564 15156
rect 1476 14244 1560 15156
rect 480 14160 1560 14244
rect 480 14120 520 14160
rect 1520 14120 1560 14160
rect 1600 15156 2680 15240
rect 1600 14244 1684 15156
rect 2596 14244 2680 15156
rect 1600 14160 2680 14244
rect 1600 14120 1640 14160
rect 2640 14120 2680 14160
rect 2720 15156 3800 15240
rect 2720 14244 2804 15156
rect 3716 14244 3800 15156
rect 2720 14160 3800 14244
rect 2720 14120 2760 14160
rect 3760 14120 3800 14160
rect 3840 15156 4920 15240
rect 3840 14244 3924 15156
rect 4836 14244 4920 15156
rect 3840 14160 4920 14244
rect 3840 14120 3880 14160
rect 4880 14120 4920 14160
rect 5680 15156 6760 15240
rect 5680 14244 5764 15156
rect 6676 14244 6760 15156
rect 5680 14160 6760 14244
rect 5680 14120 5720 14160
rect 6720 14120 6760 14160
rect 6800 15156 7880 15240
rect 6800 14244 6884 15156
rect 7796 14244 7880 15156
rect 6800 14160 7880 14244
rect 6800 14120 6840 14160
rect 7840 14120 7880 14160
rect 7920 15156 9000 15240
rect 7920 14244 8004 15156
rect 8916 14244 9000 15156
rect 7920 14160 9000 14244
rect 7920 14120 7960 14160
rect 8960 14120 9000 14160
rect 9040 15156 10120 15240
rect 9040 14244 9124 15156
rect 10036 14244 10120 15156
rect 9040 14160 10120 14244
rect 9040 14120 9080 14160
rect 10080 14120 10120 14160
rect 400 14116 10200 14120
rect 400 14084 404 14116
rect 436 14084 4964 14116
rect 4996 14084 5124 14116
rect 5156 14084 5284 14116
rect 5316 14084 5444 14116
rect 5476 14084 5604 14116
rect 5636 14084 10164 14116
rect 10196 14084 10200 14116
rect 400 14080 10200 14084
rect 0 14036 10600 14040
rect 0 14004 4 14036
rect 36 14004 324 14036
rect 356 14004 5044 14036
rect 5076 14004 5524 14036
rect 5556 14004 10244 14036
rect 10276 14004 10564 14036
rect 10596 14004 10600 14036
rect 0 14000 10600 14004
rect 0 13956 10600 13960
rect 0 13924 84 13956
rect 116 13924 244 13956
rect 276 13924 4484 13956
rect 4516 13924 4644 13956
rect 4676 13924 10324 13956
rect 10356 13924 10484 13956
rect 10516 13924 10600 13956
rect 0 13920 10600 13924
rect 0 13876 10600 13880
rect 0 13844 164 13876
rect 196 13844 4564 13876
rect 4596 13844 10404 13876
rect 10436 13844 10600 13876
rect 0 13840 10600 13844
rect 0 13796 10600 13800
rect 0 13764 84 13796
rect 116 13764 244 13796
rect 276 13764 4484 13796
rect 4516 13764 4644 13796
rect 4676 13764 10324 13796
rect 10356 13764 10484 13796
rect 10516 13764 10600 13796
rect 0 13760 10600 13764
rect 0 13716 10600 13720
rect 0 13684 4 13716
rect 36 13684 324 13716
rect 356 13684 5044 13716
rect 5076 13684 5524 13716
rect 5556 13684 10244 13716
rect 10276 13684 10564 13716
rect 10596 13684 10600 13716
rect 0 13680 10600 13684
rect 0 13636 10600 13640
rect 0 13604 4244 13636
rect 4276 13604 4404 13636
rect 4436 13604 10600 13636
rect 0 13599 10600 13604
rect 0 13481 1561 13599
rect 1679 13481 2521 13599
rect 2639 13596 7961 13599
rect 2639 13564 4244 13596
rect 4276 13564 4404 13596
rect 4436 13564 7961 13596
rect 2639 13556 7961 13564
rect 2639 13524 4244 13556
rect 4276 13524 4404 13556
rect 4436 13524 7961 13556
rect 2639 13516 7961 13524
rect 2639 13484 4244 13516
rect 4276 13484 4404 13516
rect 4436 13484 7961 13516
rect 2639 13481 7961 13484
rect 8079 13481 8921 13599
rect 9039 13481 10600 13599
rect 0 13476 10600 13481
rect 0 13444 4244 13476
rect 4276 13444 4404 13476
rect 4436 13444 10600 13476
rect 0 13440 10600 13444
rect 0 13396 10600 13400
rect 0 13364 4724 13396
rect 4756 13364 4884 13396
rect 4916 13364 5044 13396
rect 5076 13364 5524 13396
rect 5556 13364 5684 13396
rect 5716 13364 5844 13396
rect 5876 13364 6164 13396
rect 6196 13364 6324 13396
rect 6356 13364 10600 13396
rect 0 13359 10600 13364
rect 0 13241 1081 13359
rect 1199 13241 2041 13359
rect 2159 13241 3001 13359
rect 3119 13356 7481 13359
rect 3119 13324 4724 13356
rect 4756 13324 4884 13356
rect 4916 13324 5044 13356
rect 5076 13324 5524 13356
rect 5556 13324 5684 13356
rect 5716 13324 5844 13356
rect 5876 13324 6164 13356
rect 6196 13324 6324 13356
rect 6356 13324 7481 13356
rect 3119 13316 7481 13324
rect 3119 13284 4724 13316
rect 4756 13284 4884 13316
rect 4916 13284 5044 13316
rect 5076 13284 5524 13316
rect 5556 13284 5684 13316
rect 5716 13284 5844 13316
rect 5876 13284 6164 13316
rect 6196 13284 6324 13316
rect 6356 13284 7481 13316
rect 3119 13276 7481 13284
rect 3119 13244 4724 13276
rect 4756 13244 4884 13276
rect 4916 13244 5044 13276
rect 5076 13244 5524 13276
rect 5556 13244 5684 13276
rect 5716 13244 5844 13276
rect 5876 13244 6164 13276
rect 6196 13244 6324 13276
rect 6356 13244 7481 13276
rect 3119 13241 7481 13244
rect 7599 13241 8441 13359
rect 8559 13241 9401 13359
rect 9519 13241 10600 13359
rect 0 13236 10600 13241
rect 0 13204 4724 13236
rect 4756 13204 4884 13236
rect 4916 13204 5044 13236
rect 5076 13204 5524 13236
rect 5556 13204 5684 13236
rect 5716 13204 5844 13236
rect 5876 13204 6164 13236
rect 6196 13204 6324 13236
rect 6356 13204 10600 13236
rect 0 13200 10600 13204
rect 0 13156 10600 13160
rect 0 13124 4484 13156
rect 4516 13124 4644 13156
rect 4676 13124 10600 13156
rect 0 13119 10600 13124
rect 0 13001 601 13119
rect 719 13001 3481 13119
rect 3599 13116 7001 13119
rect 3599 13084 4484 13116
rect 4516 13084 4644 13116
rect 4676 13084 7001 13116
rect 3599 13076 7001 13084
rect 3599 13044 4484 13076
rect 4516 13044 4644 13076
rect 4676 13044 7001 13076
rect 3599 13036 7001 13044
rect 3599 13004 4484 13036
rect 4516 13004 4644 13036
rect 4676 13004 7001 13036
rect 3599 13001 7001 13004
rect 7119 13001 9881 13119
rect 9999 13001 10600 13119
rect 0 12996 10600 13001
rect 0 12964 4484 12996
rect 4516 12964 4644 12996
rect 4676 12964 10600 12996
rect 0 12960 10600 12964
rect 0 12916 10600 12920
rect 0 12884 5924 12916
rect 5956 12884 6084 12916
rect 6116 12884 10600 12916
rect 0 12879 10600 12884
rect 0 12761 121 12879
rect 239 12761 3961 12879
rect 4079 12876 6521 12879
rect 4079 12844 5924 12876
rect 5956 12844 6084 12876
rect 6116 12844 6521 12876
rect 4079 12836 6521 12844
rect 4079 12804 5924 12836
rect 5956 12804 6084 12836
rect 6116 12804 6521 12836
rect 4079 12796 6521 12804
rect 4079 12764 5924 12796
rect 5956 12764 6084 12796
rect 6116 12764 6521 12796
rect 4079 12761 6521 12764
rect 6639 12761 10361 12879
rect 10479 12761 10600 12879
rect 0 12756 10600 12761
rect 0 12724 5924 12756
rect 5956 12724 6084 12756
rect 6116 12724 10600 12756
rect 0 12720 10600 12724
rect 4240 12636 4440 12640
rect 4240 12604 4244 12636
rect 4276 12604 4404 12636
rect 4436 12604 4440 12636
rect 4240 12600 4440 12604
rect 4480 12636 4680 12640
rect 4480 12604 4484 12636
rect 4516 12604 4644 12636
rect 4676 12604 4680 12636
rect 4480 12600 4680 12604
rect 4720 12636 5080 12640
rect 4720 12604 4724 12636
rect 4756 12604 4884 12636
rect 4916 12604 5044 12636
rect 5076 12604 5080 12636
rect 4720 12600 5080 12604
rect 5120 12636 5480 12640
rect 5120 12604 5124 12636
rect 5156 12604 5284 12636
rect 5316 12604 5444 12636
rect 5476 12604 5480 12636
rect 5120 12600 5480 12604
rect 5520 12636 5880 12640
rect 5520 12604 5524 12636
rect 5556 12604 5684 12636
rect 5716 12604 5844 12636
rect 5876 12604 5880 12636
rect 5520 12600 5880 12604
rect 5920 12636 6120 12640
rect 5920 12604 5924 12636
rect 5956 12604 6084 12636
rect 6116 12604 6120 12636
rect 5920 12600 6120 12604
rect 6160 12636 6360 12640
rect 6160 12604 6164 12636
rect 6196 12604 6324 12636
rect 6356 12604 6360 12636
rect 6160 12600 6360 12604
rect 4240 12556 4440 12560
rect 4240 12524 4244 12556
rect 4276 12524 4404 12556
rect 4436 12524 4440 12556
rect 4240 12520 4440 12524
rect 4480 12556 4680 12560
rect 4480 12524 4484 12556
rect 4516 12524 4644 12556
rect 4676 12524 4680 12556
rect 4480 12520 4680 12524
rect 4720 12556 5080 12560
rect 4720 12524 4724 12556
rect 4756 12524 4884 12556
rect 4916 12524 5044 12556
rect 5076 12524 5080 12556
rect 4720 12520 5080 12524
rect 5120 12556 5480 12560
rect 5120 12524 5124 12556
rect 5156 12524 5284 12556
rect 5316 12524 5444 12556
rect 5476 12524 5480 12556
rect 5120 12520 5480 12524
rect 5520 12556 5880 12560
rect 5520 12524 5524 12556
rect 5556 12524 5684 12556
rect 5716 12524 5844 12556
rect 5876 12524 5880 12556
rect 5520 12520 5880 12524
rect 5920 12556 6120 12560
rect 5920 12524 5924 12556
rect 5956 12524 6084 12556
rect 6116 12524 6120 12556
rect 5920 12520 6120 12524
rect 6160 12556 6360 12560
rect 6160 12524 6164 12556
rect 6196 12524 6324 12556
rect 6356 12524 6360 12556
rect 6160 12520 6360 12524
rect 4240 12476 4440 12480
rect 4240 12444 4244 12476
rect 4276 12444 4404 12476
rect 4436 12444 4440 12476
rect 4240 12440 4440 12444
rect 4480 12476 4680 12480
rect 4480 12444 4484 12476
rect 4516 12444 4644 12476
rect 4676 12444 4680 12476
rect 4480 12440 4680 12444
rect 4720 12476 5080 12480
rect 4720 12444 4724 12476
rect 4756 12444 4884 12476
rect 4916 12444 5044 12476
rect 5076 12444 5080 12476
rect 4720 12440 5080 12444
rect 5120 12476 5480 12480
rect 5120 12444 5124 12476
rect 5156 12444 5284 12476
rect 5316 12444 5444 12476
rect 5476 12444 5480 12476
rect 5120 12440 5480 12444
rect 5520 12476 5880 12480
rect 5520 12444 5524 12476
rect 5556 12444 5684 12476
rect 5716 12444 5844 12476
rect 5876 12444 5880 12476
rect 5520 12440 5880 12444
rect 5920 12476 6120 12480
rect 5920 12444 5924 12476
rect 5956 12444 6084 12476
rect 6116 12444 6120 12476
rect 5920 12440 6120 12444
rect 6160 12476 6360 12480
rect 6160 12444 6164 12476
rect 6196 12444 6324 12476
rect 6356 12444 6360 12476
rect 6160 12440 6360 12444
rect 4240 12396 4440 12400
rect 4240 12364 4244 12396
rect 4276 12364 4404 12396
rect 4436 12364 4440 12396
rect 4240 12360 4440 12364
rect 4480 12396 4680 12400
rect 4480 12364 4484 12396
rect 4516 12364 4644 12396
rect 4676 12364 4680 12396
rect 4480 12360 4680 12364
rect 4720 12396 5080 12400
rect 4720 12364 4724 12396
rect 4756 12364 4884 12396
rect 4916 12364 5044 12396
rect 5076 12364 5080 12396
rect 4720 12360 5080 12364
rect 5120 12396 5480 12400
rect 5120 12364 5124 12396
rect 5156 12364 5284 12396
rect 5316 12364 5444 12396
rect 5476 12364 5480 12396
rect 5120 12360 5480 12364
rect 5520 12396 5880 12400
rect 5520 12364 5524 12396
rect 5556 12364 5684 12396
rect 5716 12364 5844 12396
rect 5876 12364 5880 12396
rect 5520 12360 5880 12364
rect 5920 12396 6120 12400
rect 5920 12364 5924 12396
rect 5956 12364 6084 12396
rect 6116 12364 6120 12396
rect 5920 12360 6120 12364
rect 6160 12396 6360 12400
rect 6160 12364 6164 12396
rect 6196 12364 6324 12396
rect 6356 12364 6360 12396
rect 6160 12360 6360 12364
rect 4240 12316 4440 12320
rect 4240 12284 4244 12316
rect 4276 12284 4404 12316
rect 4436 12284 4440 12316
rect 4240 12280 4440 12284
rect 4480 12316 4680 12320
rect 4480 12284 4484 12316
rect 4516 12284 4644 12316
rect 4676 12284 4680 12316
rect 4480 12280 4680 12284
rect 4720 12316 5080 12320
rect 4720 12284 4724 12316
rect 4756 12284 4884 12316
rect 4916 12284 5044 12316
rect 5076 12284 5080 12316
rect 4720 12280 5080 12284
rect 5120 12316 5480 12320
rect 5120 12284 5124 12316
rect 5156 12284 5284 12316
rect 5316 12284 5444 12316
rect 5476 12284 5480 12316
rect 5120 12280 5480 12284
rect 5520 12316 5880 12320
rect 5520 12284 5524 12316
rect 5556 12284 5684 12316
rect 5716 12284 5844 12316
rect 5876 12284 5880 12316
rect 5520 12280 5880 12284
rect 5920 12316 6120 12320
rect 5920 12284 5924 12316
rect 5956 12284 6084 12316
rect 6116 12284 6120 12316
rect 5920 12280 6120 12284
rect 6160 12316 6360 12320
rect 6160 12284 6164 12316
rect 6196 12284 6324 12316
rect 6356 12284 6360 12316
rect 6160 12280 6360 12284
rect 4240 12236 4440 12240
rect 4240 12204 4244 12236
rect 4276 12204 4404 12236
rect 4436 12204 4440 12236
rect 4240 12200 4440 12204
rect 4480 12236 4680 12240
rect 4480 12204 4484 12236
rect 4516 12204 4644 12236
rect 4676 12204 4680 12236
rect 4480 12200 4680 12204
rect 4720 12236 5080 12240
rect 4720 12204 4724 12236
rect 4756 12204 4884 12236
rect 4916 12204 5044 12236
rect 5076 12204 5080 12236
rect 4720 12200 5080 12204
rect 5120 12236 5480 12240
rect 5120 12204 5124 12236
rect 5156 12204 5284 12236
rect 5316 12204 5444 12236
rect 5476 12204 5480 12236
rect 5120 12200 5480 12204
rect 5520 12236 5880 12240
rect 5520 12204 5524 12236
rect 5556 12204 5684 12236
rect 5716 12204 5844 12236
rect 5876 12204 5880 12236
rect 5520 12200 5880 12204
rect 5920 12236 6120 12240
rect 5920 12204 5924 12236
rect 5956 12204 6084 12236
rect 6116 12204 6120 12236
rect 5920 12200 6120 12204
rect 6160 12236 6360 12240
rect 6160 12204 6164 12236
rect 6196 12204 6324 12236
rect 6356 12204 6360 12236
rect 6160 12200 6360 12204
rect 4240 12156 4440 12160
rect 4240 12124 4244 12156
rect 4276 12124 4404 12156
rect 4436 12124 4440 12156
rect 4240 12120 4440 12124
rect 4480 12156 4680 12160
rect 4480 12124 4484 12156
rect 4516 12124 4644 12156
rect 4676 12124 4680 12156
rect 4480 12120 4680 12124
rect 4720 12156 5080 12160
rect 4720 12124 4724 12156
rect 4756 12124 4884 12156
rect 4916 12124 5044 12156
rect 5076 12124 5080 12156
rect 4720 12120 5080 12124
rect 5120 12156 5480 12160
rect 5120 12124 5124 12156
rect 5156 12124 5284 12156
rect 5316 12124 5444 12156
rect 5476 12124 5480 12156
rect 5120 12120 5480 12124
rect 5520 12156 5880 12160
rect 5520 12124 5524 12156
rect 5556 12124 5684 12156
rect 5716 12124 5844 12156
rect 5876 12124 5880 12156
rect 5520 12120 5880 12124
rect 5920 12156 6120 12160
rect 5920 12124 5924 12156
rect 5956 12124 6084 12156
rect 6116 12124 6120 12156
rect 5920 12120 6120 12124
rect 6160 12156 6360 12160
rect 6160 12124 6164 12156
rect 6196 12124 6324 12156
rect 6356 12124 6360 12156
rect 6160 12120 6360 12124
rect 4240 11836 4440 11840
rect 4240 11804 4244 11836
rect 4276 11804 4404 11836
rect 4436 11804 4440 11836
rect 4240 11800 4440 11804
rect 4480 11836 4680 11840
rect 4480 11804 4484 11836
rect 4516 11804 4644 11836
rect 4676 11804 4680 11836
rect 4480 11800 4680 11804
rect 4720 11836 5080 11840
rect 4720 11804 4724 11836
rect 4756 11804 4884 11836
rect 4916 11804 5044 11836
rect 5076 11804 5080 11836
rect 4720 11800 5080 11804
rect 5120 11836 5480 11840
rect 5120 11804 5124 11836
rect 5156 11804 5284 11836
rect 5316 11804 5444 11836
rect 5476 11804 5480 11836
rect 5120 11800 5480 11804
rect 5520 11836 5880 11840
rect 5520 11804 5524 11836
rect 5556 11804 5684 11836
rect 5716 11804 5844 11836
rect 5876 11804 5880 11836
rect 5520 11800 5880 11804
rect 5920 11836 6120 11840
rect 5920 11804 5924 11836
rect 5956 11804 6084 11836
rect 6116 11804 6120 11836
rect 5920 11800 6120 11804
rect 6160 11836 6360 11840
rect 6160 11804 6164 11836
rect 6196 11804 6324 11836
rect 6356 11804 6360 11836
rect 6160 11800 6360 11804
rect 4240 11756 4440 11760
rect 4240 11724 4244 11756
rect 4276 11724 4404 11756
rect 4436 11724 4440 11756
rect 4240 11720 4440 11724
rect 4480 11756 4680 11760
rect 4480 11724 4484 11756
rect 4516 11724 4644 11756
rect 4676 11724 4680 11756
rect 4480 11720 4680 11724
rect 4720 11756 5080 11760
rect 4720 11724 4724 11756
rect 4756 11724 4884 11756
rect 4916 11724 5044 11756
rect 5076 11724 5080 11756
rect 4720 11720 5080 11724
rect 5120 11756 5480 11760
rect 5120 11724 5124 11756
rect 5156 11724 5284 11756
rect 5316 11724 5444 11756
rect 5476 11724 5480 11756
rect 5120 11720 5480 11724
rect 5520 11756 5880 11760
rect 5520 11724 5524 11756
rect 5556 11724 5684 11756
rect 5716 11724 5844 11756
rect 5876 11724 5880 11756
rect 5520 11720 5880 11724
rect 5920 11756 6120 11760
rect 5920 11724 5924 11756
rect 5956 11724 6084 11756
rect 6116 11724 6120 11756
rect 5920 11720 6120 11724
rect 6160 11756 6360 11760
rect 6160 11724 6164 11756
rect 6196 11724 6324 11756
rect 6356 11724 6360 11756
rect 6160 11720 6360 11724
rect 4240 11676 4440 11680
rect 4240 11644 4244 11676
rect 4276 11644 4404 11676
rect 4436 11644 4440 11676
rect 4240 11640 4440 11644
rect 4480 11676 4680 11680
rect 4480 11644 4484 11676
rect 4516 11644 4644 11676
rect 4676 11644 4680 11676
rect 4480 11640 4680 11644
rect 4720 11676 5080 11680
rect 4720 11644 4724 11676
rect 4756 11644 4884 11676
rect 4916 11644 5044 11676
rect 5076 11644 5080 11676
rect 4720 11640 5080 11644
rect 5120 11676 5480 11680
rect 5120 11644 5124 11676
rect 5156 11644 5284 11676
rect 5316 11644 5444 11676
rect 5476 11644 5480 11676
rect 5120 11640 5480 11644
rect 5520 11676 5880 11680
rect 5520 11644 5524 11676
rect 5556 11644 5684 11676
rect 5716 11644 5844 11676
rect 5876 11644 5880 11676
rect 5520 11640 5880 11644
rect 5920 11676 6120 11680
rect 5920 11644 5924 11676
rect 5956 11644 6084 11676
rect 6116 11644 6120 11676
rect 5920 11640 6120 11644
rect 6160 11676 6360 11680
rect 6160 11644 6164 11676
rect 6196 11644 6324 11676
rect 6356 11644 6360 11676
rect 6160 11640 6360 11644
rect 4240 11596 4440 11600
rect 4240 11564 4244 11596
rect 4276 11564 4404 11596
rect 4436 11564 4440 11596
rect 4240 11560 4440 11564
rect 4480 11596 4680 11600
rect 4480 11564 4484 11596
rect 4516 11564 4644 11596
rect 4676 11564 4680 11596
rect 4480 11560 4680 11564
rect 4720 11596 5080 11600
rect 4720 11564 4724 11596
rect 4756 11564 4884 11596
rect 4916 11564 5044 11596
rect 5076 11564 5080 11596
rect 4720 11560 5080 11564
rect 5120 11596 5480 11600
rect 5120 11564 5124 11596
rect 5156 11564 5284 11596
rect 5316 11564 5444 11596
rect 5476 11564 5480 11596
rect 5120 11560 5480 11564
rect 5520 11596 5880 11600
rect 5520 11564 5524 11596
rect 5556 11564 5684 11596
rect 5716 11564 5844 11596
rect 5876 11564 5880 11596
rect 5520 11560 5880 11564
rect 5920 11596 6120 11600
rect 5920 11564 5924 11596
rect 5956 11564 6084 11596
rect 6116 11564 6120 11596
rect 5920 11560 6120 11564
rect 6160 11596 6360 11600
rect 6160 11564 6164 11596
rect 6196 11564 6324 11596
rect 6356 11564 6360 11596
rect 6160 11560 6360 11564
rect 4240 11516 4440 11520
rect 4240 11484 4244 11516
rect 4276 11484 4404 11516
rect 4436 11484 4440 11516
rect 4240 11480 4440 11484
rect 4480 11516 4680 11520
rect 4480 11484 4484 11516
rect 4516 11484 4644 11516
rect 4676 11484 4680 11516
rect 4480 11480 4680 11484
rect 4720 11516 5080 11520
rect 4720 11484 4724 11516
rect 4756 11484 4884 11516
rect 4916 11484 5044 11516
rect 5076 11484 5080 11516
rect 4720 11480 5080 11484
rect 5120 11516 5480 11520
rect 5120 11484 5124 11516
rect 5156 11484 5284 11516
rect 5316 11484 5444 11516
rect 5476 11484 5480 11516
rect 5120 11480 5480 11484
rect 5520 11516 5880 11520
rect 5520 11484 5524 11516
rect 5556 11484 5684 11516
rect 5716 11484 5844 11516
rect 5876 11484 5880 11516
rect 5520 11480 5880 11484
rect 5920 11516 6120 11520
rect 5920 11484 5924 11516
rect 5956 11484 6084 11516
rect 6116 11484 6120 11516
rect 5920 11480 6120 11484
rect 6160 11516 6360 11520
rect 6160 11484 6164 11516
rect 6196 11484 6324 11516
rect 6356 11484 6360 11516
rect 6160 11480 6360 11484
rect 4240 11436 4440 11440
rect 4240 11404 4244 11436
rect 4276 11404 4404 11436
rect 4436 11404 4440 11436
rect 4240 11400 4440 11404
rect 4480 11436 4680 11440
rect 4480 11404 4484 11436
rect 4516 11404 4644 11436
rect 4676 11404 4680 11436
rect 4480 11400 4680 11404
rect 4720 11436 5080 11440
rect 4720 11404 4724 11436
rect 4756 11404 4884 11436
rect 4916 11404 5044 11436
rect 5076 11404 5080 11436
rect 4720 11400 5080 11404
rect 5120 11436 5480 11440
rect 5120 11404 5124 11436
rect 5156 11404 5284 11436
rect 5316 11404 5444 11436
rect 5476 11404 5480 11436
rect 5120 11400 5480 11404
rect 5520 11436 5880 11440
rect 5520 11404 5524 11436
rect 5556 11404 5684 11436
rect 5716 11404 5844 11436
rect 5876 11404 5880 11436
rect 5520 11400 5880 11404
rect 5920 11436 6120 11440
rect 5920 11404 5924 11436
rect 5956 11404 6084 11436
rect 6116 11404 6120 11436
rect 5920 11400 6120 11404
rect 6160 11436 6360 11440
rect 6160 11404 6164 11436
rect 6196 11404 6324 11436
rect 6356 11404 6360 11436
rect 6160 11400 6360 11404
rect 4240 10876 4440 10880
rect 4240 10844 4244 10876
rect 4276 10844 4404 10876
rect 4436 10844 4440 10876
rect 4240 10840 4440 10844
rect 4480 10876 4680 10880
rect 4480 10844 4484 10876
rect 4516 10844 4644 10876
rect 4676 10844 4680 10876
rect 4480 10840 4680 10844
rect 4720 10876 5080 10880
rect 4720 10844 4724 10876
rect 4756 10844 4884 10876
rect 4916 10844 5044 10876
rect 5076 10844 5080 10876
rect 4720 10840 5080 10844
rect 5120 10876 5480 10880
rect 5120 10844 5124 10876
rect 5156 10844 5284 10876
rect 5316 10844 5444 10876
rect 5476 10844 5480 10876
rect 5120 10840 5480 10844
rect 5520 10876 5880 10880
rect 5520 10844 5524 10876
rect 5556 10844 5684 10876
rect 5716 10844 5844 10876
rect 5876 10844 5880 10876
rect 5520 10840 5880 10844
rect 5920 10876 6120 10880
rect 5920 10844 5924 10876
rect 5956 10844 6084 10876
rect 6116 10844 6120 10876
rect 5920 10840 6120 10844
rect 6160 10876 6360 10880
rect 6160 10844 6164 10876
rect 6196 10844 6324 10876
rect 6356 10844 6360 10876
rect 6160 10840 6360 10844
rect 4240 10796 4440 10800
rect 4240 10764 4244 10796
rect 4276 10764 4404 10796
rect 4436 10764 4440 10796
rect 4240 10760 4440 10764
rect 4480 10796 4680 10800
rect 4480 10764 4484 10796
rect 4516 10764 4644 10796
rect 4676 10764 4680 10796
rect 4480 10760 4680 10764
rect 4720 10796 5080 10800
rect 4720 10764 4724 10796
rect 4756 10764 4884 10796
rect 4916 10764 5044 10796
rect 5076 10764 5080 10796
rect 4720 10760 5080 10764
rect 5120 10796 5480 10800
rect 5120 10764 5124 10796
rect 5156 10764 5284 10796
rect 5316 10764 5444 10796
rect 5476 10764 5480 10796
rect 5120 10760 5480 10764
rect 5520 10796 5880 10800
rect 5520 10764 5524 10796
rect 5556 10764 5684 10796
rect 5716 10764 5844 10796
rect 5876 10764 5880 10796
rect 5520 10760 5880 10764
rect 5920 10796 6120 10800
rect 5920 10764 5924 10796
rect 5956 10764 6084 10796
rect 6116 10764 6120 10796
rect 5920 10760 6120 10764
rect 6160 10796 6360 10800
rect 6160 10764 6164 10796
rect 6196 10764 6324 10796
rect 6356 10764 6360 10796
rect 6160 10760 6360 10764
rect 4240 10716 4440 10720
rect 4240 10684 4244 10716
rect 4276 10684 4404 10716
rect 4436 10684 4440 10716
rect 4240 10680 4440 10684
rect 4480 10716 4680 10720
rect 4480 10684 4484 10716
rect 4516 10684 4644 10716
rect 4676 10684 4680 10716
rect 4480 10680 4680 10684
rect 4720 10716 5080 10720
rect 4720 10684 4724 10716
rect 4756 10684 4884 10716
rect 4916 10684 5044 10716
rect 5076 10684 5080 10716
rect 4720 10680 5080 10684
rect 5120 10716 5480 10720
rect 5120 10684 5124 10716
rect 5156 10684 5284 10716
rect 5316 10684 5444 10716
rect 5476 10684 5480 10716
rect 5120 10680 5480 10684
rect 5520 10716 5880 10720
rect 5520 10684 5524 10716
rect 5556 10684 5684 10716
rect 5716 10684 5844 10716
rect 5876 10684 5880 10716
rect 5520 10680 5880 10684
rect 5920 10716 6120 10720
rect 5920 10684 5924 10716
rect 5956 10684 6084 10716
rect 6116 10684 6120 10716
rect 5920 10680 6120 10684
rect 6160 10716 6360 10720
rect 6160 10684 6164 10716
rect 6196 10684 6324 10716
rect 6356 10684 6360 10716
rect 6160 10680 6360 10684
rect 4240 10636 4440 10640
rect 4240 10604 4244 10636
rect 4276 10604 4404 10636
rect 4436 10604 4440 10636
rect 4240 10600 4440 10604
rect 4480 10636 4680 10640
rect 4480 10604 4484 10636
rect 4516 10604 4644 10636
rect 4676 10604 4680 10636
rect 4480 10600 4680 10604
rect 4720 10636 5080 10640
rect 4720 10604 4724 10636
rect 4756 10604 4884 10636
rect 4916 10604 5044 10636
rect 5076 10604 5080 10636
rect 4720 10600 5080 10604
rect 5120 10636 5480 10640
rect 5120 10604 5124 10636
rect 5156 10604 5284 10636
rect 5316 10604 5444 10636
rect 5476 10604 5480 10636
rect 5120 10600 5480 10604
rect 5520 10636 5880 10640
rect 5520 10604 5524 10636
rect 5556 10604 5684 10636
rect 5716 10604 5844 10636
rect 5876 10604 5880 10636
rect 5520 10600 5880 10604
rect 5920 10636 6120 10640
rect 5920 10604 5924 10636
rect 5956 10604 6084 10636
rect 6116 10604 6120 10636
rect 5920 10600 6120 10604
rect 6160 10636 6360 10640
rect 6160 10604 6164 10636
rect 6196 10604 6324 10636
rect 6356 10604 6360 10636
rect 6160 10600 6360 10604
rect 4240 10556 4440 10560
rect 4240 10524 4244 10556
rect 4276 10524 4404 10556
rect 4436 10524 4440 10556
rect 4240 10520 4440 10524
rect 4480 10556 4680 10560
rect 4480 10524 4484 10556
rect 4516 10524 4644 10556
rect 4676 10524 4680 10556
rect 4480 10520 4680 10524
rect 4720 10556 5080 10560
rect 4720 10524 4724 10556
rect 4756 10524 4884 10556
rect 4916 10524 5044 10556
rect 5076 10524 5080 10556
rect 4720 10520 5080 10524
rect 5120 10556 5480 10560
rect 5120 10524 5124 10556
rect 5156 10524 5284 10556
rect 5316 10524 5444 10556
rect 5476 10524 5480 10556
rect 5120 10520 5480 10524
rect 5520 10556 5880 10560
rect 5520 10524 5524 10556
rect 5556 10524 5684 10556
rect 5716 10524 5844 10556
rect 5876 10524 5880 10556
rect 5520 10520 5880 10524
rect 5920 10556 6120 10560
rect 5920 10524 5924 10556
rect 5956 10524 6084 10556
rect 6116 10524 6120 10556
rect 5920 10520 6120 10524
rect 6160 10556 6360 10560
rect 6160 10524 6164 10556
rect 6196 10524 6324 10556
rect 6356 10524 6360 10556
rect 6160 10520 6360 10524
rect 4240 10476 4440 10480
rect 4240 10444 4244 10476
rect 4276 10444 4404 10476
rect 4436 10444 4440 10476
rect 4240 10440 4440 10444
rect 4480 10476 4680 10480
rect 4480 10444 4484 10476
rect 4516 10444 4644 10476
rect 4676 10444 4680 10476
rect 4480 10440 4680 10444
rect 4720 10476 5080 10480
rect 4720 10444 4724 10476
rect 4756 10444 4884 10476
rect 4916 10444 5044 10476
rect 5076 10444 5080 10476
rect 4720 10440 5080 10444
rect 5120 10476 5480 10480
rect 5120 10444 5124 10476
rect 5156 10444 5284 10476
rect 5316 10444 5444 10476
rect 5476 10444 5480 10476
rect 5120 10440 5480 10444
rect 5520 10476 5880 10480
rect 5520 10444 5524 10476
rect 5556 10444 5684 10476
rect 5716 10444 5844 10476
rect 5876 10444 5880 10476
rect 5520 10440 5880 10444
rect 5920 10476 6120 10480
rect 5920 10444 5924 10476
rect 5956 10444 6084 10476
rect 6116 10444 6120 10476
rect 5920 10440 6120 10444
rect 6160 10476 6360 10480
rect 6160 10444 6164 10476
rect 6196 10444 6324 10476
rect 6356 10444 6360 10476
rect 6160 10440 6360 10444
rect 4240 10396 4440 10400
rect 4240 10364 4244 10396
rect 4276 10364 4404 10396
rect 4436 10364 4440 10396
rect 4240 10360 4440 10364
rect 4480 10396 4680 10400
rect 4480 10364 4484 10396
rect 4516 10364 4644 10396
rect 4676 10364 4680 10396
rect 4480 10360 4680 10364
rect 4720 10396 5080 10400
rect 4720 10364 4724 10396
rect 4756 10364 4884 10396
rect 4916 10364 5044 10396
rect 5076 10364 5080 10396
rect 4720 10360 5080 10364
rect 5120 10396 5480 10400
rect 5120 10364 5124 10396
rect 5156 10364 5284 10396
rect 5316 10364 5444 10396
rect 5476 10364 5480 10396
rect 5120 10360 5480 10364
rect 5520 10396 5880 10400
rect 5520 10364 5524 10396
rect 5556 10364 5684 10396
rect 5716 10364 5844 10396
rect 5876 10364 5880 10396
rect 5520 10360 5880 10364
rect 5920 10396 6120 10400
rect 5920 10364 5924 10396
rect 5956 10364 6084 10396
rect 6116 10364 6120 10396
rect 5920 10360 6120 10364
rect 6160 10396 6360 10400
rect 6160 10364 6164 10396
rect 6196 10364 6324 10396
rect 6356 10364 6360 10396
rect 6160 10360 6360 10364
rect 4240 10316 4440 10320
rect 4240 10284 4244 10316
rect 4276 10284 4404 10316
rect 4436 10284 4440 10316
rect 4240 10280 4440 10284
rect 4480 10316 4680 10320
rect 4480 10284 4484 10316
rect 4516 10284 4644 10316
rect 4676 10284 4680 10316
rect 4480 10280 4680 10284
rect 4720 10316 5080 10320
rect 4720 10284 4724 10316
rect 4756 10284 4884 10316
rect 4916 10284 5044 10316
rect 5076 10284 5080 10316
rect 4720 10280 5080 10284
rect 5120 10316 5480 10320
rect 5120 10284 5124 10316
rect 5156 10284 5284 10316
rect 5316 10284 5444 10316
rect 5476 10284 5480 10316
rect 5120 10280 5480 10284
rect 5520 10316 5880 10320
rect 5520 10284 5524 10316
rect 5556 10284 5684 10316
rect 5716 10284 5844 10316
rect 5876 10284 5880 10316
rect 5520 10280 5880 10284
rect 5920 10316 6120 10320
rect 5920 10284 5924 10316
rect 5956 10284 6084 10316
rect 6116 10284 6120 10316
rect 5920 10280 6120 10284
rect 6160 10316 6360 10320
rect 6160 10284 6164 10316
rect 6196 10284 6324 10316
rect 6356 10284 6360 10316
rect 6160 10280 6360 10284
rect 4240 10236 4440 10240
rect 4240 10204 4244 10236
rect 4276 10204 4404 10236
rect 4436 10204 4440 10236
rect 4240 10200 4440 10204
rect 4480 10236 4680 10240
rect 4480 10204 4484 10236
rect 4516 10204 4644 10236
rect 4676 10204 4680 10236
rect 4480 10200 4680 10204
rect 4720 10236 5080 10240
rect 4720 10204 4724 10236
rect 4756 10204 4884 10236
rect 4916 10204 5044 10236
rect 5076 10204 5080 10236
rect 4720 10200 5080 10204
rect 5120 10236 5480 10240
rect 5120 10204 5124 10236
rect 5156 10204 5284 10236
rect 5316 10204 5444 10236
rect 5476 10204 5480 10236
rect 5120 10200 5480 10204
rect 5520 10236 5880 10240
rect 5520 10204 5524 10236
rect 5556 10204 5684 10236
rect 5716 10204 5844 10236
rect 5876 10204 5880 10236
rect 5520 10200 5880 10204
rect 5920 10236 6120 10240
rect 5920 10204 5924 10236
rect 5956 10204 6084 10236
rect 6116 10204 6120 10236
rect 5920 10200 6120 10204
rect 6160 10236 6360 10240
rect 6160 10204 6164 10236
rect 6196 10204 6324 10236
rect 6356 10204 6360 10236
rect 6160 10200 6360 10204
rect 4240 10156 4440 10160
rect 4240 10124 4244 10156
rect 4276 10124 4404 10156
rect 4436 10124 4440 10156
rect 4240 10120 4440 10124
rect 4480 10156 4680 10160
rect 4480 10124 4484 10156
rect 4516 10124 4644 10156
rect 4676 10124 4680 10156
rect 4480 10120 4680 10124
rect 4720 10156 5080 10160
rect 4720 10124 4724 10156
rect 4756 10124 4884 10156
rect 4916 10124 5044 10156
rect 5076 10124 5080 10156
rect 4720 10120 5080 10124
rect 5120 10156 5480 10160
rect 5120 10124 5124 10156
rect 5156 10124 5284 10156
rect 5316 10124 5444 10156
rect 5476 10124 5480 10156
rect 5120 10120 5480 10124
rect 5520 10156 5880 10160
rect 5520 10124 5524 10156
rect 5556 10124 5684 10156
rect 5716 10124 5844 10156
rect 5876 10124 5880 10156
rect 5520 10120 5880 10124
rect 5920 10156 6120 10160
rect 5920 10124 5924 10156
rect 5956 10124 6084 10156
rect 6116 10124 6120 10156
rect 5920 10120 6120 10124
rect 6160 10156 6360 10160
rect 6160 10124 6164 10156
rect 6196 10124 6324 10156
rect 6356 10124 6360 10156
rect 6160 10120 6360 10124
rect 4240 10076 4440 10080
rect 4240 10044 4244 10076
rect 4276 10044 4404 10076
rect 4436 10044 4440 10076
rect 4240 10040 4440 10044
rect 4480 10076 4680 10080
rect 4480 10044 4484 10076
rect 4516 10044 4644 10076
rect 4676 10044 4680 10076
rect 4480 10040 4680 10044
rect 4720 10076 5080 10080
rect 4720 10044 4724 10076
rect 4756 10044 4884 10076
rect 4916 10044 5044 10076
rect 5076 10044 5080 10076
rect 4720 10040 5080 10044
rect 5120 10076 5480 10080
rect 5120 10044 5124 10076
rect 5156 10044 5284 10076
rect 5316 10044 5444 10076
rect 5476 10044 5480 10076
rect 5120 10040 5480 10044
rect 5520 10076 5880 10080
rect 5520 10044 5524 10076
rect 5556 10044 5684 10076
rect 5716 10044 5844 10076
rect 5876 10044 5880 10076
rect 5520 10040 5880 10044
rect 5920 10076 6120 10080
rect 5920 10044 5924 10076
rect 5956 10044 6084 10076
rect 6116 10044 6120 10076
rect 5920 10040 6120 10044
rect 6160 10076 6360 10080
rect 6160 10044 6164 10076
rect 6196 10044 6324 10076
rect 6356 10044 6360 10076
rect 6160 10040 6360 10044
rect 4240 9996 4440 10000
rect 4240 9964 4244 9996
rect 4276 9964 4404 9996
rect 4436 9964 4440 9996
rect 4240 9960 4440 9964
rect 4480 9996 4680 10000
rect 4480 9964 4484 9996
rect 4516 9964 4644 9996
rect 4676 9964 4680 9996
rect 4480 9960 4680 9964
rect 4720 9996 5080 10000
rect 4720 9964 4724 9996
rect 4756 9964 4884 9996
rect 4916 9964 5044 9996
rect 5076 9964 5080 9996
rect 4720 9960 5080 9964
rect 5120 9996 5480 10000
rect 5120 9964 5124 9996
rect 5156 9964 5284 9996
rect 5316 9964 5444 9996
rect 5476 9964 5480 9996
rect 5120 9960 5480 9964
rect 5520 9996 5880 10000
rect 5520 9964 5524 9996
rect 5556 9964 5684 9996
rect 5716 9964 5844 9996
rect 5876 9964 5880 9996
rect 5520 9960 5880 9964
rect 5920 9996 6120 10000
rect 5920 9964 5924 9996
rect 5956 9964 6084 9996
rect 6116 9964 6120 9996
rect 5920 9960 6120 9964
rect 6160 9996 6360 10000
rect 6160 9964 6164 9996
rect 6196 9964 6324 9996
rect 6356 9964 6360 9996
rect 6160 9960 6360 9964
rect 4240 9916 4440 9920
rect 4240 9884 4244 9916
rect 4276 9884 4404 9916
rect 4436 9884 4440 9916
rect 4240 9880 4440 9884
rect 4480 9916 4680 9920
rect 4480 9884 4484 9916
rect 4516 9884 4644 9916
rect 4676 9884 4680 9916
rect 4480 9880 4680 9884
rect 4720 9916 5080 9920
rect 4720 9884 4724 9916
rect 4756 9884 4884 9916
rect 4916 9884 5044 9916
rect 5076 9884 5080 9916
rect 4720 9880 5080 9884
rect 5120 9916 5480 9920
rect 5120 9884 5124 9916
rect 5156 9884 5284 9916
rect 5316 9884 5444 9916
rect 5476 9884 5480 9916
rect 5120 9880 5480 9884
rect 5520 9916 5880 9920
rect 5520 9884 5524 9916
rect 5556 9884 5684 9916
rect 5716 9884 5844 9916
rect 5876 9884 5880 9916
rect 5520 9880 5880 9884
rect 5920 9916 6120 9920
rect 5920 9884 5924 9916
rect 5956 9884 6084 9916
rect 6116 9884 6120 9916
rect 5920 9880 6120 9884
rect 6160 9916 6360 9920
rect 6160 9884 6164 9916
rect 6196 9884 6324 9916
rect 6356 9884 6360 9916
rect 6160 9880 6360 9884
rect 4240 9836 4440 9840
rect 4240 9804 4244 9836
rect 4276 9804 4404 9836
rect 4436 9804 4440 9836
rect 4240 9800 4440 9804
rect 4480 9836 4680 9840
rect 4480 9804 4484 9836
rect 4516 9804 4644 9836
rect 4676 9804 4680 9836
rect 4480 9800 4680 9804
rect 4720 9836 5080 9840
rect 4720 9804 4724 9836
rect 4756 9804 4884 9836
rect 4916 9804 5044 9836
rect 5076 9804 5080 9836
rect 4720 9800 5080 9804
rect 5120 9836 5480 9840
rect 5120 9804 5124 9836
rect 5156 9804 5284 9836
rect 5316 9804 5444 9836
rect 5476 9804 5480 9836
rect 5120 9800 5480 9804
rect 5520 9836 5880 9840
rect 5520 9804 5524 9836
rect 5556 9804 5684 9836
rect 5716 9804 5844 9836
rect 5876 9804 5880 9836
rect 5520 9800 5880 9804
rect 5920 9836 6120 9840
rect 5920 9804 5924 9836
rect 5956 9804 6084 9836
rect 6116 9804 6120 9836
rect 5920 9800 6120 9804
rect 6160 9836 6360 9840
rect 6160 9804 6164 9836
rect 6196 9804 6324 9836
rect 6356 9804 6360 9836
rect 6160 9800 6360 9804
rect 4240 9756 4440 9760
rect 4240 9724 4244 9756
rect 4276 9724 4404 9756
rect 4436 9724 4440 9756
rect 4240 9720 4440 9724
rect 4480 9756 4680 9760
rect 4480 9724 4484 9756
rect 4516 9724 4644 9756
rect 4676 9724 4680 9756
rect 4480 9720 4680 9724
rect 4720 9756 5080 9760
rect 4720 9724 4724 9756
rect 4756 9724 4884 9756
rect 4916 9724 5044 9756
rect 5076 9724 5080 9756
rect 4720 9720 5080 9724
rect 5120 9756 5480 9760
rect 5120 9724 5124 9756
rect 5156 9724 5284 9756
rect 5316 9724 5444 9756
rect 5476 9724 5480 9756
rect 5120 9720 5480 9724
rect 5520 9756 5880 9760
rect 5520 9724 5524 9756
rect 5556 9724 5684 9756
rect 5716 9724 5844 9756
rect 5876 9724 5880 9756
rect 5520 9720 5880 9724
rect 5920 9756 6120 9760
rect 5920 9724 5924 9756
rect 5956 9724 6084 9756
rect 6116 9724 6120 9756
rect 5920 9720 6120 9724
rect 6160 9756 6360 9760
rect 6160 9724 6164 9756
rect 6196 9724 6324 9756
rect 6356 9724 6360 9756
rect 6160 9720 6360 9724
rect 4240 9356 4440 9360
rect 4240 9324 4244 9356
rect 4276 9324 4404 9356
rect 4436 9324 4440 9356
rect 4240 9320 4440 9324
rect 4480 9356 4680 9360
rect 4480 9324 4484 9356
rect 4516 9324 4644 9356
rect 4676 9324 4680 9356
rect 4480 9320 4680 9324
rect 4720 9356 5080 9360
rect 4720 9324 4724 9356
rect 4756 9324 4884 9356
rect 4916 9324 5044 9356
rect 5076 9324 5080 9356
rect 4720 9320 5080 9324
rect 5120 9356 5480 9360
rect 5120 9324 5124 9356
rect 5156 9324 5284 9356
rect 5316 9324 5444 9356
rect 5476 9324 5480 9356
rect 5120 9320 5480 9324
rect 5520 9356 5880 9360
rect 5520 9324 5524 9356
rect 5556 9324 5684 9356
rect 5716 9324 5844 9356
rect 5876 9324 5880 9356
rect 5520 9320 5880 9324
rect 5920 9356 6120 9360
rect 5920 9324 5924 9356
rect 5956 9324 6084 9356
rect 6116 9324 6120 9356
rect 5920 9320 6120 9324
rect 6160 9356 6360 9360
rect 6160 9324 6164 9356
rect 6196 9324 6324 9356
rect 6356 9324 6360 9356
rect 6160 9320 6360 9324
rect 4240 9276 4440 9280
rect 4240 9244 4244 9276
rect 4276 9244 4404 9276
rect 4436 9244 4440 9276
rect 4240 9240 4440 9244
rect 4480 9276 4680 9280
rect 4480 9244 4484 9276
rect 4516 9244 4644 9276
rect 4676 9244 4680 9276
rect 4480 9240 4680 9244
rect 4720 9276 5080 9280
rect 4720 9244 4724 9276
rect 4756 9244 4884 9276
rect 4916 9244 5044 9276
rect 5076 9244 5080 9276
rect 4720 9240 5080 9244
rect 5120 9276 5480 9280
rect 5120 9244 5124 9276
rect 5156 9244 5284 9276
rect 5316 9244 5444 9276
rect 5476 9244 5480 9276
rect 5120 9240 5480 9244
rect 5520 9276 5880 9280
rect 5520 9244 5524 9276
rect 5556 9244 5684 9276
rect 5716 9244 5844 9276
rect 5876 9244 5880 9276
rect 5520 9240 5880 9244
rect 5920 9276 6120 9280
rect 5920 9244 5924 9276
rect 5956 9244 6084 9276
rect 6116 9244 6120 9276
rect 5920 9240 6120 9244
rect 6160 9276 6360 9280
rect 6160 9244 6164 9276
rect 6196 9244 6324 9276
rect 6356 9244 6360 9276
rect 6160 9240 6360 9244
rect 4240 9196 4440 9200
rect 4240 9164 4244 9196
rect 4276 9164 4404 9196
rect 4436 9164 4440 9196
rect 4240 9160 4440 9164
rect 4480 9196 4680 9200
rect 4480 9164 4484 9196
rect 4516 9164 4644 9196
rect 4676 9164 4680 9196
rect 4480 9160 4680 9164
rect 4720 9196 5080 9200
rect 4720 9164 4724 9196
rect 4756 9164 4884 9196
rect 4916 9164 5044 9196
rect 5076 9164 5080 9196
rect 4720 9160 5080 9164
rect 5120 9196 5480 9200
rect 5120 9164 5124 9196
rect 5156 9164 5284 9196
rect 5316 9164 5444 9196
rect 5476 9164 5480 9196
rect 5120 9160 5480 9164
rect 5520 9196 5880 9200
rect 5520 9164 5524 9196
rect 5556 9164 5684 9196
rect 5716 9164 5844 9196
rect 5876 9164 5880 9196
rect 5520 9160 5880 9164
rect 5920 9196 6120 9200
rect 5920 9164 5924 9196
rect 5956 9164 6084 9196
rect 6116 9164 6120 9196
rect 5920 9160 6120 9164
rect 6160 9196 6360 9200
rect 6160 9164 6164 9196
rect 6196 9164 6324 9196
rect 6356 9164 6360 9196
rect 6160 9160 6360 9164
rect 4240 8876 4440 8880
rect 4240 8844 4244 8876
rect 4276 8844 4404 8876
rect 4436 8844 4440 8876
rect 4240 8840 4440 8844
rect 4480 8876 4680 8880
rect 4480 8844 4484 8876
rect 4516 8844 4644 8876
rect 4676 8844 4680 8876
rect 4480 8840 4680 8844
rect 4720 8876 5080 8880
rect 4720 8844 4724 8876
rect 4756 8844 4884 8876
rect 4916 8844 5044 8876
rect 5076 8844 5080 8876
rect 4720 8840 5080 8844
rect 5120 8876 5480 8880
rect 5120 8844 5124 8876
rect 5156 8844 5284 8876
rect 5316 8844 5444 8876
rect 5476 8844 5480 8876
rect 5120 8840 5480 8844
rect 5520 8876 5880 8880
rect 5520 8844 5524 8876
rect 5556 8844 5684 8876
rect 5716 8844 5844 8876
rect 5876 8844 5880 8876
rect 5520 8840 5880 8844
rect 5920 8876 6120 8880
rect 5920 8844 5924 8876
rect 5956 8844 6084 8876
rect 6116 8844 6120 8876
rect 5920 8840 6120 8844
rect 6160 8876 6360 8880
rect 6160 8844 6164 8876
rect 6196 8844 6324 8876
rect 6356 8844 6360 8876
rect 6160 8840 6360 8844
rect 4240 8796 4440 8800
rect 4240 8764 4244 8796
rect 4276 8764 4404 8796
rect 4436 8764 4440 8796
rect 4240 8760 4440 8764
rect 4480 8796 4680 8800
rect 4480 8764 4484 8796
rect 4516 8764 4644 8796
rect 4676 8764 4680 8796
rect 4480 8760 4680 8764
rect 4720 8796 5080 8800
rect 4720 8764 4724 8796
rect 4756 8764 4884 8796
rect 4916 8764 5044 8796
rect 5076 8764 5080 8796
rect 4720 8760 5080 8764
rect 5120 8796 5480 8800
rect 5120 8764 5124 8796
rect 5156 8764 5284 8796
rect 5316 8764 5444 8796
rect 5476 8764 5480 8796
rect 5120 8760 5480 8764
rect 5520 8796 5880 8800
rect 5520 8764 5524 8796
rect 5556 8764 5684 8796
rect 5716 8764 5844 8796
rect 5876 8764 5880 8796
rect 5520 8760 5880 8764
rect 5920 8796 6120 8800
rect 5920 8764 5924 8796
rect 5956 8764 6084 8796
rect 6116 8764 6120 8796
rect 5920 8760 6120 8764
rect 6160 8796 6360 8800
rect 6160 8764 6164 8796
rect 6196 8764 6324 8796
rect 6356 8764 6360 8796
rect 6160 8760 6360 8764
rect 4240 8716 4440 8720
rect 4240 8684 4244 8716
rect 4276 8684 4404 8716
rect 4436 8684 4440 8716
rect 4240 8680 4440 8684
rect 4480 8716 4680 8720
rect 4480 8684 4484 8716
rect 4516 8684 4644 8716
rect 4676 8684 4680 8716
rect 4480 8680 4680 8684
rect 4720 8716 5080 8720
rect 4720 8684 4724 8716
rect 4756 8684 4884 8716
rect 4916 8684 5044 8716
rect 5076 8684 5080 8716
rect 4720 8680 5080 8684
rect 5120 8716 5480 8720
rect 5120 8684 5124 8716
rect 5156 8684 5284 8716
rect 5316 8684 5444 8716
rect 5476 8684 5480 8716
rect 5120 8680 5480 8684
rect 5520 8716 5880 8720
rect 5520 8684 5524 8716
rect 5556 8684 5684 8716
rect 5716 8684 5844 8716
rect 5876 8684 5880 8716
rect 5520 8680 5880 8684
rect 5920 8716 6120 8720
rect 5920 8684 5924 8716
rect 5956 8684 6084 8716
rect 6116 8684 6120 8716
rect 5920 8680 6120 8684
rect 6160 8716 6360 8720
rect 6160 8684 6164 8716
rect 6196 8684 6324 8716
rect 6356 8684 6360 8716
rect 6160 8680 6360 8684
rect 4240 8636 4440 8640
rect 4240 8604 4244 8636
rect 4276 8604 4404 8636
rect 4436 8604 4440 8636
rect 4240 8600 4440 8604
rect 4480 8636 4680 8640
rect 4480 8604 4484 8636
rect 4516 8604 4644 8636
rect 4676 8604 4680 8636
rect 4480 8600 4680 8604
rect 4720 8636 5080 8640
rect 4720 8604 4724 8636
rect 4756 8604 4884 8636
rect 4916 8604 5044 8636
rect 5076 8604 5080 8636
rect 4720 8600 5080 8604
rect 5120 8636 5480 8640
rect 5120 8604 5124 8636
rect 5156 8604 5284 8636
rect 5316 8604 5444 8636
rect 5476 8604 5480 8636
rect 5120 8600 5480 8604
rect 5520 8636 5880 8640
rect 5520 8604 5524 8636
rect 5556 8604 5684 8636
rect 5716 8604 5844 8636
rect 5876 8604 5880 8636
rect 5520 8600 5880 8604
rect 5920 8636 6120 8640
rect 5920 8604 5924 8636
rect 5956 8604 6084 8636
rect 6116 8604 6120 8636
rect 5920 8600 6120 8604
rect 6160 8636 6360 8640
rect 6160 8604 6164 8636
rect 6196 8604 6324 8636
rect 6356 8604 6360 8636
rect 6160 8600 6360 8604
rect 4240 8556 4440 8560
rect 4240 8524 4244 8556
rect 4276 8524 4404 8556
rect 4436 8524 4440 8556
rect 4240 8520 4440 8524
rect 4480 8556 4680 8560
rect 4480 8524 4484 8556
rect 4516 8524 4644 8556
rect 4676 8524 4680 8556
rect 4480 8520 4680 8524
rect 4720 8556 5080 8560
rect 4720 8524 4724 8556
rect 4756 8524 4884 8556
rect 4916 8524 5044 8556
rect 5076 8524 5080 8556
rect 4720 8520 5080 8524
rect 5120 8556 5480 8560
rect 5120 8524 5124 8556
rect 5156 8524 5284 8556
rect 5316 8524 5444 8556
rect 5476 8524 5480 8556
rect 5120 8520 5480 8524
rect 5520 8556 5880 8560
rect 5520 8524 5524 8556
rect 5556 8524 5684 8556
rect 5716 8524 5844 8556
rect 5876 8524 5880 8556
rect 5520 8520 5880 8524
rect 5920 8556 6120 8560
rect 5920 8524 5924 8556
rect 5956 8524 6084 8556
rect 6116 8524 6120 8556
rect 5920 8520 6120 8524
rect 6160 8556 6360 8560
rect 6160 8524 6164 8556
rect 6196 8524 6324 8556
rect 6356 8524 6360 8556
rect 6160 8520 6360 8524
rect 4240 7636 4440 7640
rect 4240 7604 4244 7636
rect 4276 7604 4404 7636
rect 4436 7604 4440 7636
rect 4240 7600 4440 7604
rect 4480 7636 4680 7640
rect 4480 7604 4484 7636
rect 4516 7604 4644 7636
rect 4676 7604 4680 7636
rect 4480 7600 4680 7604
rect 4720 7636 5080 7640
rect 4720 7604 4724 7636
rect 4756 7604 4884 7636
rect 4916 7604 5044 7636
rect 5076 7604 5080 7636
rect 4720 7600 5080 7604
rect 5120 7636 5480 7640
rect 5120 7604 5124 7636
rect 5156 7604 5284 7636
rect 5316 7604 5444 7636
rect 5476 7604 5480 7636
rect 5120 7600 5480 7604
rect 5520 7636 5880 7640
rect 5520 7604 5524 7636
rect 5556 7604 5684 7636
rect 5716 7604 5844 7636
rect 5876 7604 5880 7636
rect 5520 7600 5880 7604
rect 5920 7636 6120 7640
rect 5920 7604 5924 7636
rect 5956 7604 6084 7636
rect 6116 7604 6120 7636
rect 5920 7600 6120 7604
rect 6160 7636 6360 7640
rect 6160 7604 6164 7636
rect 6196 7604 6324 7636
rect 6356 7604 6360 7636
rect 6160 7600 6360 7604
rect 4240 7556 4440 7560
rect 4240 7524 4244 7556
rect 4276 7524 4404 7556
rect 4436 7524 4440 7556
rect 4240 7520 4440 7524
rect 4480 7556 4680 7560
rect 4480 7524 4484 7556
rect 4516 7524 4644 7556
rect 4676 7524 4680 7556
rect 4480 7520 4680 7524
rect 4720 7556 5080 7560
rect 4720 7524 4724 7556
rect 4756 7524 4884 7556
rect 4916 7524 5044 7556
rect 5076 7524 5080 7556
rect 4720 7520 5080 7524
rect 5120 7556 5480 7560
rect 5120 7524 5124 7556
rect 5156 7524 5284 7556
rect 5316 7524 5444 7556
rect 5476 7524 5480 7556
rect 5120 7520 5480 7524
rect 5520 7556 5880 7560
rect 5520 7524 5524 7556
rect 5556 7524 5684 7556
rect 5716 7524 5844 7556
rect 5876 7524 5880 7556
rect 5520 7520 5880 7524
rect 5920 7556 6120 7560
rect 5920 7524 5924 7556
rect 5956 7524 6084 7556
rect 6116 7524 6120 7556
rect 5920 7520 6120 7524
rect 6160 7556 6360 7560
rect 6160 7524 6164 7556
rect 6196 7524 6324 7556
rect 6356 7524 6360 7556
rect 6160 7520 6360 7524
rect 4240 7476 4440 7480
rect 4240 7444 4244 7476
rect 4276 7444 4404 7476
rect 4436 7444 4440 7476
rect 4240 7440 4440 7444
rect 4480 7476 4680 7480
rect 4480 7444 4484 7476
rect 4516 7444 4644 7476
rect 4676 7444 4680 7476
rect 4480 7440 4680 7444
rect 4720 7476 5080 7480
rect 4720 7444 4724 7476
rect 4756 7444 4884 7476
rect 4916 7444 5044 7476
rect 5076 7444 5080 7476
rect 4720 7440 5080 7444
rect 5120 7476 5480 7480
rect 5120 7444 5124 7476
rect 5156 7444 5284 7476
rect 5316 7444 5444 7476
rect 5476 7444 5480 7476
rect 5120 7440 5480 7444
rect 5520 7476 5880 7480
rect 5520 7444 5524 7476
rect 5556 7444 5684 7476
rect 5716 7444 5844 7476
rect 5876 7444 5880 7476
rect 5520 7440 5880 7444
rect 5920 7476 6120 7480
rect 5920 7444 5924 7476
rect 5956 7444 6084 7476
rect 6116 7444 6120 7476
rect 5920 7440 6120 7444
rect 6160 7476 6360 7480
rect 6160 7444 6164 7476
rect 6196 7444 6324 7476
rect 6356 7444 6360 7476
rect 6160 7440 6360 7444
rect 4240 7396 4440 7400
rect 4240 7364 4244 7396
rect 4276 7364 4404 7396
rect 4436 7364 4440 7396
rect 4240 7360 4440 7364
rect 4480 7396 4680 7400
rect 4480 7364 4484 7396
rect 4516 7364 4644 7396
rect 4676 7364 4680 7396
rect 4480 7360 4680 7364
rect 4720 7396 5080 7400
rect 4720 7364 4724 7396
rect 4756 7364 4884 7396
rect 4916 7364 5044 7396
rect 5076 7364 5080 7396
rect 4720 7360 5080 7364
rect 5120 7396 5480 7400
rect 5120 7364 5124 7396
rect 5156 7364 5284 7396
rect 5316 7364 5444 7396
rect 5476 7364 5480 7396
rect 5120 7360 5480 7364
rect 5520 7396 5880 7400
rect 5520 7364 5524 7396
rect 5556 7364 5684 7396
rect 5716 7364 5844 7396
rect 5876 7364 5880 7396
rect 5520 7360 5880 7364
rect 5920 7396 6120 7400
rect 5920 7364 5924 7396
rect 5956 7364 6084 7396
rect 6116 7364 6120 7396
rect 5920 7360 6120 7364
rect 6160 7396 6360 7400
rect 6160 7364 6164 7396
rect 6196 7364 6324 7396
rect 6356 7364 6360 7396
rect 6160 7360 6360 7364
rect 4240 7316 4440 7320
rect 4240 7284 4244 7316
rect 4276 7284 4404 7316
rect 4436 7284 4440 7316
rect 4240 7280 4440 7284
rect 4480 7316 4680 7320
rect 4480 7284 4484 7316
rect 4516 7284 4644 7316
rect 4676 7284 4680 7316
rect 4480 7280 4680 7284
rect 4720 7316 5080 7320
rect 4720 7284 4724 7316
rect 4756 7284 4884 7316
rect 4916 7284 5044 7316
rect 5076 7284 5080 7316
rect 4720 7280 5080 7284
rect 5120 7316 5480 7320
rect 5120 7284 5124 7316
rect 5156 7284 5284 7316
rect 5316 7284 5444 7316
rect 5476 7284 5480 7316
rect 5120 7280 5480 7284
rect 5520 7316 5880 7320
rect 5520 7284 5524 7316
rect 5556 7284 5684 7316
rect 5716 7284 5844 7316
rect 5876 7284 5880 7316
rect 5520 7280 5880 7284
rect 5920 7316 6120 7320
rect 5920 7284 5924 7316
rect 5956 7284 6084 7316
rect 6116 7284 6120 7316
rect 5920 7280 6120 7284
rect 6160 7316 6360 7320
rect 6160 7284 6164 7316
rect 6196 7284 6324 7316
rect 6356 7284 6360 7316
rect 6160 7280 6360 7284
rect 4240 7236 4440 7240
rect 4240 7204 4244 7236
rect 4276 7204 4404 7236
rect 4436 7204 4440 7236
rect 4240 7200 4440 7204
rect 4480 7236 4680 7240
rect 4480 7204 4484 7236
rect 4516 7204 4644 7236
rect 4676 7204 4680 7236
rect 4480 7200 4680 7204
rect 4720 7236 5080 7240
rect 4720 7204 4724 7236
rect 4756 7204 4884 7236
rect 4916 7204 5044 7236
rect 5076 7204 5080 7236
rect 4720 7200 5080 7204
rect 5120 7236 5480 7240
rect 5120 7204 5124 7236
rect 5156 7204 5284 7236
rect 5316 7204 5444 7236
rect 5476 7204 5480 7236
rect 5120 7200 5480 7204
rect 5520 7236 5880 7240
rect 5520 7204 5524 7236
rect 5556 7204 5684 7236
rect 5716 7204 5844 7236
rect 5876 7204 5880 7236
rect 5520 7200 5880 7204
rect 5920 7236 6120 7240
rect 5920 7204 5924 7236
rect 5956 7204 6084 7236
rect 6116 7204 6120 7236
rect 5920 7200 6120 7204
rect 6160 7236 6360 7240
rect 6160 7204 6164 7236
rect 6196 7204 6324 7236
rect 6356 7204 6360 7236
rect 6160 7200 6360 7204
rect 4240 7156 4440 7160
rect 4240 7124 4244 7156
rect 4276 7124 4404 7156
rect 4436 7124 4440 7156
rect 4240 7120 4440 7124
rect 4480 7156 4680 7160
rect 4480 7124 4484 7156
rect 4516 7124 4644 7156
rect 4676 7124 4680 7156
rect 4480 7120 4680 7124
rect 4720 7156 5080 7160
rect 4720 7124 4724 7156
rect 4756 7124 4884 7156
rect 4916 7124 5044 7156
rect 5076 7124 5080 7156
rect 4720 7120 5080 7124
rect 5120 7156 5480 7160
rect 5120 7124 5124 7156
rect 5156 7124 5284 7156
rect 5316 7124 5444 7156
rect 5476 7124 5480 7156
rect 5120 7120 5480 7124
rect 5520 7156 5880 7160
rect 5520 7124 5524 7156
rect 5556 7124 5684 7156
rect 5716 7124 5844 7156
rect 5876 7124 5880 7156
rect 5520 7120 5880 7124
rect 5920 7156 6120 7160
rect 5920 7124 5924 7156
rect 5956 7124 6084 7156
rect 6116 7124 6120 7156
rect 5920 7120 6120 7124
rect 6160 7156 6360 7160
rect 6160 7124 6164 7156
rect 6196 7124 6324 7156
rect 6356 7124 6360 7156
rect 6160 7120 6360 7124
rect 4240 7076 4440 7080
rect 4240 7044 4244 7076
rect 4276 7044 4404 7076
rect 4436 7044 4440 7076
rect 4240 7040 4440 7044
rect 4480 7076 4680 7080
rect 4480 7044 4484 7076
rect 4516 7044 4644 7076
rect 4676 7044 4680 7076
rect 4480 7040 4680 7044
rect 4720 7076 5080 7080
rect 4720 7044 4724 7076
rect 4756 7044 4884 7076
rect 4916 7044 5044 7076
rect 5076 7044 5080 7076
rect 4720 7040 5080 7044
rect 5120 7076 5480 7080
rect 5120 7044 5124 7076
rect 5156 7044 5284 7076
rect 5316 7044 5444 7076
rect 5476 7044 5480 7076
rect 5120 7040 5480 7044
rect 5520 7076 5880 7080
rect 5520 7044 5524 7076
rect 5556 7044 5684 7076
rect 5716 7044 5844 7076
rect 5876 7044 5880 7076
rect 5520 7040 5880 7044
rect 5920 7076 6120 7080
rect 5920 7044 5924 7076
rect 5956 7044 6084 7076
rect 6116 7044 6120 7076
rect 5920 7040 6120 7044
rect 6160 7076 6360 7080
rect 6160 7044 6164 7076
rect 6196 7044 6324 7076
rect 6356 7044 6360 7076
rect 6160 7040 6360 7044
rect 4240 6756 4440 6760
rect 4240 6724 4244 6756
rect 4276 6724 4404 6756
rect 4436 6724 4440 6756
rect 4240 6720 4440 6724
rect 4480 6756 4680 6760
rect 4480 6724 4484 6756
rect 4516 6724 4644 6756
rect 4676 6724 4680 6756
rect 4480 6720 4680 6724
rect 4720 6756 5080 6760
rect 4720 6724 4724 6756
rect 4756 6724 4884 6756
rect 4916 6724 5044 6756
rect 5076 6724 5080 6756
rect 4720 6720 5080 6724
rect 5120 6756 5480 6760
rect 5120 6724 5124 6756
rect 5156 6724 5284 6756
rect 5316 6724 5444 6756
rect 5476 6724 5480 6756
rect 5120 6720 5480 6724
rect 5520 6756 5880 6760
rect 5520 6724 5524 6756
rect 5556 6724 5684 6756
rect 5716 6724 5844 6756
rect 5876 6724 5880 6756
rect 5520 6720 5880 6724
rect 5920 6756 6120 6760
rect 5920 6724 5924 6756
rect 5956 6724 6084 6756
rect 6116 6724 6120 6756
rect 5920 6720 6120 6724
rect 6160 6756 6360 6760
rect 6160 6724 6164 6756
rect 6196 6724 6324 6756
rect 6356 6724 6360 6756
rect 6160 6720 6360 6724
rect 4240 6676 4440 6680
rect 4240 6644 4244 6676
rect 4276 6644 4404 6676
rect 4436 6644 4440 6676
rect 4240 6640 4440 6644
rect 4480 6676 4680 6680
rect 4480 6644 4484 6676
rect 4516 6644 4644 6676
rect 4676 6644 4680 6676
rect 4480 6640 4680 6644
rect 4720 6676 5080 6680
rect 4720 6644 4724 6676
rect 4756 6644 4884 6676
rect 4916 6644 5044 6676
rect 5076 6644 5080 6676
rect 4720 6640 5080 6644
rect 5120 6676 5480 6680
rect 5120 6644 5124 6676
rect 5156 6644 5284 6676
rect 5316 6644 5444 6676
rect 5476 6644 5480 6676
rect 5120 6640 5480 6644
rect 5520 6676 5880 6680
rect 5520 6644 5524 6676
rect 5556 6644 5684 6676
rect 5716 6644 5844 6676
rect 5876 6644 5880 6676
rect 5520 6640 5880 6644
rect 5920 6676 6120 6680
rect 5920 6644 5924 6676
rect 5956 6644 6084 6676
rect 6116 6644 6120 6676
rect 5920 6640 6120 6644
rect 6160 6676 6360 6680
rect 6160 6644 6164 6676
rect 6196 6644 6324 6676
rect 6356 6644 6360 6676
rect 6160 6640 6360 6644
rect 4240 6596 4440 6600
rect 4240 6564 4244 6596
rect 4276 6564 4404 6596
rect 4436 6564 4440 6596
rect 4240 6560 4440 6564
rect 4480 6596 4680 6600
rect 4480 6564 4484 6596
rect 4516 6564 4644 6596
rect 4676 6564 4680 6596
rect 4480 6560 4680 6564
rect 4720 6596 5080 6600
rect 4720 6564 4724 6596
rect 4756 6564 4884 6596
rect 4916 6564 5044 6596
rect 5076 6564 5080 6596
rect 4720 6560 5080 6564
rect 5120 6596 5480 6600
rect 5120 6564 5124 6596
rect 5156 6564 5284 6596
rect 5316 6564 5444 6596
rect 5476 6564 5480 6596
rect 5120 6560 5480 6564
rect 5520 6596 5880 6600
rect 5520 6564 5524 6596
rect 5556 6564 5684 6596
rect 5716 6564 5844 6596
rect 5876 6564 5880 6596
rect 5520 6560 5880 6564
rect 5920 6596 6120 6600
rect 5920 6564 5924 6596
rect 5956 6564 6084 6596
rect 6116 6564 6120 6596
rect 5920 6560 6120 6564
rect 6160 6596 6360 6600
rect 6160 6564 6164 6596
rect 6196 6564 6324 6596
rect 6356 6564 6360 6596
rect 6160 6560 6360 6564
rect 4240 6516 4440 6520
rect 4240 6484 4244 6516
rect 4276 6484 4404 6516
rect 4436 6484 4440 6516
rect 4240 6480 4440 6484
rect 4480 6516 4680 6520
rect 4480 6484 4484 6516
rect 4516 6484 4644 6516
rect 4676 6484 4680 6516
rect 4480 6480 4680 6484
rect 4720 6516 5080 6520
rect 4720 6484 4724 6516
rect 4756 6484 4884 6516
rect 4916 6484 5044 6516
rect 5076 6484 5080 6516
rect 4720 6480 5080 6484
rect 5120 6516 5480 6520
rect 5120 6484 5124 6516
rect 5156 6484 5284 6516
rect 5316 6484 5444 6516
rect 5476 6484 5480 6516
rect 5120 6480 5480 6484
rect 5520 6516 5880 6520
rect 5520 6484 5524 6516
rect 5556 6484 5684 6516
rect 5716 6484 5844 6516
rect 5876 6484 5880 6516
rect 5520 6480 5880 6484
rect 5920 6516 6120 6520
rect 5920 6484 5924 6516
rect 5956 6484 6084 6516
rect 6116 6484 6120 6516
rect 5920 6480 6120 6484
rect 6160 6516 6360 6520
rect 6160 6484 6164 6516
rect 6196 6484 6324 6516
rect 6356 6484 6360 6516
rect 6160 6480 6360 6484
rect 4240 6436 4440 6440
rect 4240 6404 4244 6436
rect 4276 6404 4404 6436
rect 4436 6404 4440 6436
rect 4240 6400 4440 6404
rect 4480 6436 4680 6440
rect 4480 6404 4484 6436
rect 4516 6404 4644 6436
rect 4676 6404 4680 6436
rect 4480 6400 4680 6404
rect 4720 6436 5080 6440
rect 4720 6404 4724 6436
rect 4756 6404 4884 6436
rect 4916 6404 5044 6436
rect 5076 6404 5080 6436
rect 4720 6400 5080 6404
rect 5120 6436 5480 6440
rect 5120 6404 5124 6436
rect 5156 6404 5284 6436
rect 5316 6404 5444 6436
rect 5476 6404 5480 6436
rect 5120 6400 5480 6404
rect 5520 6436 5880 6440
rect 5520 6404 5524 6436
rect 5556 6404 5684 6436
rect 5716 6404 5844 6436
rect 5876 6404 5880 6436
rect 5520 6400 5880 6404
rect 5920 6436 6120 6440
rect 5920 6404 5924 6436
rect 5956 6404 6084 6436
rect 6116 6404 6120 6436
rect 5920 6400 6120 6404
rect 6160 6436 6360 6440
rect 6160 6404 6164 6436
rect 6196 6404 6324 6436
rect 6356 6404 6360 6436
rect 6160 6400 6360 6404
rect 4240 6356 4440 6360
rect 4240 6324 4244 6356
rect 4276 6324 4404 6356
rect 4436 6324 4440 6356
rect 4240 6320 4440 6324
rect 4480 6356 4680 6360
rect 4480 6324 4484 6356
rect 4516 6324 4644 6356
rect 4676 6324 4680 6356
rect 4480 6320 4680 6324
rect 4720 6356 5080 6360
rect 4720 6324 4724 6356
rect 4756 6324 4884 6356
rect 4916 6324 5044 6356
rect 5076 6324 5080 6356
rect 4720 6320 5080 6324
rect 5120 6356 5480 6360
rect 5120 6324 5124 6356
rect 5156 6324 5284 6356
rect 5316 6324 5444 6356
rect 5476 6324 5480 6356
rect 5120 6320 5480 6324
rect 5520 6356 5880 6360
rect 5520 6324 5524 6356
rect 5556 6324 5684 6356
rect 5716 6324 5844 6356
rect 5876 6324 5880 6356
rect 5520 6320 5880 6324
rect 5920 6356 6120 6360
rect 5920 6324 5924 6356
rect 5956 6324 6084 6356
rect 6116 6324 6120 6356
rect 5920 6320 6120 6324
rect 6160 6356 6360 6360
rect 6160 6324 6164 6356
rect 6196 6324 6324 6356
rect 6356 6324 6360 6356
rect 6160 6320 6360 6324
rect 4240 5796 4440 5800
rect 4240 5764 4244 5796
rect 4276 5764 4404 5796
rect 4436 5764 4440 5796
rect 4240 5760 4440 5764
rect 4480 5796 4680 5800
rect 4480 5764 4484 5796
rect 4516 5764 4644 5796
rect 4676 5764 4680 5796
rect 4480 5760 4680 5764
rect 4720 5796 5080 5800
rect 4720 5764 4724 5796
rect 4756 5764 4884 5796
rect 4916 5764 5044 5796
rect 5076 5764 5080 5796
rect 4720 5760 5080 5764
rect 5120 5796 5480 5800
rect 5120 5764 5124 5796
rect 5156 5764 5284 5796
rect 5316 5764 5444 5796
rect 5476 5764 5480 5796
rect 5120 5760 5480 5764
rect 5520 5796 5880 5800
rect 5520 5764 5524 5796
rect 5556 5764 5684 5796
rect 5716 5764 5844 5796
rect 5876 5764 5880 5796
rect 5520 5760 5880 5764
rect 5920 5796 6120 5800
rect 5920 5764 5924 5796
rect 5956 5764 6084 5796
rect 6116 5764 6120 5796
rect 5920 5760 6120 5764
rect 6160 5796 6360 5800
rect 6160 5764 6164 5796
rect 6196 5764 6324 5796
rect 6356 5764 6360 5796
rect 6160 5760 6360 5764
rect 4240 5716 4440 5720
rect 4240 5684 4244 5716
rect 4276 5684 4404 5716
rect 4436 5684 4440 5716
rect 4240 5680 4440 5684
rect 4480 5716 4680 5720
rect 4480 5684 4484 5716
rect 4516 5684 4644 5716
rect 4676 5684 4680 5716
rect 4480 5680 4680 5684
rect 4720 5716 5080 5720
rect 4720 5684 4724 5716
rect 4756 5684 4884 5716
rect 4916 5684 5044 5716
rect 5076 5684 5080 5716
rect 4720 5680 5080 5684
rect 5120 5716 5480 5720
rect 5120 5684 5124 5716
rect 5156 5684 5284 5716
rect 5316 5684 5444 5716
rect 5476 5684 5480 5716
rect 5120 5680 5480 5684
rect 5520 5716 5880 5720
rect 5520 5684 5524 5716
rect 5556 5684 5684 5716
rect 5716 5684 5844 5716
rect 5876 5684 5880 5716
rect 5520 5680 5880 5684
rect 5920 5716 6120 5720
rect 5920 5684 5924 5716
rect 5956 5684 6084 5716
rect 6116 5684 6120 5716
rect 5920 5680 6120 5684
rect 6160 5716 6360 5720
rect 6160 5684 6164 5716
rect 6196 5684 6324 5716
rect 6356 5684 6360 5716
rect 6160 5680 6360 5684
rect 4240 5636 4440 5640
rect 4240 5604 4244 5636
rect 4276 5604 4404 5636
rect 4436 5604 4440 5636
rect 4240 5600 4440 5604
rect 4480 5636 4680 5640
rect 4480 5604 4484 5636
rect 4516 5604 4644 5636
rect 4676 5604 4680 5636
rect 4480 5600 4680 5604
rect 4720 5636 5080 5640
rect 4720 5604 4724 5636
rect 4756 5604 4884 5636
rect 4916 5604 5044 5636
rect 5076 5604 5080 5636
rect 4720 5600 5080 5604
rect 5120 5636 5480 5640
rect 5120 5604 5124 5636
rect 5156 5604 5284 5636
rect 5316 5604 5444 5636
rect 5476 5604 5480 5636
rect 5120 5600 5480 5604
rect 5520 5636 5880 5640
rect 5520 5604 5524 5636
rect 5556 5604 5684 5636
rect 5716 5604 5844 5636
rect 5876 5604 5880 5636
rect 5520 5600 5880 5604
rect 5920 5636 6120 5640
rect 5920 5604 5924 5636
rect 5956 5604 6084 5636
rect 6116 5604 6120 5636
rect 5920 5600 6120 5604
rect 6160 5636 6360 5640
rect 6160 5604 6164 5636
rect 6196 5604 6324 5636
rect 6356 5604 6360 5636
rect 6160 5600 6360 5604
rect 4240 5556 4440 5560
rect 4240 5524 4244 5556
rect 4276 5524 4404 5556
rect 4436 5524 4440 5556
rect 4240 5520 4440 5524
rect 4480 5556 4680 5560
rect 4480 5524 4484 5556
rect 4516 5524 4644 5556
rect 4676 5524 4680 5556
rect 4480 5520 4680 5524
rect 4720 5556 5080 5560
rect 4720 5524 4724 5556
rect 4756 5524 4884 5556
rect 4916 5524 5044 5556
rect 5076 5524 5080 5556
rect 4720 5520 5080 5524
rect 5120 5556 5480 5560
rect 5120 5524 5124 5556
rect 5156 5524 5284 5556
rect 5316 5524 5444 5556
rect 5476 5524 5480 5556
rect 5120 5520 5480 5524
rect 5520 5556 5880 5560
rect 5520 5524 5524 5556
rect 5556 5524 5684 5556
rect 5716 5524 5844 5556
rect 5876 5524 5880 5556
rect 5520 5520 5880 5524
rect 5920 5556 6120 5560
rect 5920 5524 5924 5556
rect 5956 5524 6084 5556
rect 6116 5524 6120 5556
rect 5920 5520 6120 5524
rect 6160 5556 6360 5560
rect 6160 5524 6164 5556
rect 6196 5524 6324 5556
rect 6356 5524 6360 5556
rect 6160 5520 6360 5524
rect 4240 5476 4440 5480
rect 4240 5444 4244 5476
rect 4276 5444 4404 5476
rect 4436 5444 4440 5476
rect 4240 5440 4440 5444
rect 4480 5476 4680 5480
rect 4480 5444 4484 5476
rect 4516 5444 4644 5476
rect 4676 5444 4680 5476
rect 4480 5440 4680 5444
rect 4720 5476 5080 5480
rect 4720 5444 4724 5476
rect 4756 5444 4884 5476
rect 4916 5444 5044 5476
rect 5076 5444 5080 5476
rect 4720 5440 5080 5444
rect 5120 5476 5480 5480
rect 5120 5444 5124 5476
rect 5156 5444 5284 5476
rect 5316 5444 5444 5476
rect 5476 5444 5480 5476
rect 5120 5440 5480 5444
rect 5520 5476 5880 5480
rect 5520 5444 5524 5476
rect 5556 5444 5684 5476
rect 5716 5444 5844 5476
rect 5876 5444 5880 5476
rect 5520 5440 5880 5444
rect 5920 5476 6120 5480
rect 5920 5444 5924 5476
rect 5956 5444 6084 5476
rect 6116 5444 6120 5476
rect 5920 5440 6120 5444
rect 6160 5476 6360 5480
rect 6160 5444 6164 5476
rect 6196 5444 6324 5476
rect 6356 5444 6360 5476
rect 6160 5440 6360 5444
rect 4240 5396 4440 5400
rect 4240 5364 4244 5396
rect 4276 5364 4404 5396
rect 4436 5364 4440 5396
rect 4240 5360 4440 5364
rect 4480 5396 4680 5400
rect 4480 5364 4484 5396
rect 4516 5364 4644 5396
rect 4676 5364 4680 5396
rect 4480 5360 4680 5364
rect 4720 5396 5080 5400
rect 4720 5364 4724 5396
rect 4756 5364 4884 5396
rect 4916 5364 5044 5396
rect 5076 5364 5080 5396
rect 4720 5360 5080 5364
rect 5120 5396 5480 5400
rect 5120 5364 5124 5396
rect 5156 5364 5284 5396
rect 5316 5364 5444 5396
rect 5476 5364 5480 5396
rect 5120 5360 5480 5364
rect 5520 5396 5880 5400
rect 5520 5364 5524 5396
rect 5556 5364 5684 5396
rect 5716 5364 5844 5396
rect 5876 5364 5880 5396
rect 5520 5360 5880 5364
rect 5920 5396 6120 5400
rect 5920 5364 5924 5396
rect 5956 5364 6084 5396
rect 6116 5364 6120 5396
rect 5920 5360 6120 5364
rect 6160 5396 6360 5400
rect 6160 5364 6164 5396
rect 6196 5364 6324 5396
rect 6356 5364 6360 5396
rect 6160 5360 6360 5364
rect 4240 5316 4440 5320
rect 4240 5284 4244 5316
rect 4276 5284 4404 5316
rect 4436 5284 4440 5316
rect 4240 5280 4440 5284
rect 4480 5316 4680 5320
rect 4480 5284 4484 5316
rect 4516 5284 4644 5316
rect 4676 5284 4680 5316
rect 4480 5280 4680 5284
rect 4720 5316 5080 5320
rect 4720 5284 4724 5316
rect 4756 5284 4884 5316
rect 4916 5284 5044 5316
rect 5076 5284 5080 5316
rect 4720 5280 5080 5284
rect 5120 5316 5480 5320
rect 5120 5284 5124 5316
rect 5156 5284 5284 5316
rect 5316 5284 5444 5316
rect 5476 5284 5480 5316
rect 5120 5280 5480 5284
rect 5520 5316 5880 5320
rect 5520 5284 5524 5316
rect 5556 5284 5684 5316
rect 5716 5284 5844 5316
rect 5876 5284 5880 5316
rect 5520 5280 5880 5284
rect 5920 5316 6120 5320
rect 5920 5284 5924 5316
rect 5956 5284 6084 5316
rect 6116 5284 6120 5316
rect 5920 5280 6120 5284
rect 6160 5316 6360 5320
rect 6160 5284 6164 5316
rect 6196 5284 6324 5316
rect 6356 5284 6360 5316
rect 6160 5280 6360 5284
rect 4240 5236 4440 5240
rect 4240 5204 4244 5236
rect 4276 5204 4404 5236
rect 4436 5204 4440 5236
rect 4240 5200 4440 5204
rect 4480 5236 4680 5240
rect 4480 5204 4484 5236
rect 4516 5204 4644 5236
rect 4676 5204 4680 5236
rect 4480 5200 4680 5204
rect 4720 5236 5080 5240
rect 4720 5204 4724 5236
rect 4756 5204 4884 5236
rect 4916 5204 5044 5236
rect 5076 5204 5080 5236
rect 4720 5200 5080 5204
rect 5120 5236 5480 5240
rect 5120 5204 5124 5236
rect 5156 5204 5284 5236
rect 5316 5204 5444 5236
rect 5476 5204 5480 5236
rect 5120 5200 5480 5204
rect 5520 5236 5880 5240
rect 5520 5204 5524 5236
rect 5556 5204 5684 5236
rect 5716 5204 5844 5236
rect 5876 5204 5880 5236
rect 5520 5200 5880 5204
rect 5920 5236 6120 5240
rect 5920 5204 5924 5236
rect 5956 5204 6084 5236
rect 6116 5204 6120 5236
rect 5920 5200 6120 5204
rect 6160 5236 6360 5240
rect 6160 5204 6164 5236
rect 6196 5204 6324 5236
rect 6356 5204 6360 5236
rect 6160 5200 6360 5204
rect 4240 5156 4440 5160
rect 4240 5124 4244 5156
rect 4276 5124 4404 5156
rect 4436 5124 4440 5156
rect 4240 5120 4440 5124
rect 4480 5156 4680 5160
rect 4480 5124 4484 5156
rect 4516 5124 4644 5156
rect 4676 5124 4680 5156
rect 4480 5120 4680 5124
rect 4720 5156 5080 5160
rect 4720 5124 4724 5156
rect 4756 5124 4884 5156
rect 4916 5124 5044 5156
rect 5076 5124 5080 5156
rect 4720 5120 5080 5124
rect 5120 5156 5480 5160
rect 5120 5124 5124 5156
rect 5156 5124 5284 5156
rect 5316 5124 5444 5156
rect 5476 5124 5480 5156
rect 5120 5120 5480 5124
rect 5520 5156 5880 5160
rect 5520 5124 5524 5156
rect 5556 5124 5684 5156
rect 5716 5124 5844 5156
rect 5876 5124 5880 5156
rect 5520 5120 5880 5124
rect 5920 5156 6120 5160
rect 5920 5124 5924 5156
rect 5956 5124 6084 5156
rect 6116 5124 6120 5156
rect 5920 5120 6120 5124
rect 6160 5156 6360 5160
rect 6160 5124 6164 5156
rect 6196 5124 6324 5156
rect 6356 5124 6360 5156
rect 6160 5120 6360 5124
rect 4240 5076 4440 5080
rect 4240 5044 4244 5076
rect 4276 5044 4404 5076
rect 4436 5044 4440 5076
rect 4240 5040 4440 5044
rect 4480 5076 4680 5080
rect 4480 5044 4484 5076
rect 4516 5044 4644 5076
rect 4676 5044 4680 5076
rect 4480 5040 4680 5044
rect 4720 5076 5080 5080
rect 4720 5044 4724 5076
rect 4756 5044 4884 5076
rect 4916 5044 5044 5076
rect 5076 5044 5080 5076
rect 4720 5040 5080 5044
rect 5120 5076 5480 5080
rect 5120 5044 5124 5076
rect 5156 5044 5284 5076
rect 5316 5044 5444 5076
rect 5476 5044 5480 5076
rect 5120 5040 5480 5044
rect 5520 5076 5880 5080
rect 5520 5044 5524 5076
rect 5556 5044 5684 5076
rect 5716 5044 5844 5076
rect 5876 5044 5880 5076
rect 5520 5040 5880 5044
rect 5920 5076 6120 5080
rect 5920 5044 5924 5076
rect 5956 5044 6084 5076
rect 6116 5044 6120 5076
rect 5920 5040 6120 5044
rect 6160 5076 6360 5080
rect 6160 5044 6164 5076
rect 6196 5044 6324 5076
rect 6356 5044 6360 5076
rect 6160 5040 6360 5044
rect 4240 4996 4440 5000
rect 4240 4964 4244 4996
rect 4276 4964 4404 4996
rect 4436 4964 4440 4996
rect 4240 4960 4440 4964
rect 4480 4996 4680 5000
rect 4480 4964 4484 4996
rect 4516 4964 4644 4996
rect 4676 4964 4680 4996
rect 4480 4960 4680 4964
rect 4720 4996 5080 5000
rect 4720 4964 4724 4996
rect 4756 4964 4884 4996
rect 4916 4964 5044 4996
rect 5076 4964 5080 4996
rect 4720 4960 5080 4964
rect 5120 4996 5480 5000
rect 5120 4964 5124 4996
rect 5156 4964 5284 4996
rect 5316 4964 5444 4996
rect 5476 4964 5480 4996
rect 5120 4960 5480 4964
rect 5520 4996 5880 5000
rect 5520 4964 5524 4996
rect 5556 4964 5684 4996
rect 5716 4964 5844 4996
rect 5876 4964 5880 4996
rect 5520 4960 5880 4964
rect 5920 4996 6120 5000
rect 5920 4964 5924 4996
rect 5956 4964 6084 4996
rect 6116 4964 6120 4996
rect 5920 4960 6120 4964
rect 6160 4996 6360 5000
rect 6160 4964 6164 4996
rect 6196 4964 6324 4996
rect 6356 4964 6360 4996
rect 6160 4960 6360 4964
rect 4240 4436 4440 4440
rect 4240 4404 4244 4436
rect 4276 4404 4404 4436
rect 4436 4404 4440 4436
rect 4240 4400 4440 4404
rect 4480 4436 4680 4440
rect 4480 4404 4484 4436
rect 4516 4404 4644 4436
rect 4676 4404 4680 4436
rect 4480 4400 4680 4404
rect 4720 4436 5080 4440
rect 4720 4404 4724 4436
rect 4756 4404 4884 4436
rect 4916 4404 5044 4436
rect 5076 4404 5080 4436
rect 4720 4400 5080 4404
rect 5120 4436 5480 4440
rect 5120 4404 5124 4436
rect 5156 4404 5284 4436
rect 5316 4404 5444 4436
rect 5476 4404 5480 4436
rect 5120 4400 5480 4404
rect 5520 4436 5880 4440
rect 5520 4404 5524 4436
rect 5556 4404 5684 4436
rect 5716 4404 5844 4436
rect 5876 4404 5880 4436
rect 5520 4400 5880 4404
rect 5920 4436 6120 4440
rect 5920 4404 5924 4436
rect 5956 4404 6084 4436
rect 6116 4404 6120 4436
rect 5920 4400 6120 4404
rect 6160 4436 6360 4440
rect 6160 4404 6164 4436
rect 6196 4404 6324 4436
rect 6356 4404 6360 4436
rect 6160 4400 6360 4404
rect 4240 4356 4440 4360
rect 4240 4324 4244 4356
rect 4276 4324 4404 4356
rect 4436 4324 4440 4356
rect 4240 4320 4440 4324
rect 4480 4356 4680 4360
rect 4480 4324 4484 4356
rect 4516 4324 4644 4356
rect 4676 4324 4680 4356
rect 4480 4320 4680 4324
rect 4720 4356 5080 4360
rect 4720 4324 4724 4356
rect 4756 4324 4884 4356
rect 4916 4324 5044 4356
rect 5076 4324 5080 4356
rect 4720 4320 5080 4324
rect 5120 4356 5480 4360
rect 5120 4324 5124 4356
rect 5156 4324 5284 4356
rect 5316 4324 5444 4356
rect 5476 4324 5480 4356
rect 5120 4320 5480 4324
rect 5520 4356 5880 4360
rect 5520 4324 5524 4356
rect 5556 4324 5684 4356
rect 5716 4324 5844 4356
rect 5876 4324 5880 4356
rect 5520 4320 5880 4324
rect 5920 4356 6120 4360
rect 5920 4324 5924 4356
rect 5956 4324 6084 4356
rect 6116 4324 6120 4356
rect 5920 4320 6120 4324
rect 6160 4356 6360 4360
rect 6160 4324 6164 4356
rect 6196 4324 6324 4356
rect 6356 4324 6360 4356
rect 6160 4320 6360 4324
rect 4240 4276 4440 4280
rect 4240 4244 4244 4276
rect 4276 4244 4404 4276
rect 4436 4244 4440 4276
rect 4240 4240 4440 4244
rect 4480 4276 4680 4280
rect 4480 4244 4484 4276
rect 4516 4244 4644 4276
rect 4676 4244 4680 4276
rect 4480 4240 4680 4244
rect 4720 4276 5080 4280
rect 4720 4244 4724 4276
rect 4756 4244 4884 4276
rect 4916 4244 5044 4276
rect 5076 4244 5080 4276
rect 4720 4240 5080 4244
rect 5120 4276 5480 4280
rect 5120 4244 5124 4276
rect 5156 4244 5284 4276
rect 5316 4244 5444 4276
rect 5476 4244 5480 4276
rect 5120 4240 5480 4244
rect 5520 4276 5880 4280
rect 5520 4244 5524 4276
rect 5556 4244 5684 4276
rect 5716 4244 5844 4276
rect 5876 4244 5880 4276
rect 5520 4240 5880 4244
rect 5920 4276 6120 4280
rect 5920 4244 5924 4276
rect 5956 4244 6084 4276
rect 6116 4244 6120 4276
rect 5920 4240 6120 4244
rect 6160 4276 6360 4280
rect 6160 4244 6164 4276
rect 6196 4244 6324 4276
rect 6356 4244 6360 4276
rect 6160 4240 6360 4244
rect 4240 4196 4440 4200
rect 4240 4164 4244 4196
rect 4276 4164 4404 4196
rect 4436 4164 4440 4196
rect 4240 4160 4440 4164
rect 4480 4196 4680 4200
rect 4480 4164 4484 4196
rect 4516 4164 4644 4196
rect 4676 4164 4680 4196
rect 4480 4160 4680 4164
rect 4720 4196 5080 4200
rect 4720 4164 4724 4196
rect 4756 4164 4884 4196
rect 4916 4164 5044 4196
rect 5076 4164 5080 4196
rect 4720 4160 5080 4164
rect 5120 4196 5480 4200
rect 5120 4164 5124 4196
rect 5156 4164 5284 4196
rect 5316 4164 5444 4196
rect 5476 4164 5480 4196
rect 5120 4160 5480 4164
rect 5520 4196 5880 4200
rect 5520 4164 5524 4196
rect 5556 4164 5684 4196
rect 5716 4164 5844 4196
rect 5876 4164 5880 4196
rect 5520 4160 5880 4164
rect 5920 4196 6120 4200
rect 5920 4164 5924 4196
rect 5956 4164 6084 4196
rect 6116 4164 6120 4196
rect 5920 4160 6120 4164
rect 6160 4196 6360 4200
rect 6160 4164 6164 4196
rect 6196 4164 6324 4196
rect 6356 4164 6360 4196
rect 6160 4160 6360 4164
rect 4240 4116 4440 4120
rect 4240 4084 4244 4116
rect 4276 4084 4404 4116
rect 4436 4084 4440 4116
rect 4240 4080 4440 4084
rect 4480 4116 4680 4120
rect 4480 4084 4484 4116
rect 4516 4084 4644 4116
rect 4676 4084 4680 4116
rect 4480 4080 4680 4084
rect 4720 4116 5080 4120
rect 4720 4084 4724 4116
rect 4756 4084 4884 4116
rect 4916 4084 5044 4116
rect 5076 4084 5080 4116
rect 4720 4080 5080 4084
rect 5120 4116 5480 4120
rect 5120 4084 5124 4116
rect 5156 4084 5284 4116
rect 5316 4084 5444 4116
rect 5476 4084 5480 4116
rect 5120 4080 5480 4084
rect 5520 4116 5880 4120
rect 5520 4084 5524 4116
rect 5556 4084 5684 4116
rect 5716 4084 5844 4116
rect 5876 4084 5880 4116
rect 5520 4080 5880 4084
rect 5920 4116 6120 4120
rect 5920 4084 5924 4116
rect 5956 4084 6084 4116
rect 6116 4084 6120 4116
rect 5920 4080 6120 4084
rect 6160 4116 6360 4120
rect 6160 4084 6164 4116
rect 6196 4084 6324 4116
rect 6356 4084 6360 4116
rect 6160 4080 6360 4084
rect 4240 4036 4440 4040
rect 4240 4004 4244 4036
rect 4276 4004 4404 4036
rect 4436 4004 4440 4036
rect 4240 4000 4440 4004
rect 4480 4036 4680 4040
rect 4480 4004 4484 4036
rect 4516 4004 4644 4036
rect 4676 4004 4680 4036
rect 4480 4000 4680 4004
rect 4720 4036 5080 4040
rect 4720 4004 4724 4036
rect 4756 4004 4884 4036
rect 4916 4004 5044 4036
rect 5076 4004 5080 4036
rect 4720 4000 5080 4004
rect 5120 4036 5480 4040
rect 5120 4004 5124 4036
rect 5156 4004 5284 4036
rect 5316 4004 5444 4036
rect 5476 4004 5480 4036
rect 5120 4000 5480 4004
rect 5520 4036 5880 4040
rect 5520 4004 5524 4036
rect 5556 4004 5684 4036
rect 5716 4004 5844 4036
rect 5876 4004 5880 4036
rect 5520 4000 5880 4004
rect 5920 4036 6120 4040
rect 5920 4004 5924 4036
rect 5956 4004 6084 4036
rect 6116 4004 6120 4036
rect 5920 4000 6120 4004
rect 6160 4036 6360 4040
rect 6160 4004 6164 4036
rect 6196 4004 6324 4036
rect 6356 4004 6360 4036
rect 6160 4000 6360 4004
rect 4240 3956 4440 3960
rect 4240 3924 4244 3956
rect 4276 3924 4404 3956
rect 4436 3924 4440 3956
rect 4240 3920 4440 3924
rect 4480 3956 4680 3960
rect 4480 3924 4484 3956
rect 4516 3924 4644 3956
rect 4676 3924 4680 3956
rect 4480 3920 4680 3924
rect 4720 3956 5080 3960
rect 4720 3924 4724 3956
rect 4756 3924 4884 3956
rect 4916 3924 5044 3956
rect 5076 3924 5080 3956
rect 4720 3920 5080 3924
rect 5120 3956 5480 3960
rect 5120 3924 5124 3956
rect 5156 3924 5284 3956
rect 5316 3924 5444 3956
rect 5476 3924 5480 3956
rect 5120 3920 5480 3924
rect 5520 3956 5880 3960
rect 5520 3924 5524 3956
rect 5556 3924 5684 3956
rect 5716 3924 5844 3956
rect 5876 3924 5880 3956
rect 5520 3920 5880 3924
rect 5920 3956 6120 3960
rect 5920 3924 5924 3956
rect 5956 3924 6084 3956
rect 6116 3924 6120 3956
rect 5920 3920 6120 3924
rect 6160 3956 6360 3960
rect 6160 3924 6164 3956
rect 6196 3924 6324 3956
rect 6356 3924 6360 3956
rect 6160 3920 6360 3924
rect 4240 3156 4440 3160
rect 4240 3124 4244 3156
rect 4276 3124 4404 3156
rect 4436 3124 4440 3156
rect 4240 3120 4440 3124
rect 4480 3156 4680 3160
rect 4480 3124 4484 3156
rect 4516 3124 4644 3156
rect 4676 3124 4680 3156
rect 4480 3120 4680 3124
rect 4720 3156 5080 3160
rect 4720 3124 4724 3156
rect 4756 3124 4884 3156
rect 4916 3124 5044 3156
rect 5076 3124 5080 3156
rect 4720 3120 5080 3124
rect 5120 3156 5480 3160
rect 5120 3124 5124 3156
rect 5156 3124 5284 3156
rect 5316 3124 5444 3156
rect 5476 3124 5480 3156
rect 5120 3120 5480 3124
rect 5520 3156 5880 3160
rect 5520 3124 5524 3156
rect 5556 3124 5684 3156
rect 5716 3124 5844 3156
rect 5876 3124 5880 3156
rect 5520 3120 5880 3124
rect 5920 3156 6120 3160
rect 5920 3124 5924 3156
rect 5956 3124 6084 3156
rect 6116 3124 6120 3156
rect 5920 3120 6120 3124
rect 6160 3156 6360 3160
rect 6160 3124 6164 3156
rect 6196 3124 6324 3156
rect 6356 3124 6360 3156
rect 6160 3120 6360 3124
rect 4240 3076 4440 3080
rect 4240 3044 4244 3076
rect 4276 3044 4404 3076
rect 4436 3044 4440 3076
rect 4240 3040 4440 3044
rect 4480 3076 4680 3080
rect 4480 3044 4484 3076
rect 4516 3044 4644 3076
rect 4676 3044 4680 3076
rect 4480 3040 4680 3044
rect 4720 3076 5080 3080
rect 4720 3044 4724 3076
rect 4756 3044 4884 3076
rect 4916 3044 5044 3076
rect 5076 3044 5080 3076
rect 4720 3040 5080 3044
rect 5120 3076 5480 3080
rect 5120 3044 5124 3076
rect 5156 3044 5284 3076
rect 5316 3044 5444 3076
rect 5476 3044 5480 3076
rect 5120 3040 5480 3044
rect 5520 3076 5880 3080
rect 5520 3044 5524 3076
rect 5556 3044 5684 3076
rect 5716 3044 5844 3076
rect 5876 3044 5880 3076
rect 5520 3040 5880 3044
rect 5920 3076 6120 3080
rect 5920 3044 5924 3076
rect 5956 3044 6084 3076
rect 6116 3044 6120 3076
rect 5920 3040 6120 3044
rect 6160 3076 6360 3080
rect 6160 3044 6164 3076
rect 6196 3044 6324 3076
rect 6356 3044 6360 3076
rect 6160 3040 6360 3044
rect 4240 2996 4440 3000
rect 4240 2964 4244 2996
rect 4276 2964 4404 2996
rect 4436 2964 4440 2996
rect 4240 2960 4440 2964
rect 4480 2996 4680 3000
rect 4480 2964 4484 2996
rect 4516 2964 4644 2996
rect 4676 2964 4680 2996
rect 4480 2960 4680 2964
rect 4720 2996 5080 3000
rect 4720 2964 4724 2996
rect 4756 2964 4884 2996
rect 4916 2964 5044 2996
rect 5076 2964 5080 2996
rect 4720 2960 5080 2964
rect 5120 2996 5480 3000
rect 5120 2964 5124 2996
rect 5156 2964 5284 2996
rect 5316 2964 5444 2996
rect 5476 2964 5480 2996
rect 5120 2960 5480 2964
rect 5520 2996 5880 3000
rect 5520 2964 5524 2996
rect 5556 2964 5684 2996
rect 5716 2964 5844 2996
rect 5876 2964 5880 2996
rect 5520 2960 5880 2964
rect 5920 2996 6120 3000
rect 5920 2964 5924 2996
rect 5956 2964 6084 2996
rect 6116 2964 6120 2996
rect 5920 2960 6120 2964
rect 6160 2996 6360 3000
rect 6160 2964 6164 2996
rect 6196 2964 6324 2996
rect 6356 2964 6360 2996
rect 6160 2960 6360 2964
rect 4240 2916 4440 2920
rect 4240 2884 4244 2916
rect 4276 2884 4404 2916
rect 4436 2884 4440 2916
rect 4240 2880 4440 2884
rect 4480 2916 4680 2920
rect 4480 2884 4484 2916
rect 4516 2884 4644 2916
rect 4676 2884 4680 2916
rect 4480 2880 4680 2884
rect 4720 2916 5080 2920
rect 4720 2884 4724 2916
rect 4756 2884 4884 2916
rect 4916 2884 5044 2916
rect 5076 2884 5080 2916
rect 4720 2880 5080 2884
rect 5120 2916 5480 2920
rect 5120 2884 5124 2916
rect 5156 2884 5284 2916
rect 5316 2884 5444 2916
rect 5476 2884 5480 2916
rect 5120 2880 5480 2884
rect 5520 2916 5880 2920
rect 5520 2884 5524 2916
rect 5556 2884 5684 2916
rect 5716 2884 5844 2916
rect 5876 2884 5880 2916
rect 5520 2880 5880 2884
rect 5920 2916 6120 2920
rect 5920 2884 5924 2916
rect 5956 2884 6084 2916
rect 6116 2884 6120 2916
rect 5920 2880 6120 2884
rect 6160 2916 6360 2920
rect 6160 2884 6164 2916
rect 6196 2884 6324 2916
rect 6356 2884 6360 2916
rect 6160 2880 6360 2884
rect 4240 2836 4440 2840
rect 4240 2804 4244 2836
rect 4276 2804 4404 2836
rect 4436 2804 4440 2836
rect 4240 2800 4440 2804
rect 4480 2836 4680 2840
rect 4480 2804 4484 2836
rect 4516 2804 4644 2836
rect 4676 2804 4680 2836
rect 4480 2800 4680 2804
rect 4720 2836 5080 2840
rect 4720 2804 4724 2836
rect 4756 2804 4884 2836
rect 4916 2804 5044 2836
rect 5076 2804 5080 2836
rect 4720 2800 5080 2804
rect 5120 2836 5480 2840
rect 5120 2804 5124 2836
rect 5156 2804 5284 2836
rect 5316 2804 5444 2836
rect 5476 2804 5480 2836
rect 5120 2800 5480 2804
rect 5520 2836 5880 2840
rect 5520 2804 5524 2836
rect 5556 2804 5684 2836
rect 5716 2804 5844 2836
rect 5876 2804 5880 2836
rect 5520 2800 5880 2804
rect 5920 2836 6120 2840
rect 5920 2804 5924 2836
rect 5956 2804 6084 2836
rect 6116 2804 6120 2836
rect 5920 2800 6120 2804
rect 6160 2836 6360 2840
rect 6160 2804 6164 2836
rect 6196 2804 6324 2836
rect 6356 2804 6360 2836
rect 6160 2800 6360 2804
rect 4240 2756 4440 2760
rect 4240 2724 4244 2756
rect 4276 2724 4404 2756
rect 4436 2724 4440 2756
rect 4240 2720 4440 2724
rect 4480 2756 4680 2760
rect 4480 2724 4484 2756
rect 4516 2724 4644 2756
rect 4676 2724 4680 2756
rect 4480 2720 4680 2724
rect 4720 2756 5080 2760
rect 4720 2724 4724 2756
rect 4756 2724 4884 2756
rect 4916 2724 5044 2756
rect 5076 2724 5080 2756
rect 4720 2720 5080 2724
rect 5120 2756 5480 2760
rect 5120 2724 5124 2756
rect 5156 2724 5284 2756
rect 5316 2724 5444 2756
rect 5476 2724 5480 2756
rect 5120 2720 5480 2724
rect 5520 2756 5880 2760
rect 5520 2724 5524 2756
rect 5556 2724 5684 2756
rect 5716 2724 5844 2756
rect 5876 2724 5880 2756
rect 5520 2720 5880 2724
rect 5920 2756 6120 2760
rect 5920 2724 5924 2756
rect 5956 2724 6084 2756
rect 6116 2724 6120 2756
rect 5920 2720 6120 2724
rect 6160 2756 6360 2760
rect 6160 2724 6164 2756
rect 6196 2724 6324 2756
rect 6356 2724 6360 2756
rect 6160 2720 6360 2724
rect 4240 2676 4440 2680
rect 4240 2644 4244 2676
rect 4276 2644 4404 2676
rect 4436 2644 4440 2676
rect 4240 2640 4440 2644
rect 4480 2676 4680 2680
rect 4480 2644 4484 2676
rect 4516 2644 4644 2676
rect 4676 2644 4680 2676
rect 4480 2640 4680 2644
rect 4720 2676 5080 2680
rect 4720 2644 4724 2676
rect 4756 2644 4884 2676
rect 4916 2644 5044 2676
rect 5076 2644 5080 2676
rect 4720 2640 5080 2644
rect 5120 2676 5480 2680
rect 5120 2644 5124 2676
rect 5156 2644 5284 2676
rect 5316 2644 5444 2676
rect 5476 2644 5480 2676
rect 5120 2640 5480 2644
rect 5520 2676 5880 2680
rect 5520 2644 5524 2676
rect 5556 2644 5684 2676
rect 5716 2644 5844 2676
rect 5876 2644 5880 2676
rect 5520 2640 5880 2644
rect 5920 2676 6120 2680
rect 5920 2644 5924 2676
rect 5956 2644 6084 2676
rect 6116 2644 6120 2676
rect 5920 2640 6120 2644
rect 6160 2676 6360 2680
rect 6160 2644 6164 2676
rect 6196 2644 6324 2676
rect 6356 2644 6360 2676
rect 6160 2640 6360 2644
rect 4240 2596 4440 2600
rect 4240 2564 4244 2596
rect 4276 2564 4404 2596
rect 4436 2564 4440 2596
rect 4240 2560 4440 2564
rect 4480 2596 4680 2600
rect 4480 2564 4484 2596
rect 4516 2564 4644 2596
rect 4676 2564 4680 2596
rect 4480 2560 4680 2564
rect 4720 2596 5080 2600
rect 4720 2564 4724 2596
rect 4756 2564 4884 2596
rect 4916 2564 5044 2596
rect 5076 2564 5080 2596
rect 4720 2560 5080 2564
rect 5120 2596 5480 2600
rect 5120 2564 5124 2596
rect 5156 2564 5284 2596
rect 5316 2564 5444 2596
rect 5476 2564 5480 2596
rect 5120 2560 5480 2564
rect 5520 2596 5880 2600
rect 5520 2564 5524 2596
rect 5556 2564 5684 2596
rect 5716 2564 5844 2596
rect 5876 2564 5880 2596
rect 5520 2560 5880 2564
rect 5920 2596 6120 2600
rect 5920 2564 5924 2596
rect 5956 2564 6084 2596
rect 6116 2564 6120 2596
rect 5920 2560 6120 2564
rect 6160 2596 6360 2600
rect 6160 2564 6164 2596
rect 6196 2564 6324 2596
rect 6356 2564 6360 2596
rect 6160 2560 6360 2564
rect 4240 2516 4440 2520
rect 4240 2484 4244 2516
rect 4276 2484 4404 2516
rect 4436 2484 4440 2516
rect 4240 2480 4440 2484
rect 4480 2516 4680 2520
rect 4480 2484 4484 2516
rect 4516 2484 4644 2516
rect 4676 2484 4680 2516
rect 4480 2480 4680 2484
rect 4720 2516 5080 2520
rect 4720 2484 4724 2516
rect 4756 2484 4884 2516
rect 4916 2484 5044 2516
rect 5076 2484 5080 2516
rect 4720 2480 5080 2484
rect 5120 2516 5480 2520
rect 5120 2484 5124 2516
rect 5156 2484 5284 2516
rect 5316 2484 5444 2516
rect 5476 2484 5480 2516
rect 5120 2480 5480 2484
rect 5520 2516 5880 2520
rect 5520 2484 5524 2516
rect 5556 2484 5684 2516
rect 5716 2484 5844 2516
rect 5876 2484 5880 2516
rect 5520 2480 5880 2484
rect 5920 2516 6120 2520
rect 5920 2484 5924 2516
rect 5956 2484 6084 2516
rect 6116 2484 6120 2516
rect 5920 2480 6120 2484
rect 6160 2516 6360 2520
rect 6160 2484 6164 2516
rect 6196 2484 6324 2516
rect 6356 2484 6360 2516
rect 6160 2480 6360 2484
rect 4240 2436 4440 2440
rect 4240 2404 4244 2436
rect 4276 2404 4404 2436
rect 4436 2404 4440 2436
rect 4240 2400 4440 2404
rect 4480 2436 4680 2440
rect 4480 2404 4484 2436
rect 4516 2404 4644 2436
rect 4676 2404 4680 2436
rect 4480 2400 4680 2404
rect 4720 2436 5080 2440
rect 4720 2404 4724 2436
rect 4756 2404 4884 2436
rect 4916 2404 5044 2436
rect 5076 2404 5080 2436
rect 4720 2400 5080 2404
rect 5120 2436 5480 2440
rect 5120 2404 5124 2436
rect 5156 2404 5284 2436
rect 5316 2404 5444 2436
rect 5476 2404 5480 2436
rect 5120 2400 5480 2404
rect 5520 2436 5880 2440
rect 5520 2404 5524 2436
rect 5556 2404 5684 2436
rect 5716 2404 5844 2436
rect 5876 2404 5880 2436
rect 5520 2400 5880 2404
rect 5920 2436 6120 2440
rect 5920 2404 5924 2436
rect 5956 2404 6084 2436
rect 6116 2404 6120 2436
rect 5920 2400 6120 2404
rect 6160 2436 6360 2440
rect 6160 2404 6164 2436
rect 6196 2404 6324 2436
rect 6356 2404 6360 2436
rect 6160 2400 6360 2404
rect 4240 2356 4440 2360
rect 4240 2324 4244 2356
rect 4276 2324 4404 2356
rect 4436 2324 4440 2356
rect 4240 2320 4440 2324
rect 4480 2356 4680 2360
rect 4480 2324 4484 2356
rect 4516 2324 4644 2356
rect 4676 2324 4680 2356
rect 4480 2320 4680 2324
rect 4720 2356 5080 2360
rect 4720 2324 4724 2356
rect 4756 2324 4884 2356
rect 4916 2324 5044 2356
rect 5076 2324 5080 2356
rect 4720 2320 5080 2324
rect 5120 2356 5480 2360
rect 5120 2324 5124 2356
rect 5156 2324 5284 2356
rect 5316 2324 5444 2356
rect 5476 2324 5480 2356
rect 5120 2320 5480 2324
rect 5520 2356 5880 2360
rect 5520 2324 5524 2356
rect 5556 2324 5684 2356
rect 5716 2324 5844 2356
rect 5876 2324 5880 2356
rect 5520 2320 5880 2324
rect 5920 2356 6120 2360
rect 5920 2324 5924 2356
rect 5956 2324 6084 2356
rect 6116 2324 6120 2356
rect 5920 2320 6120 2324
rect 6160 2356 6360 2360
rect 6160 2324 6164 2356
rect 6196 2324 6324 2356
rect 6356 2324 6360 2356
rect 6160 2320 6360 2324
rect 4240 2276 4440 2280
rect 4240 2244 4244 2276
rect 4276 2244 4404 2276
rect 4436 2244 4440 2276
rect 4240 2240 4440 2244
rect 4480 2276 4680 2280
rect 4480 2244 4484 2276
rect 4516 2244 4644 2276
rect 4676 2244 4680 2276
rect 4480 2240 4680 2244
rect 4720 2276 5080 2280
rect 4720 2244 4724 2276
rect 4756 2244 4884 2276
rect 4916 2244 5044 2276
rect 5076 2244 5080 2276
rect 4720 2240 5080 2244
rect 5120 2276 5480 2280
rect 5120 2244 5124 2276
rect 5156 2244 5284 2276
rect 5316 2244 5444 2276
rect 5476 2244 5480 2276
rect 5120 2240 5480 2244
rect 5520 2276 5880 2280
rect 5520 2244 5524 2276
rect 5556 2244 5684 2276
rect 5716 2244 5844 2276
rect 5876 2244 5880 2276
rect 5520 2240 5880 2244
rect 5920 2276 6120 2280
rect 5920 2244 5924 2276
rect 5956 2244 6084 2276
rect 6116 2244 6120 2276
rect 5920 2240 6120 2244
rect 6160 2276 6360 2280
rect 6160 2244 6164 2276
rect 6196 2244 6324 2276
rect 6356 2244 6360 2276
rect 6160 2240 6360 2244
rect 4240 2196 4440 2200
rect 4240 2164 4244 2196
rect 4276 2164 4404 2196
rect 4436 2164 4440 2196
rect 4240 2160 4440 2164
rect 4480 2196 4680 2200
rect 4480 2164 4484 2196
rect 4516 2164 4644 2196
rect 4676 2164 4680 2196
rect 4480 2160 4680 2164
rect 4720 2196 5080 2200
rect 4720 2164 4724 2196
rect 4756 2164 4884 2196
rect 4916 2164 5044 2196
rect 5076 2164 5080 2196
rect 4720 2160 5080 2164
rect 5120 2196 5480 2200
rect 5120 2164 5124 2196
rect 5156 2164 5284 2196
rect 5316 2164 5444 2196
rect 5476 2164 5480 2196
rect 5120 2160 5480 2164
rect 5520 2196 5880 2200
rect 5520 2164 5524 2196
rect 5556 2164 5684 2196
rect 5716 2164 5844 2196
rect 5876 2164 5880 2196
rect 5520 2160 5880 2164
rect 5920 2196 6120 2200
rect 5920 2164 5924 2196
rect 5956 2164 6084 2196
rect 6116 2164 6120 2196
rect 5920 2160 6120 2164
rect 6160 2196 6360 2200
rect 6160 2164 6164 2196
rect 6196 2164 6324 2196
rect 6356 2164 6360 2196
rect 6160 2160 6360 2164
rect 4240 2116 4440 2120
rect 4240 2084 4244 2116
rect 4276 2084 4404 2116
rect 4436 2084 4440 2116
rect 4240 2080 4440 2084
rect 4480 2116 4680 2120
rect 4480 2084 4484 2116
rect 4516 2084 4644 2116
rect 4676 2084 4680 2116
rect 4480 2080 4680 2084
rect 4720 2116 5080 2120
rect 4720 2084 4724 2116
rect 4756 2084 4884 2116
rect 4916 2084 5044 2116
rect 5076 2084 5080 2116
rect 4720 2080 5080 2084
rect 5120 2116 5480 2120
rect 5120 2084 5124 2116
rect 5156 2084 5284 2116
rect 5316 2084 5444 2116
rect 5476 2084 5480 2116
rect 5120 2080 5480 2084
rect 5520 2116 5880 2120
rect 5520 2084 5524 2116
rect 5556 2084 5684 2116
rect 5716 2084 5844 2116
rect 5876 2084 5880 2116
rect 5520 2080 5880 2084
rect 5920 2116 6120 2120
rect 5920 2084 5924 2116
rect 5956 2084 6084 2116
rect 6116 2084 6120 2116
rect 5920 2080 6120 2084
rect 6160 2116 6360 2120
rect 6160 2084 6164 2116
rect 6196 2084 6324 2116
rect 6356 2084 6360 2116
rect 6160 2080 6360 2084
rect 4240 2036 4440 2040
rect 4240 2004 4244 2036
rect 4276 2004 4404 2036
rect 4436 2004 4440 2036
rect 4240 2000 4440 2004
rect 4480 2036 4680 2040
rect 4480 2004 4484 2036
rect 4516 2004 4644 2036
rect 4676 2004 4680 2036
rect 4480 2000 4680 2004
rect 4720 2036 5080 2040
rect 4720 2004 4724 2036
rect 4756 2004 4884 2036
rect 4916 2004 5044 2036
rect 5076 2004 5080 2036
rect 4720 2000 5080 2004
rect 5120 2036 5480 2040
rect 5120 2004 5124 2036
rect 5156 2004 5284 2036
rect 5316 2004 5444 2036
rect 5476 2004 5480 2036
rect 5120 2000 5480 2004
rect 5520 2036 5880 2040
rect 5520 2004 5524 2036
rect 5556 2004 5684 2036
rect 5716 2004 5844 2036
rect 5876 2004 5880 2036
rect 5520 2000 5880 2004
rect 5920 2036 6120 2040
rect 5920 2004 5924 2036
rect 5956 2004 6084 2036
rect 6116 2004 6120 2036
rect 5920 2000 6120 2004
rect 6160 2036 6360 2040
rect 6160 2004 6164 2036
rect 6196 2004 6324 2036
rect 6356 2004 6360 2036
rect 6160 2000 6360 2004
rect 4240 1636 4440 1640
rect 4240 1604 4244 1636
rect 4276 1604 4404 1636
rect 4436 1604 4440 1636
rect 4240 1600 4440 1604
rect 4480 1636 4680 1640
rect 4480 1604 4484 1636
rect 4516 1604 4644 1636
rect 4676 1604 4680 1636
rect 4480 1600 4680 1604
rect 4720 1636 5080 1640
rect 4720 1604 4724 1636
rect 4756 1604 4884 1636
rect 4916 1604 5044 1636
rect 5076 1604 5080 1636
rect 4720 1600 5080 1604
rect 5120 1636 5480 1640
rect 5120 1604 5124 1636
rect 5156 1604 5284 1636
rect 5316 1604 5444 1636
rect 5476 1604 5480 1636
rect 5120 1600 5480 1604
rect 5520 1636 5880 1640
rect 5520 1604 5524 1636
rect 5556 1604 5684 1636
rect 5716 1604 5844 1636
rect 5876 1604 5880 1636
rect 5520 1600 5880 1604
rect 5920 1636 6120 1640
rect 5920 1604 5924 1636
rect 5956 1604 6084 1636
rect 6116 1604 6120 1636
rect 5920 1600 6120 1604
rect 6160 1636 6360 1640
rect 6160 1604 6164 1636
rect 6196 1604 6324 1636
rect 6356 1604 6360 1636
rect 6160 1600 6360 1604
rect 4240 1556 4440 1560
rect 4240 1524 4244 1556
rect 4276 1524 4404 1556
rect 4436 1524 4440 1556
rect 4240 1520 4440 1524
rect 4480 1556 4680 1560
rect 4480 1524 4484 1556
rect 4516 1524 4644 1556
rect 4676 1524 4680 1556
rect 4480 1520 4680 1524
rect 4720 1556 5080 1560
rect 4720 1524 4724 1556
rect 4756 1524 4884 1556
rect 4916 1524 5044 1556
rect 5076 1524 5080 1556
rect 4720 1520 5080 1524
rect 5120 1556 5480 1560
rect 5120 1524 5124 1556
rect 5156 1524 5284 1556
rect 5316 1524 5444 1556
rect 5476 1524 5480 1556
rect 5120 1520 5480 1524
rect 5520 1556 5880 1560
rect 5520 1524 5524 1556
rect 5556 1524 5684 1556
rect 5716 1524 5844 1556
rect 5876 1524 5880 1556
rect 5520 1520 5880 1524
rect 5920 1556 6120 1560
rect 5920 1524 5924 1556
rect 5956 1524 6084 1556
rect 6116 1524 6120 1556
rect 5920 1520 6120 1524
rect 6160 1556 6360 1560
rect 6160 1524 6164 1556
rect 6196 1524 6324 1556
rect 6356 1524 6360 1556
rect 6160 1520 6360 1524
rect 4240 1476 4440 1480
rect 4240 1444 4244 1476
rect 4276 1444 4404 1476
rect 4436 1444 4440 1476
rect 4240 1440 4440 1444
rect 4480 1476 4680 1480
rect 4480 1444 4484 1476
rect 4516 1444 4644 1476
rect 4676 1444 4680 1476
rect 4480 1440 4680 1444
rect 4720 1476 5080 1480
rect 4720 1444 4724 1476
rect 4756 1444 4884 1476
rect 4916 1444 5044 1476
rect 5076 1444 5080 1476
rect 4720 1440 5080 1444
rect 5120 1476 5480 1480
rect 5120 1444 5124 1476
rect 5156 1444 5284 1476
rect 5316 1444 5444 1476
rect 5476 1444 5480 1476
rect 5120 1440 5480 1444
rect 5520 1476 5880 1480
rect 5520 1444 5524 1476
rect 5556 1444 5684 1476
rect 5716 1444 5844 1476
rect 5876 1444 5880 1476
rect 5520 1440 5880 1444
rect 5920 1476 6120 1480
rect 5920 1444 5924 1476
rect 5956 1444 6084 1476
rect 6116 1444 6120 1476
rect 5920 1440 6120 1444
rect 6160 1476 6360 1480
rect 6160 1444 6164 1476
rect 6196 1444 6324 1476
rect 6356 1444 6360 1476
rect 6160 1440 6360 1444
rect 4240 1396 4440 1400
rect 4240 1364 4244 1396
rect 4276 1364 4404 1396
rect 4436 1364 4440 1396
rect 4240 1360 4440 1364
rect 4480 1396 4680 1400
rect 4480 1364 4484 1396
rect 4516 1364 4644 1396
rect 4676 1364 4680 1396
rect 4480 1360 4680 1364
rect 4720 1396 5080 1400
rect 4720 1364 4724 1396
rect 4756 1364 4884 1396
rect 4916 1364 5044 1396
rect 5076 1364 5080 1396
rect 4720 1360 5080 1364
rect 5120 1396 5480 1400
rect 5120 1364 5124 1396
rect 5156 1364 5284 1396
rect 5316 1364 5444 1396
rect 5476 1364 5480 1396
rect 5120 1360 5480 1364
rect 5520 1396 5880 1400
rect 5520 1364 5524 1396
rect 5556 1364 5684 1396
rect 5716 1364 5844 1396
rect 5876 1364 5880 1396
rect 5520 1360 5880 1364
rect 5920 1396 6120 1400
rect 5920 1364 5924 1396
rect 5956 1364 6084 1396
rect 6116 1364 6120 1396
rect 5920 1360 6120 1364
rect 6160 1396 6360 1400
rect 6160 1364 6164 1396
rect 6196 1364 6324 1396
rect 6356 1364 6360 1396
rect 6160 1360 6360 1364
rect 4240 1316 4440 1320
rect 4240 1284 4244 1316
rect 4276 1284 4404 1316
rect 4436 1284 4440 1316
rect 4240 1280 4440 1284
rect 4480 1316 4680 1320
rect 4480 1284 4484 1316
rect 4516 1284 4644 1316
rect 4676 1284 4680 1316
rect 4480 1280 4680 1284
rect 4720 1316 5080 1320
rect 4720 1284 4724 1316
rect 4756 1284 4884 1316
rect 4916 1284 5044 1316
rect 5076 1284 5080 1316
rect 4720 1280 5080 1284
rect 5120 1316 5480 1320
rect 5120 1284 5124 1316
rect 5156 1284 5284 1316
rect 5316 1284 5444 1316
rect 5476 1284 5480 1316
rect 5120 1280 5480 1284
rect 5520 1316 5880 1320
rect 5520 1284 5524 1316
rect 5556 1284 5684 1316
rect 5716 1284 5844 1316
rect 5876 1284 5880 1316
rect 5520 1280 5880 1284
rect 5920 1316 6120 1320
rect 5920 1284 5924 1316
rect 5956 1284 6084 1316
rect 6116 1284 6120 1316
rect 5920 1280 6120 1284
rect 6160 1316 6360 1320
rect 6160 1284 6164 1316
rect 6196 1284 6324 1316
rect 6356 1284 6360 1316
rect 6160 1280 6360 1284
rect 4240 1236 4440 1240
rect 4240 1204 4244 1236
rect 4276 1204 4404 1236
rect 4436 1204 4440 1236
rect 4240 1200 4440 1204
rect 4480 1236 4680 1240
rect 4480 1204 4484 1236
rect 4516 1204 4644 1236
rect 4676 1204 4680 1236
rect 4480 1200 4680 1204
rect 4720 1236 5080 1240
rect 4720 1204 4724 1236
rect 4756 1204 4884 1236
rect 4916 1204 5044 1236
rect 5076 1204 5080 1236
rect 4720 1200 5080 1204
rect 5120 1236 5480 1240
rect 5120 1204 5124 1236
rect 5156 1204 5284 1236
rect 5316 1204 5444 1236
rect 5476 1204 5480 1236
rect 5120 1200 5480 1204
rect 5520 1236 5880 1240
rect 5520 1204 5524 1236
rect 5556 1204 5684 1236
rect 5716 1204 5844 1236
rect 5876 1204 5880 1236
rect 5520 1200 5880 1204
rect 5920 1236 6120 1240
rect 5920 1204 5924 1236
rect 5956 1204 6084 1236
rect 6116 1204 6120 1236
rect 5920 1200 6120 1204
rect 6160 1236 6360 1240
rect 6160 1204 6164 1236
rect 6196 1204 6324 1236
rect 6356 1204 6360 1236
rect 6160 1200 6360 1204
rect 4240 1156 4440 1160
rect 4240 1124 4244 1156
rect 4276 1124 4404 1156
rect 4436 1124 4440 1156
rect 4240 1120 4440 1124
rect 4480 1156 4680 1160
rect 4480 1124 4484 1156
rect 4516 1124 4644 1156
rect 4676 1124 4680 1156
rect 4480 1120 4680 1124
rect 4720 1156 5080 1160
rect 4720 1124 4724 1156
rect 4756 1124 4884 1156
rect 4916 1124 5044 1156
rect 5076 1124 5080 1156
rect 4720 1120 5080 1124
rect 5120 1156 5480 1160
rect 5120 1124 5124 1156
rect 5156 1124 5284 1156
rect 5316 1124 5444 1156
rect 5476 1124 5480 1156
rect 5120 1120 5480 1124
rect 5520 1156 5880 1160
rect 5520 1124 5524 1156
rect 5556 1124 5684 1156
rect 5716 1124 5844 1156
rect 5876 1124 5880 1156
rect 5520 1120 5880 1124
rect 5920 1156 6120 1160
rect 5920 1124 5924 1156
rect 5956 1124 6084 1156
rect 6116 1124 6120 1156
rect 5920 1120 6120 1124
rect 6160 1156 6360 1160
rect 6160 1124 6164 1156
rect 6196 1124 6324 1156
rect 6356 1124 6360 1156
rect 6160 1120 6360 1124
rect 4240 1076 4440 1080
rect 4240 1044 4244 1076
rect 4276 1044 4404 1076
rect 4436 1044 4440 1076
rect 4240 1040 4440 1044
rect 4480 1076 4680 1080
rect 4480 1044 4484 1076
rect 4516 1044 4644 1076
rect 4676 1044 4680 1076
rect 4480 1040 4680 1044
rect 4720 1076 5080 1080
rect 4720 1044 4724 1076
rect 4756 1044 4884 1076
rect 4916 1044 5044 1076
rect 5076 1044 5080 1076
rect 4720 1040 5080 1044
rect 5120 1076 5480 1080
rect 5120 1044 5124 1076
rect 5156 1044 5284 1076
rect 5316 1044 5444 1076
rect 5476 1044 5480 1076
rect 5120 1040 5480 1044
rect 5520 1076 5880 1080
rect 5520 1044 5524 1076
rect 5556 1044 5684 1076
rect 5716 1044 5844 1076
rect 5876 1044 5880 1076
rect 5520 1040 5880 1044
rect 5920 1076 6120 1080
rect 5920 1044 5924 1076
rect 5956 1044 6084 1076
rect 6116 1044 6120 1076
rect 5920 1040 6120 1044
rect 6160 1076 6360 1080
rect 6160 1044 6164 1076
rect 6196 1044 6324 1076
rect 6356 1044 6360 1076
rect 6160 1040 6360 1044
rect 4240 756 4440 760
rect 4240 724 4244 756
rect 4276 724 4404 756
rect 4436 724 4440 756
rect 4240 720 4440 724
rect 4480 756 4680 760
rect 4480 724 4484 756
rect 4516 724 4644 756
rect 4676 724 4680 756
rect 4480 720 4680 724
rect 4720 756 5080 760
rect 4720 724 4724 756
rect 4756 724 4884 756
rect 4916 724 5044 756
rect 5076 724 5080 756
rect 4720 720 5080 724
rect 5120 756 5480 760
rect 5120 724 5124 756
rect 5156 724 5284 756
rect 5316 724 5444 756
rect 5476 724 5480 756
rect 5120 720 5480 724
rect 5520 756 5880 760
rect 5520 724 5524 756
rect 5556 724 5684 756
rect 5716 724 5844 756
rect 5876 724 5880 756
rect 5520 720 5880 724
rect 5920 756 6120 760
rect 5920 724 5924 756
rect 5956 724 6084 756
rect 6116 724 6120 756
rect 5920 720 6120 724
rect 6160 756 6360 760
rect 6160 724 6164 756
rect 6196 724 6324 756
rect 6356 724 6360 756
rect 6160 720 6360 724
rect 4240 676 4440 680
rect 4240 644 4244 676
rect 4276 644 4404 676
rect 4436 644 4440 676
rect 4240 640 4440 644
rect 4480 676 4680 680
rect 4480 644 4484 676
rect 4516 644 4644 676
rect 4676 644 4680 676
rect 4480 640 4680 644
rect 4720 676 5080 680
rect 4720 644 4724 676
rect 4756 644 4884 676
rect 4916 644 5044 676
rect 5076 644 5080 676
rect 4720 640 5080 644
rect 5120 676 5480 680
rect 5120 644 5124 676
rect 5156 644 5284 676
rect 5316 644 5444 676
rect 5476 644 5480 676
rect 5120 640 5480 644
rect 5520 676 5880 680
rect 5520 644 5524 676
rect 5556 644 5684 676
rect 5716 644 5844 676
rect 5876 644 5880 676
rect 5520 640 5880 644
rect 5920 676 6120 680
rect 5920 644 5924 676
rect 5956 644 6084 676
rect 6116 644 6120 676
rect 5920 640 6120 644
rect 6160 676 6360 680
rect 6160 644 6164 676
rect 6196 644 6324 676
rect 6356 644 6360 676
rect 6160 640 6360 644
rect 4240 596 4440 600
rect 4240 564 4244 596
rect 4276 564 4404 596
rect 4436 564 4440 596
rect 4240 560 4440 564
rect 4480 596 4680 600
rect 4480 564 4484 596
rect 4516 564 4644 596
rect 4676 564 4680 596
rect 4480 560 4680 564
rect 4720 596 5080 600
rect 4720 564 4724 596
rect 4756 564 4884 596
rect 4916 564 5044 596
rect 5076 564 5080 596
rect 4720 560 5080 564
rect 5120 596 5480 600
rect 5120 564 5124 596
rect 5156 564 5284 596
rect 5316 564 5444 596
rect 5476 564 5480 596
rect 5120 560 5480 564
rect 5520 596 5880 600
rect 5520 564 5524 596
rect 5556 564 5684 596
rect 5716 564 5844 596
rect 5876 564 5880 596
rect 5520 560 5880 564
rect 5920 596 6120 600
rect 5920 564 5924 596
rect 5956 564 6084 596
rect 6116 564 6120 596
rect 5920 560 6120 564
rect 6160 596 6360 600
rect 6160 564 6164 596
rect 6196 564 6324 596
rect 6356 564 6360 596
rect 6160 560 6360 564
rect 4240 196 4440 200
rect 4240 164 4244 196
rect 4276 164 4404 196
rect 4436 164 4440 196
rect 4240 160 4440 164
rect 4480 196 4680 200
rect 4480 164 4484 196
rect 4516 164 4644 196
rect 4676 164 4680 196
rect 4480 160 4680 164
rect 4720 196 5080 200
rect 4720 164 4724 196
rect 4756 164 4884 196
rect 4916 164 5044 196
rect 5076 164 5080 196
rect 4720 160 5080 164
rect 5120 196 5480 200
rect 5120 164 5124 196
rect 5156 164 5284 196
rect 5316 164 5444 196
rect 5476 164 5480 196
rect 5120 160 5480 164
rect 5520 196 5880 200
rect 5520 164 5524 196
rect 5556 164 5684 196
rect 5716 164 5844 196
rect 5876 164 5880 196
rect 5520 160 5880 164
rect 5920 196 6120 200
rect 5920 164 5924 196
rect 5956 164 6084 196
rect 6116 164 6120 196
rect 5920 160 6120 164
rect 6160 196 6360 200
rect 6160 164 6164 196
rect 6196 164 6324 196
rect 6356 164 6360 196
rect 6160 160 6360 164
rect 4240 116 4440 120
rect 4240 84 4244 116
rect 4276 84 4404 116
rect 4436 84 4440 116
rect 4240 80 4440 84
rect 4480 116 4680 120
rect 4480 84 4484 116
rect 4516 84 4644 116
rect 4676 84 4680 116
rect 4480 80 4680 84
rect 4720 116 5080 120
rect 4720 84 4724 116
rect 4756 84 4884 116
rect 4916 84 5044 116
rect 5076 84 5080 116
rect 4720 80 5080 84
rect 5120 116 5480 120
rect 5120 84 5124 116
rect 5156 84 5284 116
rect 5316 84 5444 116
rect 5476 84 5480 116
rect 5120 80 5480 84
rect 5520 116 5880 120
rect 5520 84 5524 116
rect 5556 84 5684 116
rect 5716 84 5844 116
rect 5876 84 5880 116
rect 5520 80 5880 84
rect 5920 116 6120 120
rect 5920 84 5924 116
rect 5956 84 6084 116
rect 6116 84 6120 116
rect 5920 80 6120 84
rect 6160 116 6360 120
rect 6160 84 6164 116
rect 6196 84 6324 116
rect 6356 84 6360 116
rect 6160 80 6360 84
rect 4240 36 4440 40
rect 4240 4 4244 36
rect 4276 4 4404 36
rect 4436 4 4440 36
rect 4240 0 4440 4
rect 4480 36 4680 40
rect 4480 4 4484 36
rect 4516 4 4644 36
rect 4676 4 4680 36
rect 4480 0 4680 4
rect 4720 36 5080 40
rect 4720 4 4724 36
rect 4756 4 4884 36
rect 4916 4 5044 36
rect 5076 4 5080 36
rect 4720 0 5080 4
rect 5120 36 5480 40
rect 5120 4 5124 36
rect 5156 4 5284 36
rect 5316 4 5444 36
rect 5476 4 5480 36
rect 5120 0 5480 4
rect 5520 36 5880 40
rect 5520 4 5524 36
rect 5556 4 5684 36
rect 5716 4 5844 36
rect 5876 4 5880 36
rect 5520 0 5880 4
rect 5920 36 6120 40
rect 5920 4 5924 36
rect 5956 4 6084 36
rect 6116 4 6120 36
rect 5920 0 6120 4
rect 6160 36 6360 40
rect 6160 4 6164 36
rect 6196 4 6324 36
rect 6356 4 6360 36
rect 6160 0 6360 4
<< via4 >>
rect 1561 13481 1679 13599
rect 2521 13481 2639 13599
rect 7961 13481 8079 13599
rect 8921 13481 9039 13599
rect 1081 13241 1199 13359
rect 2041 13241 2159 13359
rect 3001 13241 3119 13359
rect 7481 13241 7599 13359
rect 8441 13241 8559 13359
rect 9401 13241 9519 13359
rect 601 13001 719 13119
rect 3481 13001 3599 13119
rect 7001 13001 7119 13119
rect 9881 13001 9999 13119
rect 121 12761 239 12879
rect 3961 12761 4079 12879
rect 6521 12761 6639 12879
rect 10361 12761 10479 12879
<< metal5 >>
rect 80 12879 280 13640
rect 80 12761 121 12879
rect 239 12761 280 12879
rect 80 12680 280 12761
rect 560 13119 760 13640
rect 560 13001 601 13119
rect 719 13001 760 13119
rect 560 12680 760 13001
rect 1040 13359 1240 13640
rect 1040 13241 1081 13359
rect 1199 13241 1240 13359
rect 1040 12680 1240 13241
rect 1520 13599 1720 13640
rect 1520 13481 1561 13599
rect 1679 13481 1720 13599
rect 1520 12680 1720 13481
rect 2000 13359 2200 13640
rect 2000 13241 2041 13359
rect 2159 13241 2200 13359
rect 2000 12680 2200 13241
rect 2480 13599 2680 13640
rect 2480 13481 2521 13599
rect 2639 13481 2680 13599
rect 2480 12680 2680 13481
rect 2960 13359 3160 13640
rect 2960 13241 3001 13359
rect 3119 13241 3160 13359
rect 2960 12680 3160 13241
rect 3440 13119 3640 13640
rect 3440 13001 3481 13119
rect 3599 13001 3640 13119
rect 3440 12680 3640 13001
rect 3920 12879 4120 13640
rect 3920 12761 3961 12879
rect 4079 12761 4120 12879
rect 3920 12680 4120 12761
rect 6480 12879 6680 13640
rect 6480 12761 6521 12879
rect 6639 12761 6680 12879
rect 6480 12680 6680 12761
rect 6960 13119 7160 13640
rect 6960 13001 7001 13119
rect 7119 13001 7160 13119
rect 6960 12680 7160 13001
rect 7440 13359 7640 13640
rect 7440 13241 7481 13359
rect 7599 13241 7640 13359
rect 7440 12680 7640 13241
rect 7920 13599 8120 13640
rect 7920 13481 7961 13599
rect 8079 13481 8120 13599
rect 7920 12680 8120 13481
rect 8400 13359 8600 13640
rect 8400 13241 8441 13359
rect 8559 13241 8600 13359
rect 8400 12680 8600 13241
rect 8880 13599 9080 13640
rect 8880 13481 8921 13599
rect 9039 13481 9080 13599
rect 8880 12680 9080 13481
rect 9360 13359 9560 13640
rect 9360 13241 9401 13359
rect 9519 13241 9560 13359
rect 9360 12680 9560 13241
rect 9840 13119 10040 13640
rect 9840 13001 9881 13119
rect 9999 13001 10040 13119
rect 9840 12680 10040 13001
rect 10320 12879 10520 13640
rect 10320 12761 10361 12879
rect 10479 12761 10520 12879
rect 10320 12680 10520 12761
rect 80 10640 280 10680
rect 560 10640 760 10680
rect 1040 10640 1240 10680
rect 1520 10640 1720 10680
rect 2000 10640 2200 10680
rect 2480 10640 2680 10680
rect 2960 10640 3160 10680
rect 3440 10640 3640 10680
rect 3920 10640 4120 10680
rect 6480 10640 6680 10680
rect 6960 10640 7160 10680
rect 7440 10640 7640 10680
rect 7920 10640 8120 10680
rect 8400 10640 8600 10680
rect 8880 10640 9080 10680
rect 9360 10640 9560 10680
rect 9840 10640 10040 10680
rect 10320 10640 10520 10680
rect 80 7600 280 7640
rect 560 7600 760 7640
rect 1040 7600 1240 7640
rect 1520 7600 1720 7640
rect 2000 7600 2200 7640
rect 2480 7600 2680 7640
rect 2960 7600 3160 7640
rect 3440 7600 3640 7640
rect 3920 7600 4120 7640
rect 6480 7600 6680 7640
rect 6960 7600 7160 7640
rect 7440 7600 7640 7640
rect 7920 7600 8120 7640
rect 8400 7600 8600 7640
rect 8880 7600 9080 7640
rect 9360 7600 9560 7640
rect 9840 7600 10040 7640
rect 10320 7600 10520 7640
rect 80 5560 280 5600
rect 560 5560 760 5600
rect 1040 5560 1240 5600
rect 1520 5560 1720 5600
rect 2000 5560 2200 5600
rect 2480 5560 2680 5600
rect 2960 5560 3160 5600
rect 3440 5560 3640 5600
rect 3920 5560 4120 5600
rect 6480 5560 6680 5600
rect 6960 5560 7160 5600
rect 7440 5560 7640 5600
rect 7920 5560 8120 5600
rect 8400 5560 8600 5600
rect 8880 5560 9080 5600
rect 9360 5560 9560 5600
rect 9840 5560 10040 5600
rect 10320 5560 10520 5600
rect 80 -40 280 0
rect 560 -40 760 0
rect 1040 -40 1240 0
rect 1520 -40 1720 0
rect 2000 -40 2200 0
rect 2480 -40 2680 0
rect 2960 -40 3160 0
rect 3440 -40 3640 0
rect 3920 -40 4120 0
use invt  br
timestamp 1638148091
transform -1 0 10600 0 1 7640
box -13 -13 4213 3013
use invt  bl
timestamp 1638148091
transform 1 0 0 0 1 7640
box -13 -13 4213 3013
use inv_2_2  ar
timestamp 1638148091
transform -1 0 10600 0 1 5600
box -13 -13 4213 2013
use inv_2_2  cr
timestamp 1638148091
transform -1 0 10600 0 1 10680
box -13 -13 4213 2013
use inv_2_2  cl
timestamp 1638148091
transform 1 0 0 0 1 10680
box -13 -13 4213 2013
use inv_2_2  al
timestamp 1638148091
transform 1 0 0 0 1 5600
box -13 -13 4213 2013
use inv_bias  biasr
timestamp 1638148091
transform -1 0 10600 0 1 520
box -13 -533 4213 5053
use inv_bias  biasl
timestamp 1638148091
transform 1 0 0 0 1 520
box -13 -533 4213 5053
<< labels >>
rlabel metal3 s 4800 -40 4840 0 4 im
port 1 nsew
rlabel metal3 s 5760 -40 5800 0 4 ip
port 2 nsew
rlabel metal3 s 5120 -40 5160 0 4 out
port 3 nsew
rlabel metal3 s 4320 -40 4360 0 4 ib
port 4 nsew
rlabel metal3 s 6240 -40 6280 0 4 q
port 5 nsew
rlabel metal5 s 80 -40 280 0 4 vdda
port 6 nsew
rlabel metal3 s 4560 -40 4600 0 4 bp
port 7 nsew
rlabel metal5 s 560 -40 760 0 4 vddx
port 8 nsew
rlabel metal5 s 1040 -40 1240 0 4 gnda
port 9 nsew
rlabel metal5 s 1520 -40 1720 0 4 vssa
port 10 nsew
rlabel metal3 s 5200 -40 5240 0 4 xn
port 11 nsew
rlabel metal3 s 5360 -40 5400 0 4 xp
port 12 nsew
rlabel metal3 s 4960 -40 5000 0 4 x
port 13 nsew
rlabel metal3 s 5600 -40 5640 0 4 y
port 14 nsew
rlabel metal3 s 6000 -40 6040 0 4 z
port 15 nsew
<< end >>
