* NGSPICE file created from cap1_10_dummy.ext - technology: sky130A

.subckt cap1_10_dummy gnda vssa
X0 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X1 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X2 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X3 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X4 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X5 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1.2e+06u
X6 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X7 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X8 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X9 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X10 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X11 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1.2e+06u
X12 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
.ends

