* load testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0

.include "array.spice"
.include "load.spice"

* supply voltages
vdda	vdda 0 1.8
vgnda	gnda 0 0.9
vssa	vssa 0 0.0

* bias current
IB ib vssa 10n

* input signals
vin	in gnda dc 0 ac 1 SINE(0 5m 1 0 0 0)
einp	ip gnda in gnda  0.5
einm	im gnda in gnda -0.5

* DUT
CP ip xp 10p
CM im xm 10p
x0 xp xm ib vdda gnda vssa load3
*x0 ip im ib vdda gnda vssa load2

*eo out vssa xp xm 1

.option gmin=1e-14
.option scale=1e-6
.control
	op
	print xp xm ib
	
*	dc vin -0.9 0.9 10m
*	let iop = i(einp)
*	plot deriv(iop)
	
	
	ac DEC 10 1m 1k
	plot vdb(xp,xm)
	
	noise v(xp,xm) vin dec 10 1 100
	print inoise_total
	
.endc

.end
