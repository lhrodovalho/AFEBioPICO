magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< error_p >>
rect 8 5920 8392 5992
rect 8 5840 80 5920
rect 94 5880 8306 5906
rect 94 3960 120 5880
rect 160 5814 8240 5840
rect 160 4072 232 5814
rect 8214 4072 8240 5814
rect 160 4000 8240 4072
rect 8280 3960 8306 5880
rect 8320 4000 8392 5920
rect 94 3934 8306 3960
rect 8 3680 8392 3752
rect 8 3600 80 3680
rect 94 3640 8306 3666
rect 94 1720 120 3640
rect 160 3574 8240 3600
rect 160 1832 232 3574
rect 8214 1832 8240 3574
rect 160 1760 8240 1832
rect 8280 1720 8306 3640
rect 8320 1760 8392 3680
rect 94 1694 8306 1720
<< nwell >>
rect 120 3960 8280 5880
rect 120 1720 8280 3640
<< pwell >>
rect -26 5894 8426 6026
rect -26 3946 106 5894
rect 8294 3946 8426 5894
rect -26 3654 8426 3946
rect -26 1706 106 3654
rect 8294 1706 8426 3654
rect -26 1574 8426 1706
rect -26 934 8426 1066
rect -26 106 106 934
rect 294 106 8106 934
rect 8294 106 8426 934
rect -26 -26 8426 106
<< mvnmos >>
rect 520 560 2120 760
rect 2440 560 4040 760
rect 4360 560 5960 760
rect 6280 560 7880 760
rect 520 160 2120 360
rect 2440 160 4040 360
rect 4360 160 5960 360
rect 6280 160 7880 360
<< mvpmos >>
rect 520 5080 2120 5680
rect 2440 5080 4040 5680
rect 4360 5080 5960 5680
rect 6280 5080 7880 5680
rect 520 4320 2120 4920
rect 2440 4320 4040 4920
rect 4360 4320 5960 4920
rect 6280 4320 7880 4920
rect 520 2840 2120 3440
rect 2440 2840 4040 3440
rect 4360 2840 5960 3440
rect 6280 2840 7880 3440
rect 520 2080 2120 2680
rect 2440 2080 4040 2680
rect 4360 2080 5960 2680
rect 6280 2080 7880 2680
<< mvndiff >>
rect 320 711 520 760
rect 320 677 343 711
rect 377 677 520 711
rect 320 643 520 677
rect 320 609 343 643
rect 377 609 520 643
rect 320 560 520 609
rect 2120 711 2440 760
rect 2120 677 2263 711
rect 2297 677 2440 711
rect 2120 643 2440 677
rect 2120 609 2263 643
rect 2297 609 2440 643
rect 2120 560 2440 609
rect 4040 711 4360 760
rect 4040 677 4183 711
rect 4217 677 4360 711
rect 4040 643 4360 677
rect 4040 609 4183 643
rect 4217 609 4360 643
rect 4040 560 4360 609
rect 5960 711 6280 760
rect 5960 677 6103 711
rect 6137 677 6280 711
rect 5960 643 6280 677
rect 5960 609 6103 643
rect 6137 609 6280 643
rect 5960 560 6280 609
rect 7880 711 8080 760
rect 7880 677 8023 711
rect 8057 677 8080 711
rect 7880 643 8080 677
rect 7880 609 8023 643
rect 8057 609 8080 643
rect 7880 560 8080 609
rect 320 311 520 360
rect 320 277 343 311
rect 377 277 520 311
rect 320 243 520 277
rect 320 209 343 243
rect 377 209 520 243
rect 320 160 520 209
rect 2120 311 2440 360
rect 2120 277 2263 311
rect 2297 277 2440 311
rect 2120 243 2440 277
rect 2120 209 2263 243
rect 2297 209 2440 243
rect 2120 160 2440 209
rect 4040 311 4360 360
rect 4040 277 4183 311
rect 4217 277 4360 311
rect 4040 243 4360 277
rect 4040 209 4183 243
rect 4217 209 4360 243
rect 4040 160 4360 209
rect 5960 311 6280 360
rect 5960 277 6103 311
rect 6137 277 6280 311
rect 5960 243 6280 277
rect 5960 209 6103 243
rect 6137 209 6280 243
rect 5960 160 6280 209
rect 7880 311 8080 360
rect 7880 277 8023 311
rect 8057 277 8080 311
rect 7880 243 8080 277
rect 7880 209 8023 243
rect 8057 209 8080 243
rect 7880 160 8080 209
<< mvpdiff >>
rect 320 5635 520 5680
rect 320 5601 343 5635
rect 377 5601 520 5635
rect 320 5567 520 5601
rect 320 5533 343 5567
rect 377 5533 520 5567
rect 320 5499 520 5533
rect 320 5465 343 5499
rect 377 5465 520 5499
rect 320 5431 520 5465
rect 320 5397 343 5431
rect 377 5397 520 5431
rect 320 5363 520 5397
rect 320 5329 343 5363
rect 377 5329 520 5363
rect 320 5295 520 5329
rect 320 5261 343 5295
rect 377 5261 520 5295
rect 320 5227 520 5261
rect 320 5193 343 5227
rect 377 5193 520 5227
rect 320 5159 520 5193
rect 320 5125 343 5159
rect 377 5125 520 5159
rect 320 5080 520 5125
rect 2120 5635 2440 5680
rect 2120 5601 2263 5635
rect 2297 5601 2440 5635
rect 2120 5567 2440 5601
rect 2120 5533 2263 5567
rect 2297 5533 2440 5567
rect 2120 5499 2440 5533
rect 2120 5465 2263 5499
rect 2297 5465 2440 5499
rect 2120 5431 2440 5465
rect 2120 5397 2263 5431
rect 2297 5397 2440 5431
rect 2120 5363 2440 5397
rect 2120 5329 2263 5363
rect 2297 5329 2440 5363
rect 2120 5295 2440 5329
rect 2120 5261 2263 5295
rect 2297 5261 2440 5295
rect 2120 5227 2440 5261
rect 2120 5193 2263 5227
rect 2297 5193 2440 5227
rect 2120 5159 2440 5193
rect 2120 5125 2263 5159
rect 2297 5125 2440 5159
rect 2120 5080 2440 5125
rect 4040 5635 4360 5680
rect 4040 5601 4183 5635
rect 4217 5601 4360 5635
rect 4040 5567 4360 5601
rect 4040 5533 4183 5567
rect 4217 5533 4360 5567
rect 4040 5499 4360 5533
rect 4040 5465 4183 5499
rect 4217 5465 4360 5499
rect 4040 5431 4360 5465
rect 4040 5397 4183 5431
rect 4217 5397 4360 5431
rect 4040 5363 4360 5397
rect 4040 5329 4183 5363
rect 4217 5329 4360 5363
rect 4040 5295 4360 5329
rect 4040 5261 4183 5295
rect 4217 5261 4360 5295
rect 4040 5227 4360 5261
rect 4040 5193 4183 5227
rect 4217 5193 4360 5227
rect 4040 5159 4360 5193
rect 4040 5125 4183 5159
rect 4217 5125 4360 5159
rect 4040 5080 4360 5125
rect 5960 5635 6280 5680
rect 5960 5601 6103 5635
rect 6137 5601 6280 5635
rect 5960 5567 6280 5601
rect 5960 5533 6103 5567
rect 6137 5533 6280 5567
rect 5960 5499 6280 5533
rect 5960 5465 6103 5499
rect 6137 5465 6280 5499
rect 5960 5431 6280 5465
rect 5960 5397 6103 5431
rect 6137 5397 6280 5431
rect 5960 5363 6280 5397
rect 5960 5329 6103 5363
rect 6137 5329 6280 5363
rect 5960 5295 6280 5329
rect 5960 5261 6103 5295
rect 6137 5261 6280 5295
rect 5960 5227 6280 5261
rect 5960 5193 6103 5227
rect 6137 5193 6280 5227
rect 5960 5159 6280 5193
rect 5960 5125 6103 5159
rect 6137 5125 6280 5159
rect 5960 5080 6280 5125
rect 7880 5635 8080 5680
rect 7880 5601 8023 5635
rect 8057 5601 8080 5635
rect 7880 5567 8080 5601
rect 7880 5533 8023 5567
rect 8057 5533 8080 5567
rect 7880 5499 8080 5533
rect 7880 5465 8023 5499
rect 8057 5465 8080 5499
rect 7880 5431 8080 5465
rect 7880 5397 8023 5431
rect 8057 5397 8080 5431
rect 7880 5363 8080 5397
rect 7880 5329 8023 5363
rect 8057 5329 8080 5363
rect 7880 5295 8080 5329
rect 7880 5261 8023 5295
rect 8057 5261 8080 5295
rect 7880 5227 8080 5261
rect 7880 5193 8023 5227
rect 8057 5193 8080 5227
rect 7880 5159 8080 5193
rect 7880 5125 8023 5159
rect 8057 5125 8080 5159
rect 7880 5080 8080 5125
rect 320 4875 520 4920
rect 320 4841 343 4875
rect 377 4841 520 4875
rect 320 4807 520 4841
rect 320 4773 343 4807
rect 377 4773 520 4807
rect 320 4739 520 4773
rect 320 4705 343 4739
rect 377 4705 520 4739
rect 320 4671 520 4705
rect 320 4637 343 4671
rect 377 4637 520 4671
rect 320 4603 520 4637
rect 320 4569 343 4603
rect 377 4569 520 4603
rect 320 4535 520 4569
rect 320 4501 343 4535
rect 377 4501 520 4535
rect 320 4467 520 4501
rect 320 4433 343 4467
rect 377 4433 520 4467
rect 320 4399 520 4433
rect 320 4365 343 4399
rect 377 4365 520 4399
rect 320 4320 520 4365
rect 2120 4875 2440 4920
rect 2120 4841 2263 4875
rect 2297 4841 2440 4875
rect 2120 4807 2440 4841
rect 2120 4773 2263 4807
rect 2297 4773 2440 4807
rect 2120 4739 2440 4773
rect 2120 4705 2263 4739
rect 2297 4705 2440 4739
rect 2120 4671 2440 4705
rect 2120 4637 2263 4671
rect 2297 4637 2440 4671
rect 2120 4603 2440 4637
rect 2120 4569 2263 4603
rect 2297 4569 2440 4603
rect 2120 4535 2440 4569
rect 2120 4501 2263 4535
rect 2297 4501 2440 4535
rect 2120 4467 2440 4501
rect 2120 4433 2263 4467
rect 2297 4433 2440 4467
rect 2120 4399 2440 4433
rect 2120 4365 2263 4399
rect 2297 4365 2440 4399
rect 2120 4320 2440 4365
rect 4040 4875 4360 4920
rect 4040 4841 4183 4875
rect 4217 4841 4360 4875
rect 4040 4807 4360 4841
rect 4040 4773 4183 4807
rect 4217 4773 4360 4807
rect 4040 4739 4360 4773
rect 4040 4705 4183 4739
rect 4217 4705 4360 4739
rect 4040 4671 4360 4705
rect 4040 4637 4183 4671
rect 4217 4637 4360 4671
rect 4040 4603 4360 4637
rect 4040 4569 4183 4603
rect 4217 4569 4360 4603
rect 4040 4535 4360 4569
rect 4040 4501 4183 4535
rect 4217 4501 4360 4535
rect 4040 4467 4360 4501
rect 4040 4433 4183 4467
rect 4217 4433 4360 4467
rect 4040 4399 4360 4433
rect 4040 4365 4183 4399
rect 4217 4365 4360 4399
rect 4040 4320 4360 4365
rect 5960 4875 6280 4920
rect 5960 4841 6103 4875
rect 6137 4841 6280 4875
rect 5960 4807 6280 4841
rect 5960 4773 6103 4807
rect 6137 4773 6280 4807
rect 5960 4739 6280 4773
rect 5960 4705 6103 4739
rect 6137 4705 6280 4739
rect 5960 4671 6280 4705
rect 5960 4637 6103 4671
rect 6137 4637 6280 4671
rect 5960 4603 6280 4637
rect 5960 4569 6103 4603
rect 6137 4569 6280 4603
rect 5960 4535 6280 4569
rect 5960 4501 6103 4535
rect 6137 4501 6280 4535
rect 5960 4467 6280 4501
rect 5960 4433 6103 4467
rect 6137 4433 6280 4467
rect 5960 4399 6280 4433
rect 5960 4365 6103 4399
rect 6137 4365 6280 4399
rect 5960 4320 6280 4365
rect 7880 4875 8080 4920
rect 7880 4841 8023 4875
rect 8057 4841 8080 4875
rect 7880 4807 8080 4841
rect 7880 4773 8023 4807
rect 8057 4773 8080 4807
rect 7880 4739 8080 4773
rect 7880 4705 8023 4739
rect 8057 4705 8080 4739
rect 7880 4671 8080 4705
rect 7880 4637 8023 4671
rect 8057 4637 8080 4671
rect 7880 4603 8080 4637
rect 7880 4569 8023 4603
rect 8057 4569 8080 4603
rect 7880 4535 8080 4569
rect 7880 4501 8023 4535
rect 8057 4501 8080 4535
rect 7880 4467 8080 4501
rect 7880 4433 8023 4467
rect 8057 4433 8080 4467
rect 7880 4399 8080 4433
rect 7880 4365 8023 4399
rect 8057 4365 8080 4399
rect 7880 4320 8080 4365
rect 320 3395 520 3440
rect 320 3361 343 3395
rect 377 3361 520 3395
rect 320 3327 520 3361
rect 320 3293 343 3327
rect 377 3293 520 3327
rect 320 3259 520 3293
rect 320 3225 343 3259
rect 377 3225 520 3259
rect 320 3191 520 3225
rect 320 3157 343 3191
rect 377 3157 520 3191
rect 320 3123 520 3157
rect 320 3089 343 3123
rect 377 3089 520 3123
rect 320 3055 520 3089
rect 320 3021 343 3055
rect 377 3021 520 3055
rect 320 2987 520 3021
rect 320 2953 343 2987
rect 377 2953 520 2987
rect 320 2919 520 2953
rect 320 2885 343 2919
rect 377 2885 520 2919
rect 320 2840 520 2885
rect 2120 3395 2440 3440
rect 2120 3361 2263 3395
rect 2297 3361 2440 3395
rect 2120 3327 2440 3361
rect 2120 3293 2263 3327
rect 2297 3293 2440 3327
rect 2120 3259 2440 3293
rect 2120 3225 2263 3259
rect 2297 3225 2440 3259
rect 2120 3191 2440 3225
rect 2120 3157 2263 3191
rect 2297 3157 2440 3191
rect 2120 3123 2440 3157
rect 2120 3089 2263 3123
rect 2297 3089 2440 3123
rect 2120 3055 2440 3089
rect 2120 3021 2263 3055
rect 2297 3021 2440 3055
rect 2120 2987 2440 3021
rect 2120 2953 2263 2987
rect 2297 2953 2440 2987
rect 2120 2919 2440 2953
rect 2120 2885 2263 2919
rect 2297 2885 2440 2919
rect 2120 2840 2440 2885
rect 4040 3395 4360 3440
rect 4040 3361 4183 3395
rect 4217 3361 4360 3395
rect 4040 3327 4360 3361
rect 4040 3293 4183 3327
rect 4217 3293 4360 3327
rect 4040 3259 4360 3293
rect 4040 3225 4183 3259
rect 4217 3225 4360 3259
rect 4040 3191 4360 3225
rect 4040 3157 4183 3191
rect 4217 3157 4360 3191
rect 4040 3123 4360 3157
rect 4040 3089 4183 3123
rect 4217 3089 4360 3123
rect 4040 3055 4360 3089
rect 4040 3021 4183 3055
rect 4217 3021 4360 3055
rect 4040 2987 4360 3021
rect 4040 2953 4183 2987
rect 4217 2953 4360 2987
rect 4040 2919 4360 2953
rect 4040 2885 4183 2919
rect 4217 2885 4360 2919
rect 4040 2840 4360 2885
rect 5960 3395 6280 3440
rect 5960 3361 6103 3395
rect 6137 3361 6280 3395
rect 5960 3327 6280 3361
rect 5960 3293 6103 3327
rect 6137 3293 6280 3327
rect 5960 3259 6280 3293
rect 5960 3225 6103 3259
rect 6137 3225 6280 3259
rect 5960 3191 6280 3225
rect 5960 3157 6103 3191
rect 6137 3157 6280 3191
rect 5960 3123 6280 3157
rect 5960 3089 6103 3123
rect 6137 3089 6280 3123
rect 5960 3055 6280 3089
rect 5960 3021 6103 3055
rect 6137 3021 6280 3055
rect 5960 2987 6280 3021
rect 5960 2953 6103 2987
rect 6137 2953 6280 2987
rect 5960 2919 6280 2953
rect 5960 2885 6103 2919
rect 6137 2885 6280 2919
rect 5960 2840 6280 2885
rect 7880 3395 8080 3440
rect 7880 3361 8023 3395
rect 8057 3361 8080 3395
rect 7880 3327 8080 3361
rect 7880 3293 8023 3327
rect 8057 3293 8080 3327
rect 7880 3259 8080 3293
rect 7880 3225 8023 3259
rect 8057 3225 8080 3259
rect 7880 3191 8080 3225
rect 7880 3157 8023 3191
rect 8057 3157 8080 3191
rect 7880 3123 8080 3157
rect 7880 3089 8023 3123
rect 8057 3089 8080 3123
rect 7880 3055 8080 3089
rect 7880 3021 8023 3055
rect 8057 3021 8080 3055
rect 7880 2987 8080 3021
rect 7880 2953 8023 2987
rect 8057 2953 8080 2987
rect 7880 2919 8080 2953
rect 7880 2885 8023 2919
rect 8057 2885 8080 2919
rect 7880 2840 8080 2885
rect 320 2635 520 2680
rect 320 2601 343 2635
rect 377 2601 520 2635
rect 320 2567 520 2601
rect 320 2533 343 2567
rect 377 2533 520 2567
rect 320 2499 520 2533
rect 320 2465 343 2499
rect 377 2465 520 2499
rect 320 2431 520 2465
rect 320 2397 343 2431
rect 377 2397 520 2431
rect 320 2363 520 2397
rect 320 2329 343 2363
rect 377 2329 520 2363
rect 320 2295 520 2329
rect 320 2261 343 2295
rect 377 2261 520 2295
rect 320 2227 520 2261
rect 320 2193 343 2227
rect 377 2193 520 2227
rect 320 2159 520 2193
rect 320 2125 343 2159
rect 377 2125 520 2159
rect 320 2080 520 2125
rect 2120 2635 2440 2680
rect 2120 2601 2263 2635
rect 2297 2601 2440 2635
rect 2120 2567 2440 2601
rect 2120 2533 2263 2567
rect 2297 2533 2440 2567
rect 2120 2499 2440 2533
rect 2120 2465 2263 2499
rect 2297 2465 2440 2499
rect 2120 2431 2440 2465
rect 2120 2397 2263 2431
rect 2297 2397 2440 2431
rect 2120 2363 2440 2397
rect 2120 2329 2263 2363
rect 2297 2329 2440 2363
rect 2120 2295 2440 2329
rect 2120 2261 2263 2295
rect 2297 2261 2440 2295
rect 2120 2227 2440 2261
rect 2120 2193 2263 2227
rect 2297 2193 2440 2227
rect 2120 2159 2440 2193
rect 2120 2125 2263 2159
rect 2297 2125 2440 2159
rect 2120 2080 2440 2125
rect 4040 2635 4360 2680
rect 4040 2601 4183 2635
rect 4217 2601 4360 2635
rect 4040 2567 4360 2601
rect 4040 2533 4183 2567
rect 4217 2533 4360 2567
rect 4040 2499 4360 2533
rect 4040 2465 4183 2499
rect 4217 2465 4360 2499
rect 4040 2431 4360 2465
rect 4040 2397 4183 2431
rect 4217 2397 4360 2431
rect 4040 2363 4360 2397
rect 4040 2329 4183 2363
rect 4217 2329 4360 2363
rect 4040 2295 4360 2329
rect 4040 2261 4183 2295
rect 4217 2261 4360 2295
rect 4040 2227 4360 2261
rect 4040 2193 4183 2227
rect 4217 2193 4360 2227
rect 4040 2159 4360 2193
rect 4040 2125 4183 2159
rect 4217 2125 4360 2159
rect 4040 2080 4360 2125
rect 5960 2635 6280 2680
rect 5960 2601 6103 2635
rect 6137 2601 6280 2635
rect 5960 2567 6280 2601
rect 5960 2533 6103 2567
rect 6137 2533 6280 2567
rect 5960 2499 6280 2533
rect 5960 2465 6103 2499
rect 6137 2465 6280 2499
rect 5960 2431 6280 2465
rect 5960 2397 6103 2431
rect 6137 2397 6280 2431
rect 5960 2363 6280 2397
rect 5960 2329 6103 2363
rect 6137 2329 6280 2363
rect 5960 2295 6280 2329
rect 5960 2261 6103 2295
rect 6137 2261 6280 2295
rect 5960 2227 6280 2261
rect 5960 2193 6103 2227
rect 6137 2193 6280 2227
rect 5960 2159 6280 2193
rect 5960 2125 6103 2159
rect 6137 2125 6280 2159
rect 5960 2080 6280 2125
rect 7880 2635 8080 2680
rect 7880 2601 8023 2635
rect 8057 2601 8080 2635
rect 7880 2567 8080 2601
rect 7880 2533 8023 2567
rect 8057 2533 8080 2567
rect 7880 2499 8080 2533
rect 7880 2465 8023 2499
rect 8057 2465 8080 2499
rect 7880 2431 8080 2465
rect 7880 2397 8023 2431
rect 8057 2397 8080 2431
rect 7880 2363 8080 2397
rect 7880 2329 8023 2363
rect 8057 2329 8080 2363
rect 7880 2295 8080 2329
rect 7880 2261 8023 2295
rect 8057 2261 8080 2295
rect 7880 2227 8080 2261
rect 7880 2193 8023 2227
rect 8057 2193 8080 2227
rect 7880 2159 8080 2193
rect 7880 2125 8023 2159
rect 8057 2125 8080 2159
rect 7880 2080 8080 2125
<< mvndiffc >>
rect 343 677 377 711
rect 343 609 377 643
rect 2263 677 2297 711
rect 2263 609 2297 643
rect 4183 677 4217 711
rect 4183 609 4217 643
rect 6103 677 6137 711
rect 6103 609 6137 643
rect 8023 677 8057 711
rect 8023 609 8057 643
rect 343 277 377 311
rect 343 209 377 243
rect 2263 277 2297 311
rect 2263 209 2297 243
rect 4183 277 4217 311
rect 4183 209 4217 243
rect 6103 277 6137 311
rect 6103 209 6137 243
rect 8023 277 8057 311
rect 8023 209 8057 243
<< mvpdiffc >>
rect 343 5601 377 5635
rect 343 5533 377 5567
rect 343 5465 377 5499
rect 343 5397 377 5431
rect 343 5329 377 5363
rect 343 5261 377 5295
rect 343 5193 377 5227
rect 343 5125 377 5159
rect 2263 5601 2297 5635
rect 2263 5533 2297 5567
rect 2263 5465 2297 5499
rect 2263 5397 2297 5431
rect 2263 5329 2297 5363
rect 2263 5261 2297 5295
rect 2263 5193 2297 5227
rect 2263 5125 2297 5159
rect 4183 5601 4217 5635
rect 4183 5533 4217 5567
rect 4183 5465 4217 5499
rect 4183 5397 4217 5431
rect 4183 5329 4217 5363
rect 4183 5261 4217 5295
rect 4183 5193 4217 5227
rect 4183 5125 4217 5159
rect 6103 5601 6137 5635
rect 6103 5533 6137 5567
rect 6103 5465 6137 5499
rect 6103 5397 6137 5431
rect 6103 5329 6137 5363
rect 6103 5261 6137 5295
rect 6103 5193 6137 5227
rect 6103 5125 6137 5159
rect 8023 5601 8057 5635
rect 8023 5533 8057 5567
rect 8023 5465 8057 5499
rect 8023 5397 8057 5431
rect 8023 5329 8057 5363
rect 8023 5261 8057 5295
rect 8023 5193 8057 5227
rect 8023 5125 8057 5159
rect 343 4841 377 4875
rect 343 4773 377 4807
rect 343 4705 377 4739
rect 343 4637 377 4671
rect 343 4569 377 4603
rect 343 4501 377 4535
rect 343 4433 377 4467
rect 343 4365 377 4399
rect 2263 4841 2297 4875
rect 2263 4773 2297 4807
rect 2263 4705 2297 4739
rect 2263 4637 2297 4671
rect 2263 4569 2297 4603
rect 2263 4501 2297 4535
rect 2263 4433 2297 4467
rect 2263 4365 2297 4399
rect 4183 4841 4217 4875
rect 4183 4773 4217 4807
rect 4183 4705 4217 4739
rect 4183 4637 4217 4671
rect 4183 4569 4217 4603
rect 4183 4501 4217 4535
rect 4183 4433 4217 4467
rect 4183 4365 4217 4399
rect 6103 4841 6137 4875
rect 6103 4773 6137 4807
rect 6103 4705 6137 4739
rect 6103 4637 6137 4671
rect 6103 4569 6137 4603
rect 6103 4501 6137 4535
rect 6103 4433 6137 4467
rect 6103 4365 6137 4399
rect 8023 4841 8057 4875
rect 8023 4773 8057 4807
rect 8023 4705 8057 4739
rect 8023 4637 8057 4671
rect 8023 4569 8057 4603
rect 8023 4501 8057 4535
rect 8023 4433 8057 4467
rect 8023 4365 8057 4399
rect 343 3361 377 3395
rect 343 3293 377 3327
rect 343 3225 377 3259
rect 343 3157 377 3191
rect 343 3089 377 3123
rect 343 3021 377 3055
rect 343 2953 377 2987
rect 343 2885 377 2919
rect 2263 3361 2297 3395
rect 2263 3293 2297 3327
rect 2263 3225 2297 3259
rect 2263 3157 2297 3191
rect 2263 3089 2297 3123
rect 2263 3021 2297 3055
rect 2263 2953 2297 2987
rect 2263 2885 2297 2919
rect 4183 3361 4217 3395
rect 4183 3293 4217 3327
rect 4183 3225 4217 3259
rect 4183 3157 4217 3191
rect 4183 3089 4217 3123
rect 4183 3021 4217 3055
rect 4183 2953 4217 2987
rect 4183 2885 4217 2919
rect 6103 3361 6137 3395
rect 6103 3293 6137 3327
rect 6103 3225 6137 3259
rect 6103 3157 6137 3191
rect 6103 3089 6137 3123
rect 6103 3021 6137 3055
rect 6103 2953 6137 2987
rect 6103 2885 6137 2919
rect 8023 3361 8057 3395
rect 8023 3293 8057 3327
rect 8023 3225 8057 3259
rect 8023 3157 8057 3191
rect 8023 3089 8057 3123
rect 8023 3021 8057 3055
rect 8023 2953 8057 2987
rect 8023 2885 8057 2919
rect 343 2601 377 2635
rect 343 2533 377 2567
rect 343 2465 377 2499
rect 343 2397 377 2431
rect 343 2329 377 2363
rect 343 2261 377 2295
rect 343 2193 377 2227
rect 343 2125 377 2159
rect 2263 2601 2297 2635
rect 2263 2533 2297 2567
rect 2263 2465 2297 2499
rect 2263 2397 2297 2431
rect 2263 2329 2297 2363
rect 2263 2261 2297 2295
rect 2263 2193 2297 2227
rect 2263 2125 2297 2159
rect 4183 2601 4217 2635
rect 4183 2533 4217 2567
rect 4183 2465 4217 2499
rect 4183 2397 4217 2431
rect 4183 2329 4217 2363
rect 4183 2261 4217 2295
rect 4183 2193 4217 2227
rect 4183 2125 4217 2159
rect 6103 2601 6137 2635
rect 6103 2533 6137 2567
rect 6103 2465 6137 2499
rect 6103 2397 6137 2431
rect 6103 2329 6137 2363
rect 6103 2261 6137 2295
rect 6103 2193 6137 2227
rect 6103 2125 6137 2159
rect 8023 2601 8057 2635
rect 8023 2533 8057 2567
rect 8023 2465 8057 2499
rect 8023 2397 8057 2431
rect 8023 2329 8057 2363
rect 8023 2261 8057 2295
rect 8023 2193 8057 2227
rect 8023 2125 8057 2159
<< psubdiff >>
rect 0 5977 8400 6000
rect 0 5943 137 5977
rect 171 5943 205 5977
rect 239 5943 273 5977
rect 307 5943 341 5977
rect 375 5943 409 5977
rect 443 5943 477 5977
rect 511 5943 545 5977
rect 579 5943 613 5977
rect 647 5943 681 5977
rect 715 5943 749 5977
rect 783 5943 817 5977
rect 851 5943 885 5977
rect 919 5943 953 5977
rect 987 5943 1021 5977
rect 1055 5943 1089 5977
rect 1123 5943 1157 5977
rect 1191 5943 1225 5977
rect 1259 5943 1293 5977
rect 1327 5943 1361 5977
rect 1395 5943 1429 5977
rect 1463 5943 1497 5977
rect 1531 5943 1565 5977
rect 1599 5943 1633 5977
rect 1667 5943 1701 5977
rect 1735 5943 1769 5977
rect 1803 5943 1837 5977
rect 1871 5943 1905 5977
rect 1939 5943 1973 5977
rect 2007 5943 2041 5977
rect 2075 5943 2109 5977
rect 2143 5943 2177 5977
rect 2211 5943 2245 5977
rect 2279 5943 2313 5977
rect 2347 5943 2381 5977
rect 2415 5943 2449 5977
rect 2483 5943 2517 5977
rect 2551 5943 2585 5977
rect 2619 5943 2653 5977
rect 2687 5943 2721 5977
rect 2755 5943 2789 5977
rect 2823 5943 2857 5977
rect 2891 5943 2925 5977
rect 2959 5943 2993 5977
rect 3027 5943 3061 5977
rect 3095 5943 3129 5977
rect 3163 5943 3197 5977
rect 3231 5943 3265 5977
rect 3299 5943 3333 5977
rect 3367 5943 3401 5977
rect 3435 5943 3469 5977
rect 3503 5943 3537 5977
rect 3571 5943 3605 5977
rect 3639 5943 3673 5977
rect 3707 5943 3741 5977
rect 3775 5943 3809 5977
rect 3843 5943 3877 5977
rect 3911 5943 3945 5977
rect 3979 5943 4013 5977
rect 4047 5943 4081 5977
rect 4115 5943 4149 5977
rect 4183 5943 4217 5977
rect 4251 5943 4285 5977
rect 4319 5943 4353 5977
rect 4387 5943 4421 5977
rect 4455 5943 4489 5977
rect 4523 5943 4557 5977
rect 4591 5943 4625 5977
rect 4659 5943 4693 5977
rect 4727 5943 4761 5977
rect 4795 5943 4829 5977
rect 4863 5943 4897 5977
rect 4931 5943 4965 5977
rect 4999 5943 5033 5977
rect 5067 5943 5101 5977
rect 5135 5943 5169 5977
rect 5203 5943 5237 5977
rect 5271 5943 5305 5977
rect 5339 5943 5373 5977
rect 5407 5943 5441 5977
rect 5475 5943 5509 5977
rect 5543 5943 5577 5977
rect 5611 5943 5645 5977
rect 5679 5943 5713 5977
rect 5747 5943 5781 5977
rect 5815 5943 5849 5977
rect 5883 5943 5917 5977
rect 5951 5943 5985 5977
rect 6019 5943 6053 5977
rect 6087 5943 6121 5977
rect 6155 5943 6189 5977
rect 6223 5943 6257 5977
rect 6291 5943 6325 5977
rect 6359 5943 6393 5977
rect 6427 5943 6461 5977
rect 6495 5943 6529 5977
rect 6563 5943 6597 5977
rect 6631 5943 6665 5977
rect 6699 5943 6733 5977
rect 6767 5943 6801 5977
rect 6835 5943 6869 5977
rect 6903 5943 6937 5977
rect 6971 5943 7005 5977
rect 7039 5943 7073 5977
rect 7107 5943 7141 5977
rect 7175 5943 7209 5977
rect 7243 5943 7277 5977
rect 7311 5943 7345 5977
rect 7379 5943 7413 5977
rect 7447 5943 7481 5977
rect 7515 5943 7549 5977
rect 7583 5943 7617 5977
rect 7651 5943 7685 5977
rect 7719 5943 7753 5977
rect 7787 5943 7821 5977
rect 7855 5943 7889 5977
rect 7923 5943 7957 5977
rect 7991 5943 8025 5977
rect 8059 5943 8093 5977
rect 8127 5943 8161 5977
rect 8195 5943 8229 5977
rect 8263 5943 8400 5977
rect 0 5920 8400 5943
rect 0 5855 80 5920
rect 0 5821 23 5855
rect 57 5821 80 5855
rect 8320 5855 8400 5920
rect 0 5787 80 5821
rect 0 5753 23 5787
rect 57 5753 80 5787
rect 0 5719 80 5753
rect 0 5685 23 5719
rect 57 5685 80 5719
rect 0 5651 80 5685
rect 0 5617 23 5651
rect 57 5617 80 5651
rect 0 5583 80 5617
rect 0 5549 23 5583
rect 57 5549 80 5583
rect 0 5515 80 5549
rect 0 5481 23 5515
rect 57 5481 80 5515
rect 0 5447 80 5481
rect 0 5413 23 5447
rect 57 5413 80 5447
rect 0 5379 80 5413
rect 0 5345 23 5379
rect 57 5345 80 5379
rect 0 5311 80 5345
rect 0 5277 23 5311
rect 57 5277 80 5311
rect 0 5243 80 5277
rect 0 5209 23 5243
rect 57 5209 80 5243
rect 0 5175 80 5209
rect 0 5141 23 5175
rect 57 5141 80 5175
rect 0 5107 80 5141
rect 0 5073 23 5107
rect 57 5073 80 5107
rect 0 5039 80 5073
rect 0 5005 23 5039
rect 57 5005 80 5039
rect 0 4971 80 5005
rect 0 4937 23 4971
rect 57 4937 80 4971
rect 0 4903 80 4937
rect 0 4869 23 4903
rect 57 4869 80 4903
rect 0 4835 80 4869
rect 0 4801 23 4835
rect 57 4801 80 4835
rect 0 4767 80 4801
rect 0 4733 23 4767
rect 57 4733 80 4767
rect 0 4699 80 4733
rect 0 4665 23 4699
rect 57 4665 80 4699
rect 0 4631 80 4665
rect 0 4597 23 4631
rect 57 4597 80 4631
rect 0 4563 80 4597
rect 0 4529 23 4563
rect 57 4529 80 4563
rect 0 4495 80 4529
rect 0 4461 23 4495
rect 57 4461 80 4495
rect 0 4427 80 4461
rect 0 4393 23 4427
rect 57 4393 80 4427
rect 0 4359 80 4393
rect 0 4325 23 4359
rect 57 4325 80 4359
rect 0 4291 80 4325
rect 0 4257 23 4291
rect 57 4257 80 4291
rect 0 4223 80 4257
rect 0 4189 23 4223
rect 57 4189 80 4223
rect 0 4155 80 4189
rect 0 4121 23 4155
rect 57 4121 80 4155
rect 0 4087 80 4121
rect 0 4053 23 4087
rect 57 4053 80 4087
rect 0 4019 80 4053
rect 0 3985 23 4019
rect 57 3985 80 4019
rect 8320 5821 8343 5855
rect 8377 5821 8400 5855
rect 8320 5787 8400 5821
rect 8320 5753 8343 5787
rect 8377 5753 8400 5787
rect 8320 5719 8400 5753
rect 8320 5685 8343 5719
rect 8377 5685 8400 5719
rect 8320 5651 8400 5685
rect 8320 5617 8343 5651
rect 8377 5617 8400 5651
rect 8320 5583 8400 5617
rect 8320 5549 8343 5583
rect 8377 5549 8400 5583
rect 8320 5515 8400 5549
rect 8320 5481 8343 5515
rect 8377 5481 8400 5515
rect 8320 5447 8400 5481
rect 8320 5413 8343 5447
rect 8377 5413 8400 5447
rect 8320 5379 8400 5413
rect 8320 5345 8343 5379
rect 8377 5345 8400 5379
rect 8320 5311 8400 5345
rect 8320 5277 8343 5311
rect 8377 5277 8400 5311
rect 8320 5243 8400 5277
rect 8320 5209 8343 5243
rect 8377 5209 8400 5243
rect 8320 5175 8400 5209
rect 8320 5141 8343 5175
rect 8377 5141 8400 5175
rect 8320 5107 8400 5141
rect 8320 5073 8343 5107
rect 8377 5073 8400 5107
rect 8320 5039 8400 5073
rect 8320 5005 8343 5039
rect 8377 5005 8400 5039
rect 8320 4971 8400 5005
rect 8320 4937 8343 4971
rect 8377 4937 8400 4971
rect 8320 4903 8400 4937
rect 8320 4869 8343 4903
rect 8377 4869 8400 4903
rect 8320 4835 8400 4869
rect 8320 4801 8343 4835
rect 8377 4801 8400 4835
rect 8320 4767 8400 4801
rect 8320 4733 8343 4767
rect 8377 4733 8400 4767
rect 8320 4699 8400 4733
rect 8320 4665 8343 4699
rect 8377 4665 8400 4699
rect 8320 4631 8400 4665
rect 8320 4597 8343 4631
rect 8377 4597 8400 4631
rect 8320 4563 8400 4597
rect 8320 4529 8343 4563
rect 8377 4529 8400 4563
rect 8320 4495 8400 4529
rect 8320 4461 8343 4495
rect 8377 4461 8400 4495
rect 8320 4427 8400 4461
rect 8320 4393 8343 4427
rect 8377 4393 8400 4427
rect 8320 4359 8400 4393
rect 8320 4325 8343 4359
rect 8377 4325 8400 4359
rect 8320 4291 8400 4325
rect 8320 4257 8343 4291
rect 8377 4257 8400 4291
rect 8320 4223 8400 4257
rect 8320 4189 8343 4223
rect 8377 4189 8400 4223
rect 8320 4155 8400 4189
rect 8320 4121 8343 4155
rect 8377 4121 8400 4155
rect 8320 4087 8400 4121
rect 8320 4053 8343 4087
rect 8377 4053 8400 4087
rect 8320 4019 8400 4053
rect 0 3920 80 3985
rect 8320 3985 8343 4019
rect 8377 3985 8400 4019
rect 8320 3920 8400 3985
rect 0 3897 8400 3920
rect 0 3863 151 3897
rect 185 3863 219 3897
rect 253 3863 287 3897
rect 321 3863 355 3897
rect 389 3863 423 3897
rect 457 3863 491 3897
rect 525 3863 559 3897
rect 593 3863 627 3897
rect 661 3863 695 3897
rect 729 3863 763 3897
rect 797 3863 831 3897
rect 865 3863 899 3897
rect 933 3863 967 3897
rect 1001 3863 1035 3897
rect 1069 3863 1103 3897
rect 1137 3863 1171 3897
rect 1205 3863 1239 3897
rect 1273 3863 1307 3897
rect 1341 3863 1375 3897
rect 1409 3863 1443 3897
rect 1477 3863 1511 3897
rect 1545 3863 1579 3897
rect 1613 3863 1647 3897
rect 1681 3863 1715 3897
rect 1749 3863 1783 3897
rect 1817 3863 1851 3897
rect 1885 3863 1919 3897
rect 1953 3863 1987 3897
rect 2021 3863 2055 3897
rect 2089 3863 2123 3897
rect 2157 3863 2191 3897
rect 2225 3863 2259 3897
rect 2293 3863 2327 3897
rect 2361 3863 2395 3897
rect 2429 3863 2463 3897
rect 2497 3863 2531 3897
rect 2565 3863 2599 3897
rect 2633 3863 2667 3897
rect 2701 3863 2735 3897
rect 2769 3863 2803 3897
rect 2837 3863 2871 3897
rect 2905 3863 2939 3897
rect 2973 3863 3007 3897
rect 3041 3863 3075 3897
rect 3109 3863 3143 3897
rect 3177 3863 3211 3897
rect 3245 3863 3279 3897
rect 3313 3863 3347 3897
rect 3381 3863 3415 3897
rect 3449 3863 3483 3897
rect 3517 3863 3551 3897
rect 3585 3863 3619 3897
rect 3653 3863 3687 3897
rect 3721 3863 3755 3897
rect 3789 3863 3823 3897
rect 3857 3863 3891 3897
rect 3925 3863 3959 3897
rect 3993 3863 4027 3897
rect 4061 3863 4095 3897
rect 4129 3863 4163 3897
rect 4197 3863 4231 3897
rect 4265 3863 4299 3897
rect 4333 3863 4367 3897
rect 4401 3863 4435 3897
rect 4469 3863 4503 3897
rect 4537 3863 4571 3897
rect 4605 3863 4639 3897
rect 4673 3863 4707 3897
rect 4741 3863 4775 3897
rect 4809 3863 4843 3897
rect 4877 3863 4911 3897
rect 4945 3863 4979 3897
rect 5013 3863 5047 3897
rect 5081 3863 5115 3897
rect 5149 3863 5183 3897
rect 5217 3863 5251 3897
rect 5285 3863 5319 3897
rect 5353 3863 5387 3897
rect 5421 3863 5455 3897
rect 5489 3863 5523 3897
rect 5557 3863 5591 3897
rect 5625 3863 5659 3897
rect 5693 3863 5727 3897
rect 5761 3863 5795 3897
rect 5829 3863 5863 3897
rect 5897 3863 5931 3897
rect 5965 3863 5999 3897
rect 6033 3863 6067 3897
rect 6101 3863 6135 3897
rect 6169 3863 6203 3897
rect 6237 3863 6271 3897
rect 6305 3863 6339 3897
rect 6373 3863 6407 3897
rect 6441 3863 6475 3897
rect 6509 3863 6543 3897
rect 6577 3863 6611 3897
rect 6645 3863 6679 3897
rect 6713 3863 6747 3897
rect 6781 3863 6815 3897
rect 6849 3863 6883 3897
rect 6917 3863 6951 3897
rect 6985 3863 7019 3897
rect 7053 3863 7087 3897
rect 7121 3863 7155 3897
rect 7189 3863 7223 3897
rect 7257 3863 7291 3897
rect 7325 3863 7359 3897
rect 7393 3863 7427 3897
rect 7461 3863 7495 3897
rect 7529 3863 7563 3897
rect 7597 3863 7631 3897
rect 7665 3863 7699 3897
rect 7733 3863 7767 3897
rect 7801 3863 7835 3897
rect 7869 3863 7903 3897
rect 7937 3863 7971 3897
rect 8005 3863 8039 3897
rect 8073 3863 8107 3897
rect 8141 3863 8175 3897
rect 8209 3863 8400 3897
rect 0 3840 8400 3863
rect 0 3737 8400 3760
rect 0 3703 151 3737
rect 185 3703 219 3737
rect 253 3703 287 3737
rect 321 3703 355 3737
rect 389 3703 423 3737
rect 457 3703 491 3737
rect 525 3703 559 3737
rect 593 3703 627 3737
rect 661 3703 695 3737
rect 729 3703 763 3737
rect 797 3703 831 3737
rect 865 3703 899 3737
rect 933 3703 967 3737
rect 1001 3703 1035 3737
rect 1069 3703 1103 3737
rect 1137 3703 1171 3737
rect 1205 3703 1239 3737
rect 1273 3703 1307 3737
rect 1341 3703 1375 3737
rect 1409 3703 1443 3737
rect 1477 3703 1511 3737
rect 1545 3703 1579 3737
rect 1613 3703 1647 3737
rect 1681 3703 1715 3737
rect 1749 3703 1783 3737
rect 1817 3703 1851 3737
rect 1885 3703 1919 3737
rect 1953 3703 1987 3737
rect 2021 3703 2055 3737
rect 2089 3703 2123 3737
rect 2157 3703 2191 3737
rect 2225 3703 2259 3737
rect 2293 3703 2327 3737
rect 2361 3703 2395 3737
rect 2429 3703 2463 3737
rect 2497 3703 2531 3737
rect 2565 3703 2599 3737
rect 2633 3703 2667 3737
rect 2701 3703 2735 3737
rect 2769 3703 2803 3737
rect 2837 3703 2871 3737
rect 2905 3703 2939 3737
rect 2973 3703 3007 3737
rect 3041 3703 3075 3737
rect 3109 3703 3143 3737
rect 3177 3703 3211 3737
rect 3245 3703 3279 3737
rect 3313 3703 3347 3737
rect 3381 3703 3415 3737
rect 3449 3703 3483 3737
rect 3517 3703 3551 3737
rect 3585 3703 3619 3737
rect 3653 3703 3687 3737
rect 3721 3703 3755 3737
rect 3789 3703 3823 3737
rect 3857 3703 3891 3737
rect 3925 3703 3959 3737
rect 3993 3703 4027 3737
rect 4061 3703 4095 3737
rect 4129 3703 4163 3737
rect 4197 3703 4231 3737
rect 4265 3703 4299 3737
rect 4333 3703 4367 3737
rect 4401 3703 4435 3737
rect 4469 3703 4503 3737
rect 4537 3703 4571 3737
rect 4605 3703 4639 3737
rect 4673 3703 4707 3737
rect 4741 3703 4775 3737
rect 4809 3703 4843 3737
rect 4877 3703 4911 3737
rect 4945 3703 4979 3737
rect 5013 3703 5047 3737
rect 5081 3703 5115 3737
rect 5149 3703 5183 3737
rect 5217 3703 5251 3737
rect 5285 3703 5319 3737
rect 5353 3703 5387 3737
rect 5421 3703 5455 3737
rect 5489 3703 5523 3737
rect 5557 3703 5591 3737
rect 5625 3703 5659 3737
rect 5693 3703 5727 3737
rect 5761 3703 5795 3737
rect 5829 3703 5863 3737
rect 5897 3703 5931 3737
rect 5965 3703 5999 3737
rect 6033 3703 6067 3737
rect 6101 3703 6135 3737
rect 6169 3703 6203 3737
rect 6237 3703 6271 3737
rect 6305 3703 6339 3737
rect 6373 3703 6407 3737
rect 6441 3703 6475 3737
rect 6509 3703 6543 3737
rect 6577 3703 6611 3737
rect 6645 3703 6679 3737
rect 6713 3703 6747 3737
rect 6781 3703 6815 3737
rect 6849 3703 6883 3737
rect 6917 3703 6951 3737
rect 6985 3703 7019 3737
rect 7053 3703 7087 3737
rect 7121 3703 7155 3737
rect 7189 3703 7223 3737
rect 7257 3703 7291 3737
rect 7325 3703 7359 3737
rect 7393 3703 7427 3737
rect 7461 3703 7495 3737
rect 7529 3703 7563 3737
rect 7597 3703 7631 3737
rect 7665 3703 7699 3737
rect 7733 3703 7767 3737
rect 7801 3703 7835 3737
rect 7869 3703 7903 3737
rect 7937 3703 7971 3737
rect 8005 3703 8039 3737
rect 8073 3703 8107 3737
rect 8141 3703 8175 3737
rect 8209 3703 8400 3737
rect 0 3680 8400 3703
rect 0 3615 80 3680
rect 0 3581 23 3615
rect 57 3581 80 3615
rect 8320 3615 8400 3680
rect 0 3547 80 3581
rect 0 3513 23 3547
rect 57 3513 80 3547
rect 0 3479 80 3513
rect 0 3445 23 3479
rect 57 3445 80 3479
rect 0 3411 80 3445
rect 0 3377 23 3411
rect 57 3377 80 3411
rect 0 3343 80 3377
rect 0 3309 23 3343
rect 57 3309 80 3343
rect 0 3275 80 3309
rect 0 3241 23 3275
rect 57 3241 80 3275
rect 0 3207 80 3241
rect 0 3173 23 3207
rect 57 3173 80 3207
rect 0 3139 80 3173
rect 0 3105 23 3139
rect 57 3105 80 3139
rect 0 3071 80 3105
rect 0 3037 23 3071
rect 57 3037 80 3071
rect 0 3003 80 3037
rect 0 2969 23 3003
rect 57 2969 80 3003
rect 0 2935 80 2969
rect 0 2901 23 2935
rect 57 2901 80 2935
rect 0 2867 80 2901
rect 0 2833 23 2867
rect 57 2833 80 2867
rect 0 2799 80 2833
rect 0 2765 23 2799
rect 57 2765 80 2799
rect 0 2731 80 2765
rect 0 2697 23 2731
rect 57 2697 80 2731
rect 0 2663 80 2697
rect 0 2629 23 2663
rect 57 2629 80 2663
rect 0 2595 80 2629
rect 0 2561 23 2595
rect 57 2561 80 2595
rect 0 2527 80 2561
rect 0 2493 23 2527
rect 57 2493 80 2527
rect 0 2459 80 2493
rect 0 2425 23 2459
rect 57 2425 80 2459
rect 0 2391 80 2425
rect 0 2357 23 2391
rect 57 2357 80 2391
rect 0 2323 80 2357
rect 0 2289 23 2323
rect 57 2289 80 2323
rect 0 2255 80 2289
rect 0 2221 23 2255
rect 57 2221 80 2255
rect 0 2187 80 2221
rect 0 2153 23 2187
rect 57 2153 80 2187
rect 0 2119 80 2153
rect 0 2085 23 2119
rect 57 2085 80 2119
rect 0 2051 80 2085
rect 0 2017 23 2051
rect 57 2017 80 2051
rect 0 1983 80 2017
rect 0 1949 23 1983
rect 57 1949 80 1983
rect 0 1915 80 1949
rect 0 1881 23 1915
rect 57 1881 80 1915
rect 0 1847 80 1881
rect 0 1813 23 1847
rect 57 1813 80 1847
rect 0 1779 80 1813
rect 0 1745 23 1779
rect 57 1745 80 1779
rect 8320 3581 8343 3615
rect 8377 3581 8400 3615
rect 8320 3547 8400 3581
rect 8320 3513 8343 3547
rect 8377 3513 8400 3547
rect 8320 3479 8400 3513
rect 8320 3445 8343 3479
rect 8377 3445 8400 3479
rect 8320 3411 8400 3445
rect 8320 3377 8343 3411
rect 8377 3377 8400 3411
rect 8320 3343 8400 3377
rect 8320 3309 8343 3343
rect 8377 3309 8400 3343
rect 8320 3275 8400 3309
rect 8320 3241 8343 3275
rect 8377 3241 8400 3275
rect 8320 3207 8400 3241
rect 8320 3173 8343 3207
rect 8377 3173 8400 3207
rect 8320 3139 8400 3173
rect 8320 3105 8343 3139
rect 8377 3105 8400 3139
rect 8320 3071 8400 3105
rect 8320 3037 8343 3071
rect 8377 3037 8400 3071
rect 8320 3003 8400 3037
rect 8320 2969 8343 3003
rect 8377 2969 8400 3003
rect 8320 2935 8400 2969
rect 8320 2901 8343 2935
rect 8377 2901 8400 2935
rect 8320 2867 8400 2901
rect 8320 2833 8343 2867
rect 8377 2833 8400 2867
rect 8320 2799 8400 2833
rect 8320 2765 8343 2799
rect 8377 2765 8400 2799
rect 8320 2731 8400 2765
rect 8320 2697 8343 2731
rect 8377 2697 8400 2731
rect 8320 2663 8400 2697
rect 8320 2629 8343 2663
rect 8377 2629 8400 2663
rect 8320 2595 8400 2629
rect 8320 2561 8343 2595
rect 8377 2561 8400 2595
rect 8320 2527 8400 2561
rect 8320 2493 8343 2527
rect 8377 2493 8400 2527
rect 8320 2459 8400 2493
rect 8320 2425 8343 2459
rect 8377 2425 8400 2459
rect 8320 2391 8400 2425
rect 8320 2357 8343 2391
rect 8377 2357 8400 2391
rect 8320 2323 8400 2357
rect 8320 2289 8343 2323
rect 8377 2289 8400 2323
rect 8320 2255 8400 2289
rect 8320 2221 8343 2255
rect 8377 2221 8400 2255
rect 8320 2187 8400 2221
rect 8320 2153 8343 2187
rect 8377 2153 8400 2187
rect 8320 2119 8400 2153
rect 8320 2085 8343 2119
rect 8377 2085 8400 2119
rect 8320 2051 8400 2085
rect 8320 2017 8343 2051
rect 8377 2017 8400 2051
rect 8320 1983 8400 2017
rect 8320 1949 8343 1983
rect 8377 1949 8400 1983
rect 8320 1915 8400 1949
rect 8320 1881 8343 1915
rect 8377 1881 8400 1915
rect 8320 1847 8400 1881
rect 8320 1813 8343 1847
rect 8377 1813 8400 1847
rect 8320 1779 8400 1813
rect 0 1680 80 1745
rect 8320 1745 8343 1779
rect 8377 1745 8400 1779
rect 8320 1680 8400 1745
rect 0 1657 8400 1680
rect 0 1623 137 1657
rect 171 1623 205 1657
rect 239 1623 273 1657
rect 307 1623 341 1657
rect 375 1623 409 1657
rect 443 1623 477 1657
rect 511 1623 545 1657
rect 579 1623 613 1657
rect 647 1623 681 1657
rect 715 1623 749 1657
rect 783 1623 817 1657
rect 851 1623 885 1657
rect 919 1623 953 1657
rect 987 1623 1021 1657
rect 1055 1623 1089 1657
rect 1123 1623 1157 1657
rect 1191 1623 1225 1657
rect 1259 1623 1293 1657
rect 1327 1623 1361 1657
rect 1395 1623 1429 1657
rect 1463 1623 1497 1657
rect 1531 1623 1565 1657
rect 1599 1623 1633 1657
rect 1667 1623 1701 1657
rect 1735 1623 1769 1657
rect 1803 1623 1837 1657
rect 1871 1623 1905 1657
rect 1939 1623 1973 1657
rect 2007 1623 2041 1657
rect 2075 1623 2109 1657
rect 2143 1623 2177 1657
rect 2211 1623 2245 1657
rect 2279 1623 2313 1657
rect 2347 1623 2381 1657
rect 2415 1623 2449 1657
rect 2483 1623 2517 1657
rect 2551 1623 2585 1657
rect 2619 1623 2653 1657
rect 2687 1623 2721 1657
rect 2755 1623 2789 1657
rect 2823 1623 2857 1657
rect 2891 1623 2925 1657
rect 2959 1623 2993 1657
rect 3027 1623 3061 1657
rect 3095 1623 3129 1657
rect 3163 1623 3197 1657
rect 3231 1623 3265 1657
rect 3299 1623 3333 1657
rect 3367 1623 3401 1657
rect 3435 1623 3469 1657
rect 3503 1623 3537 1657
rect 3571 1623 3605 1657
rect 3639 1623 3673 1657
rect 3707 1623 3741 1657
rect 3775 1623 3809 1657
rect 3843 1623 3877 1657
rect 3911 1623 3945 1657
rect 3979 1623 4013 1657
rect 4047 1623 4081 1657
rect 4115 1623 4149 1657
rect 4183 1623 4217 1657
rect 4251 1623 4285 1657
rect 4319 1623 4353 1657
rect 4387 1623 4421 1657
rect 4455 1623 4489 1657
rect 4523 1623 4557 1657
rect 4591 1623 4625 1657
rect 4659 1623 4693 1657
rect 4727 1623 4761 1657
rect 4795 1623 4829 1657
rect 4863 1623 4897 1657
rect 4931 1623 4965 1657
rect 4999 1623 5033 1657
rect 5067 1623 5101 1657
rect 5135 1623 5169 1657
rect 5203 1623 5237 1657
rect 5271 1623 5305 1657
rect 5339 1623 5373 1657
rect 5407 1623 5441 1657
rect 5475 1623 5509 1657
rect 5543 1623 5577 1657
rect 5611 1623 5645 1657
rect 5679 1623 5713 1657
rect 5747 1623 5781 1657
rect 5815 1623 5849 1657
rect 5883 1623 5917 1657
rect 5951 1623 5985 1657
rect 6019 1623 6053 1657
rect 6087 1623 6121 1657
rect 6155 1623 6189 1657
rect 6223 1623 6257 1657
rect 6291 1623 6325 1657
rect 6359 1623 6393 1657
rect 6427 1623 6461 1657
rect 6495 1623 6529 1657
rect 6563 1623 6597 1657
rect 6631 1623 6665 1657
rect 6699 1623 6733 1657
rect 6767 1623 6801 1657
rect 6835 1623 6869 1657
rect 6903 1623 6937 1657
rect 6971 1623 7005 1657
rect 7039 1623 7073 1657
rect 7107 1623 7141 1657
rect 7175 1623 7209 1657
rect 7243 1623 7277 1657
rect 7311 1623 7345 1657
rect 7379 1623 7413 1657
rect 7447 1623 7481 1657
rect 7515 1623 7549 1657
rect 7583 1623 7617 1657
rect 7651 1623 7685 1657
rect 7719 1623 7753 1657
rect 7787 1623 7821 1657
rect 7855 1623 7889 1657
rect 7923 1623 7957 1657
rect 7991 1623 8025 1657
rect 8059 1623 8093 1657
rect 8127 1623 8161 1657
rect 8195 1623 8229 1657
rect 8263 1623 8400 1657
rect 0 1600 8400 1623
rect 0 1017 8400 1040
rect 0 983 137 1017
rect 171 983 205 1017
rect 239 983 273 1017
rect 307 983 341 1017
rect 375 983 409 1017
rect 443 983 477 1017
rect 511 983 545 1017
rect 579 983 613 1017
rect 647 983 681 1017
rect 715 983 749 1017
rect 783 983 817 1017
rect 851 983 885 1017
rect 919 983 953 1017
rect 987 983 1021 1017
rect 1055 983 1089 1017
rect 1123 983 1157 1017
rect 1191 983 1225 1017
rect 1259 983 1293 1017
rect 1327 983 1361 1017
rect 1395 983 1429 1017
rect 1463 983 1497 1017
rect 1531 983 1565 1017
rect 1599 983 1633 1017
rect 1667 983 1701 1017
rect 1735 983 1769 1017
rect 1803 983 1837 1017
rect 1871 983 1905 1017
rect 1939 983 1973 1017
rect 2007 983 2041 1017
rect 2075 983 2109 1017
rect 2143 983 2177 1017
rect 2211 983 2245 1017
rect 2279 983 2313 1017
rect 2347 983 2381 1017
rect 2415 983 2449 1017
rect 2483 983 2517 1017
rect 2551 983 2585 1017
rect 2619 983 2653 1017
rect 2687 983 2721 1017
rect 2755 983 2789 1017
rect 2823 983 2857 1017
rect 2891 983 2925 1017
rect 2959 983 2993 1017
rect 3027 983 3061 1017
rect 3095 983 3129 1017
rect 3163 983 3197 1017
rect 3231 983 3265 1017
rect 3299 983 3333 1017
rect 3367 983 3401 1017
rect 3435 983 3469 1017
rect 3503 983 3537 1017
rect 3571 983 3605 1017
rect 3639 983 3673 1017
rect 3707 983 3741 1017
rect 3775 983 3809 1017
rect 3843 983 3877 1017
rect 3911 983 3945 1017
rect 3979 983 4013 1017
rect 4047 983 4081 1017
rect 4115 983 4149 1017
rect 4183 983 4217 1017
rect 4251 983 4285 1017
rect 4319 983 4353 1017
rect 4387 983 4421 1017
rect 4455 983 4489 1017
rect 4523 983 4557 1017
rect 4591 983 4625 1017
rect 4659 983 4693 1017
rect 4727 983 4761 1017
rect 4795 983 4829 1017
rect 4863 983 4897 1017
rect 4931 983 4965 1017
rect 4999 983 5033 1017
rect 5067 983 5101 1017
rect 5135 983 5169 1017
rect 5203 983 5237 1017
rect 5271 983 5305 1017
rect 5339 983 5373 1017
rect 5407 983 5441 1017
rect 5475 983 5509 1017
rect 5543 983 5577 1017
rect 5611 983 5645 1017
rect 5679 983 5713 1017
rect 5747 983 5781 1017
rect 5815 983 5849 1017
rect 5883 983 5917 1017
rect 5951 983 5985 1017
rect 6019 983 6053 1017
rect 6087 983 6121 1017
rect 6155 983 6189 1017
rect 6223 983 6257 1017
rect 6291 983 6325 1017
rect 6359 983 6393 1017
rect 6427 983 6461 1017
rect 6495 983 6529 1017
rect 6563 983 6597 1017
rect 6631 983 6665 1017
rect 6699 983 6733 1017
rect 6767 983 6801 1017
rect 6835 983 6869 1017
rect 6903 983 6937 1017
rect 6971 983 7005 1017
rect 7039 983 7073 1017
rect 7107 983 7141 1017
rect 7175 983 7209 1017
rect 7243 983 7277 1017
rect 7311 983 7345 1017
rect 7379 983 7413 1017
rect 7447 983 7481 1017
rect 7515 983 7549 1017
rect 7583 983 7617 1017
rect 7651 983 7685 1017
rect 7719 983 7753 1017
rect 7787 983 7821 1017
rect 7855 983 7889 1017
rect 7923 983 7957 1017
rect 7991 983 8025 1017
rect 8059 983 8093 1017
rect 8127 983 8161 1017
rect 8195 983 8229 1017
rect 8263 983 8400 1017
rect 0 960 8400 983
rect 0 911 80 960
rect 0 877 23 911
rect 57 877 80 911
rect 8320 911 8400 960
rect 0 843 80 877
rect 0 809 23 843
rect 57 809 80 843
rect 0 775 80 809
rect 0 741 23 775
rect 57 741 80 775
rect 8320 877 8343 911
rect 8377 877 8400 911
rect 8320 843 8400 877
rect 8320 809 8343 843
rect 8377 809 8400 843
rect 8320 775 8400 809
rect 0 707 80 741
rect 0 673 23 707
rect 57 673 80 707
rect 0 639 80 673
rect 0 605 23 639
rect 57 605 80 639
rect 0 571 80 605
rect 0 537 23 571
rect 57 537 80 571
rect 8320 741 8343 775
rect 8377 741 8400 775
rect 8320 707 8400 741
rect 8320 673 8343 707
rect 8377 673 8400 707
rect 8320 639 8400 673
rect 8320 605 8343 639
rect 8377 605 8400 639
rect 8320 571 8400 605
rect 0 503 80 537
rect 0 469 23 503
rect 57 469 80 503
rect 0 435 80 469
rect 0 401 23 435
rect 57 401 80 435
rect 0 367 80 401
rect 0 333 23 367
rect 57 333 80 367
rect 8320 537 8343 571
rect 8377 537 8400 571
rect 8320 503 8400 537
rect 8320 469 8343 503
rect 8377 469 8400 503
rect 8320 435 8400 469
rect 8320 401 8343 435
rect 8377 401 8400 435
rect 8320 367 8400 401
rect 0 299 80 333
rect 0 265 23 299
rect 57 265 80 299
rect 0 231 80 265
rect 0 197 23 231
rect 57 197 80 231
rect 0 163 80 197
rect 0 129 23 163
rect 57 129 80 163
rect 8320 333 8343 367
rect 8377 333 8400 367
rect 8320 299 8400 333
rect 8320 265 8343 299
rect 8377 265 8400 299
rect 8320 231 8400 265
rect 8320 197 8343 231
rect 8377 197 8400 231
rect 8320 163 8400 197
rect 0 80 80 129
rect 8320 129 8343 163
rect 8377 129 8400 163
rect 8320 80 8400 129
rect 0 57 8400 80
rect 0 23 137 57
rect 171 23 205 57
rect 239 23 273 57
rect 307 23 341 57
rect 375 23 409 57
rect 443 23 477 57
rect 511 23 545 57
rect 579 23 613 57
rect 647 23 681 57
rect 715 23 749 57
rect 783 23 817 57
rect 851 23 885 57
rect 919 23 953 57
rect 987 23 1021 57
rect 1055 23 1089 57
rect 1123 23 1157 57
rect 1191 23 1225 57
rect 1259 23 1293 57
rect 1327 23 1361 57
rect 1395 23 1429 57
rect 1463 23 1497 57
rect 1531 23 1565 57
rect 1599 23 1633 57
rect 1667 23 1701 57
rect 1735 23 1769 57
rect 1803 23 1837 57
rect 1871 23 1905 57
rect 1939 23 1973 57
rect 2007 23 2041 57
rect 2075 23 2109 57
rect 2143 23 2177 57
rect 2211 23 2245 57
rect 2279 23 2313 57
rect 2347 23 2381 57
rect 2415 23 2449 57
rect 2483 23 2517 57
rect 2551 23 2585 57
rect 2619 23 2653 57
rect 2687 23 2721 57
rect 2755 23 2789 57
rect 2823 23 2857 57
rect 2891 23 2925 57
rect 2959 23 2993 57
rect 3027 23 3061 57
rect 3095 23 3129 57
rect 3163 23 3197 57
rect 3231 23 3265 57
rect 3299 23 3333 57
rect 3367 23 3401 57
rect 3435 23 3469 57
rect 3503 23 3537 57
rect 3571 23 3605 57
rect 3639 23 3673 57
rect 3707 23 3741 57
rect 3775 23 3809 57
rect 3843 23 3877 57
rect 3911 23 3945 57
rect 3979 23 4013 57
rect 4047 23 4081 57
rect 4115 23 4149 57
rect 4183 23 4217 57
rect 4251 23 4285 57
rect 4319 23 4353 57
rect 4387 23 4421 57
rect 4455 23 4489 57
rect 4523 23 4557 57
rect 4591 23 4625 57
rect 4659 23 4693 57
rect 4727 23 4761 57
rect 4795 23 4829 57
rect 4863 23 4897 57
rect 4931 23 4965 57
rect 4999 23 5033 57
rect 5067 23 5101 57
rect 5135 23 5169 57
rect 5203 23 5237 57
rect 5271 23 5305 57
rect 5339 23 5373 57
rect 5407 23 5441 57
rect 5475 23 5509 57
rect 5543 23 5577 57
rect 5611 23 5645 57
rect 5679 23 5713 57
rect 5747 23 5781 57
rect 5815 23 5849 57
rect 5883 23 5917 57
rect 5951 23 5985 57
rect 6019 23 6053 57
rect 6087 23 6121 57
rect 6155 23 6189 57
rect 6223 23 6257 57
rect 6291 23 6325 57
rect 6359 23 6393 57
rect 6427 23 6461 57
rect 6495 23 6529 57
rect 6563 23 6597 57
rect 6631 23 6665 57
rect 6699 23 6733 57
rect 6767 23 6801 57
rect 6835 23 6869 57
rect 6903 23 6937 57
rect 6971 23 7005 57
rect 7039 23 7073 57
rect 7107 23 7141 57
rect 7175 23 7209 57
rect 7243 23 7277 57
rect 7311 23 7345 57
rect 7379 23 7413 57
rect 7447 23 7481 57
rect 7515 23 7549 57
rect 7583 23 7617 57
rect 7651 23 7685 57
rect 7719 23 7753 57
rect 7787 23 7821 57
rect 7855 23 7889 57
rect 7923 23 7957 57
rect 7991 23 8025 57
rect 8059 23 8093 57
rect 8127 23 8161 57
rect 8195 23 8229 57
rect 8263 23 8400 57
rect 0 0 8400 23
<< mvnsubdiff >>
rect 160 5817 8240 5840
rect 160 5783 307 5817
rect 341 5783 375 5817
rect 409 5783 443 5817
rect 477 5783 511 5817
rect 545 5783 579 5817
rect 613 5783 647 5817
rect 681 5783 715 5817
rect 749 5783 783 5817
rect 817 5783 851 5817
rect 885 5783 919 5817
rect 953 5783 987 5817
rect 1021 5783 1055 5817
rect 1089 5783 1123 5817
rect 1157 5783 1191 5817
rect 1225 5783 1259 5817
rect 1293 5783 1327 5817
rect 1361 5783 1395 5817
rect 1429 5783 1463 5817
rect 1497 5783 1531 5817
rect 1565 5783 1599 5817
rect 1633 5783 1667 5817
rect 1701 5783 1735 5817
rect 1769 5783 1803 5817
rect 1837 5783 1871 5817
rect 1905 5783 1939 5817
rect 1973 5783 2007 5817
rect 2041 5783 2075 5817
rect 2109 5783 2143 5817
rect 2177 5783 2211 5817
rect 2245 5783 2279 5817
rect 2313 5783 2347 5817
rect 2381 5783 2415 5817
rect 2449 5783 2483 5817
rect 2517 5783 2551 5817
rect 2585 5783 2619 5817
rect 2653 5783 2687 5817
rect 2721 5783 2755 5817
rect 2789 5783 2823 5817
rect 2857 5783 2891 5817
rect 2925 5783 2959 5817
rect 2993 5783 3027 5817
rect 3061 5783 3095 5817
rect 3129 5783 3163 5817
rect 3197 5783 3231 5817
rect 3265 5783 3299 5817
rect 3333 5783 3367 5817
rect 3401 5783 3435 5817
rect 3469 5783 3503 5817
rect 3537 5783 3571 5817
rect 3605 5783 3639 5817
rect 3673 5783 3707 5817
rect 3741 5783 3775 5817
rect 3809 5783 3843 5817
rect 3877 5783 3911 5817
rect 3945 5783 3979 5817
rect 4013 5783 4047 5817
rect 4081 5783 4115 5817
rect 4149 5783 4183 5817
rect 4217 5783 4251 5817
rect 4285 5783 4319 5817
rect 4353 5783 4387 5817
rect 4421 5783 4455 5817
rect 4489 5783 4523 5817
rect 4557 5783 4591 5817
rect 4625 5783 4659 5817
rect 4693 5783 4727 5817
rect 4761 5783 4795 5817
rect 4829 5783 4863 5817
rect 4897 5783 4931 5817
rect 4965 5783 4999 5817
rect 5033 5783 5067 5817
rect 5101 5783 5135 5817
rect 5169 5783 5203 5817
rect 5237 5783 5271 5817
rect 5305 5783 5339 5817
rect 5373 5783 5407 5817
rect 5441 5783 5475 5817
rect 5509 5783 5543 5817
rect 5577 5783 5611 5817
rect 5645 5783 5679 5817
rect 5713 5783 5747 5817
rect 5781 5783 5815 5817
rect 5849 5783 5883 5817
rect 5917 5783 5951 5817
rect 5985 5783 6019 5817
rect 6053 5783 6087 5817
rect 6121 5783 6155 5817
rect 6189 5783 6223 5817
rect 6257 5783 6291 5817
rect 6325 5783 6359 5817
rect 6393 5783 6427 5817
rect 6461 5783 6495 5817
rect 6529 5783 6563 5817
rect 6597 5783 6631 5817
rect 6665 5783 6699 5817
rect 6733 5783 6767 5817
rect 6801 5783 6835 5817
rect 6869 5783 6903 5817
rect 6937 5783 6971 5817
rect 7005 5783 7039 5817
rect 7073 5783 7107 5817
rect 7141 5783 7175 5817
rect 7209 5783 7243 5817
rect 7277 5783 7311 5817
rect 7345 5783 7379 5817
rect 7413 5783 7447 5817
rect 7481 5783 7515 5817
rect 7549 5783 7583 5817
rect 7617 5783 7651 5817
rect 7685 5783 7719 5817
rect 7753 5783 7787 5817
rect 7821 5783 7855 5817
rect 7889 5783 7923 5817
rect 7957 5783 7991 5817
rect 8025 5783 8059 5817
rect 8093 5783 8240 5817
rect 160 5760 8240 5783
rect 160 5719 240 5760
rect 160 5685 183 5719
rect 217 5685 240 5719
rect 160 5651 240 5685
rect 8160 5719 8240 5760
rect 8160 5685 8183 5719
rect 8217 5685 8240 5719
rect 160 5617 183 5651
rect 217 5617 240 5651
rect 160 5583 240 5617
rect 160 5549 183 5583
rect 217 5549 240 5583
rect 160 5515 240 5549
rect 160 5481 183 5515
rect 217 5481 240 5515
rect 160 5447 240 5481
rect 160 5413 183 5447
rect 217 5413 240 5447
rect 160 5379 240 5413
rect 160 5345 183 5379
rect 217 5345 240 5379
rect 160 5311 240 5345
rect 160 5277 183 5311
rect 217 5277 240 5311
rect 160 5243 240 5277
rect 160 5209 183 5243
rect 217 5209 240 5243
rect 160 5175 240 5209
rect 160 5141 183 5175
rect 217 5141 240 5175
rect 160 5107 240 5141
rect 160 5073 183 5107
rect 217 5073 240 5107
rect 8160 5651 8240 5685
rect 8160 5617 8183 5651
rect 8217 5617 8240 5651
rect 8160 5583 8240 5617
rect 8160 5549 8183 5583
rect 8217 5549 8240 5583
rect 8160 5515 8240 5549
rect 8160 5481 8183 5515
rect 8217 5481 8240 5515
rect 8160 5447 8240 5481
rect 8160 5413 8183 5447
rect 8217 5413 8240 5447
rect 8160 5379 8240 5413
rect 8160 5345 8183 5379
rect 8217 5345 8240 5379
rect 8160 5311 8240 5345
rect 8160 5277 8183 5311
rect 8217 5277 8240 5311
rect 8160 5243 8240 5277
rect 8160 5209 8183 5243
rect 8217 5209 8240 5243
rect 8160 5175 8240 5209
rect 8160 5141 8183 5175
rect 8217 5141 8240 5175
rect 8160 5107 8240 5141
rect 160 5039 240 5073
rect 160 5005 183 5039
rect 217 5005 240 5039
rect 160 4971 240 5005
rect 160 4937 183 4971
rect 217 4937 240 4971
rect 160 4903 240 4937
rect 8160 5073 8183 5107
rect 8217 5073 8240 5107
rect 8160 5039 8240 5073
rect 8160 5005 8183 5039
rect 8217 5005 8240 5039
rect 8160 4971 8240 5005
rect 8160 4937 8183 4971
rect 8217 4937 8240 4971
rect 160 4869 183 4903
rect 217 4869 240 4903
rect 160 4835 240 4869
rect 160 4801 183 4835
rect 217 4801 240 4835
rect 160 4767 240 4801
rect 160 4733 183 4767
rect 217 4733 240 4767
rect 160 4699 240 4733
rect 160 4665 183 4699
rect 217 4665 240 4699
rect 160 4631 240 4665
rect 160 4597 183 4631
rect 217 4597 240 4631
rect 160 4563 240 4597
rect 160 4529 183 4563
rect 217 4529 240 4563
rect 160 4495 240 4529
rect 160 4461 183 4495
rect 217 4461 240 4495
rect 160 4427 240 4461
rect 160 4393 183 4427
rect 217 4393 240 4427
rect 160 4359 240 4393
rect 160 4325 183 4359
rect 217 4325 240 4359
rect 160 4291 240 4325
rect 8160 4903 8240 4937
rect 8160 4869 8183 4903
rect 8217 4869 8240 4903
rect 8160 4835 8240 4869
rect 8160 4801 8183 4835
rect 8217 4801 8240 4835
rect 8160 4767 8240 4801
rect 8160 4733 8183 4767
rect 8217 4733 8240 4767
rect 8160 4699 8240 4733
rect 8160 4665 8183 4699
rect 8217 4665 8240 4699
rect 8160 4631 8240 4665
rect 8160 4597 8183 4631
rect 8217 4597 8240 4631
rect 8160 4563 8240 4597
rect 8160 4529 8183 4563
rect 8217 4529 8240 4563
rect 8160 4495 8240 4529
rect 8160 4461 8183 4495
rect 8217 4461 8240 4495
rect 8160 4427 8240 4461
rect 8160 4393 8183 4427
rect 8217 4393 8240 4427
rect 8160 4359 8240 4393
rect 8160 4325 8183 4359
rect 8217 4325 8240 4359
rect 160 4257 183 4291
rect 217 4257 240 4291
rect 160 4223 240 4257
rect 160 4189 183 4223
rect 217 4189 240 4223
rect 160 4155 240 4189
rect 8160 4291 8240 4325
rect 8160 4257 8183 4291
rect 8217 4257 8240 4291
rect 8160 4223 8240 4257
rect 8160 4189 8183 4223
rect 8217 4189 8240 4223
rect 160 4121 183 4155
rect 217 4121 240 4155
rect 160 4080 240 4121
rect 8160 4155 8240 4189
rect 8160 4121 8183 4155
rect 8217 4121 8240 4155
rect 8160 4080 8240 4121
rect 160 4057 8240 4080
rect 160 4023 307 4057
rect 341 4023 375 4057
rect 409 4023 443 4057
rect 477 4023 511 4057
rect 545 4023 579 4057
rect 613 4023 647 4057
rect 681 4023 715 4057
rect 749 4023 783 4057
rect 817 4023 851 4057
rect 885 4023 919 4057
rect 953 4023 987 4057
rect 1021 4023 1055 4057
rect 1089 4023 1123 4057
rect 1157 4023 1191 4057
rect 1225 4023 1259 4057
rect 1293 4023 1327 4057
rect 1361 4023 1395 4057
rect 1429 4023 1463 4057
rect 1497 4023 1531 4057
rect 1565 4023 1599 4057
rect 1633 4023 1667 4057
rect 1701 4023 1735 4057
rect 1769 4023 1803 4057
rect 1837 4023 1871 4057
rect 1905 4023 1939 4057
rect 1973 4023 2007 4057
rect 2041 4023 2075 4057
rect 2109 4023 2143 4057
rect 2177 4023 2211 4057
rect 2245 4023 2279 4057
rect 2313 4023 2347 4057
rect 2381 4023 2415 4057
rect 2449 4023 2483 4057
rect 2517 4023 2551 4057
rect 2585 4023 2619 4057
rect 2653 4023 2687 4057
rect 2721 4023 2755 4057
rect 2789 4023 2823 4057
rect 2857 4023 2891 4057
rect 2925 4023 2959 4057
rect 2993 4023 3027 4057
rect 3061 4023 3095 4057
rect 3129 4023 3163 4057
rect 3197 4023 3231 4057
rect 3265 4023 3299 4057
rect 3333 4023 3367 4057
rect 3401 4023 3435 4057
rect 3469 4023 3503 4057
rect 3537 4023 3571 4057
rect 3605 4023 3639 4057
rect 3673 4023 3707 4057
rect 3741 4023 3775 4057
rect 3809 4023 3843 4057
rect 3877 4023 3911 4057
rect 3945 4023 3979 4057
rect 4013 4023 4047 4057
rect 4081 4023 4115 4057
rect 4149 4023 4183 4057
rect 4217 4023 4251 4057
rect 4285 4023 4319 4057
rect 4353 4023 4387 4057
rect 4421 4023 4455 4057
rect 4489 4023 4523 4057
rect 4557 4023 4591 4057
rect 4625 4023 4659 4057
rect 4693 4023 4727 4057
rect 4761 4023 4795 4057
rect 4829 4023 4863 4057
rect 4897 4023 4931 4057
rect 4965 4023 4999 4057
rect 5033 4023 5067 4057
rect 5101 4023 5135 4057
rect 5169 4023 5203 4057
rect 5237 4023 5271 4057
rect 5305 4023 5339 4057
rect 5373 4023 5407 4057
rect 5441 4023 5475 4057
rect 5509 4023 5543 4057
rect 5577 4023 5611 4057
rect 5645 4023 5679 4057
rect 5713 4023 5747 4057
rect 5781 4023 5815 4057
rect 5849 4023 5883 4057
rect 5917 4023 5951 4057
rect 5985 4023 6019 4057
rect 6053 4023 6087 4057
rect 6121 4023 6155 4057
rect 6189 4023 6223 4057
rect 6257 4023 6291 4057
rect 6325 4023 6359 4057
rect 6393 4023 6427 4057
rect 6461 4023 6495 4057
rect 6529 4023 6563 4057
rect 6597 4023 6631 4057
rect 6665 4023 6699 4057
rect 6733 4023 6767 4057
rect 6801 4023 6835 4057
rect 6869 4023 6903 4057
rect 6937 4023 6971 4057
rect 7005 4023 7039 4057
rect 7073 4023 7107 4057
rect 7141 4023 7175 4057
rect 7209 4023 7243 4057
rect 7277 4023 7311 4057
rect 7345 4023 7379 4057
rect 7413 4023 7447 4057
rect 7481 4023 7515 4057
rect 7549 4023 7583 4057
rect 7617 4023 7651 4057
rect 7685 4023 7719 4057
rect 7753 4023 7787 4057
rect 7821 4023 7855 4057
rect 7889 4023 7923 4057
rect 7957 4023 7991 4057
rect 8025 4023 8059 4057
rect 8093 4023 8240 4057
rect 160 4000 8240 4023
rect 160 3577 8240 3600
rect 160 3543 307 3577
rect 341 3543 375 3577
rect 409 3543 443 3577
rect 477 3543 511 3577
rect 545 3543 579 3577
rect 613 3543 647 3577
rect 681 3543 715 3577
rect 749 3543 783 3577
rect 817 3543 851 3577
rect 885 3543 919 3577
rect 953 3543 987 3577
rect 1021 3543 1055 3577
rect 1089 3543 1123 3577
rect 1157 3543 1191 3577
rect 1225 3543 1259 3577
rect 1293 3543 1327 3577
rect 1361 3543 1395 3577
rect 1429 3543 1463 3577
rect 1497 3543 1531 3577
rect 1565 3543 1599 3577
rect 1633 3543 1667 3577
rect 1701 3543 1735 3577
rect 1769 3543 1803 3577
rect 1837 3543 1871 3577
rect 1905 3543 1939 3577
rect 1973 3543 2007 3577
rect 2041 3543 2075 3577
rect 2109 3543 2143 3577
rect 2177 3543 2211 3577
rect 2245 3543 2279 3577
rect 2313 3543 2347 3577
rect 2381 3543 2415 3577
rect 2449 3543 2483 3577
rect 2517 3543 2551 3577
rect 2585 3543 2619 3577
rect 2653 3543 2687 3577
rect 2721 3543 2755 3577
rect 2789 3543 2823 3577
rect 2857 3543 2891 3577
rect 2925 3543 2959 3577
rect 2993 3543 3027 3577
rect 3061 3543 3095 3577
rect 3129 3543 3163 3577
rect 3197 3543 3231 3577
rect 3265 3543 3299 3577
rect 3333 3543 3367 3577
rect 3401 3543 3435 3577
rect 3469 3543 3503 3577
rect 3537 3543 3571 3577
rect 3605 3543 3639 3577
rect 3673 3543 3707 3577
rect 3741 3543 3775 3577
rect 3809 3543 3843 3577
rect 3877 3543 3911 3577
rect 3945 3543 3979 3577
rect 4013 3543 4047 3577
rect 4081 3543 4115 3577
rect 4149 3543 4183 3577
rect 4217 3543 4251 3577
rect 4285 3543 4319 3577
rect 4353 3543 4387 3577
rect 4421 3543 4455 3577
rect 4489 3543 4523 3577
rect 4557 3543 4591 3577
rect 4625 3543 4659 3577
rect 4693 3543 4727 3577
rect 4761 3543 4795 3577
rect 4829 3543 4863 3577
rect 4897 3543 4931 3577
rect 4965 3543 4999 3577
rect 5033 3543 5067 3577
rect 5101 3543 5135 3577
rect 5169 3543 5203 3577
rect 5237 3543 5271 3577
rect 5305 3543 5339 3577
rect 5373 3543 5407 3577
rect 5441 3543 5475 3577
rect 5509 3543 5543 3577
rect 5577 3543 5611 3577
rect 5645 3543 5679 3577
rect 5713 3543 5747 3577
rect 5781 3543 5815 3577
rect 5849 3543 5883 3577
rect 5917 3543 5951 3577
rect 5985 3543 6019 3577
rect 6053 3543 6087 3577
rect 6121 3543 6155 3577
rect 6189 3543 6223 3577
rect 6257 3543 6291 3577
rect 6325 3543 6359 3577
rect 6393 3543 6427 3577
rect 6461 3543 6495 3577
rect 6529 3543 6563 3577
rect 6597 3543 6631 3577
rect 6665 3543 6699 3577
rect 6733 3543 6767 3577
rect 6801 3543 6835 3577
rect 6869 3543 6903 3577
rect 6937 3543 6971 3577
rect 7005 3543 7039 3577
rect 7073 3543 7107 3577
rect 7141 3543 7175 3577
rect 7209 3543 7243 3577
rect 7277 3543 7311 3577
rect 7345 3543 7379 3577
rect 7413 3543 7447 3577
rect 7481 3543 7515 3577
rect 7549 3543 7583 3577
rect 7617 3543 7651 3577
rect 7685 3543 7719 3577
rect 7753 3543 7787 3577
rect 7821 3543 7855 3577
rect 7889 3543 7923 3577
rect 7957 3543 7991 3577
rect 8025 3543 8059 3577
rect 8093 3543 8240 3577
rect 160 3520 8240 3543
rect 160 3465 240 3520
rect 160 3431 183 3465
rect 217 3431 240 3465
rect 8160 3465 8240 3520
rect 160 3397 240 3431
rect 160 3363 183 3397
rect 217 3363 240 3397
rect 160 3329 240 3363
rect 160 3295 183 3329
rect 217 3295 240 3329
rect 160 3261 240 3295
rect 160 3227 183 3261
rect 217 3227 240 3261
rect 160 3193 240 3227
rect 160 3159 183 3193
rect 217 3159 240 3193
rect 160 3125 240 3159
rect 160 3091 183 3125
rect 217 3091 240 3125
rect 160 3057 240 3091
rect 160 3023 183 3057
rect 217 3023 240 3057
rect 160 2989 240 3023
rect 160 2955 183 2989
rect 217 2955 240 2989
rect 160 2921 240 2955
rect 160 2887 183 2921
rect 217 2887 240 2921
rect 160 2853 240 2887
rect 160 2819 183 2853
rect 217 2819 240 2853
rect 8160 3431 8183 3465
rect 8217 3431 8240 3465
rect 8160 3397 8240 3431
rect 8160 3363 8183 3397
rect 8217 3363 8240 3397
rect 8160 3329 8240 3363
rect 8160 3295 8183 3329
rect 8217 3295 8240 3329
rect 8160 3261 8240 3295
rect 8160 3227 8183 3261
rect 8217 3227 8240 3261
rect 8160 3193 8240 3227
rect 8160 3159 8183 3193
rect 8217 3159 8240 3193
rect 8160 3125 8240 3159
rect 8160 3091 8183 3125
rect 8217 3091 8240 3125
rect 8160 3057 8240 3091
rect 8160 3023 8183 3057
rect 8217 3023 8240 3057
rect 8160 2989 8240 3023
rect 8160 2955 8183 2989
rect 8217 2955 8240 2989
rect 8160 2921 8240 2955
rect 8160 2887 8183 2921
rect 8217 2887 8240 2921
rect 8160 2853 8240 2887
rect 160 2785 240 2819
rect 160 2751 183 2785
rect 217 2751 240 2785
rect 160 2717 240 2751
rect 160 2683 183 2717
rect 217 2683 240 2717
rect 160 2649 240 2683
rect 8160 2819 8183 2853
rect 8217 2819 8240 2853
rect 8160 2785 8240 2819
rect 8160 2751 8183 2785
rect 8217 2751 8240 2785
rect 8160 2717 8240 2751
rect 8160 2683 8183 2717
rect 8217 2683 8240 2717
rect 160 2615 183 2649
rect 217 2615 240 2649
rect 160 2581 240 2615
rect 160 2547 183 2581
rect 217 2547 240 2581
rect 160 2513 240 2547
rect 160 2479 183 2513
rect 217 2479 240 2513
rect 160 2445 240 2479
rect 160 2411 183 2445
rect 217 2411 240 2445
rect 160 2377 240 2411
rect 160 2343 183 2377
rect 217 2343 240 2377
rect 160 2309 240 2343
rect 160 2275 183 2309
rect 217 2275 240 2309
rect 160 2241 240 2275
rect 160 2207 183 2241
rect 217 2207 240 2241
rect 160 2173 240 2207
rect 160 2139 183 2173
rect 217 2139 240 2173
rect 160 2105 240 2139
rect 160 2071 183 2105
rect 217 2071 240 2105
rect 8160 2649 8240 2683
rect 8160 2615 8183 2649
rect 8217 2615 8240 2649
rect 8160 2581 8240 2615
rect 8160 2547 8183 2581
rect 8217 2547 8240 2581
rect 8160 2513 8240 2547
rect 8160 2479 8183 2513
rect 8217 2479 8240 2513
rect 8160 2445 8240 2479
rect 8160 2411 8183 2445
rect 8217 2411 8240 2445
rect 8160 2377 8240 2411
rect 8160 2343 8183 2377
rect 8217 2343 8240 2377
rect 8160 2309 8240 2343
rect 8160 2275 8183 2309
rect 8217 2275 8240 2309
rect 8160 2241 8240 2275
rect 8160 2207 8183 2241
rect 8217 2207 8240 2241
rect 8160 2173 8240 2207
rect 8160 2139 8183 2173
rect 8217 2139 8240 2173
rect 8160 2105 8240 2139
rect 160 2037 240 2071
rect 160 2003 183 2037
rect 217 2003 240 2037
rect 160 1969 240 2003
rect 160 1935 183 1969
rect 217 1935 240 1969
rect 160 1840 240 1935
rect 8160 2071 8183 2105
rect 8217 2071 8240 2105
rect 8160 2037 8240 2071
rect 8160 2003 8183 2037
rect 8217 2003 8240 2037
rect 8160 1969 8240 2003
rect 8160 1935 8183 1969
rect 8217 1935 8240 1969
rect 8160 1840 8240 1935
rect 160 1817 8240 1840
rect 160 1783 307 1817
rect 341 1783 375 1817
rect 409 1783 443 1817
rect 477 1783 511 1817
rect 545 1783 579 1817
rect 613 1783 647 1817
rect 681 1783 715 1817
rect 749 1783 783 1817
rect 817 1783 851 1817
rect 885 1783 919 1817
rect 953 1783 987 1817
rect 1021 1783 1055 1817
rect 1089 1783 1123 1817
rect 1157 1783 1191 1817
rect 1225 1783 1259 1817
rect 1293 1783 1327 1817
rect 1361 1783 1395 1817
rect 1429 1783 1463 1817
rect 1497 1783 1531 1817
rect 1565 1783 1599 1817
rect 1633 1783 1667 1817
rect 1701 1783 1735 1817
rect 1769 1783 1803 1817
rect 1837 1783 1871 1817
rect 1905 1783 1939 1817
rect 1973 1783 2007 1817
rect 2041 1783 2075 1817
rect 2109 1783 2143 1817
rect 2177 1783 2211 1817
rect 2245 1783 2279 1817
rect 2313 1783 2347 1817
rect 2381 1783 2415 1817
rect 2449 1783 2483 1817
rect 2517 1783 2551 1817
rect 2585 1783 2619 1817
rect 2653 1783 2687 1817
rect 2721 1783 2755 1817
rect 2789 1783 2823 1817
rect 2857 1783 2891 1817
rect 2925 1783 2959 1817
rect 2993 1783 3027 1817
rect 3061 1783 3095 1817
rect 3129 1783 3163 1817
rect 3197 1783 3231 1817
rect 3265 1783 3299 1817
rect 3333 1783 3367 1817
rect 3401 1783 3435 1817
rect 3469 1783 3503 1817
rect 3537 1783 3571 1817
rect 3605 1783 3639 1817
rect 3673 1783 3707 1817
rect 3741 1783 3775 1817
rect 3809 1783 3843 1817
rect 3877 1783 3911 1817
rect 3945 1783 3979 1817
rect 4013 1783 4047 1817
rect 4081 1783 4115 1817
rect 4149 1783 4183 1817
rect 4217 1783 4251 1817
rect 4285 1783 4319 1817
rect 4353 1783 4387 1817
rect 4421 1783 4455 1817
rect 4489 1783 4523 1817
rect 4557 1783 4591 1817
rect 4625 1783 4659 1817
rect 4693 1783 4727 1817
rect 4761 1783 4795 1817
rect 4829 1783 4863 1817
rect 4897 1783 4931 1817
rect 4965 1783 4999 1817
rect 5033 1783 5067 1817
rect 5101 1783 5135 1817
rect 5169 1783 5203 1817
rect 5237 1783 5271 1817
rect 5305 1783 5339 1817
rect 5373 1783 5407 1817
rect 5441 1783 5475 1817
rect 5509 1783 5543 1817
rect 5577 1783 5611 1817
rect 5645 1783 5679 1817
rect 5713 1783 5747 1817
rect 5781 1783 5815 1817
rect 5849 1783 5883 1817
rect 5917 1783 5951 1817
rect 5985 1783 6019 1817
rect 6053 1783 6087 1817
rect 6121 1783 6155 1817
rect 6189 1783 6223 1817
rect 6257 1783 6291 1817
rect 6325 1783 6359 1817
rect 6393 1783 6427 1817
rect 6461 1783 6495 1817
rect 6529 1783 6563 1817
rect 6597 1783 6631 1817
rect 6665 1783 6699 1817
rect 6733 1783 6767 1817
rect 6801 1783 6835 1817
rect 6869 1783 6903 1817
rect 6937 1783 6971 1817
rect 7005 1783 7039 1817
rect 7073 1783 7107 1817
rect 7141 1783 7175 1817
rect 7209 1783 7243 1817
rect 7277 1783 7311 1817
rect 7345 1783 7379 1817
rect 7413 1783 7447 1817
rect 7481 1783 7515 1817
rect 7549 1783 7583 1817
rect 7617 1783 7651 1817
rect 7685 1783 7719 1817
rect 7753 1783 7787 1817
rect 7821 1783 7855 1817
rect 7889 1783 7923 1817
rect 7957 1783 7991 1817
rect 8025 1783 8059 1817
rect 8093 1783 8240 1817
rect 160 1760 8240 1783
<< psubdiffcont >>
rect 137 5943 171 5977
rect 205 5943 239 5977
rect 273 5943 307 5977
rect 341 5943 375 5977
rect 409 5943 443 5977
rect 477 5943 511 5977
rect 545 5943 579 5977
rect 613 5943 647 5977
rect 681 5943 715 5977
rect 749 5943 783 5977
rect 817 5943 851 5977
rect 885 5943 919 5977
rect 953 5943 987 5977
rect 1021 5943 1055 5977
rect 1089 5943 1123 5977
rect 1157 5943 1191 5977
rect 1225 5943 1259 5977
rect 1293 5943 1327 5977
rect 1361 5943 1395 5977
rect 1429 5943 1463 5977
rect 1497 5943 1531 5977
rect 1565 5943 1599 5977
rect 1633 5943 1667 5977
rect 1701 5943 1735 5977
rect 1769 5943 1803 5977
rect 1837 5943 1871 5977
rect 1905 5943 1939 5977
rect 1973 5943 2007 5977
rect 2041 5943 2075 5977
rect 2109 5943 2143 5977
rect 2177 5943 2211 5977
rect 2245 5943 2279 5977
rect 2313 5943 2347 5977
rect 2381 5943 2415 5977
rect 2449 5943 2483 5977
rect 2517 5943 2551 5977
rect 2585 5943 2619 5977
rect 2653 5943 2687 5977
rect 2721 5943 2755 5977
rect 2789 5943 2823 5977
rect 2857 5943 2891 5977
rect 2925 5943 2959 5977
rect 2993 5943 3027 5977
rect 3061 5943 3095 5977
rect 3129 5943 3163 5977
rect 3197 5943 3231 5977
rect 3265 5943 3299 5977
rect 3333 5943 3367 5977
rect 3401 5943 3435 5977
rect 3469 5943 3503 5977
rect 3537 5943 3571 5977
rect 3605 5943 3639 5977
rect 3673 5943 3707 5977
rect 3741 5943 3775 5977
rect 3809 5943 3843 5977
rect 3877 5943 3911 5977
rect 3945 5943 3979 5977
rect 4013 5943 4047 5977
rect 4081 5943 4115 5977
rect 4149 5943 4183 5977
rect 4217 5943 4251 5977
rect 4285 5943 4319 5977
rect 4353 5943 4387 5977
rect 4421 5943 4455 5977
rect 4489 5943 4523 5977
rect 4557 5943 4591 5977
rect 4625 5943 4659 5977
rect 4693 5943 4727 5977
rect 4761 5943 4795 5977
rect 4829 5943 4863 5977
rect 4897 5943 4931 5977
rect 4965 5943 4999 5977
rect 5033 5943 5067 5977
rect 5101 5943 5135 5977
rect 5169 5943 5203 5977
rect 5237 5943 5271 5977
rect 5305 5943 5339 5977
rect 5373 5943 5407 5977
rect 5441 5943 5475 5977
rect 5509 5943 5543 5977
rect 5577 5943 5611 5977
rect 5645 5943 5679 5977
rect 5713 5943 5747 5977
rect 5781 5943 5815 5977
rect 5849 5943 5883 5977
rect 5917 5943 5951 5977
rect 5985 5943 6019 5977
rect 6053 5943 6087 5977
rect 6121 5943 6155 5977
rect 6189 5943 6223 5977
rect 6257 5943 6291 5977
rect 6325 5943 6359 5977
rect 6393 5943 6427 5977
rect 6461 5943 6495 5977
rect 6529 5943 6563 5977
rect 6597 5943 6631 5977
rect 6665 5943 6699 5977
rect 6733 5943 6767 5977
rect 6801 5943 6835 5977
rect 6869 5943 6903 5977
rect 6937 5943 6971 5977
rect 7005 5943 7039 5977
rect 7073 5943 7107 5977
rect 7141 5943 7175 5977
rect 7209 5943 7243 5977
rect 7277 5943 7311 5977
rect 7345 5943 7379 5977
rect 7413 5943 7447 5977
rect 7481 5943 7515 5977
rect 7549 5943 7583 5977
rect 7617 5943 7651 5977
rect 7685 5943 7719 5977
rect 7753 5943 7787 5977
rect 7821 5943 7855 5977
rect 7889 5943 7923 5977
rect 7957 5943 7991 5977
rect 8025 5943 8059 5977
rect 8093 5943 8127 5977
rect 8161 5943 8195 5977
rect 8229 5943 8263 5977
rect 23 5821 57 5855
rect 23 5753 57 5787
rect 23 5685 57 5719
rect 23 5617 57 5651
rect 23 5549 57 5583
rect 23 5481 57 5515
rect 23 5413 57 5447
rect 23 5345 57 5379
rect 23 5277 57 5311
rect 23 5209 57 5243
rect 23 5141 57 5175
rect 23 5073 57 5107
rect 23 5005 57 5039
rect 23 4937 57 4971
rect 23 4869 57 4903
rect 23 4801 57 4835
rect 23 4733 57 4767
rect 23 4665 57 4699
rect 23 4597 57 4631
rect 23 4529 57 4563
rect 23 4461 57 4495
rect 23 4393 57 4427
rect 23 4325 57 4359
rect 23 4257 57 4291
rect 23 4189 57 4223
rect 23 4121 57 4155
rect 23 4053 57 4087
rect 23 3985 57 4019
rect 8343 5821 8377 5855
rect 8343 5753 8377 5787
rect 8343 5685 8377 5719
rect 8343 5617 8377 5651
rect 8343 5549 8377 5583
rect 8343 5481 8377 5515
rect 8343 5413 8377 5447
rect 8343 5345 8377 5379
rect 8343 5277 8377 5311
rect 8343 5209 8377 5243
rect 8343 5141 8377 5175
rect 8343 5073 8377 5107
rect 8343 5005 8377 5039
rect 8343 4937 8377 4971
rect 8343 4869 8377 4903
rect 8343 4801 8377 4835
rect 8343 4733 8377 4767
rect 8343 4665 8377 4699
rect 8343 4597 8377 4631
rect 8343 4529 8377 4563
rect 8343 4461 8377 4495
rect 8343 4393 8377 4427
rect 8343 4325 8377 4359
rect 8343 4257 8377 4291
rect 8343 4189 8377 4223
rect 8343 4121 8377 4155
rect 8343 4053 8377 4087
rect 8343 3985 8377 4019
rect 151 3863 185 3897
rect 219 3863 253 3897
rect 287 3863 321 3897
rect 355 3863 389 3897
rect 423 3863 457 3897
rect 491 3863 525 3897
rect 559 3863 593 3897
rect 627 3863 661 3897
rect 695 3863 729 3897
rect 763 3863 797 3897
rect 831 3863 865 3897
rect 899 3863 933 3897
rect 967 3863 1001 3897
rect 1035 3863 1069 3897
rect 1103 3863 1137 3897
rect 1171 3863 1205 3897
rect 1239 3863 1273 3897
rect 1307 3863 1341 3897
rect 1375 3863 1409 3897
rect 1443 3863 1477 3897
rect 1511 3863 1545 3897
rect 1579 3863 1613 3897
rect 1647 3863 1681 3897
rect 1715 3863 1749 3897
rect 1783 3863 1817 3897
rect 1851 3863 1885 3897
rect 1919 3863 1953 3897
rect 1987 3863 2021 3897
rect 2055 3863 2089 3897
rect 2123 3863 2157 3897
rect 2191 3863 2225 3897
rect 2259 3863 2293 3897
rect 2327 3863 2361 3897
rect 2395 3863 2429 3897
rect 2463 3863 2497 3897
rect 2531 3863 2565 3897
rect 2599 3863 2633 3897
rect 2667 3863 2701 3897
rect 2735 3863 2769 3897
rect 2803 3863 2837 3897
rect 2871 3863 2905 3897
rect 2939 3863 2973 3897
rect 3007 3863 3041 3897
rect 3075 3863 3109 3897
rect 3143 3863 3177 3897
rect 3211 3863 3245 3897
rect 3279 3863 3313 3897
rect 3347 3863 3381 3897
rect 3415 3863 3449 3897
rect 3483 3863 3517 3897
rect 3551 3863 3585 3897
rect 3619 3863 3653 3897
rect 3687 3863 3721 3897
rect 3755 3863 3789 3897
rect 3823 3863 3857 3897
rect 3891 3863 3925 3897
rect 3959 3863 3993 3897
rect 4027 3863 4061 3897
rect 4095 3863 4129 3897
rect 4163 3863 4197 3897
rect 4231 3863 4265 3897
rect 4299 3863 4333 3897
rect 4367 3863 4401 3897
rect 4435 3863 4469 3897
rect 4503 3863 4537 3897
rect 4571 3863 4605 3897
rect 4639 3863 4673 3897
rect 4707 3863 4741 3897
rect 4775 3863 4809 3897
rect 4843 3863 4877 3897
rect 4911 3863 4945 3897
rect 4979 3863 5013 3897
rect 5047 3863 5081 3897
rect 5115 3863 5149 3897
rect 5183 3863 5217 3897
rect 5251 3863 5285 3897
rect 5319 3863 5353 3897
rect 5387 3863 5421 3897
rect 5455 3863 5489 3897
rect 5523 3863 5557 3897
rect 5591 3863 5625 3897
rect 5659 3863 5693 3897
rect 5727 3863 5761 3897
rect 5795 3863 5829 3897
rect 5863 3863 5897 3897
rect 5931 3863 5965 3897
rect 5999 3863 6033 3897
rect 6067 3863 6101 3897
rect 6135 3863 6169 3897
rect 6203 3863 6237 3897
rect 6271 3863 6305 3897
rect 6339 3863 6373 3897
rect 6407 3863 6441 3897
rect 6475 3863 6509 3897
rect 6543 3863 6577 3897
rect 6611 3863 6645 3897
rect 6679 3863 6713 3897
rect 6747 3863 6781 3897
rect 6815 3863 6849 3897
rect 6883 3863 6917 3897
rect 6951 3863 6985 3897
rect 7019 3863 7053 3897
rect 7087 3863 7121 3897
rect 7155 3863 7189 3897
rect 7223 3863 7257 3897
rect 7291 3863 7325 3897
rect 7359 3863 7393 3897
rect 7427 3863 7461 3897
rect 7495 3863 7529 3897
rect 7563 3863 7597 3897
rect 7631 3863 7665 3897
rect 7699 3863 7733 3897
rect 7767 3863 7801 3897
rect 7835 3863 7869 3897
rect 7903 3863 7937 3897
rect 7971 3863 8005 3897
rect 8039 3863 8073 3897
rect 8107 3863 8141 3897
rect 8175 3863 8209 3897
rect 151 3703 185 3737
rect 219 3703 253 3737
rect 287 3703 321 3737
rect 355 3703 389 3737
rect 423 3703 457 3737
rect 491 3703 525 3737
rect 559 3703 593 3737
rect 627 3703 661 3737
rect 695 3703 729 3737
rect 763 3703 797 3737
rect 831 3703 865 3737
rect 899 3703 933 3737
rect 967 3703 1001 3737
rect 1035 3703 1069 3737
rect 1103 3703 1137 3737
rect 1171 3703 1205 3737
rect 1239 3703 1273 3737
rect 1307 3703 1341 3737
rect 1375 3703 1409 3737
rect 1443 3703 1477 3737
rect 1511 3703 1545 3737
rect 1579 3703 1613 3737
rect 1647 3703 1681 3737
rect 1715 3703 1749 3737
rect 1783 3703 1817 3737
rect 1851 3703 1885 3737
rect 1919 3703 1953 3737
rect 1987 3703 2021 3737
rect 2055 3703 2089 3737
rect 2123 3703 2157 3737
rect 2191 3703 2225 3737
rect 2259 3703 2293 3737
rect 2327 3703 2361 3737
rect 2395 3703 2429 3737
rect 2463 3703 2497 3737
rect 2531 3703 2565 3737
rect 2599 3703 2633 3737
rect 2667 3703 2701 3737
rect 2735 3703 2769 3737
rect 2803 3703 2837 3737
rect 2871 3703 2905 3737
rect 2939 3703 2973 3737
rect 3007 3703 3041 3737
rect 3075 3703 3109 3737
rect 3143 3703 3177 3737
rect 3211 3703 3245 3737
rect 3279 3703 3313 3737
rect 3347 3703 3381 3737
rect 3415 3703 3449 3737
rect 3483 3703 3517 3737
rect 3551 3703 3585 3737
rect 3619 3703 3653 3737
rect 3687 3703 3721 3737
rect 3755 3703 3789 3737
rect 3823 3703 3857 3737
rect 3891 3703 3925 3737
rect 3959 3703 3993 3737
rect 4027 3703 4061 3737
rect 4095 3703 4129 3737
rect 4163 3703 4197 3737
rect 4231 3703 4265 3737
rect 4299 3703 4333 3737
rect 4367 3703 4401 3737
rect 4435 3703 4469 3737
rect 4503 3703 4537 3737
rect 4571 3703 4605 3737
rect 4639 3703 4673 3737
rect 4707 3703 4741 3737
rect 4775 3703 4809 3737
rect 4843 3703 4877 3737
rect 4911 3703 4945 3737
rect 4979 3703 5013 3737
rect 5047 3703 5081 3737
rect 5115 3703 5149 3737
rect 5183 3703 5217 3737
rect 5251 3703 5285 3737
rect 5319 3703 5353 3737
rect 5387 3703 5421 3737
rect 5455 3703 5489 3737
rect 5523 3703 5557 3737
rect 5591 3703 5625 3737
rect 5659 3703 5693 3737
rect 5727 3703 5761 3737
rect 5795 3703 5829 3737
rect 5863 3703 5897 3737
rect 5931 3703 5965 3737
rect 5999 3703 6033 3737
rect 6067 3703 6101 3737
rect 6135 3703 6169 3737
rect 6203 3703 6237 3737
rect 6271 3703 6305 3737
rect 6339 3703 6373 3737
rect 6407 3703 6441 3737
rect 6475 3703 6509 3737
rect 6543 3703 6577 3737
rect 6611 3703 6645 3737
rect 6679 3703 6713 3737
rect 6747 3703 6781 3737
rect 6815 3703 6849 3737
rect 6883 3703 6917 3737
rect 6951 3703 6985 3737
rect 7019 3703 7053 3737
rect 7087 3703 7121 3737
rect 7155 3703 7189 3737
rect 7223 3703 7257 3737
rect 7291 3703 7325 3737
rect 7359 3703 7393 3737
rect 7427 3703 7461 3737
rect 7495 3703 7529 3737
rect 7563 3703 7597 3737
rect 7631 3703 7665 3737
rect 7699 3703 7733 3737
rect 7767 3703 7801 3737
rect 7835 3703 7869 3737
rect 7903 3703 7937 3737
rect 7971 3703 8005 3737
rect 8039 3703 8073 3737
rect 8107 3703 8141 3737
rect 8175 3703 8209 3737
rect 23 3581 57 3615
rect 23 3513 57 3547
rect 23 3445 57 3479
rect 23 3377 57 3411
rect 23 3309 57 3343
rect 23 3241 57 3275
rect 23 3173 57 3207
rect 23 3105 57 3139
rect 23 3037 57 3071
rect 23 2969 57 3003
rect 23 2901 57 2935
rect 23 2833 57 2867
rect 23 2765 57 2799
rect 23 2697 57 2731
rect 23 2629 57 2663
rect 23 2561 57 2595
rect 23 2493 57 2527
rect 23 2425 57 2459
rect 23 2357 57 2391
rect 23 2289 57 2323
rect 23 2221 57 2255
rect 23 2153 57 2187
rect 23 2085 57 2119
rect 23 2017 57 2051
rect 23 1949 57 1983
rect 23 1881 57 1915
rect 23 1813 57 1847
rect 23 1745 57 1779
rect 8343 3581 8377 3615
rect 8343 3513 8377 3547
rect 8343 3445 8377 3479
rect 8343 3377 8377 3411
rect 8343 3309 8377 3343
rect 8343 3241 8377 3275
rect 8343 3173 8377 3207
rect 8343 3105 8377 3139
rect 8343 3037 8377 3071
rect 8343 2969 8377 3003
rect 8343 2901 8377 2935
rect 8343 2833 8377 2867
rect 8343 2765 8377 2799
rect 8343 2697 8377 2731
rect 8343 2629 8377 2663
rect 8343 2561 8377 2595
rect 8343 2493 8377 2527
rect 8343 2425 8377 2459
rect 8343 2357 8377 2391
rect 8343 2289 8377 2323
rect 8343 2221 8377 2255
rect 8343 2153 8377 2187
rect 8343 2085 8377 2119
rect 8343 2017 8377 2051
rect 8343 1949 8377 1983
rect 8343 1881 8377 1915
rect 8343 1813 8377 1847
rect 8343 1745 8377 1779
rect 137 1623 171 1657
rect 205 1623 239 1657
rect 273 1623 307 1657
rect 341 1623 375 1657
rect 409 1623 443 1657
rect 477 1623 511 1657
rect 545 1623 579 1657
rect 613 1623 647 1657
rect 681 1623 715 1657
rect 749 1623 783 1657
rect 817 1623 851 1657
rect 885 1623 919 1657
rect 953 1623 987 1657
rect 1021 1623 1055 1657
rect 1089 1623 1123 1657
rect 1157 1623 1191 1657
rect 1225 1623 1259 1657
rect 1293 1623 1327 1657
rect 1361 1623 1395 1657
rect 1429 1623 1463 1657
rect 1497 1623 1531 1657
rect 1565 1623 1599 1657
rect 1633 1623 1667 1657
rect 1701 1623 1735 1657
rect 1769 1623 1803 1657
rect 1837 1623 1871 1657
rect 1905 1623 1939 1657
rect 1973 1623 2007 1657
rect 2041 1623 2075 1657
rect 2109 1623 2143 1657
rect 2177 1623 2211 1657
rect 2245 1623 2279 1657
rect 2313 1623 2347 1657
rect 2381 1623 2415 1657
rect 2449 1623 2483 1657
rect 2517 1623 2551 1657
rect 2585 1623 2619 1657
rect 2653 1623 2687 1657
rect 2721 1623 2755 1657
rect 2789 1623 2823 1657
rect 2857 1623 2891 1657
rect 2925 1623 2959 1657
rect 2993 1623 3027 1657
rect 3061 1623 3095 1657
rect 3129 1623 3163 1657
rect 3197 1623 3231 1657
rect 3265 1623 3299 1657
rect 3333 1623 3367 1657
rect 3401 1623 3435 1657
rect 3469 1623 3503 1657
rect 3537 1623 3571 1657
rect 3605 1623 3639 1657
rect 3673 1623 3707 1657
rect 3741 1623 3775 1657
rect 3809 1623 3843 1657
rect 3877 1623 3911 1657
rect 3945 1623 3979 1657
rect 4013 1623 4047 1657
rect 4081 1623 4115 1657
rect 4149 1623 4183 1657
rect 4217 1623 4251 1657
rect 4285 1623 4319 1657
rect 4353 1623 4387 1657
rect 4421 1623 4455 1657
rect 4489 1623 4523 1657
rect 4557 1623 4591 1657
rect 4625 1623 4659 1657
rect 4693 1623 4727 1657
rect 4761 1623 4795 1657
rect 4829 1623 4863 1657
rect 4897 1623 4931 1657
rect 4965 1623 4999 1657
rect 5033 1623 5067 1657
rect 5101 1623 5135 1657
rect 5169 1623 5203 1657
rect 5237 1623 5271 1657
rect 5305 1623 5339 1657
rect 5373 1623 5407 1657
rect 5441 1623 5475 1657
rect 5509 1623 5543 1657
rect 5577 1623 5611 1657
rect 5645 1623 5679 1657
rect 5713 1623 5747 1657
rect 5781 1623 5815 1657
rect 5849 1623 5883 1657
rect 5917 1623 5951 1657
rect 5985 1623 6019 1657
rect 6053 1623 6087 1657
rect 6121 1623 6155 1657
rect 6189 1623 6223 1657
rect 6257 1623 6291 1657
rect 6325 1623 6359 1657
rect 6393 1623 6427 1657
rect 6461 1623 6495 1657
rect 6529 1623 6563 1657
rect 6597 1623 6631 1657
rect 6665 1623 6699 1657
rect 6733 1623 6767 1657
rect 6801 1623 6835 1657
rect 6869 1623 6903 1657
rect 6937 1623 6971 1657
rect 7005 1623 7039 1657
rect 7073 1623 7107 1657
rect 7141 1623 7175 1657
rect 7209 1623 7243 1657
rect 7277 1623 7311 1657
rect 7345 1623 7379 1657
rect 7413 1623 7447 1657
rect 7481 1623 7515 1657
rect 7549 1623 7583 1657
rect 7617 1623 7651 1657
rect 7685 1623 7719 1657
rect 7753 1623 7787 1657
rect 7821 1623 7855 1657
rect 7889 1623 7923 1657
rect 7957 1623 7991 1657
rect 8025 1623 8059 1657
rect 8093 1623 8127 1657
rect 8161 1623 8195 1657
rect 8229 1623 8263 1657
rect 137 983 171 1017
rect 205 983 239 1017
rect 273 983 307 1017
rect 341 983 375 1017
rect 409 983 443 1017
rect 477 983 511 1017
rect 545 983 579 1017
rect 613 983 647 1017
rect 681 983 715 1017
rect 749 983 783 1017
rect 817 983 851 1017
rect 885 983 919 1017
rect 953 983 987 1017
rect 1021 983 1055 1017
rect 1089 983 1123 1017
rect 1157 983 1191 1017
rect 1225 983 1259 1017
rect 1293 983 1327 1017
rect 1361 983 1395 1017
rect 1429 983 1463 1017
rect 1497 983 1531 1017
rect 1565 983 1599 1017
rect 1633 983 1667 1017
rect 1701 983 1735 1017
rect 1769 983 1803 1017
rect 1837 983 1871 1017
rect 1905 983 1939 1017
rect 1973 983 2007 1017
rect 2041 983 2075 1017
rect 2109 983 2143 1017
rect 2177 983 2211 1017
rect 2245 983 2279 1017
rect 2313 983 2347 1017
rect 2381 983 2415 1017
rect 2449 983 2483 1017
rect 2517 983 2551 1017
rect 2585 983 2619 1017
rect 2653 983 2687 1017
rect 2721 983 2755 1017
rect 2789 983 2823 1017
rect 2857 983 2891 1017
rect 2925 983 2959 1017
rect 2993 983 3027 1017
rect 3061 983 3095 1017
rect 3129 983 3163 1017
rect 3197 983 3231 1017
rect 3265 983 3299 1017
rect 3333 983 3367 1017
rect 3401 983 3435 1017
rect 3469 983 3503 1017
rect 3537 983 3571 1017
rect 3605 983 3639 1017
rect 3673 983 3707 1017
rect 3741 983 3775 1017
rect 3809 983 3843 1017
rect 3877 983 3911 1017
rect 3945 983 3979 1017
rect 4013 983 4047 1017
rect 4081 983 4115 1017
rect 4149 983 4183 1017
rect 4217 983 4251 1017
rect 4285 983 4319 1017
rect 4353 983 4387 1017
rect 4421 983 4455 1017
rect 4489 983 4523 1017
rect 4557 983 4591 1017
rect 4625 983 4659 1017
rect 4693 983 4727 1017
rect 4761 983 4795 1017
rect 4829 983 4863 1017
rect 4897 983 4931 1017
rect 4965 983 4999 1017
rect 5033 983 5067 1017
rect 5101 983 5135 1017
rect 5169 983 5203 1017
rect 5237 983 5271 1017
rect 5305 983 5339 1017
rect 5373 983 5407 1017
rect 5441 983 5475 1017
rect 5509 983 5543 1017
rect 5577 983 5611 1017
rect 5645 983 5679 1017
rect 5713 983 5747 1017
rect 5781 983 5815 1017
rect 5849 983 5883 1017
rect 5917 983 5951 1017
rect 5985 983 6019 1017
rect 6053 983 6087 1017
rect 6121 983 6155 1017
rect 6189 983 6223 1017
rect 6257 983 6291 1017
rect 6325 983 6359 1017
rect 6393 983 6427 1017
rect 6461 983 6495 1017
rect 6529 983 6563 1017
rect 6597 983 6631 1017
rect 6665 983 6699 1017
rect 6733 983 6767 1017
rect 6801 983 6835 1017
rect 6869 983 6903 1017
rect 6937 983 6971 1017
rect 7005 983 7039 1017
rect 7073 983 7107 1017
rect 7141 983 7175 1017
rect 7209 983 7243 1017
rect 7277 983 7311 1017
rect 7345 983 7379 1017
rect 7413 983 7447 1017
rect 7481 983 7515 1017
rect 7549 983 7583 1017
rect 7617 983 7651 1017
rect 7685 983 7719 1017
rect 7753 983 7787 1017
rect 7821 983 7855 1017
rect 7889 983 7923 1017
rect 7957 983 7991 1017
rect 8025 983 8059 1017
rect 8093 983 8127 1017
rect 8161 983 8195 1017
rect 8229 983 8263 1017
rect 23 877 57 911
rect 23 809 57 843
rect 23 741 57 775
rect 8343 877 8377 911
rect 8343 809 8377 843
rect 23 673 57 707
rect 23 605 57 639
rect 23 537 57 571
rect 8343 741 8377 775
rect 8343 673 8377 707
rect 8343 605 8377 639
rect 23 469 57 503
rect 23 401 57 435
rect 23 333 57 367
rect 8343 537 8377 571
rect 8343 469 8377 503
rect 8343 401 8377 435
rect 23 265 57 299
rect 23 197 57 231
rect 23 129 57 163
rect 8343 333 8377 367
rect 8343 265 8377 299
rect 8343 197 8377 231
rect 8343 129 8377 163
rect 137 23 171 57
rect 205 23 239 57
rect 273 23 307 57
rect 341 23 375 57
rect 409 23 443 57
rect 477 23 511 57
rect 545 23 579 57
rect 613 23 647 57
rect 681 23 715 57
rect 749 23 783 57
rect 817 23 851 57
rect 885 23 919 57
rect 953 23 987 57
rect 1021 23 1055 57
rect 1089 23 1123 57
rect 1157 23 1191 57
rect 1225 23 1259 57
rect 1293 23 1327 57
rect 1361 23 1395 57
rect 1429 23 1463 57
rect 1497 23 1531 57
rect 1565 23 1599 57
rect 1633 23 1667 57
rect 1701 23 1735 57
rect 1769 23 1803 57
rect 1837 23 1871 57
rect 1905 23 1939 57
rect 1973 23 2007 57
rect 2041 23 2075 57
rect 2109 23 2143 57
rect 2177 23 2211 57
rect 2245 23 2279 57
rect 2313 23 2347 57
rect 2381 23 2415 57
rect 2449 23 2483 57
rect 2517 23 2551 57
rect 2585 23 2619 57
rect 2653 23 2687 57
rect 2721 23 2755 57
rect 2789 23 2823 57
rect 2857 23 2891 57
rect 2925 23 2959 57
rect 2993 23 3027 57
rect 3061 23 3095 57
rect 3129 23 3163 57
rect 3197 23 3231 57
rect 3265 23 3299 57
rect 3333 23 3367 57
rect 3401 23 3435 57
rect 3469 23 3503 57
rect 3537 23 3571 57
rect 3605 23 3639 57
rect 3673 23 3707 57
rect 3741 23 3775 57
rect 3809 23 3843 57
rect 3877 23 3911 57
rect 3945 23 3979 57
rect 4013 23 4047 57
rect 4081 23 4115 57
rect 4149 23 4183 57
rect 4217 23 4251 57
rect 4285 23 4319 57
rect 4353 23 4387 57
rect 4421 23 4455 57
rect 4489 23 4523 57
rect 4557 23 4591 57
rect 4625 23 4659 57
rect 4693 23 4727 57
rect 4761 23 4795 57
rect 4829 23 4863 57
rect 4897 23 4931 57
rect 4965 23 4999 57
rect 5033 23 5067 57
rect 5101 23 5135 57
rect 5169 23 5203 57
rect 5237 23 5271 57
rect 5305 23 5339 57
rect 5373 23 5407 57
rect 5441 23 5475 57
rect 5509 23 5543 57
rect 5577 23 5611 57
rect 5645 23 5679 57
rect 5713 23 5747 57
rect 5781 23 5815 57
rect 5849 23 5883 57
rect 5917 23 5951 57
rect 5985 23 6019 57
rect 6053 23 6087 57
rect 6121 23 6155 57
rect 6189 23 6223 57
rect 6257 23 6291 57
rect 6325 23 6359 57
rect 6393 23 6427 57
rect 6461 23 6495 57
rect 6529 23 6563 57
rect 6597 23 6631 57
rect 6665 23 6699 57
rect 6733 23 6767 57
rect 6801 23 6835 57
rect 6869 23 6903 57
rect 6937 23 6971 57
rect 7005 23 7039 57
rect 7073 23 7107 57
rect 7141 23 7175 57
rect 7209 23 7243 57
rect 7277 23 7311 57
rect 7345 23 7379 57
rect 7413 23 7447 57
rect 7481 23 7515 57
rect 7549 23 7583 57
rect 7617 23 7651 57
rect 7685 23 7719 57
rect 7753 23 7787 57
rect 7821 23 7855 57
rect 7889 23 7923 57
rect 7957 23 7991 57
rect 8025 23 8059 57
rect 8093 23 8127 57
rect 8161 23 8195 57
rect 8229 23 8263 57
<< mvnsubdiffcont >>
rect 307 5783 341 5817
rect 375 5783 409 5817
rect 443 5783 477 5817
rect 511 5783 545 5817
rect 579 5783 613 5817
rect 647 5783 681 5817
rect 715 5783 749 5817
rect 783 5783 817 5817
rect 851 5783 885 5817
rect 919 5783 953 5817
rect 987 5783 1021 5817
rect 1055 5783 1089 5817
rect 1123 5783 1157 5817
rect 1191 5783 1225 5817
rect 1259 5783 1293 5817
rect 1327 5783 1361 5817
rect 1395 5783 1429 5817
rect 1463 5783 1497 5817
rect 1531 5783 1565 5817
rect 1599 5783 1633 5817
rect 1667 5783 1701 5817
rect 1735 5783 1769 5817
rect 1803 5783 1837 5817
rect 1871 5783 1905 5817
rect 1939 5783 1973 5817
rect 2007 5783 2041 5817
rect 2075 5783 2109 5817
rect 2143 5783 2177 5817
rect 2211 5783 2245 5817
rect 2279 5783 2313 5817
rect 2347 5783 2381 5817
rect 2415 5783 2449 5817
rect 2483 5783 2517 5817
rect 2551 5783 2585 5817
rect 2619 5783 2653 5817
rect 2687 5783 2721 5817
rect 2755 5783 2789 5817
rect 2823 5783 2857 5817
rect 2891 5783 2925 5817
rect 2959 5783 2993 5817
rect 3027 5783 3061 5817
rect 3095 5783 3129 5817
rect 3163 5783 3197 5817
rect 3231 5783 3265 5817
rect 3299 5783 3333 5817
rect 3367 5783 3401 5817
rect 3435 5783 3469 5817
rect 3503 5783 3537 5817
rect 3571 5783 3605 5817
rect 3639 5783 3673 5817
rect 3707 5783 3741 5817
rect 3775 5783 3809 5817
rect 3843 5783 3877 5817
rect 3911 5783 3945 5817
rect 3979 5783 4013 5817
rect 4047 5783 4081 5817
rect 4115 5783 4149 5817
rect 4183 5783 4217 5817
rect 4251 5783 4285 5817
rect 4319 5783 4353 5817
rect 4387 5783 4421 5817
rect 4455 5783 4489 5817
rect 4523 5783 4557 5817
rect 4591 5783 4625 5817
rect 4659 5783 4693 5817
rect 4727 5783 4761 5817
rect 4795 5783 4829 5817
rect 4863 5783 4897 5817
rect 4931 5783 4965 5817
rect 4999 5783 5033 5817
rect 5067 5783 5101 5817
rect 5135 5783 5169 5817
rect 5203 5783 5237 5817
rect 5271 5783 5305 5817
rect 5339 5783 5373 5817
rect 5407 5783 5441 5817
rect 5475 5783 5509 5817
rect 5543 5783 5577 5817
rect 5611 5783 5645 5817
rect 5679 5783 5713 5817
rect 5747 5783 5781 5817
rect 5815 5783 5849 5817
rect 5883 5783 5917 5817
rect 5951 5783 5985 5817
rect 6019 5783 6053 5817
rect 6087 5783 6121 5817
rect 6155 5783 6189 5817
rect 6223 5783 6257 5817
rect 6291 5783 6325 5817
rect 6359 5783 6393 5817
rect 6427 5783 6461 5817
rect 6495 5783 6529 5817
rect 6563 5783 6597 5817
rect 6631 5783 6665 5817
rect 6699 5783 6733 5817
rect 6767 5783 6801 5817
rect 6835 5783 6869 5817
rect 6903 5783 6937 5817
rect 6971 5783 7005 5817
rect 7039 5783 7073 5817
rect 7107 5783 7141 5817
rect 7175 5783 7209 5817
rect 7243 5783 7277 5817
rect 7311 5783 7345 5817
rect 7379 5783 7413 5817
rect 7447 5783 7481 5817
rect 7515 5783 7549 5817
rect 7583 5783 7617 5817
rect 7651 5783 7685 5817
rect 7719 5783 7753 5817
rect 7787 5783 7821 5817
rect 7855 5783 7889 5817
rect 7923 5783 7957 5817
rect 7991 5783 8025 5817
rect 8059 5783 8093 5817
rect 183 5685 217 5719
rect 8183 5685 8217 5719
rect 183 5617 217 5651
rect 183 5549 217 5583
rect 183 5481 217 5515
rect 183 5413 217 5447
rect 183 5345 217 5379
rect 183 5277 217 5311
rect 183 5209 217 5243
rect 183 5141 217 5175
rect 183 5073 217 5107
rect 8183 5617 8217 5651
rect 8183 5549 8217 5583
rect 8183 5481 8217 5515
rect 8183 5413 8217 5447
rect 8183 5345 8217 5379
rect 8183 5277 8217 5311
rect 8183 5209 8217 5243
rect 8183 5141 8217 5175
rect 183 5005 217 5039
rect 183 4937 217 4971
rect 8183 5073 8217 5107
rect 8183 5005 8217 5039
rect 8183 4937 8217 4971
rect 183 4869 217 4903
rect 183 4801 217 4835
rect 183 4733 217 4767
rect 183 4665 217 4699
rect 183 4597 217 4631
rect 183 4529 217 4563
rect 183 4461 217 4495
rect 183 4393 217 4427
rect 183 4325 217 4359
rect 8183 4869 8217 4903
rect 8183 4801 8217 4835
rect 8183 4733 8217 4767
rect 8183 4665 8217 4699
rect 8183 4597 8217 4631
rect 8183 4529 8217 4563
rect 8183 4461 8217 4495
rect 8183 4393 8217 4427
rect 8183 4325 8217 4359
rect 183 4257 217 4291
rect 183 4189 217 4223
rect 8183 4257 8217 4291
rect 8183 4189 8217 4223
rect 183 4121 217 4155
rect 8183 4121 8217 4155
rect 307 4023 341 4057
rect 375 4023 409 4057
rect 443 4023 477 4057
rect 511 4023 545 4057
rect 579 4023 613 4057
rect 647 4023 681 4057
rect 715 4023 749 4057
rect 783 4023 817 4057
rect 851 4023 885 4057
rect 919 4023 953 4057
rect 987 4023 1021 4057
rect 1055 4023 1089 4057
rect 1123 4023 1157 4057
rect 1191 4023 1225 4057
rect 1259 4023 1293 4057
rect 1327 4023 1361 4057
rect 1395 4023 1429 4057
rect 1463 4023 1497 4057
rect 1531 4023 1565 4057
rect 1599 4023 1633 4057
rect 1667 4023 1701 4057
rect 1735 4023 1769 4057
rect 1803 4023 1837 4057
rect 1871 4023 1905 4057
rect 1939 4023 1973 4057
rect 2007 4023 2041 4057
rect 2075 4023 2109 4057
rect 2143 4023 2177 4057
rect 2211 4023 2245 4057
rect 2279 4023 2313 4057
rect 2347 4023 2381 4057
rect 2415 4023 2449 4057
rect 2483 4023 2517 4057
rect 2551 4023 2585 4057
rect 2619 4023 2653 4057
rect 2687 4023 2721 4057
rect 2755 4023 2789 4057
rect 2823 4023 2857 4057
rect 2891 4023 2925 4057
rect 2959 4023 2993 4057
rect 3027 4023 3061 4057
rect 3095 4023 3129 4057
rect 3163 4023 3197 4057
rect 3231 4023 3265 4057
rect 3299 4023 3333 4057
rect 3367 4023 3401 4057
rect 3435 4023 3469 4057
rect 3503 4023 3537 4057
rect 3571 4023 3605 4057
rect 3639 4023 3673 4057
rect 3707 4023 3741 4057
rect 3775 4023 3809 4057
rect 3843 4023 3877 4057
rect 3911 4023 3945 4057
rect 3979 4023 4013 4057
rect 4047 4023 4081 4057
rect 4115 4023 4149 4057
rect 4183 4023 4217 4057
rect 4251 4023 4285 4057
rect 4319 4023 4353 4057
rect 4387 4023 4421 4057
rect 4455 4023 4489 4057
rect 4523 4023 4557 4057
rect 4591 4023 4625 4057
rect 4659 4023 4693 4057
rect 4727 4023 4761 4057
rect 4795 4023 4829 4057
rect 4863 4023 4897 4057
rect 4931 4023 4965 4057
rect 4999 4023 5033 4057
rect 5067 4023 5101 4057
rect 5135 4023 5169 4057
rect 5203 4023 5237 4057
rect 5271 4023 5305 4057
rect 5339 4023 5373 4057
rect 5407 4023 5441 4057
rect 5475 4023 5509 4057
rect 5543 4023 5577 4057
rect 5611 4023 5645 4057
rect 5679 4023 5713 4057
rect 5747 4023 5781 4057
rect 5815 4023 5849 4057
rect 5883 4023 5917 4057
rect 5951 4023 5985 4057
rect 6019 4023 6053 4057
rect 6087 4023 6121 4057
rect 6155 4023 6189 4057
rect 6223 4023 6257 4057
rect 6291 4023 6325 4057
rect 6359 4023 6393 4057
rect 6427 4023 6461 4057
rect 6495 4023 6529 4057
rect 6563 4023 6597 4057
rect 6631 4023 6665 4057
rect 6699 4023 6733 4057
rect 6767 4023 6801 4057
rect 6835 4023 6869 4057
rect 6903 4023 6937 4057
rect 6971 4023 7005 4057
rect 7039 4023 7073 4057
rect 7107 4023 7141 4057
rect 7175 4023 7209 4057
rect 7243 4023 7277 4057
rect 7311 4023 7345 4057
rect 7379 4023 7413 4057
rect 7447 4023 7481 4057
rect 7515 4023 7549 4057
rect 7583 4023 7617 4057
rect 7651 4023 7685 4057
rect 7719 4023 7753 4057
rect 7787 4023 7821 4057
rect 7855 4023 7889 4057
rect 7923 4023 7957 4057
rect 7991 4023 8025 4057
rect 8059 4023 8093 4057
rect 307 3543 341 3577
rect 375 3543 409 3577
rect 443 3543 477 3577
rect 511 3543 545 3577
rect 579 3543 613 3577
rect 647 3543 681 3577
rect 715 3543 749 3577
rect 783 3543 817 3577
rect 851 3543 885 3577
rect 919 3543 953 3577
rect 987 3543 1021 3577
rect 1055 3543 1089 3577
rect 1123 3543 1157 3577
rect 1191 3543 1225 3577
rect 1259 3543 1293 3577
rect 1327 3543 1361 3577
rect 1395 3543 1429 3577
rect 1463 3543 1497 3577
rect 1531 3543 1565 3577
rect 1599 3543 1633 3577
rect 1667 3543 1701 3577
rect 1735 3543 1769 3577
rect 1803 3543 1837 3577
rect 1871 3543 1905 3577
rect 1939 3543 1973 3577
rect 2007 3543 2041 3577
rect 2075 3543 2109 3577
rect 2143 3543 2177 3577
rect 2211 3543 2245 3577
rect 2279 3543 2313 3577
rect 2347 3543 2381 3577
rect 2415 3543 2449 3577
rect 2483 3543 2517 3577
rect 2551 3543 2585 3577
rect 2619 3543 2653 3577
rect 2687 3543 2721 3577
rect 2755 3543 2789 3577
rect 2823 3543 2857 3577
rect 2891 3543 2925 3577
rect 2959 3543 2993 3577
rect 3027 3543 3061 3577
rect 3095 3543 3129 3577
rect 3163 3543 3197 3577
rect 3231 3543 3265 3577
rect 3299 3543 3333 3577
rect 3367 3543 3401 3577
rect 3435 3543 3469 3577
rect 3503 3543 3537 3577
rect 3571 3543 3605 3577
rect 3639 3543 3673 3577
rect 3707 3543 3741 3577
rect 3775 3543 3809 3577
rect 3843 3543 3877 3577
rect 3911 3543 3945 3577
rect 3979 3543 4013 3577
rect 4047 3543 4081 3577
rect 4115 3543 4149 3577
rect 4183 3543 4217 3577
rect 4251 3543 4285 3577
rect 4319 3543 4353 3577
rect 4387 3543 4421 3577
rect 4455 3543 4489 3577
rect 4523 3543 4557 3577
rect 4591 3543 4625 3577
rect 4659 3543 4693 3577
rect 4727 3543 4761 3577
rect 4795 3543 4829 3577
rect 4863 3543 4897 3577
rect 4931 3543 4965 3577
rect 4999 3543 5033 3577
rect 5067 3543 5101 3577
rect 5135 3543 5169 3577
rect 5203 3543 5237 3577
rect 5271 3543 5305 3577
rect 5339 3543 5373 3577
rect 5407 3543 5441 3577
rect 5475 3543 5509 3577
rect 5543 3543 5577 3577
rect 5611 3543 5645 3577
rect 5679 3543 5713 3577
rect 5747 3543 5781 3577
rect 5815 3543 5849 3577
rect 5883 3543 5917 3577
rect 5951 3543 5985 3577
rect 6019 3543 6053 3577
rect 6087 3543 6121 3577
rect 6155 3543 6189 3577
rect 6223 3543 6257 3577
rect 6291 3543 6325 3577
rect 6359 3543 6393 3577
rect 6427 3543 6461 3577
rect 6495 3543 6529 3577
rect 6563 3543 6597 3577
rect 6631 3543 6665 3577
rect 6699 3543 6733 3577
rect 6767 3543 6801 3577
rect 6835 3543 6869 3577
rect 6903 3543 6937 3577
rect 6971 3543 7005 3577
rect 7039 3543 7073 3577
rect 7107 3543 7141 3577
rect 7175 3543 7209 3577
rect 7243 3543 7277 3577
rect 7311 3543 7345 3577
rect 7379 3543 7413 3577
rect 7447 3543 7481 3577
rect 7515 3543 7549 3577
rect 7583 3543 7617 3577
rect 7651 3543 7685 3577
rect 7719 3543 7753 3577
rect 7787 3543 7821 3577
rect 7855 3543 7889 3577
rect 7923 3543 7957 3577
rect 7991 3543 8025 3577
rect 8059 3543 8093 3577
rect 183 3431 217 3465
rect 183 3363 217 3397
rect 183 3295 217 3329
rect 183 3227 217 3261
rect 183 3159 217 3193
rect 183 3091 217 3125
rect 183 3023 217 3057
rect 183 2955 217 2989
rect 183 2887 217 2921
rect 183 2819 217 2853
rect 8183 3431 8217 3465
rect 8183 3363 8217 3397
rect 8183 3295 8217 3329
rect 8183 3227 8217 3261
rect 8183 3159 8217 3193
rect 8183 3091 8217 3125
rect 8183 3023 8217 3057
rect 8183 2955 8217 2989
rect 8183 2887 8217 2921
rect 183 2751 217 2785
rect 183 2683 217 2717
rect 8183 2819 8217 2853
rect 8183 2751 8217 2785
rect 8183 2683 8217 2717
rect 183 2615 217 2649
rect 183 2547 217 2581
rect 183 2479 217 2513
rect 183 2411 217 2445
rect 183 2343 217 2377
rect 183 2275 217 2309
rect 183 2207 217 2241
rect 183 2139 217 2173
rect 183 2071 217 2105
rect 8183 2615 8217 2649
rect 8183 2547 8217 2581
rect 8183 2479 8217 2513
rect 8183 2411 8217 2445
rect 8183 2343 8217 2377
rect 8183 2275 8217 2309
rect 8183 2207 8217 2241
rect 8183 2139 8217 2173
rect 183 2003 217 2037
rect 183 1935 217 1969
rect 8183 2071 8217 2105
rect 8183 2003 8217 2037
rect 8183 1935 8217 1969
rect 307 1783 341 1817
rect 375 1783 409 1817
rect 443 1783 477 1817
rect 511 1783 545 1817
rect 579 1783 613 1817
rect 647 1783 681 1817
rect 715 1783 749 1817
rect 783 1783 817 1817
rect 851 1783 885 1817
rect 919 1783 953 1817
rect 987 1783 1021 1817
rect 1055 1783 1089 1817
rect 1123 1783 1157 1817
rect 1191 1783 1225 1817
rect 1259 1783 1293 1817
rect 1327 1783 1361 1817
rect 1395 1783 1429 1817
rect 1463 1783 1497 1817
rect 1531 1783 1565 1817
rect 1599 1783 1633 1817
rect 1667 1783 1701 1817
rect 1735 1783 1769 1817
rect 1803 1783 1837 1817
rect 1871 1783 1905 1817
rect 1939 1783 1973 1817
rect 2007 1783 2041 1817
rect 2075 1783 2109 1817
rect 2143 1783 2177 1817
rect 2211 1783 2245 1817
rect 2279 1783 2313 1817
rect 2347 1783 2381 1817
rect 2415 1783 2449 1817
rect 2483 1783 2517 1817
rect 2551 1783 2585 1817
rect 2619 1783 2653 1817
rect 2687 1783 2721 1817
rect 2755 1783 2789 1817
rect 2823 1783 2857 1817
rect 2891 1783 2925 1817
rect 2959 1783 2993 1817
rect 3027 1783 3061 1817
rect 3095 1783 3129 1817
rect 3163 1783 3197 1817
rect 3231 1783 3265 1817
rect 3299 1783 3333 1817
rect 3367 1783 3401 1817
rect 3435 1783 3469 1817
rect 3503 1783 3537 1817
rect 3571 1783 3605 1817
rect 3639 1783 3673 1817
rect 3707 1783 3741 1817
rect 3775 1783 3809 1817
rect 3843 1783 3877 1817
rect 3911 1783 3945 1817
rect 3979 1783 4013 1817
rect 4047 1783 4081 1817
rect 4115 1783 4149 1817
rect 4183 1783 4217 1817
rect 4251 1783 4285 1817
rect 4319 1783 4353 1817
rect 4387 1783 4421 1817
rect 4455 1783 4489 1817
rect 4523 1783 4557 1817
rect 4591 1783 4625 1817
rect 4659 1783 4693 1817
rect 4727 1783 4761 1817
rect 4795 1783 4829 1817
rect 4863 1783 4897 1817
rect 4931 1783 4965 1817
rect 4999 1783 5033 1817
rect 5067 1783 5101 1817
rect 5135 1783 5169 1817
rect 5203 1783 5237 1817
rect 5271 1783 5305 1817
rect 5339 1783 5373 1817
rect 5407 1783 5441 1817
rect 5475 1783 5509 1817
rect 5543 1783 5577 1817
rect 5611 1783 5645 1817
rect 5679 1783 5713 1817
rect 5747 1783 5781 1817
rect 5815 1783 5849 1817
rect 5883 1783 5917 1817
rect 5951 1783 5985 1817
rect 6019 1783 6053 1817
rect 6087 1783 6121 1817
rect 6155 1783 6189 1817
rect 6223 1783 6257 1817
rect 6291 1783 6325 1817
rect 6359 1783 6393 1817
rect 6427 1783 6461 1817
rect 6495 1783 6529 1817
rect 6563 1783 6597 1817
rect 6631 1783 6665 1817
rect 6699 1783 6733 1817
rect 6767 1783 6801 1817
rect 6835 1783 6869 1817
rect 6903 1783 6937 1817
rect 6971 1783 7005 1817
rect 7039 1783 7073 1817
rect 7107 1783 7141 1817
rect 7175 1783 7209 1817
rect 7243 1783 7277 1817
rect 7311 1783 7345 1817
rect 7379 1783 7413 1817
rect 7447 1783 7481 1817
rect 7515 1783 7549 1817
rect 7583 1783 7617 1817
rect 7651 1783 7685 1817
rect 7719 1783 7753 1817
rect 7787 1783 7821 1817
rect 7855 1783 7889 1817
rect 7923 1783 7957 1817
rect 7991 1783 8025 1817
rect 8059 1783 8093 1817
<< poly >>
rect 520 5680 2120 5720
rect 2440 5680 4040 5720
rect 4360 5680 5960 5720
rect 6280 5680 7880 5720
rect 520 4920 2120 5080
rect 2440 4920 4040 5080
rect 4360 4920 5960 5080
rect 6280 4920 7880 5080
rect 520 4217 2120 4320
rect 520 4183 555 4217
rect 589 4183 623 4217
rect 657 4183 691 4217
rect 725 4183 759 4217
rect 793 4183 827 4217
rect 861 4183 895 4217
rect 929 4183 963 4217
rect 997 4183 1031 4217
rect 1065 4183 1099 4217
rect 1133 4183 1167 4217
rect 1201 4183 1235 4217
rect 1269 4183 1303 4217
rect 1337 4183 1371 4217
rect 1405 4183 1439 4217
rect 1473 4183 1507 4217
rect 1541 4183 1575 4217
rect 1609 4183 1643 4217
rect 1677 4183 1711 4217
rect 1745 4183 1779 4217
rect 1813 4183 1847 4217
rect 1881 4183 1915 4217
rect 1949 4183 1983 4217
rect 2017 4183 2051 4217
rect 2085 4183 2120 4217
rect 520 4160 2120 4183
rect 2440 4217 4040 4320
rect 2440 4183 2475 4217
rect 2509 4183 2543 4217
rect 2577 4183 2611 4217
rect 2645 4183 2679 4217
rect 2713 4183 2747 4217
rect 2781 4183 2815 4217
rect 2849 4183 2883 4217
rect 2917 4183 2951 4217
rect 2985 4183 3019 4217
rect 3053 4183 3087 4217
rect 3121 4183 3155 4217
rect 3189 4183 3223 4217
rect 3257 4183 3291 4217
rect 3325 4183 3359 4217
rect 3393 4183 3427 4217
rect 3461 4183 3495 4217
rect 3529 4183 3563 4217
rect 3597 4183 3631 4217
rect 3665 4183 3699 4217
rect 3733 4183 3767 4217
rect 3801 4183 3835 4217
rect 3869 4183 3903 4217
rect 3937 4183 3971 4217
rect 4005 4183 4040 4217
rect 2440 4160 4040 4183
rect 4360 4217 5960 4320
rect 4360 4183 4395 4217
rect 4429 4183 4463 4217
rect 4497 4183 4531 4217
rect 4565 4183 4599 4217
rect 4633 4183 4667 4217
rect 4701 4183 4735 4217
rect 4769 4183 4803 4217
rect 4837 4183 4871 4217
rect 4905 4183 4939 4217
rect 4973 4183 5007 4217
rect 5041 4183 5075 4217
rect 5109 4183 5143 4217
rect 5177 4183 5211 4217
rect 5245 4183 5279 4217
rect 5313 4183 5347 4217
rect 5381 4183 5415 4217
rect 5449 4183 5483 4217
rect 5517 4183 5551 4217
rect 5585 4183 5619 4217
rect 5653 4183 5687 4217
rect 5721 4183 5755 4217
rect 5789 4183 5823 4217
rect 5857 4183 5891 4217
rect 5925 4183 5960 4217
rect 4360 4160 5960 4183
rect 6280 4217 7880 4320
rect 6280 4183 6315 4217
rect 6349 4183 6383 4217
rect 6417 4183 6451 4217
rect 6485 4183 6519 4217
rect 6553 4183 6587 4217
rect 6621 4183 6655 4217
rect 6689 4183 6723 4217
rect 6757 4183 6791 4217
rect 6825 4183 6859 4217
rect 6893 4183 6927 4217
rect 6961 4183 6995 4217
rect 7029 4183 7063 4217
rect 7097 4183 7131 4217
rect 7165 4183 7199 4217
rect 7233 4183 7267 4217
rect 7301 4183 7335 4217
rect 7369 4183 7403 4217
rect 7437 4183 7471 4217
rect 7505 4183 7539 4217
rect 7573 4183 7607 4217
rect 7641 4183 7675 4217
rect 7709 4183 7743 4217
rect 7777 4183 7811 4217
rect 7845 4183 7880 4217
rect 6280 4160 7880 4183
rect 520 3440 2120 3480
rect 2440 3440 4040 3480
rect 4360 3440 5960 3480
rect 6280 3440 7880 3480
rect 520 2680 2120 2840
rect 2440 2680 4040 2840
rect 4360 2680 5960 2840
rect 6280 2680 7880 2840
rect 520 1977 2120 2080
rect 520 1943 555 1977
rect 589 1943 623 1977
rect 657 1943 691 1977
rect 725 1943 759 1977
rect 793 1943 827 1977
rect 861 1943 895 1977
rect 929 1943 963 1977
rect 997 1943 1031 1977
rect 1065 1943 1099 1977
rect 1133 1943 1167 1977
rect 1201 1943 1235 1977
rect 1269 1943 1303 1977
rect 1337 1943 1371 1977
rect 1405 1943 1439 1977
rect 1473 1943 1507 1977
rect 1541 1943 1575 1977
rect 1609 1943 1643 1977
rect 1677 1943 1711 1977
rect 1745 1943 1779 1977
rect 1813 1943 1847 1977
rect 1881 1943 1915 1977
rect 1949 1943 1983 1977
rect 2017 1943 2051 1977
rect 2085 1943 2120 1977
rect 520 1920 2120 1943
rect 2440 1977 4040 2080
rect 2440 1943 2475 1977
rect 2509 1943 2543 1977
rect 2577 1943 2611 1977
rect 2645 1943 2679 1977
rect 2713 1943 2747 1977
rect 2781 1943 2815 1977
rect 2849 1943 2883 1977
rect 2917 1943 2951 1977
rect 2985 1943 3019 1977
rect 3053 1943 3087 1977
rect 3121 1943 3155 1977
rect 3189 1943 3223 1977
rect 3257 1943 3291 1977
rect 3325 1943 3359 1977
rect 3393 1943 3427 1977
rect 3461 1943 3495 1977
rect 3529 1943 3563 1977
rect 3597 1943 3631 1977
rect 3665 1943 3699 1977
rect 3733 1943 3767 1977
rect 3801 1943 3835 1977
rect 3869 1943 3903 1977
rect 3937 1943 3971 1977
rect 4005 1943 4040 1977
rect 2440 1920 4040 1943
rect 4360 1977 5960 2080
rect 4360 1943 4395 1977
rect 4429 1943 4463 1977
rect 4497 1943 4531 1977
rect 4565 1943 4599 1977
rect 4633 1943 4667 1977
rect 4701 1943 4735 1977
rect 4769 1943 4803 1977
rect 4837 1943 4871 1977
rect 4905 1943 4939 1977
rect 4973 1943 5007 1977
rect 5041 1943 5075 1977
rect 5109 1943 5143 1977
rect 5177 1943 5211 1977
rect 5245 1943 5279 1977
rect 5313 1943 5347 1977
rect 5381 1943 5415 1977
rect 5449 1943 5483 1977
rect 5517 1943 5551 1977
rect 5585 1943 5619 1977
rect 5653 1943 5687 1977
rect 5721 1943 5755 1977
rect 5789 1943 5823 1977
rect 5857 1943 5891 1977
rect 5925 1943 5960 1977
rect 4360 1920 5960 1943
rect 6280 1977 7880 2080
rect 6280 1943 6315 1977
rect 6349 1943 6383 1977
rect 6417 1943 6451 1977
rect 6485 1943 6519 1977
rect 6553 1943 6587 1977
rect 6621 1943 6655 1977
rect 6689 1943 6723 1977
rect 6757 1943 6791 1977
rect 6825 1943 6859 1977
rect 6893 1943 6927 1977
rect 6961 1943 6995 1977
rect 7029 1943 7063 1977
rect 7097 1943 7131 1977
rect 7165 1943 7199 1977
rect 7233 1943 7267 1977
rect 7301 1943 7335 1977
rect 7369 1943 7403 1977
rect 7437 1943 7471 1977
rect 7505 1943 7539 1977
rect 7573 1943 7607 1977
rect 7641 1943 7675 1977
rect 7709 1943 7743 1977
rect 7777 1943 7811 1977
rect 7845 1943 7880 1977
rect 6280 1920 7880 1943
rect 520 857 2120 880
rect 520 823 555 857
rect 589 823 623 857
rect 657 823 691 857
rect 725 823 759 857
rect 793 823 827 857
rect 861 823 895 857
rect 929 823 963 857
rect 997 823 1031 857
rect 1065 823 1099 857
rect 1133 823 1167 857
rect 1201 823 1235 857
rect 1269 823 1303 857
rect 1337 823 1371 857
rect 1405 823 1439 857
rect 1473 823 1507 857
rect 1541 823 1575 857
rect 1609 823 1643 857
rect 1677 823 1711 857
rect 1745 823 1779 857
rect 1813 823 1847 857
rect 1881 823 1915 857
rect 1949 823 1983 857
rect 2017 823 2051 857
rect 2085 823 2120 857
rect 520 760 2120 823
rect 2440 857 4040 880
rect 2440 823 2475 857
rect 2509 823 2543 857
rect 2577 823 2611 857
rect 2645 823 2679 857
rect 2713 823 2747 857
rect 2781 823 2815 857
rect 2849 823 2883 857
rect 2917 823 2951 857
rect 2985 823 3019 857
rect 3053 823 3087 857
rect 3121 823 3155 857
rect 3189 823 3223 857
rect 3257 823 3291 857
rect 3325 823 3359 857
rect 3393 823 3427 857
rect 3461 823 3495 857
rect 3529 823 3563 857
rect 3597 823 3631 857
rect 3665 823 3699 857
rect 3733 823 3767 857
rect 3801 823 3835 857
rect 3869 823 3903 857
rect 3937 823 3971 857
rect 4005 823 4040 857
rect 2440 760 4040 823
rect 4360 857 5960 880
rect 4360 823 4395 857
rect 4429 823 4463 857
rect 4497 823 4531 857
rect 4565 823 4599 857
rect 4633 823 4667 857
rect 4701 823 4735 857
rect 4769 823 4803 857
rect 4837 823 4871 857
rect 4905 823 4939 857
rect 4973 823 5007 857
rect 5041 823 5075 857
rect 5109 823 5143 857
rect 5177 823 5211 857
rect 5245 823 5279 857
rect 5313 823 5347 857
rect 5381 823 5415 857
rect 5449 823 5483 857
rect 5517 823 5551 857
rect 5585 823 5619 857
rect 5653 823 5687 857
rect 5721 823 5755 857
rect 5789 823 5823 857
rect 5857 823 5891 857
rect 5925 823 5960 857
rect 4360 760 5960 823
rect 6280 857 7880 880
rect 6280 823 6315 857
rect 6349 823 6383 857
rect 6417 823 6451 857
rect 6485 823 6519 857
rect 6553 823 6587 857
rect 6621 823 6655 857
rect 6689 823 6723 857
rect 6757 823 6791 857
rect 6825 823 6859 857
rect 6893 823 6927 857
rect 6961 823 6995 857
rect 7029 823 7063 857
rect 7097 823 7131 857
rect 7165 823 7199 857
rect 7233 823 7267 857
rect 7301 823 7335 857
rect 7369 823 7403 857
rect 7437 823 7471 857
rect 7505 823 7539 857
rect 7573 823 7607 857
rect 7641 823 7675 857
rect 7709 823 7743 857
rect 7777 823 7811 857
rect 7845 823 7880 857
rect 6280 760 7880 823
rect 520 360 2120 560
rect 2440 360 4040 560
rect 4360 360 5960 560
rect 6280 360 7880 560
rect 520 120 2120 160
rect 2440 120 4040 160
rect 4360 120 5960 160
rect 6280 120 7880 160
<< polycont >>
rect 555 4183 589 4217
rect 623 4183 657 4217
rect 691 4183 725 4217
rect 759 4183 793 4217
rect 827 4183 861 4217
rect 895 4183 929 4217
rect 963 4183 997 4217
rect 1031 4183 1065 4217
rect 1099 4183 1133 4217
rect 1167 4183 1201 4217
rect 1235 4183 1269 4217
rect 1303 4183 1337 4217
rect 1371 4183 1405 4217
rect 1439 4183 1473 4217
rect 1507 4183 1541 4217
rect 1575 4183 1609 4217
rect 1643 4183 1677 4217
rect 1711 4183 1745 4217
rect 1779 4183 1813 4217
rect 1847 4183 1881 4217
rect 1915 4183 1949 4217
rect 1983 4183 2017 4217
rect 2051 4183 2085 4217
rect 2475 4183 2509 4217
rect 2543 4183 2577 4217
rect 2611 4183 2645 4217
rect 2679 4183 2713 4217
rect 2747 4183 2781 4217
rect 2815 4183 2849 4217
rect 2883 4183 2917 4217
rect 2951 4183 2985 4217
rect 3019 4183 3053 4217
rect 3087 4183 3121 4217
rect 3155 4183 3189 4217
rect 3223 4183 3257 4217
rect 3291 4183 3325 4217
rect 3359 4183 3393 4217
rect 3427 4183 3461 4217
rect 3495 4183 3529 4217
rect 3563 4183 3597 4217
rect 3631 4183 3665 4217
rect 3699 4183 3733 4217
rect 3767 4183 3801 4217
rect 3835 4183 3869 4217
rect 3903 4183 3937 4217
rect 3971 4183 4005 4217
rect 4395 4183 4429 4217
rect 4463 4183 4497 4217
rect 4531 4183 4565 4217
rect 4599 4183 4633 4217
rect 4667 4183 4701 4217
rect 4735 4183 4769 4217
rect 4803 4183 4837 4217
rect 4871 4183 4905 4217
rect 4939 4183 4973 4217
rect 5007 4183 5041 4217
rect 5075 4183 5109 4217
rect 5143 4183 5177 4217
rect 5211 4183 5245 4217
rect 5279 4183 5313 4217
rect 5347 4183 5381 4217
rect 5415 4183 5449 4217
rect 5483 4183 5517 4217
rect 5551 4183 5585 4217
rect 5619 4183 5653 4217
rect 5687 4183 5721 4217
rect 5755 4183 5789 4217
rect 5823 4183 5857 4217
rect 5891 4183 5925 4217
rect 6315 4183 6349 4217
rect 6383 4183 6417 4217
rect 6451 4183 6485 4217
rect 6519 4183 6553 4217
rect 6587 4183 6621 4217
rect 6655 4183 6689 4217
rect 6723 4183 6757 4217
rect 6791 4183 6825 4217
rect 6859 4183 6893 4217
rect 6927 4183 6961 4217
rect 6995 4183 7029 4217
rect 7063 4183 7097 4217
rect 7131 4183 7165 4217
rect 7199 4183 7233 4217
rect 7267 4183 7301 4217
rect 7335 4183 7369 4217
rect 7403 4183 7437 4217
rect 7471 4183 7505 4217
rect 7539 4183 7573 4217
rect 7607 4183 7641 4217
rect 7675 4183 7709 4217
rect 7743 4183 7777 4217
rect 7811 4183 7845 4217
rect 555 1943 589 1977
rect 623 1943 657 1977
rect 691 1943 725 1977
rect 759 1943 793 1977
rect 827 1943 861 1977
rect 895 1943 929 1977
rect 963 1943 997 1977
rect 1031 1943 1065 1977
rect 1099 1943 1133 1977
rect 1167 1943 1201 1977
rect 1235 1943 1269 1977
rect 1303 1943 1337 1977
rect 1371 1943 1405 1977
rect 1439 1943 1473 1977
rect 1507 1943 1541 1977
rect 1575 1943 1609 1977
rect 1643 1943 1677 1977
rect 1711 1943 1745 1977
rect 1779 1943 1813 1977
rect 1847 1943 1881 1977
rect 1915 1943 1949 1977
rect 1983 1943 2017 1977
rect 2051 1943 2085 1977
rect 2475 1943 2509 1977
rect 2543 1943 2577 1977
rect 2611 1943 2645 1977
rect 2679 1943 2713 1977
rect 2747 1943 2781 1977
rect 2815 1943 2849 1977
rect 2883 1943 2917 1977
rect 2951 1943 2985 1977
rect 3019 1943 3053 1977
rect 3087 1943 3121 1977
rect 3155 1943 3189 1977
rect 3223 1943 3257 1977
rect 3291 1943 3325 1977
rect 3359 1943 3393 1977
rect 3427 1943 3461 1977
rect 3495 1943 3529 1977
rect 3563 1943 3597 1977
rect 3631 1943 3665 1977
rect 3699 1943 3733 1977
rect 3767 1943 3801 1977
rect 3835 1943 3869 1977
rect 3903 1943 3937 1977
rect 3971 1943 4005 1977
rect 4395 1943 4429 1977
rect 4463 1943 4497 1977
rect 4531 1943 4565 1977
rect 4599 1943 4633 1977
rect 4667 1943 4701 1977
rect 4735 1943 4769 1977
rect 4803 1943 4837 1977
rect 4871 1943 4905 1977
rect 4939 1943 4973 1977
rect 5007 1943 5041 1977
rect 5075 1943 5109 1977
rect 5143 1943 5177 1977
rect 5211 1943 5245 1977
rect 5279 1943 5313 1977
rect 5347 1943 5381 1977
rect 5415 1943 5449 1977
rect 5483 1943 5517 1977
rect 5551 1943 5585 1977
rect 5619 1943 5653 1977
rect 5687 1943 5721 1977
rect 5755 1943 5789 1977
rect 5823 1943 5857 1977
rect 5891 1943 5925 1977
rect 6315 1943 6349 1977
rect 6383 1943 6417 1977
rect 6451 1943 6485 1977
rect 6519 1943 6553 1977
rect 6587 1943 6621 1977
rect 6655 1943 6689 1977
rect 6723 1943 6757 1977
rect 6791 1943 6825 1977
rect 6859 1943 6893 1977
rect 6927 1943 6961 1977
rect 6995 1943 7029 1977
rect 7063 1943 7097 1977
rect 7131 1943 7165 1977
rect 7199 1943 7233 1977
rect 7267 1943 7301 1977
rect 7335 1943 7369 1977
rect 7403 1943 7437 1977
rect 7471 1943 7505 1977
rect 7539 1943 7573 1977
rect 7607 1943 7641 1977
rect 7675 1943 7709 1977
rect 7743 1943 7777 1977
rect 7811 1943 7845 1977
rect 555 823 589 857
rect 623 823 657 857
rect 691 823 725 857
rect 759 823 793 857
rect 827 823 861 857
rect 895 823 929 857
rect 963 823 997 857
rect 1031 823 1065 857
rect 1099 823 1133 857
rect 1167 823 1201 857
rect 1235 823 1269 857
rect 1303 823 1337 857
rect 1371 823 1405 857
rect 1439 823 1473 857
rect 1507 823 1541 857
rect 1575 823 1609 857
rect 1643 823 1677 857
rect 1711 823 1745 857
rect 1779 823 1813 857
rect 1847 823 1881 857
rect 1915 823 1949 857
rect 1983 823 2017 857
rect 2051 823 2085 857
rect 2475 823 2509 857
rect 2543 823 2577 857
rect 2611 823 2645 857
rect 2679 823 2713 857
rect 2747 823 2781 857
rect 2815 823 2849 857
rect 2883 823 2917 857
rect 2951 823 2985 857
rect 3019 823 3053 857
rect 3087 823 3121 857
rect 3155 823 3189 857
rect 3223 823 3257 857
rect 3291 823 3325 857
rect 3359 823 3393 857
rect 3427 823 3461 857
rect 3495 823 3529 857
rect 3563 823 3597 857
rect 3631 823 3665 857
rect 3699 823 3733 857
rect 3767 823 3801 857
rect 3835 823 3869 857
rect 3903 823 3937 857
rect 3971 823 4005 857
rect 4395 823 4429 857
rect 4463 823 4497 857
rect 4531 823 4565 857
rect 4599 823 4633 857
rect 4667 823 4701 857
rect 4735 823 4769 857
rect 4803 823 4837 857
rect 4871 823 4905 857
rect 4939 823 4973 857
rect 5007 823 5041 857
rect 5075 823 5109 857
rect 5143 823 5177 857
rect 5211 823 5245 857
rect 5279 823 5313 857
rect 5347 823 5381 857
rect 5415 823 5449 857
rect 5483 823 5517 857
rect 5551 823 5585 857
rect 5619 823 5653 857
rect 5687 823 5721 857
rect 5755 823 5789 857
rect 5823 823 5857 857
rect 5891 823 5925 857
rect 6315 823 6349 857
rect 6383 823 6417 857
rect 6451 823 6485 857
rect 6519 823 6553 857
rect 6587 823 6621 857
rect 6655 823 6689 857
rect 6723 823 6757 857
rect 6791 823 6825 857
rect 6859 823 6893 857
rect 6927 823 6961 857
rect 6995 823 7029 857
rect 7063 823 7097 857
rect 7131 823 7165 857
rect 7199 823 7233 857
rect 7267 823 7301 857
rect 7335 823 7369 857
rect 7403 823 7437 857
rect 7471 823 7505 857
rect 7539 823 7573 857
rect 7607 823 7641 857
rect 7675 823 7709 857
rect 7743 823 7777 857
rect 7811 823 7845 857
<< locali >>
rect 0 5977 8400 6000
rect 0 5943 137 5977
rect 171 5943 205 5977
rect 239 5943 273 5977
rect 307 5943 341 5977
rect 375 5943 409 5977
rect 443 5943 477 5977
rect 511 5943 545 5977
rect 579 5943 613 5977
rect 647 5943 681 5977
rect 715 5943 749 5977
rect 783 5943 817 5977
rect 851 5943 885 5977
rect 919 5943 953 5977
rect 987 5943 1021 5977
rect 1055 5943 1089 5977
rect 1123 5943 1157 5977
rect 1191 5943 1225 5977
rect 1259 5943 1293 5977
rect 1327 5943 1361 5977
rect 1395 5943 1429 5977
rect 1463 5943 1497 5977
rect 1531 5943 1565 5977
rect 1599 5943 1633 5977
rect 1667 5943 1701 5977
rect 1735 5943 1769 5977
rect 1803 5943 1837 5977
rect 1871 5943 1905 5977
rect 1939 5943 1973 5977
rect 2007 5943 2041 5977
rect 2075 5943 2109 5977
rect 2143 5943 2177 5977
rect 2211 5943 2245 5977
rect 2279 5943 2313 5977
rect 2347 5943 2381 5977
rect 2415 5943 2449 5977
rect 2483 5943 2517 5977
rect 2551 5943 2585 5977
rect 2619 5943 2653 5977
rect 2687 5943 2721 5977
rect 2755 5943 2789 5977
rect 2823 5943 2857 5977
rect 2891 5943 2925 5977
rect 2959 5943 2993 5977
rect 3027 5943 3061 5977
rect 3095 5943 3129 5977
rect 3163 5943 3197 5977
rect 3231 5943 3265 5977
rect 3299 5943 3333 5977
rect 3367 5943 3401 5977
rect 3435 5943 3469 5977
rect 3503 5943 3537 5977
rect 3571 5943 3605 5977
rect 3639 5943 3673 5977
rect 3707 5943 3741 5977
rect 3775 5943 3809 5977
rect 3843 5943 3877 5977
rect 3911 5943 3945 5977
rect 3979 5943 4013 5977
rect 4047 5943 4081 5977
rect 4115 5943 4149 5977
rect 4183 5943 4217 5977
rect 4251 5943 4285 5977
rect 4319 5943 4353 5977
rect 4387 5943 4421 5977
rect 4455 5943 4489 5977
rect 4523 5943 4557 5977
rect 4591 5943 4625 5977
rect 4659 5943 4693 5977
rect 4727 5943 4761 5977
rect 4795 5943 4829 5977
rect 4863 5943 4897 5977
rect 4931 5943 4965 5977
rect 4999 5943 5033 5977
rect 5067 5943 5101 5977
rect 5135 5943 5169 5977
rect 5203 5943 5237 5977
rect 5271 5943 5305 5977
rect 5339 5943 5373 5977
rect 5407 5943 5441 5977
rect 5475 5943 5509 5977
rect 5543 5943 5577 5977
rect 5611 5943 5645 5977
rect 5679 5943 5713 5977
rect 5747 5943 5781 5977
rect 5815 5943 5849 5977
rect 5883 5943 5917 5977
rect 5951 5943 5985 5977
rect 6019 5943 6053 5977
rect 6087 5943 6121 5977
rect 6155 5943 6189 5977
rect 6223 5943 6257 5977
rect 6291 5943 6325 5977
rect 6359 5943 6393 5977
rect 6427 5943 6461 5977
rect 6495 5943 6529 5977
rect 6563 5943 6597 5977
rect 6631 5943 6665 5977
rect 6699 5943 6733 5977
rect 6767 5943 6801 5977
rect 6835 5943 6869 5977
rect 6903 5943 6937 5977
rect 6971 5943 7005 5977
rect 7039 5943 7073 5977
rect 7107 5943 7141 5977
rect 7175 5943 7209 5977
rect 7243 5943 7277 5977
rect 7311 5943 7345 5977
rect 7379 5943 7413 5977
rect 7447 5943 7481 5977
rect 7515 5943 7549 5977
rect 7583 5943 7617 5977
rect 7651 5943 7685 5977
rect 7719 5943 7753 5977
rect 7787 5943 7821 5977
rect 7855 5943 7889 5977
rect 7923 5943 7957 5977
rect 7991 5943 8025 5977
rect 8059 5943 8093 5977
rect 8127 5943 8161 5977
rect 8195 5943 8229 5977
rect 8263 5943 8400 5977
rect 0 5920 8400 5943
rect 0 5855 80 5920
rect 0 5821 23 5855
rect 57 5821 80 5855
rect 8320 5855 8400 5920
rect 0 5787 80 5821
rect 0 5753 23 5787
rect 57 5753 80 5787
rect 0 5719 80 5753
rect 0 5685 23 5719
rect 57 5685 80 5719
rect 0 5651 80 5685
rect 0 5617 23 5651
rect 57 5617 80 5651
rect 0 5583 80 5617
rect 0 5549 23 5583
rect 57 5549 80 5583
rect 0 5515 80 5549
rect 0 5481 23 5515
rect 57 5481 80 5515
rect 0 5447 80 5481
rect 0 5413 23 5447
rect 57 5413 80 5447
rect 0 5379 80 5413
rect 0 5345 23 5379
rect 57 5345 80 5379
rect 0 5311 80 5345
rect 0 5277 23 5311
rect 57 5277 80 5311
rect 0 5243 80 5277
rect 0 5209 23 5243
rect 57 5209 80 5243
rect 0 5175 80 5209
rect 0 5141 23 5175
rect 57 5141 80 5175
rect 0 5107 80 5141
rect 0 5073 23 5107
rect 57 5073 80 5107
rect 0 5039 80 5073
rect 0 5005 23 5039
rect 57 5005 80 5039
rect 0 4971 80 5005
rect 0 4937 23 4971
rect 57 4937 80 4971
rect 0 4903 80 4937
rect 0 4869 23 4903
rect 57 4869 80 4903
rect 0 4835 80 4869
rect 0 4801 23 4835
rect 57 4801 80 4835
rect 0 4767 80 4801
rect 0 4733 23 4767
rect 57 4733 80 4767
rect 0 4699 80 4733
rect 0 4665 23 4699
rect 57 4665 80 4699
rect 0 4631 80 4665
rect 0 4597 23 4631
rect 57 4597 80 4631
rect 0 4563 80 4597
rect 0 4529 23 4563
rect 57 4529 80 4563
rect 0 4495 80 4529
rect 0 4461 23 4495
rect 57 4461 80 4495
rect 0 4427 80 4461
rect 0 4393 23 4427
rect 57 4393 80 4427
rect 0 4359 80 4393
rect 0 4325 23 4359
rect 57 4325 80 4359
rect 0 4291 80 4325
rect 0 4257 23 4291
rect 57 4257 80 4291
rect 0 4223 80 4257
rect 0 4189 23 4223
rect 57 4189 80 4223
rect 0 4155 80 4189
rect 0 4121 23 4155
rect 57 4121 80 4155
rect 0 4087 80 4121
rect 0 4053 23 4087
rect 57 4053 80 4087
rect 0 4019 80 4053
rect 0 3985 23 4019
rect 57 3985 80 4019
rect 160 5817 8240 5840
rect 160 5783 307 5817
rect 341 5783 375 5817
rect 409 5783 443 5817
rect 477 5783 511 5817
rect 545 5783 579 5817
rect 613 5783 647 5817
rect 681 5783 715 5817
rect 749 5783 783 5817
rect 817 5783 851 5817
rect 885 5783 919 5817
rect 953 5783 987 5817
rect 1021 5783 1055 5817
rect 1089 5783 1123 5817
rect 1157 5783 1191 5817
rect 1225 5783 1259 5817
rect 1293 5783 1327 5817
rect 1361 5783 1395 5817
rect 1429 5783 1463 5817
rect 1497 5783 1531 5817
rect 1565 5783 1599 5817
rect 1633 5783 1667 5817
rect 1701 5783 1735 5817
rect 1769 5783 1803 5817
rect 1837 5783 1871 5817
rect 1905 5783 1939 5817
rect 1973 5783 2007 5817
rect 2041 5783 2075 5817
rect 2109 5783 2143 5817
rect 2177 5783 2211 5817
rect 2245 5783 2279 5817
rect 2313 5783 2347 5817
rect 2381 5783 2415 5817
rect 2449 5783 2483 5817
rect 2517 5783 2551 5817
rect 2585 5783 2619 5817
rect 2653 5783 2687 5817
rect 2721 5783 2755 5817
rect 2789 5783 2823 5817
rect 2857 5783 2891 5817
rect 2925 5783 2959 5817
rect 2993 5783 3027 5817
rect 3061 5783 3095 5817
rect 3129 5783 3163 5817
rect 3197 5783 3231 5817
rect 3265 5783 3299 5817
rect 3333 5783 3367 5817
rect 3401 5783 3435 5817
rect 3469 5783 3503 5817
rect 3537 5783 3571 5817
rect 3605 5783 3639 5817
rect 3673 5783 3707 5817
rect 3741 5783 3775 5817
rect 3809 5783 3843 5817
rect 3877 5783 3911 5817
rect 3945 5783 3979 5817
rect 4013 5783 4047 5817
rect 4081 5783 4115 5817
rect 4149 5783 4183 5817
rect 4217 5783 4251 5817
rect 4285 5783 4319 5817
rect 4353 5783 4387 5817
rect 4421 5783 4455 5817
rect 4489 5783 4523 5817
rect 4557 5783 4591 5817
rect 4625 5783 4659 5817
rect 4693 5783 4727 5817
rect 4761 5783 4795 5817
rect 4829 5783 4863 5817
rect 4897 5783 4931 5817
rect 4965 5783 4999 5817
rect 5033 5783 5067 5817
rect 5101 5783 5135 5817
rect 5169 5783 5203 5817
rect 5237 5783 5271 5817
rect 5305 5783 5339 5817
rect 5373 5783 5407 5817
rect 5441 5783 5475 5817
rect 5509 5783 5543 5817
rect 5577 5783 5611 5817
rect 5645 5783 5679 5817
rect 5713 5783 5747 5817
rect 5781 5783 5815 5817
rect 5849 5783 5883 5817
rect 5917 5783 5951 5817
rect 5985 5783 6019 5817
rect 6053 5783 6087 5817
rect 6121 5783 6155 5817
rect 6189 5783 6223 5817
rect 6257 5783 6291 5817
rect 6325 5783 6359 5817
rect 6393 5783 6427 5817
rect 6461 5783 6495 5817
rect 6529 5783 6563 5817
rect 6597 5783 6631 5817
rect 6665 5783 6699 5817
rect 6733 5783 6767 5817
rect 6801 5783 6835 5817
rect 6869 5783 6903 5817
rect 6937 5783 6971 5817
rect 7005 5783 7039 5817
rect 7073 5783 7107 5817
rect 7141 5783 7175 5817
rect 7209 5783 7243 5817
rect 7277 5783 7311 5817
rect 7345 5783 7379 5817
rect 7413 5783 7447 5817
rect 7481 5783 7515 5817
rect 7549 5783 7583 5817
rect 7617 5783 7651 5817
rect 7685 5783 7719 5817
rect 7753 5783 7787 5817
rect 7821 5783 7855 5817
rect 7889 5783 7923 5817
rect 7957 5783 7991 5817
rect 8025 5783 8059 5817
rect 8093 5783 8240 5817
rect 160 5760 8240 5783
rect 160 5719 240 5760
rect 160 5685 183 5719
rect 217 5685 240 5719
rect 160 5651 240 5685
rect 160 5617 183 5651
rect 217 5617 240 5651
rect 160 5583 240 5617
rect 160 5549 183 5583
rect 217 5549 240 5583
rect 160 5515 240 5549
rect 160 5481 183 5515
rect 217 5481 240 5515
rect 160 5447 240 5481
rect 160 5413 183 5447
rect 217 5413 240 5447
rect 160 5379 240 5413
rect 160 5345 183 5379
rect 217 5345 240 5379
rect 160 5311 240 5345
rect 160 5277 183 5311
rect 217 5277 240 5311
rect 160 5243 240 5277
rect 160 5209 183 5243
rect 217 5209 240 5243
rect 160 5175 240 5209
rect 160 5141 183 5175
rect 217 5141 240 5175
rect 160 5107 240 5141
rect 160 5073 183 5107
rect 217 5073 240 5107
rect 320 5649 400 5680
rect 320 5601 343 5649
rect 377 5601 400 5649
rect 320 5577 400 5601
rect 320 5533 343 5577
rect 377 5533 400 5577
rect 320 5505 400 5533
rect 320 5465 343 5505
rect 377 5465 400 5505
rect 320 5433 400 5465
rect 320 5397 343 5433
rect 377 5397 400 5433
rect 320 5363 400 5397
rect 320 5327 343 5363
rect 377 5327 400 5363
rect 320 5295 400 5327
rect 320 5255 343 5295
rect 377 5255 400 5295
rect 320 5227 400 5255
rect 320 5183 343 5227
rect 377 5183 400 5227
rect 320 5159 400 5183
rect 320 5111 343 5159
rect 377 5111 400 5159
rect 320 5080 400 5111
rect 2240 5649 2320 5680
rect 2240 5601 2263 5649
rect 2297 5601 2320 5649
rect 2240 5577 2320 5601
rect 2240 5533 2263 5577
rect 2297 5533 2320 5577
rect 2240 5505 2320 5533
rect 2240 5465 2263 5505
rect 2297 5465 2320 5505
rect 2240 5433 2320 5465
rect 2240 5397 2263 5433
rect 2297 5397 2320 5433
rect 2240 5363 2320 5397
rect 2240 5327 2263 5363
rect 2297 5327 2320 5363
rect 2240 5295 2320 5327
rect 2240 5255 2263 5295
rect 2297 5255 2320 5295
rect 2240 5227 2320 5255
rect 2240 5183 2263 5227
rect 2297 5183 2320 5227
rect 2240 5159 2320 5183
rect 2240 5111 2263 5159
rect 2297 5111 2320 5159
rect 2240 5080 2320 5111
rect 4160 5649 4240 5760
rect 8160 5719 8240 5760
rect 8160 5685 8183 5719
rect 8217 5685 8240 5719
rect 4160 5601 4183 5649
rect 4217 5601 4240 5649
rect 4160 5577 4240 5601
rect 4160 5533 4183 5577
rect 4217 5533 4240 5577
rect 4160 5505 4240 5533
rect 4160 5465 4183 5505
rect 4217 5465 4240 5505
rect 4160 5433 4240 5465
rect 4160 5397 4183 5433
rect 4217 5397 4240 5433
rect 4160 5363 4240 5397
rect 4160 5327 4183 5363
rect 4217 5327 4240 5363
rect 4160 5295 4240 5327
rect 4160 5255 4183 5295
rect 4217 5255 4240 5295
rect 4160 5227 4240 5255
rect 4160 5183 4183 5227
rect 4217 5183 4240 5227
rect 4160 5159 4240 5183
rect 4160 5111 4183 5159
rect 4217 5111 4240 5159
rect 160 5039 240 5073
rect 4160 5040 4240 5111
rect 6080 5649 6160 5680
rect 6080 5601 6103 5649
rect 6137 5601 6160 5649
rect 6080 5577 6160 5601
rect 6080 5533 6103 5577
rect 6137 5533 6160 5577
rect 6080 5505 6160 5533
rect 6080 5465 6103 5505
rect 6137 5465 6160 5505
rect 6080 5433 6160 5465
rect 6080 5397 6103 5433
rect 6137 5397 6160 5433
rect 6080 5363 6160 5397
rect 6080 5327 6103 5363
rect 6137 5327 6160 5363
rect 6080 5295 6160 5327
rect 6080 5255 6103 5295
rect 6137 5255 6160 5295
rect 6080 5227 6160 5255
rect 6080 5183 6103 5227
rect 6137 5183 6160 5227
rect 6080 5159 6160 5183
rect 6080 5111 6103 5159
rect 6137 5111 6160 5159
rect 6080 5080 6160 5111
rect 8000 5649 8080 5680
rect 8000 5601 8023 5649
rect 8057 5601 8080 5649
rect 8000 5577 8080 5601
rect 8000 5533 8023 5577
rect 8057 5533 8080 5577
rect 8000 5505 8080 5533
rect 8000 5465 8023 5505
rect 8057 5465 8080 5505
rect 8000 5433 8080 5465
rect 8000 5397 8023 5433
rect 8057 5397 8080 5433
rect 8000 5363 8080 5397
rect 8000 5327 8023 5363
rect 8057 5327 8080 5363
rect 8000 5295 8080 5327
rect 8000 5255 8023 5295
rect 8057 5255 8080 5295
rect 8000 5227 8080 5255
rect 8000 5183 8023 5227
rect 8057 5183 8080 5227
rect 8000 5159 8080 5183
rect 8000 5111 8023 5159
rect 8057 5111 8080 5159
rect 8000 5080 8080 5111
rect 8160 5651 8240 5685
rect 8160 5617 8183 5651
rect 8217 5617 8240 5651
rect 8160 5583 8240 5617
rect 8160 5549 8183 5583
rect 8217 5549 8240 5583
rect 8160 5515 8240 5549
rect 8160 5481 8183 5515
rect 8217 5481 8240 5515
rect 8160 5447 8240 5481
rect 8160 5413 8183 5447
rect 8217 5413 8240 5447
rect 8160 5379 8240 5413
rect 8160 5345 8183 5379
rect 8217 5345 8240 5379
rect 8160 5311 8240 5345
rect 8160 5277 8183 5311
rect 8217 5277 8240 5311
rect 8160 5243 8240 5277
rect 8160 5209 8183 5243
rect 8217 5209 8240 5243
rect 8160 5175 8240 5209
rect 8160 5141 8183 5175
rect 8217 5141 8240 5175
rect 8160 5107 8240 5141
rect 8160 5073 8183 5107
rect 8217 5073 8240 5107
rect 160 5005 183 5039
rect 217 5005 240 5039
rect 160 4971 240 5005
rect 160 4937 183 4971
rect 217 4937 240 4971
rect 160 4903 240 4937
rect 2240 4960 6160 5040
rect 160 4869 183 4903
rect 217 4869 240 4903
rect 160 4835 240 4869
rect 160 4801 183 4835
rect 217 4801 240 4835
rect 160 4767 240 4801
rect 160 4733 183 4767
rect 217 4733 240 4767
rect 160 4699 240 4733
rect 160 4665 183 4699
rect 217 4665 240 4699
rect 160 4631 240 4665
rect 160 4597 183 4631
rect 217 4597 240 4631
rect 160 4563 240 4597
rect 160 4529 183 4563
rect 217 4529 240 4563
rect 160 4495 240 4529
rect 160 4461 183 4495
rect 217 4461 240 4495
rect 160 4427 240 4461
rect 160 4393 183 4427
rect 217 4393 240 4427
rect 160 4359 240 4393
rect 160 4325 183 4359
rect 217 4325 240 4359
rect 160 4291 240 4325
rect 320 4889 400 4920
rect 320 4841 343 4889
rect 377 4841 400 4889
rect 320 4817 400 4841
rect 320 4773 343 4817
rect 377 4773 400 4817
rect 320 4745 400 4773
rect 320 4705 343 4745
rect 377 4705 400 4745
rect 320 4673 400 4705
rect 320 4637 343 4673
rect 377 4637 400 4673
rect 320 4603 400 4637
rect 320 4567 343 4603
rect 377 4567 400 4603
rect 320 4535 400 4567
rect 320 4495 343 4535
rect 377 4495 400 4535
rect 320 4467 400 4495
rect 320 4423 343 4467
rect 377 4423 400 4467
rect 320 4399 400 4423
rect 320 4351 343 4399
rect 377 4351 400 4399
rect 320 4320 400 4351
rect 2240 4889 2320 4960
rect 2240 4841 2263 4889
rect 2297 4841 2320 4889
rect 2240 4817 2320 4841
rect 2240 4773 2263 4817
rect 2297 4773 2320 4817
rect 2240 4745 2320 4773
rect 2240 4705 2263 4745
rect 2297 4705 2320 4745
rect 2240 4673 2320 4705
rect 2240 4637 2263 4673
rect 2297 4637 2320 4673
rect 2240 4603 2320 4637
rect 2240 4567 2263 4603
rect 2297 4567 2320 4603
rect 2240 4535 2320 4567
rect 2240 4495 2263 4535
rect 2297 4495 2320 4535
rect 2240 4467 2320 4495
rect 2240 4423 2263 4467
rect 2297 4423 2320 4467
rect 2240 4399 2320 4423
rect 2240 4351 2263 4399
rect 2297 4351 2320 4399
rect 2240 4320 2320 4351
rect 4160 4889 4240 4920
rect 4160 4841 4183 4889
rect 4217 4841 4240 4889
rect 4160 4817 4240 4841
rect 4160 4773 4183 4817
rect 4217 4773 4240 4817
rect 4160 4745 4240 4773
rect 4160 4705 4183 4745
rect 4217 4705 4240 4745
rect 4160 4673 4240 4705
rect 4160 4637 4183 4673
rect 4217 4637 4240 4673
rect 4160 4603 4240 4637
rect 4160 4567 4183 4603
rect 4217 4567 4240 4603
rect 4160 4535 4240 4567
rect 4160 4495 4183 4535
rect 4217 4495 4240 4535
rect 4160 4467 4240 4495
rect 4160 4423 4183 4467
rect 4217 4423 4240 4467
rect 4160 4399 4240 4423
rect 4160 4351 4183 4399
rect 4217 4351 4240 4399
rect 4160 4320 4240 4351
rect 6080 4889 6160 4960
rect 8160 5039 8240 5073
rect 8160 5005 8183 5039
rect 8217 5005 8240 5039
rect 8160 4971 8240 5005
rect 8160 4937 8183 4971
rect 8217 4937 8240 4971
rect 6080 4841 6103 4889
rect 6137 4841 6160 4889
rect 6080 4817 6160 4841
rect 6080 4773 6103 4817
rect 6137 4773 6160 4817
rect 6080 4745 6160 4773
rect 6080 4705 6103 4745
rect 6137 4705 6160 4745
rect 6080 4673 6160 4705
rect 6080 4637 6103 4673
rect 6137 4637 6160 4673
rect 6080 4603 6160 4637
rect 6080 4567 6103 4603
rect 6137 4567 6160 4603
rect 6080 4535 6160 4567
rect 6080 4495 6103 4535
rect 6137 4495 6160 4535
rect 6080 4467 6160 4495
rect 6080 4423 6103 4467
rect 6137 4423 6160 4467
rect 6080 4399 6160 4423
rect 6080 4351 6103 4399
rect 6137 4351 6160 4399
rect 6080 4320 6160 4351
rect 8000 4889 8080 4920
rect 8000 4841 8023 4889
rect 8057 4841 8080 4889
rect 8000 4817 8080 4841
rect 8000 4773 8023 4817
rect 8057 4773 8080 4817
rect 8000 4745 8080 4773
rect 8000 4705 8023 4745
rect 8057 4705 8080 4745
rect 8000 4673 8080 4705
rect 8000 4637 8023 4673
rect 8057 4637 8080 4673
rect 8000 4603 8080 4637
rect 8000 4567 8023 4603
rect 8057 4567 8080 4603
rect 8000 4535 8080 4567
rect 8000 4495 8023 4535
rect 8057 4495 8080 4535
rect 8000 4467 8080 4495
rect 8000 4423 8023 4467
rect 8057 4423 8080 4467
rect 8000 4399 8080 4423
rect 8000 4351 8023 4399
rect 8057 4351 8080 4399
rect 8000 4320 8080 4351
rect 8160 4903 8240 4937
rect 8160 4869 8183 4903
rect 8217 4869 8240 4903
rect 8160 4835 8240 4869
rect 8160 4801 8183 4835
rect 8217 4801 8240 4835
rect 8160 4767 8240 4801
rect 8160 4733 8183 4767
rect 8217 4733 8240 4767
rect 8160 4699 8240 4733
rect 8160 4665 8183 4699
rect 8217 4665 8240 4699
rect 8160 4631 8240 4665
rect 8160 4597 8183 4631
rect 8217 4597 8240 4631
rect 8160 4563 8240 4597
rect 8160 4529 8183 4563
rect 8217 4529 8240 4563
rect 8160 4495 8240 4529
rect 8160 4461 8183 4495
rect 8217 4461 8240 4495
rect 8160 4427 8240 4461
rect 8160 4393 8183 4427
rect 8217 4393 8240 4427
rect 8160 4359 8240 4393
rect 8160 4325 8183 4359
rect 8217 4325 8240 4359
rect 160 4257 183 4291
rect 217 4257 240 4291
rect 160 4223 240 4257
rect 8160 4291 8240 4325
rect 8160 4257 8183 4291
rect 8217 4257 8240 4291
rect 160 4189 183 4223
rect 217 4189 240 4223
rect 160 4155 240 4189
rect 520 4217 2120 4240
rect 520 4183 547 4217
rect 589 4183 619 4217
rect 657 4183 691 4217
rect 725 4183 759 4217
rect 797 4183 827 4217
rect 869 4183 895 4217
rect 941 4183 963 4217
rect 1013 4183 1031 4217
rect 1085 4183 1099 4217
rect 1157 4183 1167 4217
rect 1229 4183 1235 4217
rect 1301 4183 1303 4217
rect 1337 4183 1339 4217
rect 1405 4183 1411 4217
rect 1473 4183 1483 4217
rect 1541 4183 1555 4217
rect 1609 4183 1627 4217
rect 1677 4183 1699 4217
rect 1745 4183 1771 4217
rect 1813 4183 1843 4217
rect 1881 4183 1915 4217
rect 1949 4183 1983 4217
rect 2021 4183 2051 4217
rect 2093 4183 2120 4217
rect 520 4160 2120 4183
rect 2440 4217 4040 4240
rect 2440 4183 2467 4217
rect 2509 4183 2539 4217
rect 2577 4183 2611 4217
rect 2645 4183 2679 4217
rect 2717 4183 2747 4217
rect 2789 4183 2815 4217
rect 2861 4183 2883 4217
rect 2933 4183 2951 4217
rect 3005 4183 3019 4217
rect 3077 4183 3087 4217
rect 3149 4183 3155 4217
rect 3221 4183 3223 4217
rect 3257 4183 3259 4217
rect 3325 4183 3331 4217
rect 3393 4183 3403 4217
rect 3461 4183 3475 4217
rect 3529 4183 3547 4217
rect 3597 4183 3619 4217
rect 3665 4183 3691 4217
rect 3733 4183 3763 4217
rect 3801 4183 3835 4217
rect 3869 4183 3903 4217
rect 3941 4183 3971 4217
rect 4013 4183 4040 4217
rect 2440 4160 4040 4183
rect 4360 4217 5960 4240
rect 4360 4183 4387 4217
rect 4429 4183 4459 4217
rect 4497 4183 4531 4217
rect 4565 4183 4599 4217
rect 4637 4183 4667 4217
rect 4709 4183 4735 4217
rect 4781 4183 4803 4217
rect 4853 4183 4871 4217
rect 4925 4183 4939 4217
rect 4997 4183 5007 4217
rect 5069 4183 5075 4217
rect 5141 4183 5143 4217
rect 5177 4183 5179 4217
rect 5245 4183 5251 4217
rect 5313 4183 5323 4217
rect 5381 4183 5395 4217
rect 5449 4183 5467 4217
rect 5517 4183 5539 4217
rect 5585 4183 5611 4217
rect 5653 4183 5683 4217
rect 5721 4183 5755 4217
rect 5789 4183 5823 4217
rect 5861 4183 5891 4217
rect 5933 4183 5960 4217
rect 4360 4160 5960 4183
rect 6280 4217 7880 4240
rect 6280 4183 6307 4217
rect 6349 4183 6379 4217
rect 6417 4183 6451 4217
rect 6485 4183 6519 4217
rect 6557 4183 6587 4217
rect 6629 4183 6655 4217
rect 6701 4183 6723 4217
rect 6773 4183 6791 4217
rect 6845 4183 6859 4217
rect 6917 4183 6927 4217
rect 6989 4183 6995 4217
rect 7061 4183 7063 4217
rect 7097 4183 7099 4217
rect 7165 4183 7171 4217
rect 7233 4183 7243 4217
rect 7301 4183 7315 4217
rect 7369 4183 7387 4217
rect 7437 4183 7459 4217
rect 7505 4183 7531 4217
rect 7573 4183 7603 4217
rect 7641 4183 7675 4217
rect 7709 4183 7743 4217
rect 7781 4183 7811 4217
rect 7853 4183 7880 4217
rect 6280 4160 7880 4183
rect 8160 4223 8240 4257
rect 8160 4189 8183 4223
rect 8217 4189 8240 4223
rect 160 4121 183 4155
rect 217 4121 240 4155
rect 160 4080 240 4121
rect 8160 4155 8240 4189
rect 8160 4121 8183 4155
rect 8217 4121 8240 4155
rect 8160 4080 8240 4121
rect 160 4057 8240 4080
rect 160 4023 307 4057
rect 341 4023 375 4057
rect 409 4023 443 4057
rect 477 4023 511 4057
rect 545 4023 579 4057
rect 613 4023 647 4057
rect 681 4023 715 4057
rect 749 4023 783 4057
rect 817 4023 851 4057
rect 885 4023 919 4057
rect 953 4023 987 4057
rect 1021 4023 1055 4057
rect 1089 4023 1123 4057
rect 1157 4023 1191 4057
rect 1225 4023 1259 4057
rect 1293 4023 1327 4057
rect 1361 4023 1395 4057
rect 1429 4023 1463 4057
rect 1497 4023 1531 4057
rect 1565 4023 1599 4057
rect 1633 4023 1667 4057
rect 1701 4023 1735 4057
rect 1769 4023 1803 4057
rect 1837 4023 1871 4057
rect 1905 4023 1939 4057
rect 1973 4023 2007 4057
rect 2041 4023 2075 4057
rect 2109 4023 2143 4057
rect 2177 4023 2211 4057
rect 2245 4023 2279 4057
rect 2313 4023 2347 4057
rect 2381 4023 2415 4057
rect 2449 4023 2483 4057
rect 2517 4023 2551 4057
rect 2585 4023 2619 4057
rect 2653 4023 2687 4057
rect 2721 4023 2755 4057
rect 2789 4023 2823 4057
rect 2857 4023 2891 4057
rect 2925 4023 2959 4057
rect 2993 4023 3027 4057
rect 3061 4023 3095 4057
rect 3129 4023 3163 4057
rect 3197 4023 3231 4057
rect 3265 4023 3299 4057
rect 3333 4023 3367 4057
rect 3401 4023 3435 4057
rect 3469 4023 3503 4057
rect 3537 4023 3571 4057
rect 3605 4023 3639 4057
rect 3673 4023 3707 4057
rect 3741 4023 3775 4057
rect 3809 4023 3843 4057
rect 3877 4023 3911 4057
rect 3945 4023 3979 4057
rect 4013 4023 4047 4057
rect 4081 4023 4115 4057
rect 4149 4023 4183 4057
rect 4217 4023 4251 4057
rect 4285 4023 4319 4057
rect 4353 4023 4387 4057
rect 4421 4023 4455 4057
rect 4489 4023 4523 4057
rect 4557 4023 4591 4057
rect 4625 4023 4659 4057
rect 4693 4023 4727 4057
rect 4761 4023 4795 4057
rect 4829 4023 4863 4057
rect 4897 4023 4931 4057
rect 4965 4023 4999 4057
rect 5033 4023 5067 4057
rect 5101 4023 5135 4057
rect 5169 4023 5203 4057
rect 5237 4023 5271 4057
rect 5305 4023 5339 4057
rect 5373 4023 5407 4057
rect 5441 4023 5475 4057
rect 5509 4023 5543 4057
rect 5577 4023 5611 4057
rect 5645 4023 5679 4057
rect 5713 4023 5747 4057
rect 5781 4023 5815 4057
rect 5849 4023 5883 4057
rect 5917 4023 5951 4057
rect 5985 4023 6019 4057
rect 6053 4023 6087 4057
rect 6121 4023 6155 4057
rect 6189 4023 6223 4057
rect 6257 4023 6291 4057
rect 6325 4023 6359 4057
rect 6393 4023 6427 4057
rect 6461 4023 6495 4057
rect 6529 4023 6563 4057
rect 6597 4023 6631 4057
rect 6665 4023 6699 4057
rect 6733 4023 6767 4057
rect 6801 4023 6835 4057
rect 6869 4023 6903 4057
rect 6937 4023 6971 4057
rect 7005 4023 7039 4057
rect 7073 4023 7107 4057
rect 7141 4023 7175 4057
rect 7209 4023 7243 4057
rect 7277 4023 7311 4057
rect 7345 4023 7379 4057
rect 7413 4023 7447 4057
rect 7481 4023 7515 4057
rect 7549 4023 7583 4057
rect 7617 4023 7651 4057
rect 7685 4023 7719 4057
rect 7753 4023 7787 4057
rect 7821 4023 7855 4057
rect 7889 4023 7923 4057
rect 7957 4023 7991 4057
rect 8025 4023 8059 4057
rect 8093 4023 8240 4057
rect 160 4000 8240 4023
rect 8320 5821 8343 5855
rect 8377 5821 8400 5855
rect 8320 5787 8400 5821
rect 8320 5753 8343 5787
rect 8377 5753 8400 5787
rect 8320 5719 8400 5753
rect 8320 5685 8343 5719
rect 8377 5685 8400 5719
rect 8320 5651 8400 5685
rect 8320 5617 8343 5651
rect 8377 5617 8400 5651
rect 8320 5583 8400 5617
rect 8320 5549 8343 5583
rect 8377 5549 8400 5583
rect 8320 5515 8400 5549
rect 8320 5481 8343 5515
rect 8377 5481 8400 5515
rect 8320 5447 8400 5481
rect 8320 5413 8343 5447
rect 8377 5413 8400 5447
rect 8320 5379 8400 5413
rect 8320 5345 8343 5379
rect 8377 5345 8400 5379
rect 8320 5311 8400 5345
rect 8320 5277 8343 5311
rect 8377 5277 8400 5311
rect 8320 5243 8400 5277
rect 8320 5209 8343 5243
rect 8377 5209 8400 5243
rect 8320 5175 8400 5209
rect 8320 5141 8343 5175
rect 8377 5141 8400 5175
rect 8320 5107 8400 5141
rect 8320 5073 8343 5107
rect 8377 5073 8400 5107
rect 8320 5039 8400 5073
rect 8320 5005 8343 5039
rect 8377 5005 8400 5039
rect 8320 4971 8400 5005
rect 8320 4937 8343 4971
rect 8377 4937 8400 4971
rect 8320 4903 8400 4937
rect 8320 4869 8343 4903
rect 8377 4869 8400 4903
rect 8320 4835 8400 4869
rect 8320 4801 8343 4835
rect 8377 4801 8400 4835
rect 8320 4767 8400 4801
rect 8320 4733 8343 4767
rect 8377 4733 8400 4767
rect 8320 4699 8400 4733
rect 8320 4665 8343 4699
rect 8377 4665 8400 4699
rect 8320 4631 8400 4665
rect 8320 4597 8343 4631
rect 8377 4597 8400 4631
rect 8320 4563 8400 4597
rect 8320 4529 8343 4563
rect 8377 4529 8400 4563
rect 8320 4495 8400 4529
rect 8320 4461 8343 4495
rect 8377 4461 8400 4495
rect 8320 4427 8400 4461
rect 8320 4393 8343 4427
rect 8377 4393 8400 4427
rect 8320 4359 8400 4393
rect 8320 4325 8343 4359
rect 8377 4325 8400 4359
rect 8320 4291 8400 4325
rect 8320 4257 8343 4291
rect 8377 4257 8400 4291
rect 8320 4223 8400 4257
rect 8320 4189 8343 4223
rect 8377 4189 8400 4223
rect 8320 4155 8400 4189
rect 8320 4121 8343 4155
rect 8377 4121 8400 4155
rect 8320 4087 8400 4121
rect 8320 4053 8343 4087
rect 8377 4053 8400 4087
rect 8320 4019 8400 4053
rect 0 3920 80 3985
rect 8320 3985 8343 4019
rect 8377 3985 8400 4019
rect 8320 3920 8400 3985
rect 0 3897 8400 3920
rect 0 3863 151 3897
rect 185 3863 219 3897
rect 253 3863 287 3897
rect 321 3863 355 3897
rect 389 3863 423 3897
rect 457 3863 491 3897
rect 525 3863 559 3897
rect 593 3863 627 3897
rect 661 3863 695 3897
rect 729 3863 763 3897
rect 797 3863 831 3897
rect 865 3863 899 3897
rect 933 3863 967 3897
rect 1001 3863 1035 3897
rect 1069 3863 1103 3897
rect 1137 3863 1171 3897
rect 1205 3863 1239 3897
rect 1273 3863 1307 3897
rect 1341 3863 1375 3897
rect 1409 3863 1443 3897
rect 1477 3863 1511 3897
rect 1545 3863 1579 3897
rect 1613 3863 1647 3897
rect 1681 3863 1715 3897
rect 1749 3863 1783 3897
rect 1817 3863 1851 3897
rect 1885 3863 1919 3897
rect 1953 3863 1987 3897
rect 2021 3863 2055 3897
rect 2089 3863 2123 3897
rect 2157 3863 2191 3897
rect 2225 3863 2259 3897
rect 2293 3863 2327 3897
rect 2361 3863 2395 3897
rect 2429 3863 2463 3897
rect 2497 3863 2531 3897
rect 2565 3863 2599 3897
rect 2633 3863 2667 3897
rect 2701 3863 2735 3897
rect 2769 3863 2803 3897
rect 2837 3863 2871 3897
rect 2905 3863 2939 3897
rect 2973 3863 3007 3897
rect 3041 3863 3075 3897
rect 3109 3863 3143 3897
rect 3177 3863 3211 3897
rect 3245 3863 3279 3897
rect 3313 3863 3347 3897
rect 3381 3863 3415 3897
rect 3449 3863 3483 3897
rect 3517 3863 3551 3897
rect 3585 3863 3619 3897
rect 3653 3863 3687 3897
rect 3721 3863 3755 3897
rect 3789 3863 3823 3897
rect 3857 3863 3891 3897
rect 3925 3863 3959 3897
rect 3993 3863 4027 3897
rect 4061 3863 4095 3897
rect 4129 3863 4163 3897
rect 4197 3863 4231 3897
rect 4265 3863 4299 3897
rect 4333 3863 4367 3897
rect 4401 3863 4435 3897
rect 4469 3863 4503 3897
rect 4537 3863 4571 3897
rect 4605 3863 4639 3897
rect 4673 3863 4707 3897
rect 4741 3863 4775 3897
rect 4809 3863 4843 3897
rect 4877 3863 4911 3897
rect 4945 3863 4979 3897
rect 5013 3863 5047 3897
rect 5081 3863 5115 3897
rect 5149 3863 5183 3897
rect 5217 3863 5251 3897
rect 5285 3863 5319 3897
rect 5353 3863 5387 3897
rect 5421 3863 5455 3897
rect 5489 3863 5523 3897
rect 5557 3863 5591 3897
rect 5625 3863 5659 3897
rect 5693 3863 5727 3897
rect 5761 3863 5795 3897
rect 5829 3863 5863 3897
rect 5897 3863 5931 3897
rect 5965 3863 5999 3897
rect 6033 3863 6067 3897
rect 6101 3863 6135 3897
rect 6169 3863 6203 3897
rect 6237 3863 6271 3897
rect 6305 3863 6339 3897
rect 6373 3863 6407 3897
rect 6441 3863 6475 3897
rect 6509 3863 6543 3897
rect 6577 3863 6611 3897
rect 6645 3863 6679 3897
rect 6713 3863 6747 3897
rect 6781 3863 6815 3897
rect 6849 3863 6883 3897
rect 6917 3863 6951 3897
rect 6985 3863 7019 3897
rect 7053 3863 7087 3897
rect 7121 3863 7155 3897
rect 7189 3863 7223 3897
rect 7257 3863 7291 3897
rect 7325 3863 7359 3897
rect 7393 3863 7427 3897
rect 7461 3863 7495 3897
rect 7529 3863 7563 3897
rect 7597 3863 7631 3897
rect 7665 3863 7699 3897
rect 7733 3863 7767 3897
rect 7801 3863 7835 3897
rect 7869 3863 7903 3897
rect 7937 3863 7971 3897
rect 8005 3863 8039 3897
rect 8073 3863 8107 3897
rect 8141 3863 8175 3897
rect 8209 3863 8400 3897
rect 0 3840 8400 3863
rect 0 3760 80 3840
rect 8320 3760 8400 3840
rect 0 3737 8400 3760
rect 0 3703 151 3737
rect 185 3703 219 3737
rect 253 3703 287 3737
rect 321 3703 355 3737
rect 389 3703 423 3737
rect 457 3703 491 3737
rect 525 3703 559 3737
rect 593 3703 627 3737
rect 661 3703 695 3737
rect 729 3703 763 3737
rect 797 3703 831 3737
rect 865 3703 899 3737
rect 933 3703 967 3737
rect 1001 3703 1035 3737
rect 1069 3703 1103 3737
rect 1137 3703 1171 3737
rect 1205 3703 1239 3737
rect 1273 3703 1307 3737
rect 1341 3703 1375 3737
rect 1409 3703 1443 3737
rect 1477 3703 1511 3737
rect 1545 3703 1579 3737
rect 1613 3703 1647 3737
rect 1681 3703 1715 3737
rect 1749 3703 1783 3737
rect 1817 3703 1851 3737
rect 1885 3703 1919 3737
rect 1953 3703 1987 3737
rect 2021 3703 2055 3737
rect 2089 3703 2123 3737
rect 2157 3703 2191 3737
rect 2225 3703 2259 3737
rect 2293 3703 2327 3737
rect 2361 3703 2395 3737
rect 2429 3703 2463 3737
rect 2497 3703 2531 3737
rect 2565 3703 2599 3737
rect 2633 3703 2667 3737
rect 2701 3703 2735 3737
rect 2769 3703 2803 3737
rect 2837 3703 2871 3737
rect 2905 3703 2939 3737
rect 2973 3703 3007 3737
rect 3041 3703 3075 3737
rect 3109 3703 3143 3737
rect 3177 3703 3211 3737
rect 3245 3703 3279 3737
rect 3313 3703 3347 3737
rect 3381 3703 3415 3737
rect 3449 3703 3483 3737
rect 3517 3703 3551 3737
rect 3585 3703 3619 3737
rect 3653 3703 3687 3737
rect 3721 3703 3755 3737
rect 3789 3703 3823 3737
rect 3857 3703 3891 3737
rect 3925 3703 3959 3737
rect 3993 3703 4027 3737
rect 4061 3703 4095 3737
rect 4129 3703 4163 3737
rect 4197 3703 4231 3737
rect 4265 3703 4299 3737
rect 4333 3703 4367 3737
rect 4401 3703 4435 3737
rect 4469 3703 4503 3737
rect 4537 3703 4571 3737
rect 4605 3703 4639 3737
rect 4673 3703 4707 3737
rect 4741 3703 4775 3737
rect 4809 3703 4843 3737
rect 4877 3703 4911 3737
rect 4945 3703 4979 3737
rect 5013 3703 5047 3737
rect 5081 3703 5115 3737
rect 5149 3703 5183 3737
rect 5217 3703 5251 3737
rect 5285 3703 5319 3737
rect 5353 3703 5387 3737
rect 5421 3703 5455 3737
rect 5489 3703 5523 3737
rect 5557 3703 5591 3737
rect 5625 3703 5659 3737
rect 5693 3703 5727 3737
rect 5761 3703 5795 3737
rect 5829 3703 5863 3737
rect 5897 3703 5931 3737
rect 5965 3703 5999 3737
rect 6033 3703 6067 3737
rect 6101 3703 6135 3737
rect 6169 3703 6203 3737
rect 6237 3703 6271 3737
rect 6305 3703 6339 3737
rect 6373 3703 6407 3737
rect 6441 3703 6475 3737
rect 6509 3703 6543 3737
rect 6577 3703 6611 3737
rect 6645 3703 6679 3737
rect 6713 3703 6747 3737
rect 6781 3703 6815 3737
rect 6849 3703 6883 3737
rect 6917 3703 6951 3737
rect 6985 3703 7019 3737
rect 7053 3703 7087 3737
rect 7121 3703 7155 3737
rect 7189 3703 7223 3737
rect 7257 3703 7291 3737
rect 7325 3703 7359 3737
rect 7393 3703 7427 3737
rect 7461 3703 7495 3737
rect 7529 3703 7563 3737
rect 7597 3703 7631 3737
rect 7665 3703 7699 3737
rect 7733 3703 7767 3737
rect 7801 3703 7835 3737
rect 7869 3703 7903 3737
rect 7937 3703 7971 3737
rect 8005 3703 8039 3737
rect 8073 3703 8107 3737
rect 8141 3703 8175 3737
rect 8209 3703 8400 3737
rect 0 3680 8400 3703
rect 0 3615 80 3680
rect 0 3581 23 3615
rect 57 3581 80 3615
rect 8320 3615 8400 3680
rect 0 3547 80 3581
rect 0 3513 23 3547
rect 57 3513 80 3547
rect 0 3479 80 3513
rect 0 3445 23 3479
rect 57 3445 80 3479
rect 0 3411 80 3445
rect 0 3377 23 3411
rect 57 3377 80 3411
rect 0 3343 80 3377
rect 0 3309 23 3343
rect 57 3309 80 3343
rect 0 3275 80 3309
rect 0 3241 23 3275
rect 57 3241 80 3275
rect 0 3207 80 3241
rect 0 3173 23 3207
rect 57 3173 80 3207
rect 0 3139 80 3173
rect 0 3105 23 3139
rect 57 3105 80 3139
rect 0 3071 80 3105
rect 0 3037 23 3071
rect 57 3037 80 3071
rect 0 3003 80 3037
rect 0 2969 23 3003
rect 57 2969 80 3003
rect 0 2935 80 2969
rect 0 2901 23 2935
rect 57 2901 80 2935
rect 0 2867 80 2901
rect 0 2833 23 2867
rect 57 2833 80 2867
rect 0 2799 80 2833
rect 0 2765 23 2799
rect 57 2765 80 2799
rect 0 2731 80 2765
rect 0 2697 23 2731
rect 57 2697 80 2731
rect 0 2663 80 2697
rect 0 2629 23 2663
rect 57 2629 80 2663
rect 0 2595 80 2629
rect 0 2561 23 2595
rect 57 2561 80 2595
rect 0 2527 80 2561
rect 0 2493 23 2527
rect 57 2493 80 2527
rect 0 2459 80 2493
rect 0 2425 23 2459
rect 57 2425 80 2459
rect 0 2391 80 2425
rect 0 2357 23 2391
rect 57 2357 80 2391
rect 0 2323 80 2357
rect 0 2289 23 2323
rect 57 2289 80 2323
rect 0 2255 80 2289
rect 0 2221 23 2255
rect 57 2221 80 2255
rect 0 2187 80 2221
rect 0 2153 23 2187
rect 57 2153 80 2187
rect 0 2119 80 2153
rect 0 2085 23 2119
rect 57 2085 80 2119
rect 0 2051 80 2085
rect 0 2017 23 2051
rect 57 2017 80 2051
rect 0 1983 80 2017
rect 0 1949 23 1983
rect 57 1949 80 1983
rect 0 1915 80 1949
rect 0 1881 23 1915
rect 57 1881 80 1915
rect 0 1847 80 1881
rect 0 1813 23 1847
rect 57 1813 80 1847
rect 0 1779 80 1813
rect 0 1745 23 1779
rect 57 1745 80 1779
rect 160 3577 8240 3600
rect 160 3543 307 3577
rect 341 3543 375 3577
rect 409 3543 443 3577
rect 477 3543 511 3577
rect 545 3543 579 3577
rect 613 3543 647 3577
rect 681 3543 715 3577
rect 749 3543 783 3577
rect 817 3543 851 3577
rect 885 3543 919 3577
rect 953 3543 987 3577
rect 1021 3543 1055 3577
rect 1089 3543 1123 3577
rect 1157 3543 1191 3577
rect 1225 3543 1259 3577
rect 1293 3543 1327 3577
rect 1361 3543 1395 3577
rect 1429 3543 1463 3577
rect 1497 3543 1531 3577
rect 1565 3543 1599 3577
rect 1633 3543 1667 3577
rect 1701 3543 1735 3577
rect 1769 3543 1803 3577
rect 1837 3543 1871 3577
rect 1905 3543 1939 3577
rect 1973 3543 2007 3577
rect 2041 3543 2075 3577
rect 2109 3543 2143 3577
rect 2177 3543 2211 3577
rect 2245 3543 2279 3577
rect 2313 3543 2347 3577
rect 2381 3543 2415 3577
rect 2449 3543 2483 3577
rect 2517 3543 2551 3577
rect 2585 3543 2619 3577
rect 2653 3543 2687 3577
rect 2721 3543 2755 3577
rect 2789 3543 2823 3577
rect 2857 3543 2891 3577
rect 2925 3543 2959 3577
rect 2993 3543 3027 3577
rect 3061 3543 3095 3577
rect 3129 3543 3163 3577
rect 3197 3543 3231 3577
rect 3265 3543 3299 3577
rect 3333 3543 3367 3577
rect 3401 3543 3435 3577
rect 3469 3543 3503 3577
rect 3537 3543 3571 3577
rect 3605 3543 3639 3577
rect 3673 3543 3707 3577
rect 3741 3543 3775 3577
rect 3809 3543 3843 3577
rect 3877 3543 3911 3577
rect 3945 3543 3979 3577
rect 4013 3543 4047 3577
rect 4081 3543 4115 3577
rect 4149 3543 4183 3577
rect 4217 3543 4251 3577
rect 4285 3543 4319 3577
rect 4353 3543 4387 3577
rect 4421 3543 4455 3577
rect 4489 3543 4523 3577
rect 4557 3543 4591 3577
rect 4625 3543 4659 3577
rect 4693 3543 4727 3577
rect 4761 3543 4795 3577
rect 4829 3543 4863 3577
rect 4897 3543 4931 3577
rect 4965 3543 4999 3577
rect 5033 3543 5067 3577
rect 5101 3543 5135 3577
rect 5169 3543 5203 3577
rect 5237 3543 5271 3577
rect 5305 3543 5339 3577
rect 5373 3543 5407 3577
rect 5441 3543 5475 3577
rect 5509 3543 5543 3577
rect 5577 3543 5611 3577
rect 5645 3543 5679 3577
rect 5713 3543 5747 3577
rect 5781 3543 5815 3577
rect 5849 3543 5883 3577
rect 5917 3543 5951 3577
rect 5985 3543 6019 3577
rect 6053 3543 6087 3577
rect 6121 3543 6155 3577
rect 6189 3543 6223 3577
rect 6257 3543 6291 3577
rect 6325 3543 6359 3577
rect 6393 3543 6427 3577
rect 6461 3543 6495 3577
rect 6529 3543 6563 3577
rect 6597 3543 6631 3577
rect 6665 3543 6699 3577
rect 6733 3543 6767 3577
rect 6801 3543 6835 3577
rect 6869 3543 6903 3577
rect 6937 3543 6971 3577
rect 7005 3543 7039 3577
rect 7073 3543 7107 3577
rect 7141 3543 7175 3577
rect 7209 3543 7243 3577
rect 7277 3543 7311 3577
rect 7345 3543 7379 3577
rect 7413 3543 7447 3577
rect 7481 3543 7515 3577
rect 7549 3543 7583 3577
rect 7617 3543 7651 3577
rect 7685 3543 7719 3577
rect 7753 3543 7787 3577
rect 7821 3543 7855 3577
rect 7889 3543 7923 3577
rect 7957 3543 7991 3577
rect 8025 3543 8059 3577
rect 8093 3543 8240 3577
rect 160 3520 8240 3543
rect 160 3465 240 3520
rect 160 3431 183 3465
rect 217 3431 240 3465
rect 160 3397 240 3431
rect 160 3363 183 3397
rect 217 3363 240 3397
rect 160 3329 240 3363
rect 160 3295 183 3329
rect 217 3295 240 3329
rect 160 3261 240 3295
rect 160 3227 183 3261
rect 217 3227 240 3261
rect 160 3193 240 3227
rect 160 3159 183 3193
rect 217 3159 240 3193
rect 160 3125 240 3159
rect 160 3091 183 3125
rect 217 3091 240 3125
rect 160 3057 240 3091
rect 160 3023 183 3057
rect 217 3023 240 3057
rect 160 2989 240 3023
rect 160 2955 183 2989
rect 217 2955 240 2989
rect 160 2921 240 2955
rect 160 2887 183 2921
rect 217 2887 240 2921
rect 160 2853 240 2887
rect 160 2819 183 2853
rect 217 2819 240 2853
rect 320 3409 400 3520
rect 320 3361 343 3409
rect 377 3361 400 3409
rect 320 3337 400 3361
rect 320 3293 343 3337
rect 377 3293 400 3337
rect 320 3265 400 3293
rect 320 3225 343 3265
rect 377 3225 400 3265
rect 320 3193 400 3225
rect 320 3157 343 3193
rect 377 3157 400 3193
rect 320 3123 400 3157
rect 320 3087 343 3123
rect 377 3087 400 3123
rect 320 3055 400 3087
rect 320 3015 343 3055
rect 377 3015 400 3055
rect 320 2987 400 3015
rect 320 2943 343 2987
rect 377 2943 400 2987
rect 320 2919 400 2943
rect 320 2871 343 2919
rect 377 2871 400 2919
rect 320 2840 400 2871
rect 2240 3409 2320 3440
rect 2240 3361 2263 3409
rect 2297 3361 2320 3409
rect 2240 3337 2320 3361
rect 2240 3293 2263 3337
rect 2297 3293 2320 3337
rect 2240 3265 2320 3293
rect 2240 3225 2263 3265
rect 2297 3225 2320 3265
rect 2240 3193 2320 3225
rect 2240 3157 2263 3193
rect 2297 3157 2320 3193
rect 2240 3123 2320 3157
rect 2240 3087 2263 3123
rect 2297 3087 2320 3123
rect 2240 3055 2320 3087
rect 2240 3015 2263 3055
rect 2297 3015 2320 3055
rect 2240 2987 2320 3015
rect 2240 2943 2263 2987
rect 2297 2943 2320 2987
rect 2240 2919 2320 2943
rect 2240 2871 2263 2919
rect 2297 2871 2320 2919
rect 2240 2840 2320 2871
rect 4160 3409 4240 3440
rect 4160 3361 4183 3409
rect 4217 3361 4240 3409
rect 4160 3337 4240 3361
rect 4160 3293 4183 3337
rect 4217 3293 4240 3337
rect 4160 3265 4240 3293
rect 4160 3225 4183 3265
rect 4217 3225 4240 3265
rect 4160 3193 4240 3225
rect 4160 3157 4183 3193
rect 4217 3157 4240 3193
rect 4160 3123 4240 3157
rect 4160 3087 4183 3123
rect 4217 3087 4240 3123
rect 4160 3055 4240 3087
rect 4160 3015 4183 3055
rect 4217 3015 4240 3055
rect 4160 2987 4240 3015
rect 4160 2943 4183 2987
rect 4217 2943 4240 2987
rect 4160 2919 4240 2943
rect 4160 2871 4183 2919
rect 4217 2871 4240 2919
rect 160 2785 240 2819
rect 4160 2800 4240 2871
rect 6080 3409 6160 3440
rect 6080 3361 6103 3409
rect 6137 3361 6160 3409
rect 6080 3337 6160 3361
rect 6080 3293 6103 3337
rect 6137 3293 6160 3337
rect 6080 3265 6160 3293
rect 6080 3225 6103 3265
rect 6137 3225 6160 3265
rect 6080 3193 6160 3225
rect 6080 3157 6103 3193
rect 6137 3157 6160 3193
rect 6080 3123 6160 3157
rect 6080 3087 6103 3123
rect 6137 3087 6160 3123
rect 6080 3055 6160 3087
rect 6080 3015 6103 3055
rect 6137 3015 6160 3055
rect 6080 2987 6160 3015
rect 6080 2943 6103 2987
rect 6137 2943 6160 2987
rect 6080 2919 6160 2943
rect 6080 2871 6103 2919
rect 6137 2871 6160 2919
rect 6080 2840 6160 2871
rect 8000 3409 8080 3520
rect 8000 3361 8023 3409
rect 8057 3361 8080 3409
rect 8000 3337 8080 3361
rect 8000 3293 8023 3337
rect 8057 3293 8080 3337
rect 8000 3265 8080 3293
rect 8000 3225 8023 3265
rect 8057 3225 8080 3265
rect 8000 3193 8080 3225
rect 8000 3157 8023 3193
rect 8057 3157 8080 3193
rect 8000 3123 8080 3157
rect 8000 3087 8023 3123
rect 8057 3087 8080 3123
rect 8000 3055 8080 3087
rect 8000 3015 8023 3055
rect 8057 3015 8080 3055
rect 8000 2987 8080 3015
rect 8000 2943 8023 2987
rect 8057 2943 8080 2987
rect 8000 2919 8080 2943
rect 8000 2871 8023 2919
rect 8057 2871 8080 2919
rect 8000 2840 8080 2871
rect 8160 3465 8240 3520
rect 8160 3431 8183 3465
rect 8217 3431 8240 3465
rect 8160 3397 8240 3431
rect 8160 3363 8183 3397
rect 8217 3363 8240 3397
rect 8160 3329 8240 3363
rect 8160 3295 8183 3329
rect 8217 3295 8240 3329
rect 8160 3261 8240 3295
rect 8160 3227 8183 3261
rect 8217 3227 8240 3261
rect 8160 3193 8240 3227
rect 8160 3159 8183 3193
rect 8217 3159 8240 3193
rect 8160 3125 8240 3159
rect 8160 3091 8183 3125
rect 8217 3091 8240 3125
rect 8160 3057 8240 3091
rect 8160 3023 8183 3057
rect 8217 3023 8240 3057
rect 8160 2989 8240 3023
rect 8160 2955 8183 2989
rect 8217 2955 8240 2989
rect 8160 2921 8240 2955
rect 8160 2887 8183 2921
rect 8217 2887 8240 2921
rect 8160 2853 8240 2887
rect 8160 2819 8183 2853
rect 8217 2819 8240 2853
rect 160 2751 183 2785
rect 217 2751 240 2785
rect 160 2717 240 2751
rect 160 2683 183 2717
rect 217 2683 240 2717
rect 160 2649 240 2683
rect 2240 2720 6160 2800
rect 160 2615 183 2649
rect 217 2615 240 2649
rect 160 2581 240 2615
rect 160 2547 183 2581
rect 217 2547 240 2581
rect 160 2513 240 2547
rect 160 2479 183 2513
rect 217 2479 240 2513
rect 160 2445 240 2479
rect 160 2411 183 2445
rect 217 2411 240 2445
rect 160 2377 240 2411
rect 160 2343 183 2377
rect 217 2343 240 2377
rect 160 2309 240 2343
rect 160 2275 183 2309
rect 217 2275 240 2309
rect 160 2241 240 2275
rect 160 2207 183 2241
rect 217 2207 240 2241
rect 160 2173 240 2207
rect 160 2139 183 2173
rect 217 2139 240 2173
rect 160 2105 240 2139
rect 160 2071 183 2105
rect 217 2071 240 2105
rect 320 2649 400 2680
rect 320 2601 343 2649
rect 377 2601 400 2649
rect 320 2577 400 2601
rect 320 2533 343 2577
rect 377 2533 400 2577
rect 320 2505 400 2533
rect 320 2465 343 2505
rect 377 2465 400 2505
rect 320 2433 400 2465
rect 320 2397 343 2433
rect 377 2397 400 2433
rect 320 2363 400 2397
rect 320 2327 343 2363
rect 377 2327 400 2363
rect 320 2295 400 2327
rect 320 2255 343 2295
rect 377 2255 400 2295
rect 320 2227 400 2255
rect 320 2183 343 2227
rect 377 2183 400 2227
rect 320 2159 400 2183
rect 320 2111 343 2159
rect 377 2111 400 2159
rect 320 2080 400 2111
rect 2240 2649 2320 2720
rect 2240 2601 2263 2649
rect 2297 2601 2320 2649
rect 2240 2577 2320 2601
rect 2240 2533 2263 2577
rect 2297 2533 2320 2577
rect 2240 2505 2320 2533
rect 2240 2465 2263 2505
rect 2297 2465 2320 2505
rect 2240 2433 2320 2465
rect 2240 2397 2263 2433
rect 2297 2397 2320 2433
rect 2240 2363 2320 2397
rect 2240 2327 2263 2363
rect 2297 2327 2320 2363
rect 2240 2295 2320 2327
rect 2240 2255 2263 2295
rect 2297 2255 2320 2295
rect 2240 2227 2320 2255
rect 2240 2183 2263 2227
rect 2297 2183 2320 2227
rect 2240 2159 2320 2183
rect 2240 2111 2263 2159
rect 2297 2111 2320 2159
rect 2240 2080 2320 2111
rect 4160 2649 4240 2680
rect 4160 2601 4183 2649
rect 4217 2601 4240 2649
rect 4160 2577 4240 2601
rect 4160 2533 4183 2577
rect 4217 2533 4240 2577
rect 4160 2505 4240 2533
rect 4160 2465 4183 2505
rect 4217 2465 4240 2505
rect 4160 2433 4240 2465
rect 4160 2397 4183 2433
rect 4217 2397 4240 2433
rect 4160 2363 4240 2397
rect 4160 2327 4183 2363
rect 4217 2327 4240 2363
rect 4160 2295 4240 2327
rect 4160 2255 4183 2295
rect 4217 2255 4240 2295
rect 4160 2227 4240 2255
rect 4160 2183 4183 2227
rect 4217 2183 4240 2227
rect 4160 2159 4240 2183
rect 4160 2111 4183 2159
rect 4217 2111 4240 2159
rect 4160 2080 4240 2111
rect 6080 2649 6160 2720
rect 8160 2785 8240 2819
rect 8160 2751 8183 2785
rect 8217 2751 8240 2785
rect 8160 2717 8240 2751
rect 8160 2683 8183 2717
rect 8217 2683 8240 2717
rect 6080 2601 6103 2649
rect 6137 2601 6160 2649
rect 6080 2577 6160 2601
rect 6080 2533 6103 2577
rect 6137 2533 6160 2577
rect 6080 2505 6160 2533
rect 6080 2465 6103 2505
rect 6137 2465 6160 2505
rect 6080 2433 6160 2465
rect 6080 2397 6103 2433
rect 6137 2397 6160 2433
rect 6080 2363 6160 2397
rect 6080 2327 6103 2363
rect 6137 2327 6160 2363
rect 6080 2295 6160 2327
rect 6080 2255 6103 2295
rect 6137 2255 6160 2295
rect 6080 2227 6160 2255
rect 6080 2183 6103 2227
rect 6137 2183 6160 2227
rect 6080 2159 6160 2183
rect 6080 2111 6103 2159
rect 6137 2111 6160 2159
rect 6080 2080 6160 2111
rect 8000 2649 8080 2680
rect 8000 2601 8023 2649
rect 8057 2601 8080 2649
rect 8000 2577 8080 2601
rect 8000 2533 8023 2577
rect 8057 2533 8080 2577
rect 8000 2505 8080 2533
rect 8000 2465 8023 2505
rect 8057 2465 8080 2505
rect 8000 2433 8080 2465
rect 8000 2397 8023 2433
rect 8057 2397 8080 2433
rect 8000 2363 8080 2397
rect 8000 2327 8023 2363
rect 8057 2327 8080 2363
rect 8000 2295 8080 2327
rect 8000 2255 8023 2295
rect 8057 2255 8080 2295
rect 8000 2227 8080 2255
rect 8000 2183 8023 2227
rect 8057 2183 8080 2227
rect 8000 2159 8080 2183
rect 8000 2111 8023 2159
rect 8057 2111 8080 2159
rect 8000 2080 8080 2111
rect 8160 2649 8240 2683
rect 8160 2615 8183 2649
rect 8217 2615 8240 2649
rect 8160 2581 8240 2615
rect 8160 2547 8183 2581
rect 8217 2547 8240 2581
rect 8160 2513 8240 2547
rect 8160 2479 8183 2513
rect 8217 2479 8240 2513
rect 8160 2445 8240 2479
rect 8160 2411 8183 2445
rect 8217 2411 8240 2445
rect 8160 2377 8240 2411
rect 8160 2343 8183 2377
rect 8217 2343 8240 2377
rect 8160 2309 8240 2343
rect 8160 2275 8183 2309
rect 8217 2275 8240 2309
rect 8160 2241 8240 2275
rect 8160 2207 8183 2241
rect 8217 2207 8240 2241
rect 8160 2173 8240 2207
rect 8160 2139 8183 2173
rect 8217 2139 8240 2173
rect 8160 2105 8240 2139
rect 160 2037 240 2071
rect 160 2003 183 2037
rect 217 2003 240 2037
rect 160 1969 240 2003
rect 8160 2071 8183 2105
rect 8217 2071 8240 2105
rect 8160 2037 8240 2071
rect 8160 2003 8183 2037
rect 8217 2003 8240 2037
rect 160 1935 183 1969
rect 217 1935 240 1969
rect 160 1840 240 1935
rect 520 1977 2120 2000
rect 520 1943 547 1977
rect 589 1943 619 1977
rect 657 1943 691 1977
rect 725 1943 759 1977
rect 797 1943 827 1977
rect 869 1943 895 1977
rect 941 1943 963 1977
rect 1013 1943 1031 1977
rect 1085 1943 1099 1977
rect 1157 1943 1167 1977
rect 1229 1943 1235 1977
rect 1301 1943 1303 1977
rect 1337 1943 1339 1977
rect 1405 1943 1411 1977
rect 1473 1943 1483 1977
rect 1541 1943 1555 1977
rect 1609 1943 1627 1977
rect 1677 1943 1699 1977
rect 1745 1943 1771 1977
rect 1813 1943 1843 1977
rect 1881 1943 1915 1977
rect 1949 1943 1983 1977
rect 2021 1943 2051 1977
rect 2093 1943 2120 1977
rect 520 1920 2120 1943
rect 2440 1977 4040 2000
rect 2440 1943 2467 1977
rect 2509 1943 2539 1977
rect 2577 1943 2611 1977
rect 2645 1943 2679 1977
rect 2717 1943 2747 1977
rect 2789 1943 2815 1977
rect 2861 1943 2883 1977
rect 2933 1943 2951 1977
rect 3005 1943 3019 1977
rect 3077 1943 3087 1977
rect 3149 1943 3155 1977
rect 3221 1943 3223 1977
rect 3257 1943 3259 1977
rect 3325 1943 3331 1977
rect 3393 1943 3403 1977
rect 3461 1943 3475 1977
rect 3529 1943 3547 1977
rect 3597 1943 3619 1977
rect 3665 1943 3691 1977
rect 3733 1943 3763 1977
rect 3801 1943 3835 1977
rect 3869 1943 3903 1977
rect 3941 1943 3971 1977
rect 4013 1943 4040 1977
rect 2440 1920 4040 1943
rect 4360 1977 5960 2000
rect 4360 1943 4387 1977
rect 4429 1943 4459 1977
rect 4497 1943 4531 1977
rect 4565 1943 4599 1977
rect 4637 1943 4667 1977
rect 4709 1943 4735 1977
rect 4781 1943 4803 1977
rect 4853 1943 4871 1977
rect 4925 1943 4939 1977
rect 4997 1943 5007 1977
rect 5069 1943 5075 1977
rect 5141 1943 5143 1977
rect 5177 1943 5179 1977
rect 5245 1943 5251 1977
rect 5313 1943 5323 1977
rect 5381 1943 5395 1977
rect 5449 1943 5467 1977
rect 5517 1943 5539 1977
rect 5585 1943 5611 1977
rect 5653 1943 5683 1977
rect 5721 1943 5755 1977
rect 5789 1943 5823 1977
rect 5861 1943 5891 1977
rect 5933 1943 5960 1977
rect 4360 1920 5960 1943
rect 6280 1977 7880 2000
rect 6280 1943 6307 1977
rect 6349 1943 6379 1977
rect 6417 1943 6451 1977
rect 6485 1943 6519 1977
rect 6557 1943 6587 1977
rect 6629 1943 6655 1977
rect 6701 1943 6723 1977
rect 6773 1943 6791 1977
rect 6845 1943 6859 1977
rect 6917 1943 6927 1977
rect 6989 1943 6995 1977
rect 7061 1943 7063 1977
rect 7097 1943 7099 1977
rect 7165 1943 7171 1977
rect 7233 1943 7243 1977
rect 7301 1943 7315 1977
rect 7369 1943 7387 1977
rect 7437 1943 7459 1977
rect 7505 1943 7531 1977
rect 7573 1943 7603 1977
rect 7641 1943 7675 1977
rect 7709 1943 7743 1977
rect 7781 1943 7811 1977
rect 7853 1943 7880 1977
rect 6280 1920 7880 1943
rect 8160 1969 8240 2003
rect 8160 1935 8183 1969
rect 8217 1935 8240 1969
rect 8160 1840 8240 1935
rect 160 1817 8240 1840
rect 160 1783 307 1817
rect 341 1783 375 1817
rect 409 1783 443 1817
rect 477 1783 511 1817
rect 545 1783 579 1817
rect 613 1783 647 1817
rect 681 1783 715 1817
rect 749 1783 783 1817
rect 817 1783 851 1817
rect 885 1783 919 1817
rect 953 1783 987 1817
rect 1021 1783 1055 1817
rect 1089 1783 1123 1817
rect 1157 1783 1191 1817
rect 1225 1783 1259 1817
rect 1293 1783 1327 1817
rect 1361 1783 1395 1817
rect 1429 1783 1463 1817
rect 1497 1783 1531 1817
rect 1565 1783 1599 1817
rect 1633 1783 1667 1817
rect 1701 1783 1735 1817
rect 1769 1783 1803 1817
rect 1837 1783 1871 1817
rect 1905 1783 1939 1817
rect 1973 1783 2007 1817
rect 2041 1783 2075 1817
rect 2109 1783 2143 1817
rect 2177 1783 2211 1817
rect 2245 1783 2279 1817
rect 2313 1783 2347 1817
rect 2381 1783 2415 1817
rect 2449 1783 2483 1817
rect 2517 1783 2551 1817
rect 2585 1783 2619 1817
rect 2653 1783 2687 1817
rect 2721 1783 2755 1817
rect 2789 1783 2823 1817
rect 2857 1783 2891 1817
rect 2925 1783 2959 1817
rect 2993 1783 3027 1817
rect 3061 1783 3095 1817
rect 3129 1783 3163 1817
rect 3197 1783 3231 1817
rect 3265 1783 3299 1817
rect 3333 1783 3367 1817
rect 3401 1783 3435 1817
rect 3469 1783 3503 1817
rect 3537 1783 3571 1817
rect 3605 1783 3639 1817
rect 3673 1783 3707 1817
rect 3741 1783 3775 1817
rect 3809 1783 3843 1817
rect 3877 1783 3911 1817
rect 3945 1783 3979 1817
rect 4013 1783 4047 1817
rect 4081 1783 4115 1817
rect 4149 1783 4183 1817
rect 4217 1783 4251 1817
rect 4285 1783 4319 1817
rect 4353 1783 4387 1817
rect 4421 1783 4455 1817
rect 4489 1783 4523 1817
rect 4557 1783 4591 1817
rect 4625 1783 4659 1817
rect 4693 1783 4727 1817
rect 4761 1783 4795 1817
rect 4829 1783 4863 1817
rect 4897 1783 4931 1817
rect 4965 1783 4999 1817
rect 5033 1783 5067 1817
rect 5101 1783 5135 1817
rect 5169 1783 5203 1817
rect 5237 1783 5271 1817
rect 5305 1783 5339 1817
rect 5373 1783 5407 1817
rect 5441 1783 5475 1817
rect 5509 1783 5543 1817
rect 5577 1783 5611 1817
rect 5645 1783 5679 1817
rect 5713 1783 5747 1817
rect 5781 1783 5815 1817
rect 5849 1783 5883 1817
rect 5917 1783 5951 1817
rect 5985 1783 6019 1817
rect 6053 1783 6087 1817
rect 6121 1783 6155 1817
rect 6189 1783 6223 1817
rect 6257 1783 6291 1817
rect 6325 1783 6359 1817
rect 6393 1783 6427 1817
rect 6461 1783 6495 1817
rect 6529 1783 6563 1817
rect 6597 1783 6631 1817
rect 6665 1783 6699 1817
rect 6733 1783 6767 1817
rect 6801 1783 6835 1817
rect 6869 1783 6903 1817
rect 6937 1783 6971 1817
rect 7005 1783 7039 1817
rect 7073 1783 7107 1817
rect 7141 1783 7175 1817
rect 7209 1783 7243 1817
rect 7277 1783 7311 1817
rect 7345 1783 7379 1817
rect 7413 1783 7447 1817
rect 7481 1783 7515 1817
rect 7549 1783 7583 1817
rect 7617 1783 7651 1817
rect 7685 1783 7719 1817
rect 7753 1783 7787 1817
rect 7821 1783 7855 1817
rect 7889 1783 7923 1817
rect 7957 1783 7991 1817
rect 8025 1783 8059 1817
rect 8093 1783 8240 1817
rect 160 1760 8240 1783
rect 8320 3581 8343 3615
rect 8377 3581 8400 3615
rect 8320 3547 8400 3581
rect 8320 3513 8343 3547
rect 8377 3513 8400 3547
rect 8320 3479 8400 3513
rect 8320 3445 8343 3479
rect 8377 3445 8400 3479
rect 8320 3411 8400 3445
rect 8320 3377 8343 3411
rect 8377 3377 8400 3411
rect 8320 3343 8400 3377
rect 8320 3309 8343 3343
rect 8377 3309 8400 3343
rect 8320 3275 8400 3309
rect 8320 3241 8343 3275
rect 8377 3241 8400 3275
rect 8320 3207 8400 3241
rect 8320 3173 8343 3207
rect 8377 3173 8400 3207
rect 8320 3139 8400 3173
rect 8320 3105 8343 3139
rect 8377 3105 8400 3139
rect 8320 3071 8400 3105
rect 8320 3037 8343 3071
rect 8377 3037 8400 3071
rect 8320 3003 8400 3037
rect 8320 2969 8343 3003
rect 8377 2969 8400 3003
rect 8320 2935 8400 2969
rect 8320 2901 8343 2935
rect 8377 2901 8400 2935
rect 8320 2867 8400 2901
rect 8320 2833 8343 2867
rect 8377 2833 8400 2867
rect 8320 2799 8400 2833
rect 8320 2765 8343 2799
rect 8377 2765 8400 2799
rect 8320 2731 8400 2765
rect 8320 2697 8343 2731
rect 8377 2697 8400 2731
rect 8320 2663 8400 2697
rect 8320 2629 8343 2663
rect 8377 2629 8400 2663
rect 8320 2595 8400 2629
rect 8320 2561 8343 2595
rect 8377 2561 8400 2595
rect 8320 2527 8400 2561
rect 8320 2493 8343 2527
rect 8377 2493 8400 2527
rect 8320 2459 8400 2493
rect 8320 2425 8343 2459
rect 8377 2425 8400 2459
rect 8320 2391 8400 2425
rect 8320 2357 8343 2391
rect 8377 2357 8400 2391
rect 8320 2323 8400 2357
rect 8320 2289 8343 2323
rect 8377 2289 8400 2323
rect 8320 2255 8400 2289
rect 8320 2221 8343 2255
rect 8377 2221 8400 2255
rect 8320 2187 8400 2221
rect 8320 2153 8343 2187
rect 8377 2153 8400 2187
rect 8320 2119 8400 2153
rect 8320 2085 8343 2119
rect 8377 2085 8400 2119
rect 8320 2051 8400 2085
rect 8320 2017 8343 2051
rect 8377 2017 8400 2051
rect 8320 1983 8400 2017
rect 8320 1949 8343 1983
rect 8377 1949 8400 1983
rect 8320 1915 8400 1949
rect 8320 1881 8343 1915
rect 8377 1881 8400 1915
rect 8320 1847 8400 1881
rect 8320 1813 8343 1847
rect 8377 1813 8400 1847
rect 8320 1779 8400 1813
rect 0 1680 80 1745
rect 8320 1745 8343 1779
rect 8377 1745 8400 1779
rect 8320 1680 8400 1745
rect 0 1657 8400 1680
rect 0 1623 137 1657
rect 171 1623 205 1657
rect 239 1623 273 1657
rect 307 1623 341 1657
rect 375 1623 409 1657
rect 443 1623 477 1657
rect 511 1623 545 1657
rect 579 1623 613 1657
rect 647 1623 681 1657
rect 715 1623 749 1657
rect 783 1623 817 1657
rect 851 1623 885 1657
rect 919 1623 953 1657
rect 987 1623 1021 1657
rect 1055 1623 1089 1657
rect 1123 1623 1157 1657
rect 1191 1623 1225 1657
rect 1259 1623 1293 1657
rect 1327 1623 1361 1657
rect 1395 1623 1429 1657
rect 1463 1623 1497 1657
rect 1531 1623 1565 1657
rect 1599 1623 1633 1657
rect 1667 1623 1701 1657
rect 1735 1623 1769 1657
rect 1803 1623 1837 1657
rect 1871 1623 1905 1657
rect 1939 1623 1973 1657
rect 2007 1623 2041 1657
rect 2075 1623 2109 1657
rect 2143 1623 2177 1657
rect 2211 1623 2245 1657
rect 2279 1623 2313 1657
rect 2347 1623 2381 1657
rect 2415 1623 2449 1657
rect 2483 1623 2517 1657
rect 2551 1623 2585 1657
rect 2619 1623 2653 1657
rect 2687 1623 2721 1657
rect 2755 1623 2789 1657
rect 2823 1623 2857 1657
rect 2891 1623 2925 1657
rect 2959 1623 2993 1657
rect 3027 1623 3061 1657
rect 3095 1623 3129 1657
rect 3163 1623 3197 1657
rect 3231 1623 3265 1657
rect 3299 1623 3333 1657
rect 3367 1623 3401 1657
rect 3435 1623 3469 1657
rect 3503 1623 3537 1657
rect 3571 1623 3605 1657
rect 3639 1623 3673 1657
rect 3707 1623 3741 1657
rect 3775 1623 3809 1657
rect 3843 1623 3877 1657
rect 3911 1623 3945 1657
rect 3979 1623 4013 1657
rect 4047 1623 4081 1657
rect 4115 1623 4149 1657
rect 4183 1623 4217 1657
rect 4251 1623 4285 1657
rect 4319 1623 4353 1657
rect 4387 1623 4421 1657
rect 4455 1623 4489 1657
rect 4523 1623 4557 1657
rect 4591 1623 4625 1657
rect 4659 1623 4693 1657
rect 4727 1623 4761 1657
rect 4795 1623 4829 1657
rect 4863 1623 4897 1657
rect 4931 1623 4965 1657
rect 4999 1623 5033 1657
rect 5067 1623 5101 1657
rect 5135 1623 5169 1657
rect 5203 1623 5237 1657
rect 5271 1623 5305 1657
rect 5339 1623 5373 1657
rect 5407 1623 5441 1657
rect 5475 1623 5509 1657
rect 5543 1623 5577 1657
rect 5611 1623 5645 1657
rect 5679 1623 5713 1657
rect 5747 1623 5781 1657
rect 5815 1623 5849 1657
rect 5883 1623 5917 1657
rect 5951 1623 5985 1657
rect 6019 1623 6053 1657
rect 6087 1623 6121 1657
rect 6155 1623 6189 1657
rect 6223 1623 6257 1657
rect 6291 1623 6325 1657
rect 6359 1623 6393 1657
rect 6427 1623 6461 1657
rect 6495 1623 6529 1657
rect 6563 1623 6597 1657
rect 6631 1623 6665 1657
rect 6699 1623 6733 1657
rect 6767 1623 6801 1657
rect 6835 1623 6869 1657
rect 6903 1623 6937 1657
rect 6971 1623 7005 1657
rect 7039 1623 7073 1657
rect 7107 1623 7141 1657
rect 7175 1623 7209 1657
rect 7243 1623 7277 1657
rect 7311 1623 7345 1657
rect 7379 1623 7413 1657
rect 7447 1623 7481 1657
rect 7515 1623 7549 1657
rect 7583 1623 7617 1657
rect 7651 1623 7685 1657
rect 7719 1623 7753 1657
rect 7787 1623 7821 1657
rect 7855 1623 7889 1657
rect 7923 1623 7957 1657
rect 7991 1623 8025 1657
rect 8059 1623 8093 1657
rect 8127 1623 8161 1657
rect 8195 1623 8229 1657
rect 8263 1623 8400 1657
rect 0 1600 8400 1623
rect 0 1040 80 1600
rect 160 1337 240 1520
rect 160 1303 183 1337
rect 217 1303 240 1337
rect 160 1120 240 1303
rect 480 1337 560 1520
rect 480 1303 503 1337
rect 537 1303 560 1337
rect 480 1120 560 1303
rect 640 1337 720 1520
rect 640 1303 663 1337
rect 697 1303 720 1337
rect 640 1120 720 1303
rect 800 1337 880 1520
rect 800 1303 823 1337
rect 857 1303 880 1337
rect 800 1120 880 1303
rect 960 1337 1040 1520
rect 960 1303 983 1337
rect 1017 1303 1040 1337
rect 960 1120 1040 1303
rect 1120 1337 1200 1520
rect 1120 1303 1143 1337
rect 1177 1303 1200 1337
rect 1120 1120 1200 1303
rect 1440 1337 1520 1520
rect 1440 1303 1463 1337
rect 1497 1303 1520 1337
rect 1440 1120 1520 1303
rect 1600 1337 1680 1520
rect 1600 1303 1623 1337
rect 1657 1303 1680 1337
rect 1600 1120 1680 1303
rect 1760 1337 1840 1520
rect 1760 1303 1783 1337
rect 1817 1303 1840 1337
rect 1760 1120 1840 1303
rect 1920 1337 2000 1520
rect 1920 1303 1943 1337
rect 1977 1303 2000 1337
rect 1920 1120 2000 1303
rect 2080 1337 2160 1520
rect 2080 1303 2103 1337
rect 2137 1303 2160 1337
rect 2080 1120 2160 1303
rect 2240 1337 2320 1520
rect 2240 1303 2263 1337
rect 2297 1303 2320 1337
rect 2240 1120 2320 1303
rect 2400 1337 2480 1520
rect 2400 1303 2423 1337
rect 2457 1303 2480 1337
rect 2400 1120 2480 1303
rect 2560 1337 2640 1520
rect 2560 1303 2583 1337
rect 2617 1303 2640 1337
rect 2560 1120 2640 1303
rect 2720 1337 2800 1520
rect 2720 1303 2743 1337
rect 2777 1303 2800 1337
rect 2720 1120 2800 1303
rect 2880 1337 2960 1520
rect 2880 1303 2903 1337
rect 2937 1303 2960 1337
rect 2880 1120 2960 1303
rect 3040 1337 3120 1520
rect 3040 1303 3063 1337
rect 3097 1303 3120 1337
rect 3040 1120 3120 1303
rect 3360 1337 3440 1520
rect 3360 1303 3383 1337
rect 3417 1303 3440 1337
rect 3360 1120 3440 1303
rect 3520 1337 3600 1520
rect 3520 1303 3543 1337
rect 3577 1303 3600 1337
rect 3520 1120 3600 1303
rect 3680 1337 3760 1520
rect 3680 1303 3703 1337
rect 3737 1303 3760 1337
rect 3680 1120 3760 1303
rect 3840 1337 3920 1520
rect 3840 1303 3863 1337
rect 3897 1303 3920 1337
rect 3840 1120 3920 1303
rect 4000 1337 4080 1520
rect 4000 1303 4023 1337
rect 4057 1303 4080 1337
rect 4000 1120 4080 1303
rect 4320 1337 4400 1520
rect 4320 1303 4343 1337
rect 4377 1303 4400 1337
rect 4320 1120 4400 1303
rect 4480 1337 4560 1520
rect 4480 1303 4503 1337
rect 4537 1303 4560 1337
rect 4480 1120 4560 1303
rect 4640 1337 4720 1520
rect 4640 1303 4663 1337
rect 4697 1303 4720 1337
rect 4640 1120 4720 1303
rect 4800 1337 4880 1520
rect 4800 1303 4823 1337
rect 4857 1303 4880 1337
rect 4800 1120 4880 1303
rect 4960 1337 5040 1520
rect 4960 1303 4983 1337
rect 5017 1303 5040 1337
rect 4960 1120 5040 1303
rect 5280 1337 5360 1520
rect 5280 1303 5303 1337
rect 5337 1303 5360 1337
rect 5280 1120 5360 1303
rect 5440 1337 5520 1520
rect 5440 1303 5463 1337
rect 5497 1303 5520 1337
rect 5440 1120 5520 1303
rect 5600 1337 5680 1520
rect 5600 1303 5623 1337
rect 5657 1303 5680 1337
rect 5600 1120 5680 1303
rect 5760 1337 5840 1520
rect 5760 1303 5783 1337
rect 5817 1303 5840 1337
rect 5760 1120 5840 1303
rect 5920 1337 6000 1520
rect 5920 1303 5943 1337
rect 5977 1303 6000 1337
rect 5920 1120 6000 1303
rect 6080 1337 6160 1520
rect 6080 1303 6103 1337
rect 6137 1303 6160 1337
rect 6080 1120 6160 1303
rect 6240 1337 6320 1520
rect 6240 1303 6263 1337
rect 6297 1303 6320 1337
rect 6240 1120 6320 1303
rect 6400 1337 6480 1520
rect 6400 1303 6423 1337
rect 6457 1303 6480 1337
rect 6400 1120 6480 1303
rect 6560 1337 6640 1520
rect 6560 1303 6583 1337
rect 6617 1303 6640 1337
rect 6560 1120 6640 1303
rect 6720 1337 6800 1520
rect 6720 1303 6743 1337
rect 6777 1303 6800 1337
rect 6720 1120 6800 1303
rect 6880 1337 6960 1520
rect 6880 1303 6903 1337
rect 6937 1303 6960 1337
rect 6880 1120 6960 1303
rect 7200 1337 7280 1520
rect 7200 1303 7223 1337
rect 7257 1303 7280 1337
rect 7200 1120 7280 1303
rect 7360 1337 7440 1520
rect 7360 1303 7383 1337
rect 7417 1303 7440 1337
rect 7360 1120 7440 1303
rect 7520 1337 7600 1520
rect 7520 1303 7543 1337
rect 7577 1303 7600 1337
rect 7520 1120 7600 1303
rect 7680 1337 7760 1520
rect 7680 1303 7703 1337
rect 7737 1303 7760 1337
rect 7680 1120 7760 1303
rect 7840 1337 7920 1520
rect 7840 1303 7863 1337
rect 7897 1303 7920 1337
rect 7840 1120 7920 1303
rect 8160 1337 8240 1520
rect 8160 1303 8183 1337
rect 8217 1303 8240 1337
rect 8160 1120 8240 1303
rect 8320 1040 8400 1600
rect 0 1017 8400 1040
rect 0 983 137 1017
rect 171 983 205 1017
rect 239 983 273 1017
rect 307 983 341 1017
rect 375 983 409 1017
rect 443 983 477 1017
rect 511 983 545 1017
rect 579 983 613 1017
rect 647 983 681 1017
rect 715 983 749 1017
rect 783 983 817 1017
rect 851 983 885 1017
rect 919 983 953 1017
rect 987 983 1021 1017
rect 1055 983 1089 1017
rect 1123 983 1157 1017
rect 1191 983 1225 1017
rect 1259 983 1293 1017
rect 1327 983 1361 1017
rect 1395 983 1429 1017
rect 1463 983 1497 1017
rect 1531 983 1565 1017
rect 1599 983 1633 1017
rect 1667 983 1701 1017
rect 1735 983 1769 1017
rect 1803 983 1837 1017
rect 1871 983 1905 1017
rect 1939 983 1973 1017
rect 2007 983 2041 1017
rect 2075 983 2109 1017
rect 2143 983 2177 1017
rect 2211 983 2245 1017
rect 2279 983 2313 1017
rect 2347 983 2381 1017
rect 2415 983 2449 1017
rect 2483 983 2517 1017
rect 2551 983 2585 1017
rect 2619 983 2653 1017
rect 2687 983 2721 1017
rect 2755 983 2789 1017
rect 2823 983 2857 1017
rect 2891 983 2925 1017
rect 2959 983 2993 1017
rect 3027 983 3061 1017
rect 3095 983 3129 1017
rect 3163 983 3197 1017
rect 3231 983 3265 1017
rect 3299 983 3333 1017
rect 3367 983 3401 1017
rect 3435 983 3469 1017
rect 3503 983 3537 1017
rect 3571 983 3605 1017
rect 3639 983 3673 1017
rect 3707 983 3741 1017
rect 3775 983 3809 1017
rect 3843 983 3877 1017
rect 3911 983 3945 1017
rect 3979 983 4013 1017
rect 4047 983 4081 1017
rect 4115 983 4149 1017
rect 4183 983 4217 1017
rect 4251 983 4285 1017
rect 4319 983 4353 1017
rect 4387 983 4421 1017
rect 4455 983 4489 1017
rect 4523 983 4557 1017
rect 4591 983 4625 1017
rect 4659 983 4693 1017
rect 4727 983 4761 1017
rect 4795 983 4829 1017
rect 4863 983 4897 1017
rect 4931 983 4965 1017
rect 4999 983 5033 1017
rect 5067 983 5101 1017
rect 5135 983 5169 1017
rect 5203 983 5237 1017
rect 5271 983 5305 1017
rect 5339 983 5373 1017
rect 5407 983 5441 1017
rect 5475 983 5509 1017
rect 5543 983 5577 1017
rect 5611 983 5645 1017
rect 5679 983 5713 1017
rect 5747 983 5781 1017
rect 5815 983 5849 1017
rect 5883 983 5917 1017
rect 5951 983 5985 1017
rect 6019 983 6053 1017
rect 6087 983 6121 1017
rect 6155 983 6189 1017
rect 6223 983 6257 1017
rect 6291 983 6325 1017
rect 6359 983 6393 1017
rect 6427 983 6461 1017
rect 6495 983 6529 1017
rect 6563 983 6597 1017
rect 6631 983 6665 1017
rect 6699 983 6733 1017
rect 6767 983 6801 1017
rect 6835 983 6869 1017
rect 6903 983 6937 1017
rect 6971 983 7005 1017
rect 7039 983 7073 1017
rect 7107 983 7141 1017
rect 7175 983 7209 1017
rect 7243 983 7277 1017
rect 7311 983 7345 1017
rect 7379 983 7413 1017
rect 7447 983 7481 1017
rect 7515 983 7549 1017
rect 7583 983 7617 1017
rect 7651 983 7685 1017
rect 7719 983 7753 1017
rect 7787 983 7821 1017
rect 7855 983 7889 1017
rect 7923 983 7957 1017
rect 7991 983 8025 1017
rect 8059 983 8093 1017
rect 8127 983 8161 1017
rect 8195 983 8229 1017
rect 8263 983 8400 1017
rect 0 960 8400 983
rect 0 911 80 960
rect 0 877 23 911
rect 57 877 80 911
rect 8320 911 8400 960
rect 0 843 80 877
rect 0 809 23 843
rect 57 809 80 843
rect 0 775 80 809
rect 520 857 2120 880
rect 520 823 547 857
rect 589 823 619 857
rect 657 823 691 857
rect 725 823 759 857
rect 797 823 827 857
rect 869 823 895 857
rect 941 823 963 857
rect 1013 823 1031 857
rect 1085 823 1099 857
rect 1157 823 1167 857
rect 1229 823 1235 857
rect 1301 823 1303 857
rect 1337 823 1339 857
rect 1405 823 1411 857
rect 1473 823 1483 857
rect 1541 823 1555 857
rect 1609 823 1627 857
rect 1677 823 1699 857
rect 1745 823 1771 857
rect 1813 823 1843 857
rect 1881 823 1915 857
rect 1949 823 1983 857
rect 2021 823 2051 857
rect 2093 823 2120 857
rect 520 800 2120 823
rect 2440 857 4040 880
rect 2440 823 2467 857
rect 2509 823 2539 857
rect 2577 823 2611 857
rect 2645 823 2679 857
rect 2717 823 2747 857
rect 2789 823 2815 857
rect 2861 823 2883 857
rect 2933 823 2951 857
rect 3005 823 3019 857
rect 3077 823 3087 857
rect 3149 823 3155 857
rect 3221 823 3223 857
rect 3257 823 3259 857
rect 3325 823 3331 857
rect 3393 823 3403 857
rect 3461 823 3475 857
rect 3529 823 3547 857
rect 3597 823 3619 857
rect 3665 823 3691 857
rect 3733 823 3763 857
rect 3801 823 3835 857
rect 3869 823 3903 857
rect 3941 823 3971 857
rect 4013 823 4040 857
rect 2440 800 4040 823
rect 4360 857 5960 880
rect 4360 823 4387 857
rect 4429 823 4459 857
rect 4497 823 4531 857
rect 4565 823 4599 857
rect 4637 823 4667 857
rect 4709 823 4735 857
rect 4781 823 4803 857
rect 4853 823 4871 857
rect 4925 823 4939 857
rect 4997 823 5007 857
rect 5069 823 5075 857
rect 5141 823 5143 857
rect 5177 823 5179 857
rect 5245 823 5251 857
rect 5313 823 5323 857
rect 5381 823 5395 857
rect 5449 823 5467 857
rect 5517 823 5539 857
rect 5585 823 5611 857
rect 5653 823 5683 857
rect 5721 823 5755 857
rect 5789 823 5823 857
rect 5861 823 5891 857
rect 5933 823 5960 857
rect 4360 800 5960 823
rect 6280 857 7880 880
rect 6280 823 6307 857
rect 6349 823 6379 857
rect 6417 823 6451 857
rect 6485 823 6519 857
rect 6557 823 6587 857
rect 6629 823 6655 857
rect 6701 823 6723 857
rect 6773 823 6791 857
rect 6845 823 6859 857
rect 6917 823 6927 857
rect 6989 823 6995 857
rect 7061 823 7063 857
rect 7097 823 7099 857
rect 7165 823 7171 857
rect 7233 823 7243 857
rect 7301 823 7315 857
rect 7369 823 7387 857
rect 7437 823 7459 857
rect 7505 823 7531 857
rect 7573 823 7603 857
rect 7641 823 7675 857
rect 7709 823 7743 857
rect 7781 823 7811 857
rect 7853 823 7880 857
rect 6280 800 7880 823
rect 8320 877 8343 911
rect 8377 877 8400 911
rect 8320 843 8400 877
rect 8320 809 8343 843
rect 8377 809 8400 843
rect 0 741 23 775
rect 57 741 80 775
rect 8320 775 8400 809
rect 0 707 80 741
rect 0 673 23 707
rect 57 673 80 707
rect 0 639 80 673
rect 0 605 23 639
rect 57 605 80 639
rect 0 571 80 605
rect 0 537 23 571
rect 57 537 80 571
rect 320 713 400 760
rect 320 677 343 713
rect 377 677 400 713
rect 320 643 400 677
rect 320 607 343 643
rect 377 607 400 643
rect 320 560 400 607
rect 2240 713 2320 760
rect 2240 677 2263 713
rect 2297 677 2320 713
rect 2240 643 2320 677
rect 2240 607 2263 643
rect 2297 607 2320 643
rect 0 503 80 537
rect 0 469 23 503
rect 57 469 80 503
rect 0 435 80 469
rect 0 401 23 435
rect 57 401 80 435
rect 0 367 80 401
rect 2240 480 2320 607
rect 4160 713 4240 760
rect 4160 677 4183 713
rect 4217 677 4240 713
rect 4160 643 4240 677
rect 4160 607 4183 643
rect 4217 607 4240 643
rect 4160 560 4240 607
rect 6080 713 6160 760
rect 6080 677 6103 713
rect 6137 677 6160 713
rect 6080 643 6160 677
rect 6080 607 6103 643
rect 6137 607 6160 643
rect 6080 480 6160 607
rect 8000 713 8080 760
rect 8000 677 8023 713
rect 8057 677 8080 713
rect 8000 643 8080 677
rect 8000 607 8023 643
rect 8057 607 8080 643
rect 8000 560 8080 607
rect 8320 741 8343 775
rect 8377 741 8400 775
rect 8320 707 8400 741
rect 8320 673 8343 707
rect 8377 673 8400 707
rect 8320 639 8400 673
rect 8320 605 8343 639
rect 8377 605 8400 639
rect 8320 571 8400 605
rect 2240 400 6160 480
rect 8320 537 8343 571
rect 8377 537 8400 571
rect 8320 503 8400 537
rect 8320 469 8343 503
rect 8377 469 8400 503
rect 8320 435 8400 469
rect 8320 401 8343 435
rect 8377 401 8400 435
rect 0 333 23 367
rect 57 333 80 367
rect 0 299 80 333
rect 0 265 23 299
rect 57 265 80 299
rect 0 231 80 265
rect 0 197 23 231
rect 57 197 80 231
rect 0 163 80 197
rect 0 129 23 163
rect 57 129 80 163
rect 0 80 80 129
rect 320 313 400 360
rect 320 277 343 313
rect 377 277 400 313
rect 320 243 400 277
rect 320 207 343 243
rect 377 207 400 243
rect 320 80 400 207
rect 2240 313 2320 360
rect 2240 277 2263 313
rect 2297 277 2320 313
rect 2240 243 2320 277
rect 2240 207 2263 243
rect 2297 207 2320 243
rect 2240 160 2320 207
rect 4160 313 4240 400
rect 8320 367 8400 401
rect 4160 277 4183 313
rect 4217 277 4240 313
rect 4160 243 4240 277
rect 4160 207 4183 243
rect 4217 207 4240 243
rect 4160 160 4240 207
rect 6080 313 6160 360
rect 6080 277 6103 313
rect 6137 277 6160 313
rect 6080 243 6160 277
rect 6080 207 6103 243
rect 6137 207 6160 243
rect 6080 160 6160 207
rect 8000 313 8080 360
rect 8000 277 8023 313
rect 8057 277 8080 313
rect 8000 243 8080 277
rect 8000 207 8023 243
rect 8057 207 8080 243
rect 8000 80 8080 207
rect 8320 333 8343 367
rect 8377 333 8400 367
rect 8320 299 8400 333
rect 8320 265 8343 299
rect 8377 265 8400 299
rect 8320 231 8400 265
rect 8320 197 8343 231
rect 8377 197 8400 231
rect 8320 163 8400 197
rect 8320 129 8343 163
rect 8377 129 8400 163
rect 8320 80 8400 129
rect 0 57 8400 80
rect 0 23 137 57
rect 171 23 205 57
rect 239 23 273 57
rect 307 23 341 57
rect 375 23 409 57
rect 443 23 477 57
rect 511 23 545 57
rect 579 23 613 57
rect 647 23 681 57
rect 715 23 749 57
rect 783 23 817 57
rect 851 23 885 57
rect 919 23 953 57
rect 987 23 1021 57
rect 1055 23 1089 57
rect 1123 23 1157 57
rect 1191 23 1225 57
rect 1259 23 1293 57
rect 1327 23 1361 57
rect 1395 23 1429 57
rect 1463 23 1497 57
rect 1531 23 1565 57
rect 1599 23 1633 57
rect 1667 23 1701 57
rect 1735 23 1769 57
rect 1803 23 1837 57
rect 1871 23 1905 57
rect 1939 23 1973 57
rect 2007 23 2041 57
rect 2075 23 2109 57
rect 2143 23 2177 57
rect 2211 23 2245 57
rect 2279 23 2313 57
rect 2347 23 2381 57
rect 2415 23 2449 57
rect 2483 23 2517 57
rect 2551 23 2585 57
rect 2619 23 2653 57
rect 2687 23 2721 57
rect 2755 23 2789 57
rect 2823 23 2857 57
rect 2891 23 2925 57
rect 2959 23 2993 57
rect 3027 23 3061 57
rect 3095 23 3129 57
rect 3163 23 3197 57
rect 3231 23 3265 57
rect 3299 23 3333 57
rect 3367 23 3401 57
rect 3435 23 3469 57
rect 3503 23 3537 57
rect 3571 23 3605 57
rect 3639 23 3673 57
rect 3707 23 3741 57
rect 3775 23 3809 57
rect 3843 23 3877 57
rect 3911 23 3945 57
rect 3979 23 4013 57
rect 4047 23 4081 57
rect 4115 23 4149 57
rect 4183 23 4217 57
rect 4251 23 4285 57
rect 4319 23 4353 57
rect 4387 23 4421 57
rect 4455 23 4489 57
rect 4523 23 4557 57
rect 4591 23 4625 57
rect 4659 23 4693 57
rect 4727 23 4761 57
rect 4795 23 4829 57
rect 4863 23 4897 57
rect 4931 23 4965 57
rect 4999 23 5033 57
rect 5067 23 5101 57
rect 5135 23 5169 57
rect 5203 23 5237 57
rect 5271 23 5305 57
rect 5339 23 5373 57
rect 5407 23 5441 57
rect 5475 23 5509 57
rect 5543 23 5577 57
rect 5611 23 5645 57
rect 5679 23 5713 57
rect 5747 23 5781 57
rect 5815 23 5849 57
rect 5883 23 5917 57
rect 5951 23 5985 57
rect 6019 23 6053 57
rect 6087 23 6121 57
rect 6155 23 6189 57
rect 6223 23 6257 57
rect 6291 23 6325 57
rect 6359 23 6393 57
rect 6427 23 6461 57
rect 6495 23 6529 57
rect 6563 23 6597 57
rect 6631 23 6665 57
rect 6699 23 6733 57
rect 6767 23 6801 57
rect 6835 23 6869 57
rect 6903 23 6937 57
rect 6971 23 7005 57
rect 7039 23 7073 57
rect 7107 23 7141 57
rect 7175 23 7209 57
rect 7243 23 7277 57
rect 7311 23 7345 57
rect 7379 23 7413 57
rect 7447 23 7481 57
rect 7515 23 7549 57
rect 7583 23 7617 57
rect 7651 23 7685 57
rect 7719 23 7753 57
rect 7787 23 7821 57
rect 7855 23 7889 57
rect 7923 23 7957 57
rect 7991 23 8025 57
rect 8059 23 8093 57
rect 8127 23 8161 57
rect 8195 23 8229 57
rect 8263 23 8400 57
rect 0 0 8400 23
<< viali >>
rect 343 5635 377 5649
rect 343 5615 377 5635
rect 343 5567 377 5577
rect 343 5543 377 5567
rect 343 5499 377 5505
rect 343 5471 377 5499
rect 343 5431 377 5433
rect 343 5399 377 5431
rect 343 5329 377 5361
rect 343 5327 377 5329
rect 343 5261 377 5289
rect 343 5255 377 5261
rect 343 5193 377 5217
rect 343 5183 377 5193
rect 343 5125 377 5145
rect 343 5111 377 5125
rect 2263 5635 2297 5649
rect 2263 5615 2297 5635
rect 2263 5567 2297 5577
rect 2263 5543 2297 5567
rect 2263 5499 2297 5505
rect 2263 5471 2297 5499
rect 2263 5431 2297 5433
rect 2263 5399 2297 5431
rect 2263 5329 2297 5361
rect 2263 5327 2297 5329
rect 2263 5261 2297 5289
rect 2263 5255 2297 5261
rect 2263 5193 2297 5217
rect 2263 5183 2297 5193
rect 2263 5125 2297 5145
rect 2263 5111 2297 5125
rect 4183 5635 4217 5649
rect 4183 5615 4217 5635
rect 4183 5567 4217 5577
rect 4183 5543 4217 5567
rect 4183 5499 4217 5505
rect 4183 5471 4217 5499
rect 4183 5431 4217 5433
rect 4183 5399 4217 5431
rect 4183 5329 4217 5361
rect 4183 5327 4217 5329
rect 4183 5261 4217 5289
rect 4183 5255 4217 5261
rect 4183 5193 4217 5217
rect 4183 5183 4217 5193
rect 4183 5125 4217 5145
rect 4183 5111 4217 5125
rect 6103 5635 6137 5649
rect 6103 5615 6137 5635
rect 6103 5567 6137 5577
rect 6103 5543 6137 5567
rect 6103 5499 6137 5505
rect 6103 5471 6137 5499
rect 6103 5431 6137 5433
rect 6103 5399 6137 5431
rect 6103 5329 6137 5361
rect 6103 5327 6137 5329
rect 6103 5261 6137 5289
rect 6103 5255 6137 5261
rect 6103 5193 6137 5217
rect 6103 5183 6137 5193
rect 6103 5125 6137 5145
rect 6103 5111 6137 5125
rect 8023 5635 8057 5649
rect 8023 5615 8057 5635
rect 8023 5567 8057 5577
rect 8023 5543 8057 5567
rect 8023 5499 8057 5505
rect 8023 5471 8057 5499
rect 8023 5431 8057 5433
rect 8023 5399 8057 5431
rect 8023 5329 8057 5361
rect 8023 5327 8057 5329
rect 8023 5261 8057 5289
rect 8023 5255 8057 5261
rect 8023 5193 8057 5217
rect 8023 5183 8057 5193
rect 8023 5125 8057 5145
rect 8023 5111 8057 5125
rect 343 4875 377 4889
rect 343 4855 377 4875
rect 343 4807 377 4817
rect 343 4783 377 4807
rect 343 4739 377 4745
rect 343 4711 377 4739
rect 343 4671 377 4673
rect 343 4639 377 4671
rect 343 4569 377 4601
rect 343 4567 377 4569
rect 343 4501 377 4529
rect 343 4495 377 4501
rect 343 4433 377 4457
rect 343 4423 377 4433
rect 343 4365 377 4385
rect 343 4351 377 4365
rect 2263 4875 2297 4889
rect 2263 4855 2297 4875
rect 2263 4807 2297 4817
rect 2263 4783 2297 4807
rect 2263 4739 2297 4745
rect 2263 4711 2297 4739
rect 2263 4671 2297 4673
rect 2263 4639 2297 4671
rect 2263 4569 2297 4601
rect 2263 4567 2297 4569
rect 2263 4501 2297 4529
rect 2263 4495 2297 4501
rect 2263 4433 2297 4457
rect 2263 4423 2297 4433
rect 2263 4365 2297 4385
rect 2263 4351 2297 4365
rect 4183 4875 4217 4889
rect 4183 4855 4217 4875
rect 4183 4807 4217 4817
rect 4183 4783 4217 4807
rect 4183 4739 4217 4745
rect 4183 4711 4217 4739
rect 4183 4671 4217 4673
rect 4183 4639 4217 4671
rect 4183 4569 4217 4601
rect 4183 4567 4217 4569
rect 4183 4501 4217 4529
rect 4183 4495 4217 4501
rect 4183 4433 4217 4457
rect 4183 4423 4217 4433
rect 4183 4365 4217 4385
rect 4183 4351 4217 4365
rect 6103 4875 6137 4889
rect 6103 4855 6137 4875
rect 6103 4807 6137 4817
rect 6103 4783 6137 4807
rect 6103 4739 6137 4745
rect 6103 4711 6137 4739
rect 6103 4671 6137 4673
rect 6103 4639 6137 4671
rect 6103 4569 6137 4601
rect 6103 4567 6137 4569
rect 6103 4501 6137 4529
rect 6103 4495 6137 4501
rect 6103 4433 6137 4457
rect 6103 4423 6137 4433
rect 6103 4365 6137 4385
rect 6103 4351 6137 4365
rect 8023 4875 8057 4889
rect 8023 4855 8057 4875
rect 8023 4807 8057 4817
rect 8023 4783 8057 4807
rect 8023 4739 8057 4745
rect 8023 4711 8057 4739
rect 8023 4671 8057 4673
rect 8023 4639 8057 4671
rect 8023 4569 8057 4601
rect 8023 4567 8057 4569
rect 8023 4501 8057 4529
rect 8023 4495 8057 4501
rect 8023 4433 8057 4457
rect 8023 4423 8057 4433
rect 8023 4365 8057 4385
rect 8023 4351 8057 4365
rect 547 4183 555 4217
rect 555 4183 581 4217
rect 619 4183 623 4217
rect 623 4183 653 4217
rect 691 4183 725 4217
rect 763 4183 793 4217
rect 793 4183 797 4217
rect 835 4183 861 4217
rect 861 4183 869 4217
rect 907 4183 929 4217
rect 929 4183 941 4217
rect 979 4183 997 4217
rect 997 4183 1013 4217
rect 1051 4183 1065 4217
rect 1065 4183 1085 4217
rect 1123 4183 1133 4217
rect 1133 4183 1157 4217
rect 1195 4183 1201 4217
rect 1201 4183 1229 4217
rect 1267 4183 1269 4217
rect 1269 4183 1301 4217
rect 1339 4183 1371 4217
rect 1371 4183 1373 4217
rect 1411 4183 1439 4217
rect 1439 4183 1445 4217
rect 1483 4183 1507 4217
rect 1507 4183 1517 4217
rect 1555 4183 1575 4217
rect 1575 4183 1589 4217
rect 1627 4183 1643 4217
rect 1643 4183 1661 4217
rect 1699 4183 1711 4217
rect 1711 4183 1733 4217
rect 1771 4183 1779 4217
rect 1779 4183 1805 4217
rect 1843 4183 1847 4217
rect 1847 4183 1877 4217
rect 1915 4183 1949 4217
rect 1987 4183 2017 4217
rect 2017 4183 2021 4217
rect 2059 4183 2085 4217
rect 2085 4183 2093 4217
rect 2467 4183 2475 4217
rect 2475 4183 2501 4217
rect 2539 4183 2543 4217
rect 2543 4183 2573 4217
rect 2611 4183 2645 4217
rect 2683 4183 2713 4217
rect 2713 4183 2717 4217
rect 2755 4183 2781 4217
rect 2781 4183 2789 4217
rect 2827 4183 2849 4217
rect 2849 4183 2861 4217
rect 2899 4183 2917 4217
rect 2917 4183 2933 4217
rect 2971 4183 2985 4217
rect 2985 4183 3005 4217
rect 3043 4183 3053 4217
rect 3053 4183 3077 4217
rect 3115 4183 3121 4217
rect 3121 4183 3149 4217
rect 3187 4183 3189 4217
rect 3189 4183 3221 4217
rect 3259 4183 3291 4217
rect 3291 4183 3293 4217
rect 3331 4183 3359 4217
rect 3359 4183 3365 4217
rect 3403 4183 3427 4217
rect 3427 4183 3437 4217
rect 3475 4183 3495 4217
rect 3495 4183 3509 4217
rect 3547 4183 3563 4217
rect 3563 4183 3581 4217
rect 3619 4183 3631 4217
rect 3631 4183 3653 4217
rect 3691 4183 3699 4217
rect 3699 4183 3725 4217
rect 3763 4183 3767 4217
rect 3767 4183 3797 4217
rect 3835 4183 3869 4217
rect 3907 4183 3937 4217
rect 3937 4183 3941 4217
rect 3979 4183 4005 4217
rect 4005 4183 4013 4217
rect 4387 4183 4395 4217
rect 4395 4183 4421 4217
rect 4459 4183 4463 4217
rect 4463 4183 4493 4217
rect 4531 4183 4565 4217
rect 4603 4183 4633 4217
rect 4633 4183 4637 4217
rect 4675 4183 4701 4217
rect 4701 4183 4709 4217
rect 4747 4183 4769 4217
rect 4769 4183 4781 4217
rect 4819 4183 4837 4217
rect 4837 4183 4853 4217
rect 4891 4183 4905 4217
rect 4905 4183 4925 4217
rect 4963 4183 4973 4217
rect 4973 4183 4997 4217
rect 5035 4183 5041 4217
rect 5041 4183 5069 4217
rect 5107 4183 5109 4217
rect 5109 4183 5141 4217
rect 5179 4183 5211 4217
rect 5211 4183 5213 4217
rect 5251 4183 5279 4217
rect 5279 4183 5285 4217
rect 5323 4183 5347 4217
rect 5347 4183 5357 4217
rect 5395 4183 5415 4217
rect 5415 4183 5429 4217
rect 5467 4183 5483 4217
rect 5483 4183 5501 4217
rect 5539 4183 5551 4217
rect 5551 4183 5573 4217
rect 5611 4183 5619 4217
rect 5619 4183 5645 4217
rect 5683 4183 5687 4217
rect 5687 4183 5717 4217
rect 5755 4183 5789 4217
rect 5827 4183 5857 4217
rect 5857 4183 5861 4217
rect 5899 4183 5925 4217
rect 5925 4183 5933 4217
rect 6307 4183 6315 4217
rect 6315 4183 6341 4217
rect 6379 4183 6383 4217
rect 6383 4183 6413 4217
rect 6451 4183 6485 4217
rect 6523 4183 6553 4217
rect 6553 4183 6557 4217
rect 6595 4183 6621 4217
rect 6621 4183 6629 4217
rect 6667 4183 6689 4217
rect 6689 4183 6701 4217
rect 6739 4183 6757 4217
rect 6757 4183 6773 4217
rect 6811 4183 6825 4217
rect 6825 4183 6845 4217
rect 6883 4183 6893 4217
rect 6893 4183 6917 4217
rect 6955 4183 6961 4217
rect 6961 4183 6989 4217
rect 7027 4183 7029 4217
rect 7029 4183 7061 4217
rect 7099 4183 7131 4217
rect 7131 4183 7133 4217
rect 7171 4183 7199 4217
rect 7199 4183 7205 4217
rect 7243 4183 7267 4217
rect 7267 4183 7277 4217
rect 7315 4183 7335 4217
rect 7335 4183 7349 4217
rect 7387 4183 7403 4217
rect 7403 4183 7421 4217
rect 7459 4183 7471 4217
rect 7471 4183 7493 4217
rect 7531 4183 7539 4217
rect 7539 4183 7565 4217
rect 7603 4183 7607 4217
rect 7607 4183 7637 4217
rect 7675 4183 7709 4217
rect 7747 4183 7777 4217
rect 7777 4183 7781 4217
rect 7819 4183 7845 4217
rect 7845 4183 7853 4217
rect 343 3395 377 3409
rect 343 3375 377 3395
rect 343 3327 377 3337
rect 343 3303 377 3327
rect 343 3259 377 3265
rect 343 3231 377 3259
rect 343 3191 377 3193
rect 343 3159 377 3191
rect 343 3089 377 3121
rect 343 3087 377 3089
rect 343 3021 377 3049
rect 343 3015 377 3021
rect 343 2953 377 2977
rect 343 2943 377 2953
rect 343 2885 377 2905
rect 343 2871 377 2885
rect 2263 3395 2297 3409
rect 2263 3375 2297 3395
rect 2263 3327 2297 3337
rect 2263 3303 2297 3327
rect 2263 3259 2297 3265
rect 2263 3231 2297 3259
rect 2263 3191 2297 3193
rect 2263 3159 2297 3191
rect 2263 3089 2297 3121
rect 2263 3087 2297 3089
rect 2263 3021 2297 3049
rect 2263 3015 2297 3021
rect 2263 2953 2297 2977
rect 2263 2943 2297 2953
rect 2263 2885 2297 2905
rect 2263 2871 2297 2885
rect 4183 3395 4217 3409
rect 4183 3375 4217 3395
rect 4183 3327 4217 3337
rect 4183 3303 4217 3327
rect 4183 3259 4217 3265
rect 4183 3231 4217 3259
rect 4183 3191 4217 3193
rect 4183 3159 4217 3191
rect 4183 3089 4217 3121
rect 4183 3087 4217 3089
rect 4183 3021 4217 3049
rect 4183 3015 4217 3021
rect 4183 2953 4217 2977
rect 4183 2943 4217 2953
rect 4183 2885 4217 2905
rect 4183 2871 4217 2885
rect 6103 3395 6137 3409
rect 6103 3375 6137 3395
rect 6103 3327 6137 3337
rect 6103 3303 6137 3327
rect 6103 3259 6137 3265
rect 6103 3231 6137 3259
rect 6103 3191 6137 3193
rect 6103 3159 6137 3191
rect 6103 3089 6137 3121
rect 6103 3087 6137 3089
rect 6103 3021 6137 3049
rect 6103 3015 6137 3021
rect 6103 2953 6137 2977
rect 6103 2943 6137 2953
rect 6103 2885 6137 2905
rect 6103 2871 6137 2885
rect 8023 3395 8057 3409
rect 8023 3375 8057 3395
rect 8023 3327 8057 3337
rect 8023 3303 8057 3327
rect 8023 3259 8057 3265
rect 8023 3231 8057 3259
rect 8023 3191 8057 3193
rect 8023 3159 8057 3191
rect 8023 3089 8057 3121
rect 8023 3087 8057 3089
rect 8023 3021 8057 3049
rect 8023 3015 8057 3021
rect 8023 2953 8057 2977
rect 8023 2943 8057 2953
rect 8023 2885 8057 2905
rect 8023 2871 8057 2885
rect 343 2635 377 2649
rect 343 2615 377 2635
rect 343 2567 377 2577
rect 343 2543 377 2567
rect 343 2499 377 2505
rect 343 2471 377 2499
rect 343 2431 377 2433
rect 343 2399 377 2431
rect 343 2329 377 2361
rect 343 2327 377 2329
rect 343 2261 377 2289
rect 343 2255 377 2261
rect 343 2193 377 2217
rect 343 2183 377 2193
rect 343 2125 377 2145
rect 343 2111 377 2125
rect 2263 2635 2297 2649
rect 2263 2615 2297 2635
rect 2263 2567 2297 2577
rect 2263 2543 2297 2567
rect 2263 2499 2297 2505
rect 2263 2471 2297 2499
rect 2263 2431 2297 2433
rect 2263 2399 2297 2431
rect 2263 2329 2297 2361
rect 2263 2327 2297 2329
rect 2263 2261 2297 2289
rect 2263 2255 2297 2261
rect 2263 2193 2297 2217
rect 2263 2183 2297 2193
rect 2263 2125 2297 2145
rect 2263 2111 2297 2125
rect 4183 2635 4217 2649
rect 4183 2615 4217 2635
rect 4183 2567 4217 2577
rect 4183 2543 4217 2567
rect 4183 2499 4217 2505
rect 4183 2471 4217 2499
rect 4183 2431 4217 2433
rect 4183 2399 4217 2431
rect 4183 2329 4217 2361
rect 4183 2327 4217 2329
rect 4183 2261 4217 2289
rect 4183 2255 4217 2261
rect 4183 2193 4217 2217
rect 4183 2183 4217 2193
rect 4183 2125 4217 2145
rect 4183 2111 4217 2125
rect 6103 2635 6137 2649
rect 6103 2615 6137 2635
rect 6103 2567 6137 2577
rect 6103 2543 6137 2567
rect 6103 2499 6137 2505
rect 6103 2471 6137 2499
rect 6103 2431 6137 2433
rect 6103 2399 6137 2431
rect 6103 2329 6137 2361
rect 6103 2327 6137 2329
rect 6103 2261 6137 2289
rect 6103 2255 6137 2261
rect 6103 2193 6137 2217
rect 6103 2183 6137 2193
rect 6103 2125 6137 2145
rect 6103 2111 6137 2125
rect 8023 2635 8057 2649
rect 8023 2615 8057 2635
rect 8023 2567 8057 2577
rect 8023 2543 8057 2567
rect 8023 2499 8057 2505
rect 8023 2471 8057 2499
rect 8023 2431 8057 2433
rect 8023 2399 8057 2431
rect 8023 2329 8057 2361
rect 8023 2327 8057 2329
rect 8023 2261 8057 2289
rect 8023 2255 8057 2261
rect 8023 2193 8057 2217
rect 8023 2183 8057 2193
rect 8023 2125 8057 2145
rect 8023 2111 8057 2125
rect 547 1943 555 1977
rect 555 1943 581 1977
rect 619 1943 623 1977
rect 623 1943 653 1977
rect 691 1943 725 1977
rect 763 1943 793 1977
rect 793 1943 797 1977
rect 835 1943 861 1977
rect 861 1943 869 1977
rect 907 1943 929 1977
rect 929 1943 941 1977
rect 979 1943 997 1977
rect 997 1943 1013 1977
rect 1051 1943 1065 1977
rect 1065 1943 1085 1977
rect 1123 1943 1133 1977
rect 1133 1943 1157 1977
rect 1195 1943 1201 1977
rect 1201 1943 1229 1977
rect 1267 1943 1269 1977
rect 1269 1943 1301 1977
rect 1339 1943 1371 1977
rect 1371 1943 1373 1977
rect 1411 1943 1439 1977
rect 1439 1943 1445 1977
rect 1483 1943 1507 1977
rect 1507 1943 1517 1977
rect 1555 1943 1575 1977
rect 1575 1943 1589 1977
rect 1627 1943 1643 1977
rect 1643 1943 1661 1977
rect 1699 1943 1711 1977
rect 1711 1943 1733 1977
rect 1771 1943 1779 1977
rect 1779 1943 1805 1977
rect 1843 1943 1847 1977
rect 1847 1943 1877 1977
rect 1915 1943 1949 1977
rect 1987 1943 2017 1977
rect 2017 1943 2021 1977
rect 2059 1943 2085 1977
rect 2085 1943 2093 1977
rect 2467 1943 2475 1977
rect 2475 1943 2501 1977
rect 2539 1943 2543 1977
rect 2543 1943 2573 1977
rect 2611 1943 2645 1977
rect 2683 1943 2713 1977
rect 2713 1943 2717 1977
rect 2755 1943 2781 1977
rect 2781 1943 2789 1977
rect 2827 1943 2849 1977
rect 2849 1943 2861 1977
rect 2899 1943 2917 1977
rect 2917 1943 2933 1977
rect 2971 1943 2985 1977
rect 2985 1943 3005 1977
rect 3043 1943 3053 1977
rect 3053 1943 3077 1977
rect 3115 1943 3121 1977
rect 3121 1943 3149 1977
rect 3187 1943 3189 1977
rect 3189 1943 3221 1977
rect 3259 1943 3291 1977
rect 3291 1943 3293 1977
rect 3331 1943 3359 1977
rect 3359 1943 3365 1977
rect 3403 1943 3427 1977
rect 3427 1943 3437 1977
rect 3475 1943 3495 1977
rect 3495 1943 3509 1977
rect 3547 1943 3563 1977
rect 3563 1943 3581 1977
rect 3619 1943 3631 1977
rect 3631 1943 3653 1977
rect 3691 1943 3699 1977
rect 3699 1943 3725 1977
rect 3763 1943 3767 1977
rect 3767 1943 3797 1977
rect 3835 1943 3869 1977
rect 3907 1943 3937 1977
rect 3937 1943 3941 1977
rect 3979 1943 4005 1977
rect 4005 1943 4013 1977
rect 4387 1943 4395 1977
rect 4395 1943 4421 1977
rect 4459 1943 4463 1977
rect 4463 1943 4493 1977
rect 4531 1943 4565 1977
rect 4603 1943 4633 1977
rect 4633 1943 4637 1977
rect 4675 1943 4701 1977
rect 4701 1943 4709 1977
rect 4747 1943 4769 1977
rect 4769 1943 4781 1977
rect 4819 1943 4837 1977
rect 4837 1943 4853 1977
rect 4891 1943 4905 1977
rect 4905 1943 4925 1977
rect 4963 1943 4973 1977
rect 4973 1943 4997 1977
rect 5035 1943 5041 1977
rect 5041 1943 5069 1977
rect 5107 1943 5109 1977
rect 5109 1943 5141 1977
rect 5179 1943 5211 1977
rect 5211 1943 5213 1977
rect 5251 1943 5279 1977
rect 5279 1943 5285 1977
rect 5323 1943 5347 1977
rect 5347 1943 5357 1977
rect 5395 1943 5415 1977
rect 5415 1943 5429 1977
rect 5467 1943 5483 1977
rect 5483 1943 5501 1977
rect 5539 1943 5551 1977
rect 5551 1943 5573 1977
rect 5611 1943 5619 1977
rect 5619 1943 5645 1977
rect 5683 1943 5687 1977
rect 5687 1943 5717 1977
rect 5755 1943 5789 1977
rect 5827 1943 5857 1977
rect 5857 1943 5861 1977
rect 5899 1943 5925 1977
rect 5925 1943 5933 1977
rect 6307 1943 6315 1977
rect 6315 1943 6341 1977
rect 6379 1943 6383 1977
rect 6383 1943 6413 1977
rect 6451 1943 6485 1977
rect 6523 1943 6553 1977
rect 6553 1943 6557 1977
rect 6595 1943 6621 1977
rect 6621 1943 6629 1977
rect 6667 1943 6689 1977
rect 6689 1943 6701 1977
rect 6739 1943 6757 1977
rect 6757 1943 6773 1977
rect 6811 1943 6825 1977
rect 6825 1943 6845 1977
rect 6883 1943 6893 1977
rect 6893 1943 6917 1977
rect 6955 1943 6961 1977
rect 6961 1943 6989 1977
rect 7027 1943 7029 1977
rect 7029 1943 7061 1977
rect 7099 1943 7131 1977
rect 7131 1943 7133 1977
rect 7171 1943 7199 1977
rect 7199 1943 7205 1977
rect 7243 1943 7267 1977
rect 7267 1943 7277 1977
rect 7315 1943 7335 1977
rect 7335 1943 7349 1977
rect 7387 1943 7403 1977
rect 7403 1943 7421 1977
rect 7459 1943 7471 1977
rect 7471 1943 7493 1977
rect 7531 1943 7539 1977
rect 7539 1943 7565 1977
rect 7603 1943 7607 1977
rect 7607 1943 7637 1977
rect 7675 1943 7709 1977
rect 7747 1943 7777 1977
rect 7777 1943 7781 1977
rect 7819 1943 7845 1977
rect 7845 1943 7853 1977
rect 183 1303 217 1337
rect 503 1303 537 1337
rect 663 1303 697 1337
rect 823 1303 857 1337
rect 983 1303 1017 1337
rect 1143 1303 1177 1337
rect 1463 1303 1497 1337
rect 1623 1303 1657 1337
rect 1783 1303 1817 1337
rect 1943 1303 1977 1337
rect 2103 1303 2137 1337
rect 2263 1303 2297 1337
rect 2423 1303 2457 1337
rect 2583 1303 2617 1337
rect 2743 1303 2777 1337
rect 2903 1303 2937 1337
rect 3063 1303 3097 1337
rect 3383 1303 3417 1337
rect 3543 1303 3577 1337
rect 3703 1303 3737 1337
rect 3863 1303 3897 1337
rect 4023 1303 4057 1337
rect 4343 1303 4377 1337
rect 4503 1303 4537 1337
rect 4663 1303 4697 1337
rect 4823 1303 4857 1337
rect 4983 1303 5017 1337
rect 5303 1303 5337 1337
rect 5463 1303 5497 1337
rect 5623 1303 5657 1337
rect 5783 1303 5817 1337
rect 5943 1303 5977 1337
rect 6103 1303 6137 1337
rect 6263 1303 6297 1337
rect 6423 1303 6457 1337
rect 6583 1303 6617 1337
rect 6743 1303 6777 1337
rect 6903 1303 6937 1337
rect 7223 1303 7257 1337
rect 7383 1303 7417 1337
rect 7543 1303 7577 1337
rect 7703 1303 7737 1337
rect 7863 1303 7897 1337
rect 8183 1303 8217 1337
rect 547 823 555 857
rect 555 823 581 857
rect 619 823 623 857
rect 623 823 653 857
rect 691 823 725 857
rect 763 823 793 857
rect 793 823 797 857
rect 835 823 861 857
rect 861 823 869 857
rect 907 823 929 857
rect 929 823 941 857
rect 979 823 997 857
rect 997 823 1013 857
rect 1051 823 1065 857
rect 1065 823 1085 857
rect 1123 823 1133 857
rect 1133 823 1157 857
rect 1195 823 1201 857
rect 1201 823 1229 857
rect 1267 823 1269 857
rect 1269 823 1301 857
rect 1339 823 1371 857
rect 1371 823 1373 857
rect 1411 823 1439 857
rect 1439 823 1445 857
rect 1483 823 1507 857
rect 1507 823 1517 857
rect 1555 823 1575 857
rect 1575 823 1589 857
rect 1627 823 1643 857
rect 1643 823 1661 857
rect 1699 823 1711 857
rect 1711 823 1733 857
rect 1771 823 1779 857
rect 1779 823 1805 857
rect 1843 823 1847 857
rect 1847 823 1877 857
rect 1915 823 1949 857
rect 1987 823 2017 857
rect 2017 823 2021 857
rect 2059 823 2085 857
rect 2085 823 2093 857
rect 2467 823 2475 857
rect 2475 823 2501 857
rect 2539 823 2543 857
rect 2543 823 2573 857
rect 2611 823 2645 857
rect 2683 823 2713 857
rect 2713 823 2717 857
rect 2755 823 2781 857
rect 2781 823 2789 857
rect 2827 823 2849 857
rect 2849 823 2861 857
rect 2899 823 2917 857
rect 2917 823 2933 857
rect 2971 823 2985 857
rect 2985 823 3005 857
rect 3043 823 3053 857
rect 3053 823 3077 857
rect 3115 823 3121 857
rect 3121 823 3149 857
rect 3187 823 3189 857
rect 3189 823 3221 857
rect 3259 823 3291 857
rect 3291 823 3293 857
rect 3331 823 3359 857
rect 3359 823 3365 857
rect 3403 823 3427 857
rect 3427 823 3437 857
rect 3475 823 3495 857
rect 3495 823 3509 857
rect 3547 823 3563 857
rect 3563 823 3581 857
rect 3619 823 3631 857
rect 3631 823 3653 857
rect 3691 823 3699 857
rect 3699 823 3725 857
rect 3763 823 3767 857
rect 3767 823 3797 857
rect 3835 823 3869 857
rect 3907 823 3937 857
rect 3937 823 3941 857
rect 3979 823 4005 857
rect 4005 823 4013 857
rect 4387 823 4395 857
rect 4395 823 4421 857
rect 4459 823 4463 857
rect 4463 823 4493 857
rect 4531 823 4565 857
rect 4603 823 4633 857
rect 4633 823 4637 857
rect 4675 823 4701 857
rect 4701 823 4709 857
rect 4747 823 4769 857
rect 4769 823 4781 857
rect 4819 823 4837 857
rect 4837 823 4853 857
rect 4891 823 4905 857
rect 4905 823 4925 857
rect 4963 823 4973 857
rect 4973 823 4997 857
rect 5035 823 5041 857
rect 5041 823 5069 857
rect 5107 823 5109 857
rect 5109 823 5141 857
rect 5179 823 5211 857
rect 5211 823 5213 857
rect 5251 823 5279 857
rect 5279 823 5285 857
rect 5323 823 5347 857
rect 5347 823 5357 857
rect 5395 823 5415 857
rect 5415 823 5429 857
rect 5467 823 5483 857
rect 5483 823 5501 857
rect 5539 823 5551 857
rect 5551 823 5573 857
rect 5611 823 5619 857
rect 5619 823 5645 857
rect 5683 823 5687 857
rect 5687 823 5717 857
rect 5755 823 5789 857
rect 5827 823 5857 857
rect 5857 823 5861 857
rect 5899 823 5925 857
rect 5925 823 5933 857
rect 6307 823 6315 857
rect 6315 823 6341 857
rect 6379 823 6383 857
rect 6383 823 6413 857
rect 6451 823 6485 857
rect 6523 823 6553 857
rect 6553 823 6557 857
rect 6595 823 6621 857
rect 6621 823 6629 857
rect 6667 823 6689 857
rect 6689 823 6701 857
rect 6739 823 6757 857
rect 6757 823 6773 857
rect 6811 823 6825 857
rect 6825 823 6845 857
rect 6883 823 6893 857
rect 6893 823 6917 857
rect 6955 823 6961 857
rect 6961 823 6989 857
rect 7027 823 7029 857
rect 7029 823 7061 857
rect 7099 823 7131 857
rect 7131 823 7133 857
rect 7171 823 7199 857
rect 7199 823 7205 857
rect 7243 823 7267 857
rect 7267 823 7277 857
rect 7315 823 7335 857
rect 7335 823 7349 857
rect 7387 823 7403 857
rect 7403 823 7421 857
rect 7459 823 7471 857
rect 7471 823 7493 857
rect 7531 823 7539 857
rect 7539 823 7565 857
rect 7603 823 7607 857
rect 7607 823 7637 857
rect 7675 823 7709 857
rect 7747 823 7777 857
rect 7777 823 7781 857
rect 7819 823 7845 857
rect 7845 823 7853 857
rect 343 711 377 713
rect 343 679 377 711
rect 343 609 377 641
rect 343 607 377 609
rect 2263 711 2297 713
rect 2263 679 2297 711
rect 2263 609 2297 641
rect 2263 607 2297 609
rect 4183 711 4217 713
rect 4183 679 4217 711
rect 4183 609 4217 641
rect 4183 607 4217 609
rect 6103 711 6137 713
rect 6103 679 6137 711
rect 6103 609 6137 641
rect 6103 607 6137 609
rect 8023 711 8057 713
rect 8023 679 8057 711
rect 8023 609 8057 641
rect 8023 607 8057 609
rect 343 311 377 313
rect 343 279 377 311
rect 343 209 377 241
rect 343 207 377 209
rect 2263 311 2297 313
rect 2263 279 2297 311
rect 2263 209 2297 241
rect 2263 207 2297 209
rect 4183 311 4217 313
rect 4183 279 4217 311
rect 4183 209 4217 241
rect 4183 207 4217 209
rect 6103 311 6137 313
rect 6103 279 6137 311
rect 6103 209 6137 241
rect 6103 207 6137 209
rect 8023 311 8057 313
rect 8023 279 8057 311
rect 8023 209 8057 241
rect 8023 207 8057 209
<< metal1 >>
rect 320 5649 400 5680
rect 320 5615 343 5649
rect 377 5615 400 5649
rect 320 5577 400 5615
rect 320 5543 343 5577
rect 377 5543 400 5577
rect 320 5505 400 5543
rect 320 5471 343 5505
rect 377 5471 400 5505
rect 320 5433 400 5471
rect 320 5399 343 5433
rect 377 5399 400 5433
rect 320 5361 400 5399
rect 320 5327 343 5361
rect 377 5327 400 5361
rect 320 5289 400 5327
rect 320 5255 343 5289
rect 377 5255 400 5289
rect 320 5217 400 5255
rect 320 5183 343 5217
rect 377 5183 400 5217
rect 320 5145 400 5183
rect 320 5111 343 5145
rect 377 5111 400 5145
rect 320 4889 400 5111
rect 2240 5649 2320 5680
rect 2240 5615 2263 5649
rect 2297 5615 2320 5649
rect 2240 5577 2320 5615
rect 2240 5543 2263 5577
rect 2297 5543 2320 5577
rect 2240 5505 2320 5543
rect 2240 5471 2263 5505
rect 2297 5471 2320 5505
rect 2240 5433 2320 5471
rect 2240 5399 2263 5433
rect 2297 5399 2320 5433
rect 2240 5361 2320 5399
rect 2240 5327 2263 5361
rect 2297 5327 2320 5361
rect 2240 5289 2320 5327
rect 2240 5255 2263 5289
rect 2297 5255 2320 5289
rect 2240 5217 2320 5255
rect 2240 5183 2263 5217
rect 2297 5183 2320 5217
rect 2240 5145 2320 5183
rect 2240 5111 2263 5145
rect 2297 5111 2320 5145
rect 2240 5080 2320 5111
rect 4160 5649 4240 5680
rect 4160 5634 4183 5649
rect 4217 5634 4240 5649
rect 4160 5582 4174 5634
rect 4226 5582 4240 5634
rect 4160 5577 4240 5582
rect 4160 5570 4183 5577
rect 4217 5570 4240 5577
rect 4160 5518 4174 5570
rect 4226 5518 4240 5570
rect 4160 5506 4240 5518
rect 4160 5454 4174 5506
rect 4226 5454 4240 5506
rect 4160 5442 4240 5454
rect 4160 5390 4174 5442
rect 4226 5390 4240 5442
rect 4160 5378 4240 5390
rect 4160 5326 4174 5378
rect 4226 5326 4240 5378
rect 4160 5289 4240 5326
rect 4160 5255 4183 5289
rect 4217 5255 4240 5289
rect 4160 5217 4240 5255
rect 4160 5183 4183 5217
rect 4217 5183 4240 5217
rect 4160 5145 4240 5183
rect 4160 5111 4183 5145
rect 4217 5111 4240 5145
rect 4160 5080 4240 5111
rect 6080 5649 6160 5680
rect 6080 5615 6103 5649
rect 6137 5615 6160 5649
rect 6080 5577 6160 5615
rect 6080 5543 6103 5577
rect 6137 5543 6160 5577
rect 6080 5505 6160 5543
rect 6080 5471 6103 5505
rect 6137 5471 6160 5505
rect 6080 5433 6160 5471
rect 6080 5399 6103 5433
rect 6137 5399 6160 5433
rect 6080 5361 6160 5399
rect 6080 5327 6103 5361
rect 6137 5327 6160 5361
rect 6080 5289 6160 5327
rect 6080 5255 6103 5289
rect 6137 5255 6160 5289
rect 6080 5217 6160 5255
rect 6080 5183 6103 5217
rect 6137 5183 6160 5217
rect 6080 5145 6160 5183
rect 6080 5111 6103 5145
rect 6137 5111 6160 5145
rect 6080 5080 6160 5111
rect 8000 5649 8080 5680
rect 8000 5615 8023 5649
rect 8057 5615 8080 5649
rect 8000 5577 8080 5615
rect 8000 5543 8023 5577
rect 8057 5543 8080 5577
rect 8000 5505 8080 5543
rect 8000 5471 8023 5505
rect 8057 5471 8080 5505
rect 8000 5433 8080 5471
rect 8000 5399 8023 5433
rect 8057 5399 8080 5433
rect 8000 5361 8080 5399
rect 8000 5327 8023 5361
rect 8057 5327 8080 5361
rect 8000 5289 8080 5327
rect 8000 5255 8023 5289
rect 8057 5255 8080 5289
rect 8000 5217 8080 5255
rect 8000 5183 8023 5217
rect 8057 5183 8080 5217
rect 8000 5145 8080 5183
rect 8000 5111 8023 5145
rect 8057 5111 8080 5145
rect 320 4855 343 4889
rect 377 4855 400 4889
rect 320 4817 400 4855
rect 320 4783 343 4817
rect 377 4783 400 4817
rect 320 4745 400 4783
rect 320 4711 343 4745
rect 377 4711 400 4745
rect 320 4673 400 4711
rect 320 4639 343 4673
rect 377 4639 400 4673
rect 320 4601 400 4639
rect 320 4567 343 4601
rect 377 4567 400 4601
rect 320 4529 400 4567
rect 320 4495 343 4529
rect 377 4495 400 4529
rect 320 4457 400 4495
rect 320 4423 343 4457
rect 377 4423 400 4457
rect 320 4385 400 4423
rect 320 4351 343 4385
rect 377 4351 400 4385
rect 0 3986 80 4000
rect 0 3934 14 3986
rect 66 3934 80 3986
rect 0 3666 80 3934
rect 0 3614 14 3666
rect 66 3614 80 3666
rect 0 3600 80 3614
rect 160 3986 240 4000
rect 160 3934 174 3986
rect 226 3934 240 3986
rect 160 3666 240 3934
rect 160 3614 174 3666
rect 226 3614 240 3666
rect 160 3600 240 3614
rect 320 3986 400 4351
rect 2240 4889 2320 4920
rect 2240 4855 2263 4889
rect 2297 4855 2320 4889
rect 2240 4817 2320 4855
rect 2240 4783 2263 4817
rect 2297 4783 2320 4817
rect 2240 4745 2320 4783
rect 2240 4711 2263 4745
rect 2297 4711 2320 4745
rect 2240 4673 2320 4711
rect 2240 4639 2263 4673
rect 2297 4639 2320 4673
rect 2240 4601 2320 4639
rect 2240 4567 2263 4601
rect 2297 4567 2320 4601
rect 2240 4529 2320 4567
rect 2240 4495 2263 4529
rect 2297 4495 2320 4529
rect 2240 4457 2320 4495
rect 2240 4423 2263 4457
rect 2297 4423 2320 4457
rect 2240 4385 2320 4423
rect 2240 4351 2263 4385
rect 2297 4351 2320 4385
rect 2240 4320 2320 4351
rect 4160 4889 4240 4920
rect 4160 4855 4183 4889
rect 4217 4855 4240 4889
rect 4160 4817 4240 4855
rect 4160 4783 4183 4817
rect 4217 4783 4240 4817
rect 4160 4745 4240 4783
rect 4160 4711 4183 4745
rect 4217 4711 4240 4745
rect 4160 4673 4240 4711
rect 4160 4639 4183 4673
rect 4217 4639 4240 4673
rect 4160 4601 4240 4639
rect 4160 4567 4183 4601
rect 4217 4567 4240 4601
rect 4160 4529 4240 4567
rect 4160 4495 4183 4529
rect 4217 4495 4240 4529
rect 4160 4457 4240 4495
rect 4160 4423 4183 4457
rect 4217 4423 4240 4457
rect 4160 4385 4240 4423
rect 4160 4351 4183 4385
rect 4217 4351 4240 4385
rect 520 4217 2120 4240
rect 520 4183 547 4217
rect 581 4183 619 4217
rect 653 4183 691 4217
rect 725 4183 763 4217
rect 797 4183 835 4217
rect 869 4183 907 4217
rect 941 4183 979 4217
rect 1013 4183 1051 4217
rect 1085 4183 1123 4217
rect 1157 4183 1195 4217
rect 1229 4183 1267 4217
rect 1301 4183 1339 4217
rect 1373 4183 1411 4217
rect 1445 4183 1483 4217
rect 1517 4183 1555 4217
rect 1589 4183 1627 4217
rect 1661 4183 1699 4217
rect 1733 4183 1771 4217
rect 1805 4183 1843 4217
rect 1877 4183 1915 4217
rect 1949 4183 1987 4217
rect 2021 4183 2059 4217
rect 2093 4183 2120 4217
rect 520 4160 2120 4183
rect 2440 4217 4040 4240
rect 2440 4183 2467 4217
rect 2501 4183 2539 4217
rect 2573 4183 2611 4217
rect 2645 4183 2683 4217
rect 2717 4183 2755 4217
rect 2789 4183 2827 4217
rect 2861 4183 2899 4217
rect 2933 4183 2971 4217
rect 3005 4183 3043 4217
rect 3077 4183 3115 4217
rect 3149 4183 3187 4217
rect 3221 4183 3259 4217
rect 3293 4183 3331 4217
rect 3365 4183 3403 4217
rect 3437 4183 3475 4217
rect 3509 4183 3547 4217
rect 3581 4183 3619 4217
rect 3653 4183 3691 4217
rect 3725 4183 3763 4217
rect 3797 4183 3835 4217
rect 3869 4183 3907 4217
rect 3941 4183 3979 4217
rect 4013 4183 4040 4217
rect 2440 4160 4040 4183
rect 320 3934 334 3986
rect 386 3934 400 3986
rect 320 3666 400 3934
rect 320 3614 334 3666
rect 386 3614 400 3666
rect 320 3409 400 3614
rect 480 3986 560 4000
rect 480 3934 494 3986
rect 546 3934 560 3986
rect 480 3666 560 3934
rect 480 3614 494 3666
rect 546 3614 560 3666
rect 480 3600 560 3614
rect 640 3986 720 4000
rect 640 3934 654 3986
rect 706 3934 720 3986
rect 640 3666 720 3934
rect 640 3614 654 3666
rect 706 3614 720 3666
rect 640 3600 720 3614
rect 800 3986 880 4000
rect 800 3934 814 3986
rect 866 3934 880 3986
rect 800 3666 880 3934
rect 800 3614 814 3666
rect 866 3614 880 3666
rect 800 3600 880 3614
rect 960 3986 1040 4000
rect 960 3934 974 3986
rect 1026 3934 1040 3986
rect 960 3666 1040 3934
rect 960 3614 974 3666
rect 1026 3614 1040 3666
rect 960 3600 1040 3614
rect 1120 3986 1200 4000
rect 1120 3934 1134 3986
rect 1186 3934 1200 3986
rect 1120 3666 1200 3934
rect 1280 3826 1360 4160
rect 1280 3774 1294 3826
rect 1346 3774 1360 3826
rect 1280 3760 1360 3774
rect 1440 3986 1520 4000
rect 1440 3934 1454 3986
rect 1506 3934 1520 3986
rect 1120 3614 1134 3666
rect 1186 3614 1200 3666
rect 1120 3600 1200 3614
rect 1440 3666 1520 3934
rect 1440 3614 1454 3666
rect 1506 3614 1520 3666
rect 1440 3600 1520 3614
rect 1600 3986 1680 4000
rect 1600 3934 1614 3986
rect 1666 3934 1680 3986
rect 1600 3666 1680 3934
rect 1600 3614 1614 3666
rect 1666 3614 1680 3666
rect 1600 3600 1680 3614
rect 1760 3986 1840 4000
rect 1760 3934 1774 3986
rect 1826 3934 1840 3986
rect 1760 3666 1840 3934
rect 1760 3614 1774 3666
rect 1826 3614 1840 3666
rect 1760 3600 1840 3614
rect 1920 3986 2000 4000
rect 1920 3934 1934 3986
rect 1986 3934 2000 3986
rect 1920 3666 2000 3934
rect 1920 3614 1934 3666
rect 1986 3614 2000 3666
rect 1920 3600 2000 3614
rect 2080 3986 2160 4000
rect 2080 3934 2094 3986
rect 2146 3934 2160 3986
rect 2080 3666 2160 3934
rect 2080 3614 2094 3666
rect 2146 3614 2160 3666
rect 2080 3600 2160 3614
rect 2240 3986 2320 4000
rect 2240 3934 2254 3986
rect 2306 3934 2320 3986
rect 2240 3666 2320 3934
rect 2240 3614 2254 3666
rect 2306 3614 2320 3666
rect 2240 3600 2320 3614
rect 2400 3986 2480 4000
rect 2400 3934 2414 3986
rect 2466 3934 2480 3986
rect 2400 3666 2480 3934
rect 2400 3614 2414 3666
rect 2466 3614 2480 3666
rect 2400 3600 2480 3614
rect 2560 3986 2640 4000
rect 2560 3934 2574 3986
rect 2626 3934 2640 3986
rect 2560 3666 2640 3934
rect 2560 3614 2574 3666
rect 2626 3614 2640 3666
rect 2560 3600 2640 3614
rect 2720 3986 2800 4000
rect 2720 3934 2734 3986
rect 2786 3934 2800 3986
rect 2720 3666 2800 3934
rect 2720 3614 2734 3666
rect 2786 3614 2800 3666
rect 2720 3600 2800 3614
rect 2880 3986 2960 4000
rect 2880 3934 2894 3986
rect 2946 3934 2960 3986
rect 2880 3666 2960 3934
rect 2880 3614 2894 3666
rect 2946 3614 2960 3666
rect 2880 3600 2960 3614
rect 3040 3986 3120 4000
rect 3040 3934 3054 3986
rect 3106 3934 3120 3986
rect 3040 3666 3120 3934
rect 3200 3826 3280 4160
rect 3200 3774 3214 3826
rect 3266 3774 3280 3826
rect 3200 3760 3280 3774
rect 3360 3986 3440 4000
rect 3360 3934 3374 3986
rect 3426 3934 3440 3986
rect 3040 3614 3054 3666
rect 3106 3614 3120 3666
rect 3040 3600 3120 3614
rect 3360 3666 3440 3934
rect 3360 3614 3374 3666
rect 3426 3614 3440 3666
rect 3360 3600 3440 3614
rect 3520 3986 3600 4000
rect 3520 3934 3534 3986
rect 3586 3934 3600 3986
rect 3520 3666 3600 3934
rect 3520 3614 3534 3666
rect 3586 3614 3600 3666
rect 3520 3600 3600 3614
rect 3680 3986 3760 4000
rect 3680 3934 3694 3986
rect 3746 3934 3760 3986
rect 3680 3666 3760 3934
rect 3680 3614 3694 3666
rect 3746 3614 3760 3666
rect 3680 3600 3760 3614
rect 3840 3986 3920 4000
rect 3840 3934 3854 3986
rect 3906 3934 3920 3986
rect 3840 3666 3920 3934
rect 3840 3614 3854 3666
rect 3906 3614 3920 3666
rect 3840 3600 3920 3614
rect 4000 3986 4080 4000
rect 4000 3934 4014 3986
rect 4066 3934 4080 3986
rect 4000 3666 4080 3934
rect 4000 3614 4014 3666
rect 4066 3614 4080 3666
rect 4000 3600 4080 3614
rect 4160 3986 4240 4351
rect 6080 4889 6160 4920
rect 6080 4855 6103 4889
rect 6137 4855 6160 4889
rect 6080 4817 6160 4855
rect 6080 4783 6103 4817
rect 6137 4783 6160 4817
rect 6080 4745 6160 4783
rect 6080 4711 6103 4745
rect 6137 4711 6160 4745
rect 6080 4673 6160 4711
rect 6080 4639 6103 4673
rect 6137 4639 6160 4673
rect 6080 4601 6160 4639
rect 6080 4567 6103 4601
rect 6137 4567 6160 4601
rect 6080 4529 6160 4567
rect 6080 4495 6103 4529
rect 6137 4495 6160 4529
rect 6080 4457 6160 4495
rect 6080 4423 6103 4457
rect 6137 4423 6160 4457
rect 6080 4385 6160 4423
rect 6080 4351 6103 4385
rect 6137 4351 6160 4385
rect 6080 4320 6160 4351
rect 8000 4889 8080 5111
rect 8000 4855 8023 4889
rect 8057 4855 8080 4889
rect 8000 4817 8080 4855
rect 8000 4783 8023 4817
rect 8057 4783 8080 4817
rect 8000 4745 8080 4783
rect 8000 4711 8023 4745
rect 8057 4711 8080 4745
rect 8000 4673 8080 4711
rect 8000 4639 8023 4673
rect 8057 4639 8080 4673
rect 8000 4601 8080 4639
rect 8000 4567 8023 4601
rect 8057 4567 8080 4601
rect 8000 4529 8080 4567
rect 8000 4495 8023 4529
rect 8057 4495 8080 4529
rect 8000 4457 8080 4495
rect 8000 4423 8023 4457
rect 8057 4423 8080 4457
rect 8000 4385 8080 4423
rect 8000 4351 8023 4385
rect 8057 4351 8080 4385
rect 4360 4217 5960 4240
rect 4360 4183 4387 4217
rect 4421 4183 4459 4217
rect 4493 4183 4531 4217
rect 4565 4183 4603 4217
rect 4637 4183 4675 4217
rect 4709 4183 4747 4217
rect 4781 4183 4819 4217
rect 4853 4183 4891 4217
rect 4925 4183 4963 4217
rect 4997 4183 5035 4217
rect 5069 4183 5107 4217
rect 5141 4183 5179 4217
rect 5213 4183 5251 4217
rect 5285 4183 5323 4217
rect 5357 4183 5395 4217
rect 5429 4183 5467 4217
rect 5501 4183 5539 4217
rect 5573 4183 5611 4217
rect 5645 4183 5683 4217
rect 5717 4183 5755 4217
rect 5789 4183 5827 4217
rect 5861 4183 5899 4217
rect 5933 4183 5960 4217
rect 4360 4160 5960 4183
rect 6280 4217 7880 4240
rect 6280 4183 6307 4217
rect 6341 4183 6379 4217
rect 6413 4183 6451 4217
rect 6485 4183 6523 4217
rect 6557 4183 6595 4217
rect 6629 4183 6667 4217
rect 6701 4183 6739 4217
rect 6773 4183 6811 4217
rect 6845 4183 6883 4217
rect 6917 4183 6955 4217
rect 6989 4183 7027 4217
rect 7061 4183 7099 4217
rect 7133 4183 7171 4217
rect 7205 4183 7243 4217
rect 7277 4183 7315 4217
rect 7349 4183 7387 4217
rect 7421 4183 7459 4217
rect 7493 4183 7531 4217
rect 7565 4183 7603 4217
rect 7637 4183 7675 4217
rect 7709 4183 7747 4217
rect 7781 4183 7819 4217
rect 7853 4183 7880 4217
rect 6280 4160 7880 4183
rect 4160 3934 4174 3986
rect 4226 3934 4240 3986
rect 4160 3666 4240 3934
rect 4160 3614 4174 3666
rect 4226 3614 4240 3666
rect 4160 3600 4240 3614
rect 4320 3986 4400 4000
rect 4320 3934 4334 3986
rect 4386 3934 4400 3986
rect 4320 3666 4400 3934
rect 4320 3614 4334 3666
rect 4386 3614 4400 3666
rect 4320 3600 4400 3614
rect 4480 3986 4560 4000
rect 4480 3934 4494 3986
rect 4546 3934 4560 3986
rect 4480 3666 4560 3934
rect 4480 3614 4494 3666
rect 4546 3614 4560 3666
rect 4480 3600 4560 3614
rect 4640 3986 4720 4000
rect 4640 3934 4654 3986
rect 4706 3934 4720 3986
rect 4640 3666 4720 3934
rect 4640 3614 4654 3666
rect 4706 3614 4720 3666
rect 4640 3600 4720 3614
rect 4800 3986 4880 4000
rect 4800 3934 4814 3986
rect 4866 3934 4880 3986
rect 4800 3666 4880 3934
rect 4800 3614 4814 3666
rect 4866 3614 4880 3666
rect 4800 3600 4880 3614
rect 4960 3986 5040 4000
rect 4960 3934 4974 3986
rect 5026 3934 5040 3986
rect 4960 3666 5040 3934
rect 5120 3826 5200 4160
rect 5120 3774 5134 3826
rect 5186 3774 5200 3826
rect 5120 3760 5200 3774
rect 5280 3986 5360 4000
rect 5280 3934 5294 3986
rect 5346 3934 5360 3986
rect 4960 3614 4974 3666
rect 5026 3614 5040 3666
rect 4960 3600 5040 3614
rect 5280 3666 5360 3934
rect 5280 3614 5294 3666
rect 5346 3614 5360 3666
rect 5280 3600 5360 3614
rect 5440 3986 5520 4000
rect 5440 3934 5454 3986
rect 5506 3934 5520 3986
rect 5440 3666 5520 3934
rect 5440 3614 5454 3666
rect 5506 3614 5520 3666
rect 5440 3600 5520 3614
rect 5600 3986 5680 4000
rect 5600 3934 5614 3986
rect 5666 3934 5680 3986
rect 5600 3666 5680 3934
rect 5600 3614 5614 3666
rect 5666 3614 5680 3666
rect 5600 3600 5680 3614
rect 5760 3986 5840 4000
rect 5760 3934 5774 3986
rect 5826 3934 5840 3986
rect 5760 3666 5840 3934
rect 5760 3614 5774 3666
rect 5826 3614 5840 3666
rect 5760 3600 5840 3614
rect 5920 3986 6000 4000
rect 5920 3934 5934 3986
rect 5986 3934 6000 3986
rect 5920 3666 6000 3934
rect 5920 3614 5934 3666
rect 5986 3614 6000 3666
rect 5920 3600 6000 3614
rect 6080 3986 6160 4000
rect 6080 3934 6094 3986
rect 6146 3934 6160 3986
rect 6080 3666 6160 3934
rect 6080 3614 6094 3666
rect 6146 3614 6160 3666
rect 6080 3600 6160 3614
rect 6240 3986 6320 4000
rect 6240 3934 6254 3986
rect 6306 3934 6320 3986
rect 6240 3666 6320 3934
rect 6240 3614 6254 3666
rect 6306 3614 6320 3666
rect 6240 3600 6320 3614
rect 6400 3986 6480 4000
rect 6400 3934 6414 3986
rect 6466 3934 6480 3986
rect 6400 3666 6480 3934
rect 6400 3614 6414 3666
rect 6466 3614 6480 3666
rect 6400 3600 6480 3614
rect 6560 3986 6640 4000
rect 6560 3934 6574 3986
rect 6626 3934 6640 3986
rect 6560 3666 6640 3934
rect 6560 3614 6574 3666
rect 6626 3614 6640 3666
rect 6560 3600 6640 3614
rect 6720 3986 6800 4000
rect 6720 3934 6734 3986
rect 6786 3934 6800 3986
rect 6720 3666 6800 3934
rect 6720 3614 6734 3666
rect 6786 3614 6800 3666
rect 6720 3600 6800 3614
rect 6880 3986 6960 4000
rect 6880 3934 6894 3986
rect 6946 3934 6960 3986
rect 6880 3666 6960 3934
rect 7040 3826 7120 4160
rect 7040 3774 7054 3826
rect 7106 3774 7120 3826
rect 7040 3760 7120 3774
rect 7200 3986 7280 4000
rect 7200 3934 7214 3986
rect 7266 3934 7280 3986
rect 6880 3614 6894 3666
rect 6946 3614 6960 3666
rect 6880 3600 6960 3614
rect 7200 3666 7280 3934
rect 7200 3614 7214 3666
rect 7266 3614 7280 3666
rect 7200 3600 7280 3614
rect 7360 3986 7440 4000
rect 7360 3934 7374 3986
rect 7426 3934 7440 3986
rect 7360 3666 7440 3934
rect 7360 3614 7374 3666
rect 7426 3614 7440 3666
rect 7360 3600 7440 3614
rect 7520 3986 7600 4000
rect 7520 3934 7534 3986
rect 7586 3934 7600 3986
rect 7520 3666 7600 3934
rect 7520 3614 7534 3666
rect 7586 3614 7600 3666
rect 7520 3600 7600 3614
rect 7680 3986 7760 4000
rect 7680 3934 7694 3986
rect 7746 3934 7760 3986
rect 7680 3666 7760 3934
rect 7680 3614 7694 3666
rect 7746 3614 7760 3666
rect 7680 3600 7760 3614
rect 7840 3986 7920 4000
rect 7840 3934 7854 3986
rect 7906 3934 7920 3986
rect 7840 3666 7920 3934
rect 7840 3614 7854 3666
rect 7906 3614 7920 3666
rect 7840 3600 7920 3614
rect 8000 3986 8080 4351
rect 8000 3934 8014 3986
rect 8066 3934 8080 3986
rect 8000 3666 8080 3934
rect 8000 3614 8014 3666
rect 8066 3614 8080 3666
rect 320 3375 343 3409
rect 377 3375 400 3409
rect 320 3337 400 3375
rect 320 3303 343 3337
rect 377 3303 400 3337
rect 320 3265 400 3303
rect 320 3231 343 3265
rect 377 3231 400 3265
rect 320 3193 400 3231
rect 320 3159 343 3193
rect 377 3159 400 3193
rect 320 3121 400 3159
rect 320 3087 343 3121
rect 377 3087 400 3121
rect 320 3049 400 3087
rect 320 3015 343 3049
rect 377 3015 400 3049
rect 320 2977 400 3015
rect 320 2943 343 2977
rect 377 2943 400 2977
rect 320 2905 400 2943
rect 320 2871 343 2905
rect 377 2871 400 2905
rect 320 2840 400 2871
rect 2240 3409 2320 3440
rect 2240 3375 2263 3409
rect 2297 3375 2320 3409
rect 2240 3337 2320 3375
rect 2240 3303 2263 3337
rect 2297 3303 2320 3337
rect 2240 3265 2320 3303
rect 2240 3231 2263 3265
rect 2297 3231 2320 3265
rect 2240 3193 2320 3231
rect 2240 3159 2263 3193
rect 2297 3159 2320 3193
rect 2240 3121 2320 3159
rect 2240 3087 2263 3121
rect 2297 3087 2320 3121
rect 2240 3049 2320 3087
rect 2240 3015 2263 3049
rect 2297 3015 2320 3049
rect 2240 2977 2320 3015
rect 2240 2943 2263 2977
rect 2297 2943 2320 2977
rect 2240 2905 2320 2943
rect 2240 2871 2263 2905
rect 2297 2871 2320 2905
rect 2240 2840 2320 2871
rect 4160 3409 4240 3440
rect 4160 3375 4183 3409
rect 4217 3375 4240 3409
rect 4160 3337 4240 3375
rect 4160 3303 4183 3337
rect 4217 3303 4240 3337
rect 4160 3265 4240 3303
rect 4160 3231 4183 3265
rect 4217 3231 4240 3265
rect 4160 3193 4240 3231
rect 4160 3159 4183 3193
rect 4217 3159 4240 3193
rect 4160 3121 4240 3159
rect 4160 3087 4183 3121
rect 4217 3087 4240 3121
rect 4160 3049 4240 3087
rect 4160 3015 4183 3049
rect 4217 3015 4240 3049
rect 4160 2977 4240 3015
rect 4160 2943 4183 2977
rect 4217 2943 4240 2977
rect 4160 2905 4240 2943
rect 4160 2871 4183 2905
rect 4217 2871 4240 2905
rect 4160 2800 4240 2871
rect 6080 3409 6160 3440
rect 6080 3375 6103 3409
rect 6137 3375 6160 3409
rect 6080 3337 6160 3375
rect 6080 3303 6103 3337
rect 6137 3303 6160 3337
rect 6080 3265 6160 3303
rect 6080 3231 6103 3265
rect 6137 3231 6160 3265
rect 6080 3193 6160 3231
rect 6080 3159 6103 3193
rect 6137 3159 6160 3193
rect 6080 3121 6160 3159
rect 6080 3087 6103 3121
rect 6137 3087 6160 3121
rect 6080 3049 6160 3087
rect 6080 3015 6103 3049
rect 6137 3015 6160 3049
rect 6080 2977 6160 3015
rect 6080 2943 6103 2977
rect 6137 2943 6160 2977
rect 6080 2905 6160 2943
rect 6080 2871 6103 2905
rect 6137 2871 6160 2905
rect 6080 2840 6160 2871
rect 8000 3409 8080 3614
rect 8160 3986 8240 4000
rect 8160 3934 8174 3986
rect 8226 3934 8240 3986
rect 8160 3666 8240 3934
rect 8160 3614 8174 3666
rect 8226 3614 8240 3666
rect 8160 3600 8240 3614
rect 8320 3986 8400 4000
rect 8320 3934 8334 3986
rect 8386 3934 8400 3986
rect 8320 3666 8400 3934
rect 8320 3614 8334 3666
rect 8386 3614 8400 3666
rect 8320 3600 8400 3614
rect 8000 3375 8023 3409
rect 8057 3375 8080 3409
rect 8000 3337 8080 3375
rect 8000 3303 8023 3337
rect 8057 3303 8080 3337
rect 8000 3265 8080 3303
rect 8000 3231 8023 3265
rect 8057 3231 8080 3265
rect 8000 3193 8080 3231
rect 8000 3159 8023 3193
rect 8057 3159 8080 3193
rect 8000 3121 8080 3159
rect 8000 3087 8023 3121
rect 8057 3087 8080 3121
rect 8000 3049 8080 3087
rect 8000 3015 8023 3049
rect 8057 3015 8080 3049
rect 8000 2977 8080 3015
rect 8000 2943 8023 2977
rect 8057 2943 8080 2977
rect 8000 2905 8080 2943
rect 8000 2871 8023 2905
rect 8057 2871 8080 2905
rect 8000 2840 8080 2871
rect 2240 2786 2320 2800
rect 2240 2734 2254 2786
rect 2306 2734 2320 2786
rect 320 2649 400 2680
rect 320 2615 343 2649
rect 377 2615 400 2649
rect 320 2577 400 2615
rect 320 2543 343 2577
rect 377 2543 400 2577
rect 320 2505 400 2543
rect 320 2471 343 2505
rect 377 2471 400 2505
rect 320 2433 400 2471
rect 320 2399 343 2433
rect 377 2399 400 2433
rect 320 2361 400 2399
rect 320 2327 343 2361
rect 377 2327 400 2361
rect 320 2289 400 2327
rect 320 2255 343 2289
rect 377 2255 400 2289
rect 320 2217 400 2255
rect 320 2183 343 2217
rect 377 2183 400 2217
rect 320 2145 400 2183
rect 320 2111 343 2145
rect 377 2111 400 2145
rect 160 1337 240 1360
rect 160 1303 183 1337
rect 217 1303 240 1337
rect 160 1280 240 1303
rect 320 1186 400 2111
rect 2240 2649 2320 2734
rect 6080 2786 6160 2800
rect 6080 2734 6094 2786
rect 6146 2734 6160 2786
rect 2240 2615 2263 2649
rect 2297 2615 2320 2649
rect 2240 2577 2320 2615
rect 2240 2543 2263 2577
rect 2297 2543 2320 2577
rect 2240 2505 2320 2543
rect 2240 2471 2263 2505
rect 2297 2471 2320 2505
rect 2240 2433 2320 2471
rect 2240 2399 2263 2433
rect 2297 2399 2320 2433
rect 2240 2361 2320 2399
rect 2240 2327 2263 2361
rect 2297 2327 2320 2361
rect 2240 2289 2320 2327
rect 2240 2255 2263 2289
rect 2297 2255 2320 2289
rect 2240 2217 2320 2255
rect 2240 2183 2263 2217
rect 2297 2183 2320 2217
rect 2240 2145 2320 2183
rect 2240 2111 2263 2145
rect 2297 2111 2320 2145
rect 2240 2080 2320 2111
rect 4160 2649 4240 2680
rect 4160 2615 4183 2649
rect 4217 2615 4240 2649
rect 4160 2577 4240 2615
rect 4160 2543 4183 2577
rect 4217 2543 4240 2577
rect 4160 2505 4240 2543
rect 4160 2471 4183 2505
rect 4217 2471 4240 2505
rect 4160 2433 4240 2471
rect 4160 2399 4183 2433
rect 4217 2399 4240 2433
rect 4160 2361 4240 2399
rect 4160 2327 4183 2361
rect 4217 2327 4240 2361
rect 4160 2289 4240 2327
rect 4160 2255 4183 2289
rect 4217 2255 4240 2289
rect 4160 2217 4240 2255
rect 4160 2183 4183 2217
rect 4217 2183 4240 2217
rect 4160 2145 4240 2183
rect 4160 2111 4183 2145
rect 4217 2111 4240 2145
rect 520 1977 2120 2000
rect 520 1943 547 1977
rect 581 1943 619 1977
rect 653 1943 691 1977
rect 725 1943 763 1977
rect 797 1943 835 1977
rect 869 1943 907 1977
rect 941 1943 979 1977
rect 1013 1943 1051 1977
rect 1085 1943 1123 1977
rect 1157 1943 1195 1977
rect 1229 1943 1267 1977
rect 1301 1943 1339 1977
rect 1373 1943 1411 1977
rect 1445 1943 1483 1977
rect 1517 1943 1555 1977
rect 1589 1943 1627 1977
rect 1661 1943 1699 1977
rect 1733 1943 1771 1977
rect 1805 1943 1843 1977
rect 1877 1943 1915 1977
rect 1949 1943 1987 1977
rect 2021 1943 2059 1977
rect 2093 1943 2120 1977
rect 520 1920 2120 1943
rect 2440 1977 4040 2000
rect 2440 1943 2467 1977
rect 2501 1943 2539 1977
rect 2573 1943 2611 1977
rect 2645 1943 2683 1977
rect 2717 1943 2755 1977
rect 2789 1943 2827 1977
rect 2861 1943 2899 1977
rect 2933 1943 2971 1977
rect 3005 1943 3043 1977
rect 3077 1943 3115 1977
rect 3149 1943 3187 1977
rect 3221 1943 3259 1977
rect 3293 1943 3331 1977
rect 3365 1943 3403 1977
rect 3437 1943 3475 1977
rect 3509 1943 3547 1977
rect 3581 1943 3619 1977
rect 3653 1943 3691 1977
rect 3725 1943 3763 1977
rect 3797 1943 3835 1977
rect 3869 1943 3907 1977
rect 3941 1943 3979 1977
rect 4013 1943 4040 1977
rect 2440 1920 4040 1943
rect 1280 1506 1360 1920
rect 1280 1454 1294 1506
rect 1346 1454 1360 1506
rect 480 1337 560 1360
rect 480 1303 503 1337
rect 537 1303 560 1337
rect 480 1280 560 1303
rect 640 1337 720 1360
rect 640 1303 663 1337
rect 697 1303 720 1337
rect 640 1280 720 1303
rect 800 1337 880 1360
rect 800 1303 823 1337
rect 857 1303 880 1337
rect 800 1280 880 1303
rect 960 1337 1040 1360
rect 960 1303 983 1337
rect 1017 1303 1040 1337
rect 960 1280 1040 1303
rect 1120 1337 1200 1360
rect 1120 1303 1143 1337
rect 1177 1303 1200 1337
rect 1120 1280 1200 1303
rect 320 1134 334 1186
rect 386 1134 400 1186
rect 320 713 400 1134
rect 1280 880 1360 1454
rect 3200 1506 3280 1920
rect 3200 1454 3214 1506
rect 3266 1454 3280 1506
rect 1440 1337 1520 1360
rect 1440 1303 1463 1337
rect 1497 1303 1520 1337
rect 1440 1280 1520 1303
rect 1600 1337 1680 1360
rect 1600 1303 1623 1337
rect 1657 1303 1680 1337
rect 1600 1280 1680 1303
rect 1760 1337 1840 1360
rect 1760 1303 1783 1337
rect 1817 1303 1840 1337
rect 1760 1280 1840 1303
rect 1920 1337 2000 1360
rect 1920 1303 1943 1337
rect 1977 1303 2000 1337
rect 1920 1280 2000 1303
rect 2080 1337 2160 1360
rect 2080 1303 2103 1337
rect 2137 1303 2160 1337
rect 2080 1280 2160 1303
rect 2240 1337 2320 1360
rect 2240 1303 2263 1337
rect 2297 1303 2320 1337
rect 2240 1280 2320 1303
rect 2400 1337 2480 1360
rect 2400 1303 2423 1337
rect 2457 1303 2480 1337
rect 2400 1280 2480 1303
rect 2560 1337 2640 1360
rect 2560 1303 2583 1337
rect 2617 1303 2640 1337
rect 2560 1280 2640 1303
rect 2720 1337 2800 1360
rect 2720 1303 2743 1337
rect 2777 1303 2800 1337
rect 2720 1280 2800 1303
rect 2880 1337 2960 1360
rect 2880 1303 2903 1337
rect 2937 1303 2960 1337
rect 2880 1280 2960 1303
rect 3040 1337 3120 1360
rect 3040 1303 3063 1337
rect 3097 1303 3120 1337
rect 3040 1280 3120 1303
rect 3200 880 3280 1454
rect 3360 1337 3440 1360
rect 3360 1303 3383 1337
rect 3417 1303 3440 1337
rect 3360 1280 3440 1303
rect 3520 1337 3600 1360
rect 3520 1303 3543 1337
rect 3577 1303 3600 1337
rect 3520 1280 3600 1303
rect 3680 1337 3760 1360
rect 3680 1303 3703 1337
rect 3737 1303 3760 1337
rect 3680 1280 3760 1303
rect 3840 1337 3920 1360
rect 3840 1303 3863 1337
rect 3897 1303 3920 1337
rect 3840 1280 3920 1303
rect 4000 1337 4080 1360
rect 4000 1303 4023 1337
rect 4057 1303 4080 1337
rect 4000 1280 4080 1303
rect 4160 1186 4240 2111
rect 6080 2649 6160 2734
rect 6080 2615 6103 2649
rect 6137 2615 6160 2649
rect 6080 2577 6160 2615
rect 6080 2543 6103 2577
rect 6137 2543 6160 2577
rect 6080 2505 6160 2543
rect 6080 2471 6103 2505
rect 6137 2471 6160 2505
rect 6080 2433 6160 2471
rect 6080 2399 6103 2433
rect 6137 2399 6160 2433
rect 6080 2361 6160 2399
rect 6080 2327 6103 2361
rect 6137 2327 6160 2361
rect 6080 2289 6160 2327
rect 6080 2255 6103 2289
rect 6137 2255 6160 2289
rect 6080 2217 6160 2255
rect 6080 2183 6103 2217
rect 6137 2183 6160 2217
rect 6080 2145 6160 2183
rect 6080 2111 6103 2145
rect 6137 2111 6160 2145
rect 6080 2080 6160 2111
rect 8000 2649 8080 2680
rect 8000 2615 8023 2649
rect 8057 2615 8080 2649
rect 8000 2577 8080 2615
rect 8000 2543 8023 2577
rect 8057 2543 8080 2577
rect 8000 2505 8080 2543
rect 8000 2471 8023 2505
rect 8057 2471 8080 2505
rect 8000 2433 8080 2471
rect 8000 2399 8023 2433
rect 8057 2399 8080 2433
rect 8000 2361 8080 2399
rect 8000 2327 8023 2361
rect 8057 2327 8080 2361
rect 8000 2289 8080 2327
rect 8000 2255 8023 2289
rect 8057 2255 8080 2289
rect 8000 2217 8080 2255
rect 8000 2183 8023 2217
rect 8057 2183 8080 2217
rect 8000 2145 8080 2183
rect 8000 2111 8023 2145
rect 8057 2111 8080 2145
rect 4360 1977 5960 2000
rect 4360 1943 4387 1977
rect 4421 1943 4459 1977
rect 4493 1943 4531 1977
rect 4565 1943 4603 1977
rect 4637 1943 4675 1977
rect 4709 1943 4747 1977
rect 4781 1943 4819 1977
rect 4853 1943 4891 1977
rect 4925 1943 4963 1977
rect 4997 1943 5035 1977
rect 5069 1943 5107 1977
rect 5141 1943 5179 1977
rect 5213 1943 5251 1977
rect 5285 1943 5323 1977
rect 5357 1943 5395 1977
rect 5429 1943 5467 1977
rect 5501 1943 5539 1977
rect 5573 1943 5611 1977
rect 5645 1943 5683 1977
rect 5717 1943 5755 1977
rect 5789 1943 5827 1977
rect 5861 1943 5899 1977
rect 5933 1943 5960 1977
rect 4360 1920 5960 1943
rect 6280 1977 7880 2000
rect 6280 1943 6307 1977
rect 6341 1943 6379 1977
rect 6413 1943 6451 1977
rect 6485 1943 6523 1977
rect 6557 1943 6595 1977
rect 6629 1943 6667 1977
rect 6701 1943 6739 1977
rect 6773 1943 6811 1977
rect 6845 1943 6883 1977
rect 6917 1943 6955 1977
rect 6989 1943 7027 1977
rect 7061 1943 7099 1977
rect 7133 1943 7171 1977
rect 7205 1943 7243 1977
rect 7277 1943 7315 1977
rect 7349 1943 7387 1977
rect 7421 1943 7459 1977
rect 7493 1943 7531 1977
rect 7565 1943 7603 1977
rect 7637 1943 7675 1977
rect 7709 1943 7747 1977
rect 7781 1943 7819 1977
rect 7853 1943 7880 1977
rect 6280 1920 7880 1943
rect 5120 1506 5200 1920
rect 5120 1454 5134 1506
rect 5186 1454 5200 1506
rect 4320 1337 4400 1360
rect 4320 1303 4343 1337
rect 4377 1303 4400 1337
rect 4320 1280 4400 1303
rect 4480 1337 4560 1360
rect 4480 1303 4503 1337
rect 4537 1303 4560 1337
rect 4480 1280 4560 1303
rect 4640 1337 4720 1360
rect 4640 1303 4663 1337
rect 4697 1303 4720 1337
rect 4640 1280 4720 1303
rect 4800 1337 4880 1360
rect 4800 1303 4823 1337
rect 4857 1303 4880 1337
rect 4800 1280 4880 1303
rect 4960 1337 5040 1360
rect 4960 1303 4983 1337
rect 5017 1303 5040 1337
rect 4960 1280 5040 1303
rect 4160 1134 4174 1186
rect 4226 1134 4240 1186
rect 520 857 2120 880
rect 520 823 547 857
rect 581 823 619 857
rect 653 823 691 857
rect 725 823 763 857
rect 797 823 835 857
rect 869 823 907 857
rect 941 823 979 857
rect 1013 823 1051 857
rect 1085 823 1123 857
rect 1157 823 1195 857
rect 1229 823 1267 857
rect 1301 823 1339 857
rect 1373 823 1411 857
rect 1445 823 1483 857
rect 1517 823 1555 857
rect 1589 823 1627 857
rect 1661 823 1699 857
rect 1733 823 1771 857
rect 1805 823 1843 857
rect 1877 823 1915 857
rect 1949 823 1987 857
rect 2021 823 2059 857
rect 2093 823 2120 857
rect 520 800 2120 823
rect 2440 857 4040 880
rect 2440 823 2467 857
rect 2501 823 2539 857
rect 2573 823 2611 857
rect 2645 823 2683 857
rect 2717 823 2755 857
rect 2789 823 2827 857
rect 2861 823 2899 857
rect 2933 823 2971 857
rect 3005 823 3043 857
rect 3077 823 3115 857
rect 3149 823 3187 857
rect 3221 823 3259 857
rect 3293 823 3331 857
rect 3365 823 3403 857
rect 3437 823 3475 857
rect 3509 823 3547 857
rect 3581 823 3619 857
rect 3653 823 3691 857
rect 3725 823 3763 857
rect 3797 823 3835 857
rect 3869 823 3907 857
rect 3941 823 3979 857
rect 4013 823 4040 857
rect 2440 800 4040 823
rect 320 679 343 713
rect 377 679 400 713
rect 320 641 400 679
rect 320 607 343 641
rect 377 607 400 641
rect 320 560 400 607
rect 2240 713 2320 760
rect 2240 679 2263 713
rect 2297 679 2320 713
rect 2240 641 2320 679
rect 2240 607 2263 641
rect 2297 607 2320 641
rect 2240 546 2320 607
rect 4160 713 4240 1134
rect 5120 880 5200 1454
rect 7040 1506 7120 1920
rect 7040 1454 7054 1506
rect 7106 1454 7120 1506
rect 5280 1337 5360 1360
rect 5280 1303 5303 1337
rect 5337 1303 5360 1337
rect 5280 1280 5360 1303
rect 5440 1337 5520 1360
rect 5440 1303 5463 1337
rect 5497 1303 5520 1337
rect 5440 1280 5520 1303
rect 5600 1337 5680 1360
rect 5600 1303 5623 1337
rect 5657 1303 5680 1337
rect 5600 1280 5680 1303
rect 5760 1337 5840 1360
rect 5760 1303 5783 1337
rect 5817 1303 5840 1337
rect 5760 1280 5840 1303
rect 5920 1337 6000 1360
rect 5920 1303 5943 1337
rect 5977 1303 6000 1337
rect 5920 1280 6000 1303
rect 6080 1337 6160 1360
rect 6080 1303 6103 1337
rect 6137 1303 6160 1337
rect 6080 1280 6160 1303
rect 6240 1337 6320 1360
rect 6240 1303 6263 1337
rect 6297 1303 6320 1337
rect 6240 1280 6320 1303
rect 6400 1337 6480 1360
rect 6400 1303 6423 1337
rect 6457 1303 6480 1337
rect 6400 1280 6480 1303
rect 6560 1337 6640 1360
rect 6560 1303 6583 1337
rect 6617 1303 6640 1337
rect 6560 1280 6640 1303
rect 6720 1337 6800 1360
rect 6720 1303 6743 1337
rect 6777 1303 6800 1337
rect 6720 1280 6800 1303
rect 6880 1337 6960 1360
rect 6880 1303 6903 1337
rect 6937 1303 6960 1337
rect 6880 1280 6960 1303
rect 7040 880 7120 1454
rect 7200 1337 7280 1360
rect 7200 1303 7223 1337
rect 7257 1303 7280 1337
rect 7200 1280 7280 1303
rect 7360 1337 7440 1360
rect 7360 1303 7383 1337
rect 7417 1303 7440 1337
rect 7360 1280 7440 1303
rect 7520 1337 7600 1360
rect 7520 1303 7543 1337
rect 7577 1303 7600 1337
rect 7520 1280 7600 1303
rect 7680 1337 7760 1360
rect 7680 1303 7703 1337
rect 7737 1303 7760 1337
rect 7680 1280 7760 1303
rect 7840 1337 7920 1360
rect 7840 1303 7863 1337
rect 7897 1303 7920 1337
rect 7840 1280 7920 1303
rect 8000 1186 8080 2111
rect 8160 1337 8240 1360
rect 8160 1303 8183 1337
rect 8217 1303 8240 1337
rect 8160 1280 8240 1303
rect 8000 1134 8014 1186
rect 8066 1134 8080 1186
rect 4360 857 5960 880
rect 4360 823 4387 857
rect 4421 823 4459 857
rect 4493 823 4531 857
rect 4565 823 4603 857
rect 4637 823 4675 857
rect 4709 823 4747 857
rect 4781 823 4819 857
rect 4853 823 4891 857
rect 4925 823 4963 857
rect 4997 823 5035 857
rect 5069 823 5107 857
rect 5141 823 5179 857
rect 5213 823 5251 857
rect 5285 823 5323 857
rect 5357 823 5395 857
rect 5429 823 5467 857
rect 5501 823 5539 857
rect 5573 823 5611 857
rect 5645 823 5683 857
rect 5717 823 5755 857
rect 5789 823 5827 857
rect 5861 823 5899 857
rect 5933 823 5960 857
rect 4360 800 5960 823
rect 6280 857 7880 880
rect 6280 823 6307 857
rect 6341 823 6379 857
rect 6413 823 6451 857
rect 6485 823 6523 857
rect 6557 823 6595 857
rect 6629 823 6667 857
rect 6701 823 6739 857
rect 6773 823 6811 857
rect 6845 823 6883 857
rect 6917 823 6955 857
rect 6989 823 7027 857
rect 7061 823 7099 857
rect 7133 823 7171 857
rect 7205 823 7243 857
rect 7277 823 7315 857
rect 7349 823 7387 857
rect 7421 823 7459 857
rect 7493 823 7531 857
rect 7565 823 7603 857
rect 7637 823 7675 857
rect 7709 823 7747 857
rect 7781 823 7819 857
rect 7853 823 7880 857
rect 6280 800 7880 823
rect 4160 679 4183 713
rect 4217 679 4240 713
rect 4160 641 4240 679
rect 4160 607 4183 641
rect 4217 607 4240 641
rect 4160 560 4240 607
rect 6080 713 6160 760
rect 6080 679 6103 713
rect 6137 679 6160 713
rect 6080 641 6160 679
rect 6080 607 6103 641
rect 6137 607 6160 641
rect 2240 494 2254 546
rect 2306 494 2320 546
rect 2240 480 2320 494
rect 6080 546 6160 607
rect 8000 713 8080 1134
rect 8000 679 8023 713
rect 8057 679 8080 713
rect 8000 641 8080 679
rect 8000 607 8023 641
rect 8057 607 8080 641
rect 8000 560 8080 607
rect 6080 494 6094 546
rect 6146 494 6160 546
rect 6080 480 6160 494
rect 320 318 400 360
rect 320 266 334 318
rect 386 266 400 318
rect 320 254 400 266
rect 320 202 334 254
rect 386 202 400 254
rect 320 160 400 202
rect 2240 313 2320 360
rect 2240 279 2263 313
rect 2297 279 2320 313
rect 2240 241 2320 279
rect 2240 207 2263 241
rect 2297 207 2320 241
rect 2240 160 2320 207
rect 4160 313 4240 400
rect 4160 279 4183 313
rect 4217 279 4240 313
rect 4160 241 4240 279
rect 4160 207 4183 241
rect 4217 207 4240 241
rect 4160 160 4240 207
rect 6080 313 6160 360
rect 6080 279 6103 313
rect 6137 279 6160 313
rect 6080 241 6160 279
rect 6080 207 6103 241
rect 6137 207 6160 241
rect 6080 160 6160 207
rect 8000 318 8080 360
rect 8000 266 8014 318
rect 8066 266 8080 318
rect 8000 254 8080 266
rect 8000 202 8014 254
rect 8066 202 8080 254
rect 8000 160 8080 202
<< via1 >>
rect 4174 5615 4183 5634
rect 4183 5615 4217 5634
rect 4217 5615 4226 5634
rect 4174 5582 4226 5615
rect 4174 5543 4183 5570
rect 4183 5543 4217 5570
rect 4217 5543 4226 5570
rect 4174 5518 4226 5543
rect 4174 5505 4226 5506
rect 4174 5471 4183 5505
rect 4183 5471 4217 5505
rect 4217 5471 4226 5505
rect 4174 5454 4226 5471
rect 4174 5433 4226 5442
rect 4174 5399 4183 5433
rect 4183 5399 4217 5433
rect 4217 5399 4226 5433
rect 4174 5390 4226 5399
rect 4174 5361 4226 5378
rect 4174 5327 4183 5361
rect 4183 5327 4217 5361
rect 4217 5327 4226 5361
rect 4174 5326 4226 5327
rect 14 3934 66 3986
rect 14 3614 66 3666
rect 174 3934 226 3986
rect 174 3614 226 3666
rect 334 3934 386 3986
rect 334 3614 386 3666
rect 494 3934 546 3986
rect 494 3614 546 3666
rect 654 3934 706 3986
rect 654 3614 706 3666
rect 814 3934 866 3986
rect 814 3614 866 3666
rect 974 3934 1026 3986
rect 974 3614 1026 3666
rect 1134 3934 1186 3986
rect 1294 3774 1346 3826
rect 1454 3934 1506 3986
rect 1134 3614 1186 3666
rect 1454 3614 1506 3666
rect 1614 3934 1666 3986
rect 1614 3614 1666 3666
rect 1774 3934 1826 3986
rect 1774 3614 1826 3666
rect 1934 3934 1986 3986
rect 1934 3614 1986 3666
rect 2094 3934 2146 3986
rect 2094 3614 2146 3666
rect 2254 3934 2306 3986
rect 2254 3614 2306 3666
rect 2414 3934 2466 3986
rect 2414 3614 2466 3666
rect 2574 3934 2626 3986
rect 2574 3614 2626 3666
rect 2734 3934 2786 3986
rect 2734 3614 2786 3666
rect 2894 3934 2946 3986
rect 2894 3614 2946 3666
rect 3054 3934 3106 3986
rect 3214 3774 3266 3826
rect 3374 3934 3426 3986
rect 3054 3614 3106 3666
rect 3374 3614 3426 3666
rect 3534 3934 3586 3986
rect 3534 3614 3586 3666
rect 3694 3934 3746 3986
rect 3694 3614 3746 3666
rect 3854 3934 3906 3986
rect 3854 3614 3906 3666
rect 4014 3934 4066 3986
rect 4014 3614 4066 3666
rect 4174 3934 4226 3986
rect 4174 3614 4226 3666
rect 4334 3934 4386 3986
rect 4334 3614 4386 3666
rect 4494 3934 4546 3986
rect 4494 3614 4546 3666
rect 4654 3934 4706 3986
rect 4654 3614 4706 3666
rect 4814 3934 4866 3986
rect 4814 3614 4866 3666
rect 4974 3934 5026 3986
rect 5134 3774 5186 3826
rect 5294 3934 5346 3986
rect 4974 3614 5026 3666
rect 5294 3614 5346 3666
rect 5454 3934 5506 3986
rect 5454 3614 5506 3666
rect 5614 3934 5666 3986
rect 5614 3614 5666 3666
rect 5774 3934 5826 3986
rect 5774 3614 5826 3666
rect 5934 3934 5986 3986
rect 5934 3614 5986 3666
rect 6094 3934 6146 3986
rect 6094 3614 6146 3666
rect 6254 3934 6306 3986
rect 6254 3614 6306 3666
rect 6414 3934 6466 3986
rect 6414 3614 6466 3666
rect 6574 3934 6626 3986
rect 6574 3614 6626 3666
rect 6734 3934 6786 3986
rect 6734 3614 6786 3666
rect 6894 3934 6946 3986
rect 7054 3774 7106 3826
rect 7214 3934 7266 3986
rect 6894 3614 6946 3666
rect 7214 3614 7266 3666
rect 7374 3934 7426 3986
rect 7374 3614 7426 3666
rect 7534 3934 7586 3986
rect 7534 3614 7586 3666
rect 7694 3934 7746 3986
rect 7694 3614 7746 3666
rect 7854 3934 7906 3986
rect 7854 3614 7906 3666
rect 8014 3934 8066 3986
rect 8014 3614 8066 3666
rect 8174 3934 8226 3986
rect 8174 3614 8226 3666
rect 8334 3934 8386 3986
rect 8334 3614 8386 3666
rect 2254 2734 2306 2786
rect 6094 2734 6146 2786
rect 1294 1454 1346 1506
rect 334 1134 386 1186
rect 3214 1454 3266 1506
rect 5134 1454 5186 1506
rect 4174 1134 4226 1186
rect 7054 1454 7106 1506
rect 8014 1134 8066 1186
rect 2254 494 2306 546
rect 6094 494 6146 546
rect 334 313 386 318
rect 334 279 343 313
rect 343 279 377 313
rect 377 279 386 313
rect 334 266 386 279
rect 334 241 386 254
rect 334 207 343 241
rect 343 207 377 241
rect 377 207 386 241
rect 334 202 386 207
rect 8014 313 8066 318
rect 8014 279 8023 313
rect 8023 279 8057 313
rect 8057 279 8066 313
rect 8014 266 8066 279
rect 8014 241 8066 254
rect 8014 207 8023 241
rect 8023 207 8057 241
rect 8057 207 8066 241
rect 8014 202 8066 207
<< metal2 >>
rect 4160 5634 4240 5680
rect 4160 5628 4174 5634
rect 4226 5628 4240 5634
rect 4160 5572 4172 5628
rect 4228 5572 4240 5628
rect 4160 5570 4240 5572
rect 4160 5548 4174 5570
rect 4226 5548 4240 5570
rect 4160 5492 4172 5548
rect 4228 5492 4240 5548
rect 4160 5468 4174 5492
rect 4226 5468 4240 5492
rect 4160 5412 4172 5468
rect 4228 5412 4240 5468
rect 4160 5390 4174 5412
rect 4226 5390 4240 5412
rect 4160 5388 4240 5390
rect 4160 5332 4172 5388
rect 4228 5332 4240 5388
rect 4160 5326 4174 5332
rect 4226 5326 4240 5332
rect 4160 5280 4240 5326
rect 0 3988 8400 4000
rect 0 3932 12 3988
rect 68 3932 172 3988
rect 228 3932 332 3988
rect 388 3932 492 3988
rect 548 3932 652 3988
rect 708 3932 812 3988
rect 868 3932 972 3988
rect 1028 3932 1132 3988
rect 1188 3932 1452 3988
rect 1508 3932 1612 3988
rect 1668 3932 1772 3988
rect 1828 3932 1932 3988
rect 1988 3932 2092 3988
rect 2148 3932 2252 3988
rect 2308 3932 2412 3988
rect 2468 3932 2572 3988
rect 2628 3932 2732 3988
rect 2788 3932 2892 3988
rect 2948 3932 3052 3988
rect 3108 3932 3372 3988
rect 3428 3932 3532 3988
rect 3588 3932 3692 3988
rect 3748 3932 3852 3988
rect 3908 3932 4012 3988
rect 4068 3932 4172 3988
rect 4228 3932 4332 3988
rect 4388 3932 4492 3988
rect 4548 3932 4652 3988
rect 4708 3932 4812 3988
rect 4868 3932 4972 3988
rect 5028 3932 5292 3988
rect 5348 3932 5452 3988
rect 5508 3932 5612 3988
rect 5668 3932 5772 3988
rect 5828 3932 5932 3988
rect 5988 3932 6092 3988
rect 6148 3932 6252 3988
rect 6308 3932 6412 3988
rect 6468 3932 6572 3988
rect 6628 3932 6732 3988
rect 6788 3932 6892 3988
rect 6948 3932 7212 3988
rect 7268 3932 7372 3988
rect 7428 3932 7532 3988
rect 7588 3932 7692 3988
rect 7748 3932 7852 3988
rect 7908 3932 8012 3988
rect 8068 3932 8172 3988
rect 8228 3932 8332 3988
rect 8388 3932 8400 3988
rect 0 3920 8400 3932
rect 0 3826 8400 3840
rect 0 3774 1294 3826
rect 1346 3774 3214 3826
rect 3266 3774 5134 3826
rect 5186 3774 7054 3826
rect 7106 3774 8400 3826
rect 0 3760 8400 3774
rect 0 3668 8400 3680
rect 0 3612 12 3668
rect 68 3612 172 3668
rect 228 3612 332 3668
rect 388 3612 492 3668
rect 548 3612 652 3668
rect 708 3612 812 3668
rect 868 3612 972 3668
rect 1028 3612 1132 3668
rect 1188 3612 1452 3668
rect 1508 3612 1612 3668
rect 1668 3612 1772 3668
rect 1828 3612 1932 3668
rect 1988 3612 2092 3668
rect 2148 3612 2252 3668
rect 2308 3612 2412 3668
rect 2468 3612 2572 3668
rect 2628 3612 2732 3668
rect 2788 3612 2892 3668
rect 2948 3612 3052 3668
rect 3108 3612 3372 3668
rect 3428 3612 3532 3668
rect 3588 3612 3692 3668
rect 3748 3612 3852 3668
rect 3908 3612 4012 3668
rect 4068 3612 4172 3668
rect 4228 3612 4332 3668
rect 4388 3612 4492 3668
rect 4548 3612 4652 3668
rect 4708 3612 4812 3668
rect 4868 3612 4972 3668
rect 5028 3612 5292 3668
rect 5348 3612 5452 3668
rect 5508 3612 5612 3668
rect 5668 3612 5772 3668
rect 5828 3612 5932 3668
rect 5988 3612 6092 3668
rect 6148 3612 6252 3668
rect 6308 3612 6412 3668
rect 6468 3612 6572 3668
rect 6628 3612 6732 3668
rect 6788 3612 6892 3668
rect 6948 3612 7212 3668
rect 7268 3612 7372 3668
rect 7428 3612 7532 3668
rect 7588 3612 7692 3668
rect 7748 3612 7852 3668
rect 7908 3612 8012 3668
rect 8068 3612 8172 3668
rect 8228 3612 8332 3668
rect 8388 3612 8400 3668
rect 0 3600 8400 3612
rect 0 2786 8400 2800
rect 0 2734 2254 2786
rect 2306 2734 6094 2786
rect 6146 2734 8400 2786
rect 0 2720 8400 2734
rect 0 1668 8400 1680
rect 0 1612 172 1668
rect 228 1612 492 1668
rect 548 1612 652 1668
rect 708 1612 812 1668
rect 868 1612 972 1668
rect 1028 1612 1132 1668
rect 1188 1612 1452 1668
rect 1508 1612 1612 1668
rect 1668 1612 1772 1668
rect 1828 1612 1932 1668
rect 1988 1612 2092 1668
rect 2148 1612 2252 1668
rect 2308 1612 2412 1668
rect 2468 1612 2572 1668
rect 2628 1612 2732 1668
rect 2788 1612 2892 1668
rect 2948 1612 3052 1668
rect 3108 1612 3372 1668
rect 3428 1612 3532 1668
rect 3588 1612 3692 1668
rect 3748 1612 3852 1668
rect 3908 1612 4012 1668
rect 4068 1612 4332 1668
rect 4388 1612 4492 1668
rect 4548 1612 4652 1668
rect 4708 1612 4812 1668
rect 4868 1612 4972 1668
rect 5028 1612 5292 1668
rect 5348 1612 5452 1668
rect 5508 1612 5612 1668
rect 5668 1612 5772 1668
rect 5828 1612 5932 1668
rect 5988 1612 6092 1668
rect 6148 1612 6252 1668
rect 6308 1612 6412 1668
rect 6468 1612 6572 1668
rect 6628 1612 6732 1668
rect 6788 1612 6892 1668
rect 6948 1612 7212 1668
rect 7268 1612 7372 1668
rect 7428 1612 7532 1668
rect 7588 1612 7692 1668
rect 7748 1612 7852 1668
rect 7908 1612 8172 1668
rect 8228 1612 8400 1668
rect 0 1600 8400 1612
rect 0 1506 8400 1520
rect 0 1454 1294 1506
rect 1346 1454 3214 1506
rect 3266 1454 5134 1506
rect 5186 1454 7054 1506
rect 7106 1454 8400 1506
rect 0 1440 8400 1454
rect 0 1348 8400 1360
rect 0 1292 172 1348
rect 228 1292 492 1348
rect 548 1292 652 1348
rect 708 1292 812 1348
rect 868 1292 972 1348
rect 1028 1292 1132 1348
rect 1188 1292 1452 1348
rect 1508 1292 1612 1348
rect 1668 1292 1772 1348
rect 1828 1292 1932 1348
rect 1988 1292 2092 1348
rect 2148 1292 2252 1348
rect 2308 1292 2412 1348
rect 2468 1292 2572 1348
rect 2628 1292 2732 1348
rect 2788 1292 2892 1348
rect 2948 1292 3052 1348
rect 3108 1292 3372 1348
rect 3428 1292 3532 1348
rect 3588 1292 3692 1348
rect 3748 1292 3852 1348
rect 3908 1292 4012 1348
rect 4068 1292 4332 1348
rect 4388 1292 4492 1348
rect 4548 1292 4652 1348
rect 4708 1292 4812 1348
rect 4868 1292 4972 1348
rect 5028 1292 5292 1348
rect 5348 1292 5452 1348
rect 5508 1292 5612 1348
rect 5668 1292 5772 1348
rect 5828 1292 5932 1348
rect 5988 1292 6092 1348
rect 6148 1292 6252 1348
rect 6308 1292 6412 1348
rect 6468 1292 6572 1348
rect 6628 1292 6732 1348
rect 6788 1292 6892 1348
rect 6948 1292 7212 1348
rect 7268 1292 7372 1348
rect 7428 1292 7532 1348
rect 7588 1292 7692 1348
rect 7748 1292 7852 1348
rect 7908 1292 8172 1348
rect 8228 1292 8400 1348
rect 0 1280 8400 1292
rect 0 1186 8400 1200
rect 0 1134 334 1186
rect 386 1134 4174 1186
rect 4226 1134 8014 1186
rect 8066 1134 8400 1186
rect 0 1120 8400 1134
rect 0 1028 8400 1040
rect 0 972 172 1028
rect 228 972 492 1028
rect 548 972 652 1028
rect 708 972 812 1028
rect 868 972 972 1028
rect 1028 972 1132 1028
rect 1188 972 1452 1028
rect 1508 972 1612 1028
rect 1668 972 1772 1028
rect 1828 972 1932 1028
rect 1988 972 2092 1028
rect 2148 972 2252 1028
rect 2308 972 2412 1028
rect 2468 972 2572 1028
rect 2628 972 2732 1028
rect 2788 972 2892 1028
rect 2948 972 3052 1028
rect 3108 972 3372 1028
rect 3428 972 3532 1028
rect 3588 972 3692 1028
rect 3748 972 3852 1028
rect 3908 972 4012 1028
rect 4068 972 4332 1028
rect 4388 972 4492 1028
rect 4548 972 4652 1028
rect 4708 972 4812 1028
rect 4868 972 4972 1028
rect 5028 972 5292 1028
rect 5348 972 5452 1028
rect 5508 972 5612 1028
rect 5668 972 5772 1028
rect 5828 972 5932 1028
rect 5988 972 6092 1028
rect 6148 972 6252 1028
rect 6308 972 6412 1028
rect 6468 972 6572 1028
rect 6628 972 6732 1028
rect 6788 972 6892 1028
rect 6948 972 7212 1028
rect 7268 972 7372 1028
rect 7428 972 7532 1028
rect 7588 972 7692 1028
rect 7748 972 7852 1028
rect 7908 972 8172 1028
rect 8228 972 8400 1028
rect 0 960 8400 972
rect 0 546 8400 560
rect 0 494 2254 546
rect 2306 494 6094 546
rect 6146 494 8400 546
rect 0 480 8400 494
rect 320 328 400 360
rect 320 272 332 328
rect 388 272 400 328
rect 320 266 334 272
rect 386 266 400 272
rect 320 254 400 266
rect 320 248 334 254
rect 386 248 400 254
rect 320 192 332 248
rect 388 192 400 248
rect 320 160 400 192
rect 8000 328 8080 360
rect 8000 272 8012 328
rect 8068 272 8080 328
rect 8000 266 8014 272
rect 8066 266 8080 272
rect 8000 254 8080 266
rect 8000 248 8014 254
rect 8066 248 8080 254
rect 8000 192 8012 248
rect 8068 192 8080 248
rect 8000 160 8080 192
<< via2 >>
rect 4172 5582 4174 5628
rect 4174 5582 4226 5628
rect 4226 5582 4228 5628
rect 4172 5572 4228 5582
rect 4172 5518 4174 5548
rect 4174 5518 4226 5548
rect 4226 5518 4228 5548
rect 4172 5506 4228 5518
rect 4172 5492 4174 5506
rect 4174 5492 4226 5506
rect 4226 5492 4228 5506
rect 4172 5454 4174 5468
rect 4174 5454 4226 5468
rect 4226 5454 4228 5468
rect 4172 5442 4228 5454
rect 4172 5412 4174 5442
rect 4174 5412 4226 5442
rect 4226 5412 4228 5442
rect 4172 5378 4228 5388
rect 4172 5332 4174 5378
rect 4174 5332 4226 5378
rect 4226 5332 4228 5378
rect 12 3986 68 3988
rect 12 3934 14 3986
rect 14 3934 66 3986
rect 66 3934 68 3986
rect 12 3932 68 3934
rect 172 3986 228 3988
rect 172 3934 174 3986
rect 174 3934 226 3986
rect 226 3934 228 3986
rect 172 3932 228 3934
rect 332 3986 388 3988
rect 332 3934 334 3986
rect 334 3934 386 3986
rect 386 3934 388 3986
rect 332 3932 388 3934
rect 492 3986 548 3988
rect 492 3934 494 3986
rect 494 3934 546 3986
rect 546 3934 548 3986
rect 492 3932 548 3934
rect 652 3986 708 3988
rect 652 3934 654 3986
rect 654 3934 706 3986
rect 706 3934 708 3986
rect 652 3932 708 3934
rect 812 3986 868 3988
rect 812 3934 814 3986
rect 814 3934 866 3986
rect 866 3934 868 3986
rect 812 3932 868 3934
rect 972 3986 1028 3988
rect 972 3934 974 3986
rect 974 3934 1026 3986
rect 1026 3934 1028 3986
rect 972 3932 1028 3934
rect 1132 3986 1188 3988
rect 1132 3934 1134 3986
rect 1134 3934 1186 3986
rect 1186 3934 1188 3986
rect 1132 3932 1188 3934
rect 1452 3986 1508 3988
rect 1452 3934 1454 3986
rect 1454 3934 1506 3986
rect 1506 3934 1508 3986
rect 1452 3932 1508 3934
rect 1612 3986 1668 3988
rect 1612 3934 1614 3986
rect 1614 3934 1666 3986
rect 1666 3934 1668 3986
rect 1612 3932 1668 3934
rect 1772 3986 1828 3988
rect 1772 3934 1774 3986
rect 1774 3934 1826 3986
rect 1826 3934 1828 3986
rect 1772 3932 1828 3934
rect 1932 3986 1988 3988
rect 1932 3934 1934 3986
rect 1934 3934 1986 3986
rect 1986 3934 1988 3986
rect 1932 3932 1988 3934
rect 2092 3986 2148 3988
rect 2092 3934 2094 3986
rect 2094 3934 2146 3986
rect 2146 3934 2148 3986
rect 2092 3932 2148 3934
rect 2252 3986 2308 3988
rect 2252 3934 2254 3986
rect 2254 3934 2306 3986
rect 2306 3934 2308 3986
rect 2252 3932 2308 3934
rect 2412 3986 2468 3988
rect 2412 3934 2414 3986
rect 2414 3934 2466 3986
rect 2466 3934 2468 3986
rect 2412 3932 2468 3934
rect 2572 3986 2628 3988
rect 2572 3934 2574 3986
rect 2574 3934 2626 3986
rect 2626 3934 2628 3986
rect 2572 3932 2628 3934
rect 2732 3986 2788 3988
rect 2732 3934 2734 3986
rect 2734 3934 2786 3986
rect 2786 3934 2788 3986
rect 2732 3932 2788 3934
rect 2892 3986 2948 3988
rect 2892 3934 2894 3986
rect 2894 3934 2946 3986
rect 2946 3934 2948 3986
rect 2892 3932 2948 3934
rect 3052 3986 3108 3988
rect 3052 3934 3054 3986
rect 3054 3934 3106 3986
rect 3106 3934 3108 3986
rect 3052 3932 3108 3934
rect 3372 3986 3428 3988
rect 3372 3934 3374 3986
rect 3374 3934 3426 3986
rect 3426 3934 3428 3986
rect 3372 3932 3428 3934
rect 3532 3986 3588 3988
rect 3532 3934 3534 3986
rect 3534 3934 3586 3986
rect 3586 3934 3588 3986
rect 3532 3932 3588 3934
rect 3692 3986 3748 3988
rect 3692 3934 3694 3986
rect 3694 3934 3746 3986
rect 3746 3934 3748 3986
rect 3692 3932 3748 3934
rect 3852 3986 3908 3988
rect 3852 3934 3854 3986
rect 3854 3934 3906 3986
rect 3906 3934 3908 3986
rect 3852 3932 3908 3934
rect 4012 3986 4068 3988
rect 4012 3934 4014 3986
rect 4014 3934 4066 3986
rect 4066 3934 4068 3986
rect 4012 3932 4068 3934
rect 4172 3986 4228 3988
rect 4172 3934 4174 3986
rect 4174 3934 4226 3986
rect 4226 3934 4228 3986
rect 4172 3932 4228 3934
rect 4332 3986 4388 3988
rect 4332 3934 4334 3986
rect 4334 3934 4386 3986
rect 4386 3934 4388 3986
rect 4332 3932 4388 3934
rect 4492 3986 4548 3988
rect 4492 3934 4494 3986
rect 4494 3934 4546 3986
rect 4546 3934 4548 3986
rect 4492 3932 4548 3934
rect 4652 3986 4708 3988
rect 4652 3934 4654 3986
rect 4654 3934 4706 3986
rect 4706 3934 4708 3986
rect 4652 3932 4708 3934
rect 4812 3986 4868 3988
rect 4812 3934 4814 3986
rect 4814 3934 4866 3986
rect 4866 3934 4868 3986
rect 4812 3932 4868 3934
rect 4972 3986 5028 3988
rect 4972 3934 4974 3986
rect 4974 3934 5026 3986
rect 5026 3934 5028 3986
rect 4972 3932 5028 3934
rect 5292 3986 5348 3988
rect 5292 3934 5294 3986
rect 5294 3934 5346 3986
rect 5346 3934 5348 3986
rect 5292 3932 5348 3934
rect 5452 3986 5508 3988
rect 5452 3934 5454 3986
rect 5454 3934 5506 3986
rect 5506 3934 5508 3986
rect 5452 3932 5508 3934
rect 5612 3986 5668 3988
rect 5612 3934 5614 3986
rect 5614 3934 5666 3986
rect 5666 3934 5668 3986
rect 5612 3932 5668 3934
rect 5772 3986 5828 3988
rect 5772 3934 5774 3986
rect 5774 3934 5826 3986
rect 5826 3934 5828 3986
rect 5772 3932 5828 3934
rect 5932 3986 5988 3988
rect 5932 3934 5934 3986
rect 5934 3934 5986 3986
rect 5986 3934 5988 3986
rect 5932 3932 5988 3934
rect 6092 3986 6148 3988
rect 6092 3934 6094 3986
rect 6094 3934 6146 3986
rect 6146 3934 6148 3986
rect 6092 3932 6148 3934
rect 6252 3986 6308 3988
rect 6252 3934 6254 3986
rect 6254 3934 6306 3986
rect 6306 3934 6308 3986
rect 6252 3932 6308 3934
rect 6412 3986 6468 3988
rect 6412 3934 6414 3986
rect 6414 3934 6466 3986
rect 6466 3934 6468 3986
rect 6412 3932 6468 3934
rect 6572 3986 6628 3988
rect 6572 3934 6574 3986
rect 6574 3934 6626 3986
rect 6626 3934 6628 3986
rect 6572 3932 6628 3934
rect 6732 3986 6788 3988
rect 6732 3934 6734 3986
rect 6734 3934 6786 3986
rect 6786 3934 6788 3986
rect 6732 3932 6788 3934
rect 6892 3986 6948 3988
rect 6892 3934 6894 3986
rect 6894 3934 6946 3986
rect 6946 3934 6948 3986
rect 6892 3932 6948 3934
rect 7212 3986 7268 3988
rect 7212 3934 7214 3986
rect 7214 3934 7266 3986
rect 7266 3934 7268 3986
rect 7212 3932 7268 3934
rect 7372 3986 7428 3988
rect 7372 3934 7374 3986
rect 7374 3934 7426 3986
rect 7426 3934 7428 3986
rect 7372 3932 7428 3934
rect 7532 3986 7588 3988
rect 7532 3934 7534 3986
rect 7534 3934 7586 3986
rect 7586 3934 7588 3986
rect 7532 3932 7588 3934
rect 7692 3986 7748 3988
rect 7692 3934 7694 3986
rect 7694 3934 7746 3986
rect 7746 3934 7748 3986
rect 7692 3932 7748 3934
rect 7852 3986 7908 3988
rect 7852 3934 7854 3986
rect 7854 3934 7906 3986
rect 7906 3934 7908 3986
rect 7852 3932 7908 3934
rect 8012 3986 8068 3988
rect 8012 3934 8014 3986
rect 8014 3934 8066 3986
rect 8066 3934 8068 3986
rect 8012 3932 8068 3934
rect 8172 3986 8228 3988
rect 8172 3934 8174 3986
rect 8174 3934 8226 3986
rect 8226 3934 8228 3986
rect 8172 3932 8228 3934
rect 8332 3986 8388 3988
rect 8332 3934 8334 3986
rect 8334 3934 8386 3986
rect 8386 3934 8388 3986
rect 8332 3932 8388 3934
rect 12 3666 68 3668
rect 12 3614 14 3666
rect 14 3614 66 3666
rect 66 3614 68 3666
rect 12 3612 68 3614
rect 172 3666 228 3668
rect 172 3614 174 3666
rect 174 3614 226 3666
rect 226 3614 228 3666
rect 172 3612 228 3614
rect 332 3666 388 3668
rect 332 3614 334 3666
rect 334 3614 386 3666
rect 386 3614 388 3666
rect 332 3612 388 3614
rect 492 3666 548 3668
rect 492 3614 494 3666
rect 494 3614 546 3666
rect 546 3614 548 3666
rect 492 3612 548 3614
rect 652 3666 708 3668
rect 652 3614 654 3666
rect 654 3614 706 3666
rect 706 3614 708 3666
rect 652 3612 708 3614
rect 812 3666 868 3668
rect 812 3614 814 3666
rect 814 3614 866 3666
rect 866 3614 868 3666
rect 812 3612 868 3614
rect 972 3666 1028 3668
rect 972 3614 974 3666
rect 974 3614 1026 3666
rect 1026 3614 1028 3666
rect 972 3612 1028 3614
rect 1132 3666 1188 3668
rect 1132 3614 1134 3666
rect 1134 3614 1186 3666
rect 1186 3614 1188 3666
rect 1132 3612 1188 3614
rect 1452 3666 1508 3668
rect 1452 3614 1454 3666
rect 1454 3614 1506 3666
rect 1506 3614 1508 3666
rect 1452 3612 1508 3614
rect 1612 3666 1668 3668
rect 1612 3614 1614 3666
rect 1614 3614 1666 3666
rect 1666 3614 1668 3666
rect 1612 3612 1668 3614
rect 1772 3666 1828 3668
rect 1772 3614 1774 3666
rect 1774 3614 1826 3666
rect 1826 3614 1828 3666
rect 1772 3612 1828 3614
rect 1932 3666 1988 3668
rect 1932 3614 1934 3666
rect 1934 3614 1986 3666
rect 1986 3614 1988 3666
rect 1932 3612 1988 3614
rect 2092 3666 2148 3668
rect 2092 3614 2094 3666
rect 2094 3614 2146 3666
rect 2146 3614 2148 3666
rect 2092 3612 2148 3614
rect 2252 3666 2308 3668
rect 2252 3614 2254 3666
rect 2254 3614 2306 3666
rect 2306 3614 2308 3666
rect 2252 3612 2308 3614
rect 2412 3666 2468 3668
rect 2412 3614 2414 3666
rect 2414 3614 2466 3666
rect 2466 3614 2468 3666
rect 2412 3612 2468 3614
rect 2572 3666 2628 3668
rect 2572 3614 2574 3666
rect 2574 3614 2626 3666
rect 2626 3614 2628 3666
rect 2572 3612 2628 3614
rect 2732 3666 2788 3668
rect 2732 3614 2734 3666
rect 2734 3614 2786 3666
rect 2786 3614 2788 3666
rect 2732 3612 2788 3614
rect 2892 3666 2948 3668
rect 2892 3614 2894 3666
rect 2894 3614 2946 3666
rect 2946 3614 2948 3666
rect 2892 3612 2948 3614
rect 3052 3666 3108 3668
rect 3052 3614 3054 3666
rect 3054 3614 3106 3666
rect 3106 3614 3108 3666
rect 3052 3612 3108 3614
rect 3372 3666 3428 3668
rect 3372 3614 3374 3666
rect 3374 3614 3426 3666
rect 3426 3614 3428 3666
rect 3372 3612 3428 3614
rect 3532 3666 3588 3668
rect 3532 3614 3534 3666
rect 3534 3614 3586 3666
rect 3586 3614 3588 3666
rect 3532 3612 3588 3614
rect 3692 3666 3748 3668
rect 3692 3614 3694 3666
rect 3694 3614 3746 3666
rect 3746 3614 3748 3666
rect 3692 3612 3748 3614
rect 3852 3666 3908 3668
rect 3852 3614 3854 3666
rect 3854 3614 3906 3666
rect 3906 3614 3908 3666
rect 3852 3612 3908 3614
rect 4012 3666 4068 3668
rect 4012 3614 4014 3666
rect 4014 3614 4066 3666
rect 4066 3614 4068 3666
rect 4012 3612 4068 3614
rect 4172 3666 4228 3668
rect 4172 3614 4174 3666
rect 4174 3614 4226 3666
rect 4226 3614 4228 3666
rect 4172 3612 4228 3614
rect 4332 3666 4388 3668
rect 4332 3614 4334 3666
rect 4334 3614 4386 3666
rect 4386 3614 4388 3666
rect 4332 3612 4388 3614
rect 4492 3666 4548 3668
rect 4492 3614 4494 3666
rect 4494 3614 4546 3666
rect 4546 3614 4548 3666
rect 4492 3612 4548 3614
rect 4652 3666 4708 3668
rect 4652 3614 4654 3666
rect 4654 3614 4706 3666
rect 4706 3614 4708 3666
rect 4652 3612 4708 3614
rect 4812 3666 4868 3668
rect 4812 3614 4814 3666
rect 4814 3614 4866 3666
rect 4866 3614 4868 3666
rect 4812 3612 4868 3614
rect 4972 3666 5028 3668
rect 4972 3614 4974 3666
rect 4974 3614 5026 3666
rect 5026 3614 5028 3666
rect 4972 3612 5028 3614
rect 5292 3666 5348 3668
rect 5292 3614 5294 3666
rect 5294 3614 5346 3666
rect 5346 3614 5348 3666
rect 5292 3612 5348 3614
rect 5452 3666 5508 3668
rect 5452 3614 5454 3666
rect 5454 3614 5506 3666
rect 5506 3614 5508 3666
rect 5452 3612 5508 3614
rect 5612 3666 5668 3668
rect 5612 3614 5614 3666
rect 5614 3614 5666 3666
rect 5666 3614 5668 3666
rect 5612 3612 5668 3614
rect 5772 3666 5828 3668
rect 5772 3614 5774 3666
rect 5774 3614 5826 3666
rect 5826 3614 5828 3666
rect 5772 3612 5828 3614
rect 5932 3666 5988 3668
rect 5932 3614 5934 3666
rect 5934 3614 5986 3666
rect 5986 3614 5988 3666
rect 5932 3612 5988 3614
rect 6092 3666 6148 3668
rect 6092 3614 6094 3666
rect 6094 3614 6146 3666
rect 6146 3614 6148 3666
rect 6092 3612 6148 3614
rect 6252 3666 6308 3668
rect 6252 3614 6254 3666
rect 6254 3614 6306 3666
rect 6306 3614 6308 3666
rect 6252 3612 6308 3614
rect 6412 3666 6468 3668
rect 6412 3614 6414 3666
rect 6414 3614 6466 3666
rect 6466 3614 6468 3666
rect 6412 3612 6468 3614
rect 6572 3666 6628 3668
rect 6572 3614 6574 3666
rect 6574 3614 6626 3666
rect 6626 3614 6628 3666
rect 6572 3612 6628 3614
rect 6732 3666 6788 3668
rect 6732 3614 6734 3666
rect 6734 3614 6786 3666
rect 6786 3614 6788 3666
rect 6732 3612 6788 3614
rect 6892 3666 6948 3668
rect 6892 3614 6894 3666
rect 6894 3614 6946 3666
rect 6946 3614 6948 3666
rect 6892 3612 6948 3614
rect 7212 3666 7268 3668
rect 7212 3614 7214 3666
rect 7214 3614 7266 3666
rect 7266 3614 7268 3666
rect 7212 3612 7268 3614
rect 7372 3666 7428 3668
rect 7372 3614 7374 3666
rect 7374 3614 7426 3666
rect 7426 3614 7428 3666
rect 7372 3612 7428 3614
rect 7532 3666 7588 3668
rect 7532 3614 7534 3666
rect 7534 3614 7586 3666
rect 7586 3614 7588 3666
rect 7532 3612 7588 3614
rect 7692 3666 7748 3668
rect 7692 3614 7694 3666
rect 7694 3614 7746 3666
rect 7746 3614 7748 3666
rect 7692 3612 7748 3614
rect 7852 3666 7908 3668
rect 7852 3614 7854 3666
rect 7854 3614 7906 3666
rect 7906 3614 7908 3666
rect 7852 3612 7908 3614
rect 8012 3666 8068 3668
rect 8012 3614 8014 3666
rect 8014 3614 8066 3666
rect 8066 3614 8068 3666
rect 8012 3612 8068 3614
rect 8172 3666 8228 3668
rect 8172 3614 8174 3666
rect 8174 3614 8226 3666
rect 8226 3614 8228 3666
rect 8172 3612 8228 3614
rect 8332 3666 8388 3668
rect 8332 3614 8334 3666
rect 8334 3614 8386 3666
rect 8386 3614 8388 3666
rect 8332 3612 8388 3614
rect 172 1612 228 1668
rect 492 1612 548 1668
rect 652 1612 708 1668
rect 812 1612 868 1668
rect 972 1612 1028 1668
rect 1132 1612 1188 1668
rect 1452 1612 1508 1668
rect 1612 1612 1668 1668
rect 1772 1612 1828 1668
rect 1932 1612 1988 1668
rect 2092 1612 2148 1668
rect 2252 1612 2308 1668
rect 2412 1612 2468 1668
rect 2572 1612 2628 1668
rect 2732 1612 2788 1668
rect 2892 1612 2948 1668
rect 3052 1612 3108 1668
rect 3372 1612 3428 1668
rect 3532 1612 3588 1668
rect 3692 1612 3748 1668
rect 3852 1612 3908 1668
rect 4012 1612 4068 1668
rect 4332 1612 4388 1668
rect 4492 1612 4548 1668
rect 4652 1612 4708 1668
rect 4812 1612 4868 1668
rect 4972 1612 5028 1668
rect 5292 1612 5348 1668
rect 5452 1612 5508 1668
rect 5612 1612 5668 1668
rect 5772 1612 5828 1668
rect 5932 1612 5988 1668
rect 6092 1612 6148 1668
rect 6252 1612 6308 1668
rect 6412 1612 6468 1668
rect 6572 1612 6628 1668
rect 6732 1612 6788 1668
rect 6892 1612 6948 1668
rect 7212 1612 7268 1668
rect 7372 1612 7428 1668
rect 7532 1612 7588 1668
rect 7692 1612 7748 1668
rect 7852 1612 7908 1668
rect 8172 1612 8228 1668
rect 172 1292 228 1348
rect 492 1292 548 1348
rect 652 1292 708 1348
rect 812 1292 868 1348
rect 972 1292 1028 1348
rect 1132 1292 1188 1348
rect 1452 1292 1508 1348
rect 1612 1292 1668 1348
rect 1772 1292 1828 1348
rect 1932 1292 1988 1348
rect 2092 1292 2148 1348
rect 2252 1292 2308 1348
rect 2412 1292 2468 1348
rect 2572 1292 2628 1348
rect 2732 1292 2788 1348
rect 2892 1292 2948 1348
rect 3052 1292 3108 1348
rect 3372 1292 3428 1348
rect 3532 1292 3588 1348
rect 3692 1292 3748 1348
rect 3852 1292 3908 1348
rect 4012 1292 4068 1348
rect 4332 1292 4388 1348
rect 4492 1292 4548 1348
rect 4652 1292 4708 1348
rect 4812 1292 4868 1348
rect 4972 1292 5028 1348
rect 5292 1292 5348 1348
rect 5452 1292 5508 1348
rect 5612 1292 5668 1348
rect 5772 1292 5828 1348
rect 5932 1292 5988 1348
rect 6092 1292 6148 1348
rect 6252 1292 6308 1348
rect 6412 1292 6468 1348
rect 6572 1292 6628 1348
rect 6732 1292 6788 1348
rect 6892 1292 6948 1348
rect 7212 1292 7268 1348
rect 7372 1292 7428 1348
rect 7532 1292 7588 1348
rect 7692 1292 7748 1348
rect 7852 1292 7908 1348
rect 8172 1292 8228 1348
rect 172 972 228 1028
rect 492 972 548 1028
rect 652 972 708 1028
rect 812 972 868 1028
rect 972 972 1028 1028
rect 1132 972 1188 1028
rect 1452 972 1508 1028
rect 1612 972 1668 1028
rect 1772 972 1828 1028
rect 1932 972 1988 1028
rect 2092 972 2148 1028
rect 2252 972 2308 1028
rect 2412 972 2468 1028
rect 2572 972 2628 1028
rect 2732 972 2788 1028
rect 2892 972 2948 1028
rect 3052 972 3108 1028
rect 3372 972 3428 1028
rect 3532 972 3588 1028
rect 3692 972 3748 1028
rect 3852 972 3908 1028
rect 4012 972 4068 1028
rect 4332 972 4388 1028
rect 4492 972 4548 1028
rect 4652 972 4708 1028
rect 4812 972 4868 1028
rect 4972 972 5028 1028
rect 5292 972 5348 1028
rect 5452 972 5508 1028
rect 5612 972 5668 1028
rect 5772 972 5828 1028
rect 5932 972 5988 1028
rect 6092 972 6148 1028
rect 6252 972 6308 1028
rect 6412 972 6468 1028
rect 6572 972 6628 1028
rect 6732 972 6788 1028
rect 6892 972 6948 1028
rect 7212 972 7268 1028
rect 7372 972 7428 1028
rect 7532 972 7588 1028
rect 7692 972 7748 1028
rect 7852 972 7908 1028
rect 8172 972 8228 1028
rect 332 318 388 328
rect 332 272 334 318
rect 334 272 386 318
rect 386 272 388 318
rect 332 202 334 248
rect 334 202 386 248
rect 386 202 388 248
rect 332 192 388 202
rect 8012 318 8068 328
rect 8012 272 8014 318
rect 8014 272 8066 318
rect 8066 272 8068 318
rect 8012 202 8014 248
rect 8014 202 8066 248
rect 8066 202 8068 248
rect 8012 192 8068 202
<< metal3 >>
rect 4160 5632 4240 5680
rect 4160 5568 4168 5632
rect 4232 5568 4240 5632
rect 4160 5552 4240 5568
rect 4160 5488 4168 5552
rect 4232 5488 4240 5552
rect 4160 5472 4240 5488
rect 4160 5408 4168 5472
rect 4232 5408 4240 5472
rect 4160 5392 4240 5408
rect 4160 5328 4168 5392
rect 4232 5328 4240 5392
rect 4160 5280 4240 5328
rect 0 3992 80 4000
rect 0 3928 8 3992
rect 72 3928 80 3992
rect 0 3672 80 3928
rect 0 3608 8 3672
rect 72 3608 80 3672
rect 0 3600 80 3608
rect 160 3992 240 4000
rect 160 3928 168 3992
rect 232 3928 240 3992
rect 160 3672 240 3928
rect 160 3608 168 3672
rect 232 3608 240 3672
rect 160 3600 240 3608
rect 320 3992 400 4000
rect 320 3928 328 3992
rect 392 3928 400 3992
rect 320 3672 400 3928
rect 320 3608 328 3672
rect 392 3608 400 3672
rect 320 3600 400 3608
rect 480 3992 560 4000
rect 480 3928 488 3992
rect 552 3928 560 3992
rect 480 3672 560 3928
rect 480 3608 488 3672
rect 552 3608 560 3672
rect 480 3600 560 3608
rect 640 3992 720 4000
rect 640 3928 648 3992
rect 712 3928 720 3992
rect 640 3672 720 3928
rect 640 3608 648 3672
rect 712 3608 720 3672
rect 640 3600 720 3608
rect 800 3992 880 4000
rect 800 3928 808 3992
rect 872 3928 880 3992
rect 800 3672 880 3928
rect 800 3608 808 3672
rect 872 3608 880 3672
rect 800 3600 880 3608
rect 960 3992 1040 4000
rect 960 3928 968 3992
rect 1032 3928 1040 3992
rect 960 3672 1040 3928
rect 960 3608 968 3672
rect 1032 3608 1040 3672
rect 960 3600 1040 3608
rect 1120 3992 1200 4000
rect 1120 3928 1128 3992
rect 1192 3928 1200 3992
rect 1120 3672 1200 3928
rect 1120 3608 1128 3672
rect 1192 3608 1200 3672
rect 1120 3600 1200 3608
rect 1440 3992 1520 4000
rect 1440 3928 1448 3992
rect 1512 3928 1520 3992
rect 1440 3672 1520 3928
rect 1440 3608 1448 3672
rect 1512 3608 1520 3672
rect 1440 3600 1520 3608
rect 1600 3992 1680 4000
rect 1600 3928 1608 3992
rect 1672 3928 1680 3992
rect 1600 3672 1680 3928
rect 1600 3608 1608 3672
rect 1672 3608 1680 3672
rect 1600 3600 1680 3608
rect 1760 3992 1840 4000
rect 1760 3928 1768 3992
rect 1832 3928 1840 3992
rect 1760 3672 1840 3928
rect 1760 3608 1768 3672
rect 1832 3608 1840 3672
rect 1760 3600 1840 3608
rect 1920 3992 2000 4000
rect 1920 3928 1928 3992
rect 1992 3928 2000 3992
rect 1920 3672 2000 3928
rect 1920 3608 1928 3672
rect 1992 3608 2000 3672
rect 1920 3600 2000 3608
rect 2080 3992 2160 4000
rect 2080 3928 2088 3992
rect 2152 3928 2160 3992
rect 2080 3672 2160 3928
rect 2080 3608 2088 3672
rect 2152 3608 2160 3672
rect 2080 3600 2160 3608
rect 2240 3992 2320 4000
rect 2240 3928 2248 3992
rect 2312 3928 2320 3992
rect 2240 3672 2320 3928
rect 2240 3608 2248 3672
rect 2312 3608 2320 3672
rect 2240 3600 2320 3608
rect 2400 3992 2480 4000
rect 2400 3928 2408 3992
rect 2472 3928 2480 3992
rect 2400 3672 2480 3928
rect 2400 3608 2408 3672
rect 2472 3608 2480 3672
rect 2400 3600 2480 3608
rect 2560 3992 2640 4000
rect 2560 3928 2568 3992
rect 2632 3928 2640 3992
rect 2560 3672 2640 3928
rect 2560 3608 2568 3672
rect 2632 3608 2640 3672
rect 2560 3600 2640 3608
rect 2720 3992 2800 4000
rect 2720 3928 2728 3992
rect 2792 3928 2800 3992
rect 2720 3672 2800 3928
rect 2720 3608 2728 3672
rect 2792 3608 2800 3672
rect 2720 3600 2800 3608
rect 2880 3992 2960 4000
rect 2880 3928 2888 3992
rect 2952 3928 2960 3992
rect 2880 3672 2960 3928
rect 2880 3608 2888 3672
rect 2952 3608 2960 3672
rect 2880 3600 2960 3608
rect 3040 3992 3120 4000
rect 3040 3928 3048 3992
rect 3112 3928 3120 3992
rect 3040 3672 3120 3928
rect 3040 3608 3048 3672
rect 3112 3608 3120 3672
rect 3040 3600 3120 3608
rect 3360 3992 3440 4000
rect 3360 3928 3368 3992
rect 3432 3928 3440 3992
rect 3360 3672 3440 3928
rect 3360 3608 3368 3672
rect 3432 3608 3440 3672
rect 3360 3600 3440 3608
rect 3520 3992 3600 4000
rect 3520 3928 3528 3992
rect 3592 3928 3600 3992
rect 3520 3672 3600 3928
rect 3520 3608 3528 3672
rect 3592 3608 3600 3672
rect 3520 3600 3600 3608
rect 3680 3992 3760 4000
rect 3680 3928 3688 3992
rect 3752 3928 3760 3992
rect 3680 3672 3760 3928
rect 3680 3608 3688 3672
rect 3752 3608 3760 3672
rect 3680 3600 3760 3608
rect 3840 3992 3920 4000
rect 3840 3928 3848 3992
rect 3912 3928 3920 3992
rect 3840 3672 3920 3928
rect 3840 3608 3848 3672
rect 3912 3608 3920 3672
rect 3840 3600 3920 3608
rect 4000 3992 4080 4000
rect 4000 3928 4008 3992
rect 4072 3928 4080 3992
rect 4000 3672 4080 3928
rect 4000 3608 4008 3672
rect 4072 3608 4080 3672
rect 4000 3600 4080 3608
rect 4160 3992 4240 4000
rect 4160 3928 4168 3992
rect 4232 3928 4240 3992
rect 4160 3672 4240 3928
rect 4160 3608 4168 3672
rect 4232 3608 4240 3672
rect 4160 3600 4240 3608
rect 4320 3992 4400 4000
rect 4320 3928 4328 3992
rect 4392 3928 4400 3992
rect 4320 3672 4400 3928
rect 4320 3608 4328 3672
rect 4392 3608 4400 3672
rect 4320 3600 4400 3608
rect 4480 3992 4560 4000
rect 4480 3928 4488 3992
rect 4552 3928 4560 3992
rect 4480 3672 4560 3928
rect 4480 3608 4488 3672
rect 4552 3608 4560 3672
rect 4480 3600 4560 3608
rect 4640 3992 4720 4000
rect 4640 3928 4648 3992
rect 4712 3928 4720 3992
rect 4640 3672 4720 3928
rect 4640 3608 4648 3672
rect 4712 3608 4720 3672
rect 4640 3600 4720 3608
rect 4800 3992 4880 4000
rect 4800 3928 4808 3992
rect 4872 3928 4880 3992
rect 4800 3672 4880 3928
rect 4800 3608 4808 3672
rect 4872 3608 4880 3672
rect 4800 3600 4880 3608
rect 4960 3992 5040 4000
rect 4960 3928 4968 3992
rect 5032 3928 5040 3992
rect 4960 3672 5040 3928
rect 4960 3608 4968 3672
rect 5032 3608 5040 3672
rect 4960 3600 5040 3608
rect 5280 3992 5360 4000
rect 5280 3928 5288 3992
rect 5352 3928 5360 3992
rect 5280 3672 5360 3928
rect 5280 3608 5288 3672
rect 5352 3608 5360 3672
rect 5280 3600 5360 3608
rect 5440 3992 5520 4000
rect 5440 3928 5448 3992
rect 5512 3928 5520 3992
rect 5440 3672 5520 3928
rect 5440 3608 5448 3672
rect 5512 3608 5520 3672
rect 5440 3600 5520 3608
rect 5600 3992 5680 4000
rect 5600 3928 5608 3992
rect 5672 3928 5680 3992
rect 5600 3672 5680 3928
rect 5600 3608 5608 3672
rect 5672 3608 5680 3672
rect 5600 3600 5680 3608
rect 5760 3992 5840 4000
rect 5760 3928 5768 3992
rect 5832 3928 5840 3992
rect 5760 3672 5840 3928
rect 5760 3608 5768 3672
rect 5832 3608 5840 3672
rect 5760 3600 5840 3608
rect 5920 3992 6000 4000
rect 5920 3928 5928 3992
rect 5992 3928 6000 3992
rect 5920 3672 6000 3928
rect 5920 3608 5928 3672
rect 5992 3608 6000 3672
rect 5920 3600 6000 3608
rect 6080 3992 6160 4000
rect 6080 3928 6088 3992
rect 6152 3928 6160 3992
rect 6080 3672 6160 3928
rect 6080 3608 6088 3672
rect 6152 3608 6160 3672
rect 6080 3600 6160 3608
rect 6240 3992 6320 4000
rect 6240 3928 6248 3992
rect 6312 3928 6320 3992
rect 6240 3672 6320 3928
rect 6240 3608 6248 3672
rect 6312 3608 6320 3672
rect 6240 3600 6320 3608
rect 6400 3992 6480 4000
rect 6400 3928 6408 3992
rect 6472 3928 6480 3992
rect 6400 3672 6480 3928
rect 6400 3608 6408 3672
rect 6472 3608 6480 3672
rect 6400 3600 6480 3608
rect 6560 3992 6640 4000
rect 6560 3928 6568 3992
rect 6632 3928 6640 3992
rect 6560 3672 6640 3928
rect 6560 3608 6568 3672
rect 6632 3608 6640 3672
rect 6560 3600 6640 3608
rect 6720 3992 6800 4000
rect 6720 3928 6728 3992
rect 6792 3928 6800 3992
rect 6720 3672 6800 3928
rect 6720 3608 6728 3672
rect 6792 3608 6800 3672
rect 6720 3600 6800 3608
rect 6880 3992 6960 4000
rect 6880 3928 6888 3992
rect 6952 3928 6960 3992
rect 6880 3672 6960 3928
rect 6880 3608 6888 3672
rect 6952 3608 6960 3672
rect 6880 3600 6960 3608
rect 7200 3992 7280 4000
rect 7200 3928 7208 3992
rect 7272 3928 7280 3992
rect 7200 3672 7280 3928
rect 7200 3608 7208 3672
rect 7272 3608 7280 3672
rect 7200 3600 7280 3608
rect 7360 3992 7440 4000
rect 7360 3928 7368 3992
rect 7432 3928 7440 3992
rect 7360 3672 7440 3928
rect 7360 3608 7368 3672
rect 7432 3608 7440 3672
rect 7360 3600 7440 3608
rect 7520 3992 7600 4000
rect 7520 3928 7528 3992
rect 7592 3928 7600 3992
rect 7520 3672 7600 3928
rect 7520 3608 7528 3672
rect 7592 3608 7600 3672
rect 7520 3600 7600 3608
rect 7680 3992 7760 4000
rect 7680 3928 7688 3992
rect 7752 3928 7760 3992
rect 7680 3672 7760 3928
rect 7680 3608 7688 3672
rect 7752 3608 7760 3672
rect 7680 3600 7760 3608
rect 7840 3992 7920 4000
rect 7840 3928 7848 3992
rect 7912 3928 7920 3992
rect 7840 3672 7920 3928
rect 7840 3608 7848 3672
rect 7912 3608 7920 3672
rect 7840 3600 7920 3608
rect 8000 3992 8080 4000
rect 8000 3928 8008 3992
rect 8072 3928 8080 3992
rect 8000 3672 8080 3928
rect 8000 3608 8008 3672
rect 8072 3608 8080 3672
rect 8000 3600 8080 3608
rect 8160 3992 8240 4000
rect 8160 3928 8168 3992
rect 8232 3928 8240 3992
rect 8160 3672 8240 3928
rect 8160 3608 8168 3672
rect 8232 3608 8240 3672
rect 8160 3600 8240 3608
rect 8320 3992 8400 4000
rect 8320 3928 8328 3992
rect 8392 3928 8400 3992
rect 8320 3672 8400 3928
rect 8320 3608 8328 3672
rect 8392 3608 8400 3672
rect 8320 3600 8400 3608
rect 160 1668 240 1680
rect 160 1612 172 1668
rect 228 1612 240 1668
rect 160 1352 240 1612
rect 160 1288 168 1352
rect 232 1288 240 1352
rect 160 1028 240 1288
rect 160 972 172 1028
rect 228 972 240 1028
rect 160 960 240 972
rect 480 1668 560 1680
rect 480 1612 492 1668
rect 548 1612 560 1668
rect 480 1348 560 1612
rect 480 1292 492 1348
rect 548 1292 560 1348
rect 480 1028 560 1292
rect 480 972 492 1028
rect 548 972 560 1028
rect 480 960 560 972
rect 640 1668 720 1680
rect 640 1612 652 1668
rect 708 1612 720 1668
rect 640 1348 720 1612
rect 640 1292 652 1348
rect 708 1292 720 1348
rect 640 1028 720 1292
rect 640 972 652 1028
rect 708 972 720 1028
rect 640 960 720 972
rect 800 1668 880 1680
rect 800 1612 812 1668
rect 868 1612 880 1668
rect 800 1348 880 1612
rect 800 1292 812 1348
rect 868 1292 880 1348
rect 800 1028 880 1292
rect 800 972 812 1028
rect 868 972 880 1028
rect 800 960 880 972
rect 960 1668 1040 1680
rect 960 1612 972 1668
rect 1028 1612 1040 1668
rect 960 1348 1040 1612
rect 960 1292 972 1348
rect 1028 1292 1040 1348
rect 960 1028 1040 1292
rect 960 972 972 1028
rect 1028 972 1040 1028
rect 960 960 1040 972
rect 1120 1668 1200 1680
rect 1120 1612 1132 1668
rect 1188 1612 1200 1668
rect 1120 1348 1200 1612
rect 1120 1292 1132 1348
rect 1188 1292 1200 1348
rect 1120 1028 1200 1292
rect 1120 972 1132 1028
rect 1188 972 1200 1028
rect 1120 960 1200 972
rect 1440 1668 1520 1680
rect 1440 1612 1452 1668
rect 1508 1612 1520 1668
rect 1440 1348 1520 1612
rect 1440 1292 1452 1348
rect 1508 1292 1520 1348
rect 1440 1028 1520 1292
rect 1440 972 1452 1028
rect 1508 972 1520 1028
rect 1440 960 1520 972
rect 1600 1668 1680 1680
rect 1600 1612 1612 1668
rect 1668 1612 1680 1668
rect 1600 1348 1680 1612
rect 1600 1292 1612 1348
rect 1668 1292 1680 1348
rect 1600 1028 1680 1292
rect 1600 972 1612 1028
rect 1668 972 1680 1028
rect 1600 960 1680 972
rect 1760 1668 1840 1680
rect 1760 1612 1772 1668
rect 1828 1612 1840 1668
rect 1760 1348 1840 1612
rect 1760 1292 1772 1348
rect 1828 1292 1840 1348
rect 1760 1028 1840 1292
rect 1760 972 1772 1028
rect 1828 972 1840 1028
rect 1760 960 1840 972
rect 1920 1668 2000 1680
rect 1920 1612 1932 1668
rect 1988 1612 2000 1668
rect 1920 1348 2000 1612
rect 1920 1292 1932 1348
rect 1988 1292 2000 1348
rect 1920 1028 2000 1292
rect 1920 972 1932 1028
rect 1988 972 2000 1028
rect 1920 960 2000 972
rect 2080 1668 2160 1680
rect 2080 1612 2092 1668
rect 2148 1612 2160 1668
rect 2080 1348 2160 1612
rect 2080 1292 2092 1348
rect 2148 1292 2160 1348
rect 2080 1028 2160 1292
rect 2080 972 2092 1028
rect 2148 972 2160 1028
rect 2080 960 2160 972
rect 2240 1668 2320 1680
rect 2240 1612 2252 1668
rect 2308 1612 2320 1668
rect 2240 1348 2320 1612
rect 2240 1292 2252 1348
rect 2308 1292 2320 1348
rect 2240 1028 2320 1292
rect 2240 972 2252 1028
rect 2308 972 2320 1028
rect 2240 960 2320 972
rect 2400 1668 2480 1680
rect 2400 1612 2412 1668
rect 2468 1612 2480 1668
rect 2400 1348 2480 1612
rect 2400 1292 2412 1348
rect 2468 1292 2480 1348
rect 2400 1028 2480 1292
rect 2400 972 2412 1028
rect 2468 972 2480 1028
rect 2400 960 2480 972
rect 2560 1668 2640 1680
rect 2560 1612 2572 1668
rect 2628 1612 2640 1668
rect 2560 1348 2640 1612
rect 2560 1292 2572 1348
rect 2628 1292 2640 1348
rect 2560 1028 2640 1292
rect 2560 972 2572 1028
rect 2628 972 2640 1028
rect 2560 960 2640 972
rect 2720 1668 2800 1680
rect 2720 1612 2732 1668
rect 2788 1612 2800 1668
rect 2720 1348 2800 1612
rect 2720 1292 2732 1348
rect 2788 1292 2800 1348
rect 2720 1028 2800 1292
rect 2720 972 2732 1028
rect 2788 972 2800 1028
rect 2720 960 2800 972
rect 2880 1668 2960 1680
rect 2880 1612 2892 1668
rect 2948 1612 2960 1668
rect 2880 1348 2960 1612
rect 2880 1292 2892 1348
rect 2948 1292 2960 1348
rect 2880 1028 2960 1292
rect 2880 972 2892 1028
rect 2948 972 2960 1028
rect 2880 960 2960 972
rect 3040 1668 3120 1680
rect 3040 1612 3052 1668
rect 3108 1612 3120 1668
rect 3040 1348 3120 1612
rect 3040 1292 3052 1348
rect 3108 1292 3120 1348
rect 3040 1028 3120 1292
rect 3040 972 3052 1028
rect 3108 972 3120 1028
rect 3040 960 3120 972
rect 3360 1668 3440 1680
rect 3360 1612 3372 1668
rect 3428 1612 3440 1668
rect 3360 1348 3440 1612
rect 3360 1292 3372 1348
rect 3428 1292 3440 1348
rect 3360 1028 3440 1292
rect 3360 972 3372 1028
rect 3428 972 3440 1028
rect 3360 960 3440 972
rect 3520 1668 3600 1680
rect 3520 1612 3532 1668
rect 3588 1612 3600 1668
rect 3520 1348 3600 1612
rect 3520 1292 3532 1348
rect 3588 1292 3600 1348
rect 3520 1028 3600 1292
rect 3520 972 3532 1028
rect 3588 972 3600 1028
rect 3520 960 3600 972
rect 3680 1668 3760 1680
rect 3680 1612 3692 1668
rect 3748 1612 3760 1668
rect 3680 1348 3760 1612
rect 3680 1292 3692 1348
rect 3748 1292 3760 1348
rect 3680 1028 3760 1292
rect 3680 972 3692 1028
rect 3748 972 3760 1028
rect 3680 960 3760 972
rect 3840 1668 3920 1680
rect 3840 1612 3852 1668
rect 3908 1612 3920 1668
rect 3840 1348 3920 1612
rect 3840 1292 3852 1348
rect 3908 1292 3920 1348
rect 3840 1028 3920 1292
rect 3840 972 3852 1028
rect 3908 972 3920 1028
rect 3840 960 3920 972
rect 4000 1668 4080 1680
rect 4000 1612 4012 1668
rect 4068 1612 4080 1668
rect 4000 1348 4080 1612
rect 4000 1292 4012 1348
rect 4068 1292 4080 1348
rect 4000 1028 4080 1292
rect 4000 972 4012 1028
rect 4068 972 4080 1028
rect 4000 960 4080 972
rect 4320 1668 4400 1680
rect 4320 1612 4332 1668
rect 4388 1612 4400 1668
rect 4320 1348 4400 1612
rect 4320 1292 4332 1348
rect 4388 1292 4400 1348
rect 4320 1028 4400 1292
rect 4320 972 4332 1028
rect 4388 972 4400 1028
rect 4320 960 4400 972
rect 4480 1668 4560 1680
rect 4480 1612 4492 1668
rect 4548 1612 4560 1668
rect 4480 1348 4560 1612
rect 4480 1292 4492 1348
rect 4548 1292 4560 1348
rect 4480 1028 4560 1292
rect 4480 972 4492 1028
rect 4548 972 4560 1028
rect 4480 960 4560 972
rect 4640 1668 4720 1680
rect 4640 1612 4652 1668
rect 4708 1612 4720 1668
rect 4640 1348 4720 1612
rect 4640 1292 4652 1348
rect 4708 1292 4720 1348
rect 4640 1028 4720 1292
rect 4640 972 4652 1028
rect 4708 972 4720 1028
rect 4640 960 4720 972
rect 4800 1668 4880 1680
rect 4800 1612 4812 1668
rect 4868 1612 4880 1668
rect 4800 1348 4880 1612
rect 4800 1292 4812 1348
rect 4868 1292 4880 1348
rect 4800 1028 4880 1292
rect 4800 972 4812 1028
rect 4868 972 4880 1028
rect 4800 960 4880 972
rect 4960 1668 5040 1680
rect 4960 1612 4972 1668
rect 5028 1612 5040 1668
rect 4960 1348 5040 1612
rect 4960 1292 4972 1348
rect 5028 1292 5040 1348
rect 4960 1028 5040 1292
rect 4960 972 4972 1028
rect 5028 972 5040 1028
rect 4960 960 5040 972
rect 5280 1668 5360 1680
rect 5280 1612 5292 1668
rect 5348 1612 5360 1668
rect 5280 1348 5360 1612
rect 5280 1292 5292 1348
rect 5348 1292 5360 1348
rect 5280 1028 5360 1292
rect 5280 972 5292 1028
rect 5348 972 5360 1028
rect 5280 960 5360 972
rect 5440 1668 5520 1680
rect 5440 1612 5452 1668
rect 5508 1612 5520 1668
rect 5440 1348 5520 1612
rect 5440 1292 5452 1348
rect 5508 1292 5520 1348
rect 5440 1028 5520 1292
rect 5440 972 5452 1028
rect 5508 972 5520 1028
rect 5440 960 5520 972
rect 5600 1668 5680 1680
rect 5600 1612 5612 1668
rect 5668 1612 5680 1668
rect 5600 1348 5680 1612
rect 5600 1292 5612 1348
rect 5668 1292 5680 1348
rect 5600 1028 5680 1292
rect 5600 972 5612 1028
rect 5668 972 5680 1028
rect 5600 960 5680 972
rect 5760 1668 5840 1680
rect 5760 1612 5772 1668
rect 5828 1612 5840 1668
rect 5760 1348 5840 1612
rect 5760 1292 5772 1348
rect 5828 1292 5840 1348
rect 5760 1028 5840 1292
rect 5760 972 5772 1028
rect 5828 972 5840 1028
rect 5760 960 5840 972
rect 5920 1668 6000 1680
rect 5920 1612 5932 1668
rect 5988 1612 6000 1668
rect 5920 1348 6000 1612
rect 5920 1292 5932 1348
rect 5988 1292 6000 1348
rect 5920 1028 6000 1292
rect 5920 972 5932 1028
rect 5988 972 6000 1028
rect 5920 960 6000 972
rect 6080 1668 6160 1680
rect 6080 1612 6092 1668
rect 6148 1612 6160 1668
rect 6080 1348 6160 1612
rect 6080 1292 6092 1348
rect 6148 1292 6160 1348
rect 6080 1028 6160 1292
rect 6080 972 6092 1028
rect 6148 972 6160 1028
rect 6080 960 6160 972
rect 6240 1668 6320 1680
rect 6240 1612 6252 1668
rect 6308 1612 6320 1668
rect 6240 1348 6320 1612
rect 6240 1292 6252 1348
rect 6308 1292 6320 1348
rect 6240 1028 6320 1292
rect 6240 972 6252 1028
rect 6308 972 6320 1028
rect 6240 960 6320 972
rect 6400 1668 6480 1680
rect 6400 1612 6412 1668
rect 6468 1612 6480 1668
rect 6400 1348 6480 1612
rect 6400 1292 6412 1348
rect 6468 1292 6480 1348
rect 6400 1028 6480 1292
rect 6400 972 6412 1028
rect 6468 972 6480 1028
rect 6400 960 6480 972
rect 6560 1668 6640 1680
rect 6560 1612 6572 1668
rect 6628 1612 6640 1668
rect 6560 1348 6640 1612
rect 6560 1292 6572 1348
rect 6628 1292 6640 1348
rect 6560 1028 6640 1292
rect 6560 972 6572 1028
rect 6628 972 6640 1028
rect 6560 960 6640 972
rect 6720 1668 6800 1680
rect 6720 1612 6732 1668
rect 6788 1612 6800 1668
rect 6720 1348 6800 1612
rect 6720 1292 6732 1348
rect 6788 1292 6800 1348
rect 6720 1028 6800 1292
rect 6720 972 6732 1028
rect 6788 972 6800 1028
rect 6720 960 6800 972
rect 6880 1668 6960 1680
rect 6880 1612 6892 1668
rect 6948 1612 6960 1668
rect 6880 1348 6960 1612
rect 6880 1292 6892 1348
rect 6948 1292 6960 1348
rect 6880 1028 6960 1292
rect 6880 972 6892 1028
rect 6948 972 6960 1028
rect 6880 960 6960 972
rect 7200 1668 7280 1680
rect 7200 1612 7212 1668
rect 7268 1612 7280 1668
rect 7200 1348 7280 1612
rect 7200 1292 7212 1348
rect 7268 1292 7280 1348
rect 7200 1028 7280 1292
rect 7200 972 7212 1028
rect 7268 972 7280 1028
rect 7200 960 7280 972
rect 7360 1668 7440 1680
rect 7360 1612 7372 1668
rect 7428 1612 7440 1668
rect 7360 1348 7440 1612
rect 7360 1292 7372 1348
rect 7428 1292 7440 1348
rect 7360 1028 7440 1292
rect 7360 972 7372 1028
rect 7428 972 7440 1028
rect 7360 960 7440 972
rect 7520 1668 7600 1680
rect 7520 1612 7532 1668
rect 7588 1612 7600 1668
rect 7520 1348 7600 1612
rect 7520 1292 7532 1348
rect 7588 1292 7600 1348
rect 7520 1028 7600 1292
rect 7520 972 7532 1028
rect 7588 972 7600 1028
rect 7520 960 7600 972
rect 7680 1668 7760 1680
rect 7680 1612 7692 1668
rect 7748 1612 7760 1668
rect 7680 1348 7760 1612
rect 7680 1292 7692 1348
rect 7748 1292 7760 1348
rect 7680 1028 7760 1292
rect 7680 972 7692 1028
rect 7748 972 7760 1028
rect 7680 960 7760 972
rect 7840 1668 7920 1680
rect 7840 1612 7852 1668
rect 7908 1612 7920 1668
rect 7840 1348 7920 1612
rect 7840 1292 7852 1348
rect 7908 1292 7920 1348
rect 7840 1028 7920 1292
rect 7840 972 7852 1028
rect 7908 972 7920 1028
rect 7840 960 7920 972
rect 8160 1668 8240 1680
rect 8160 1612 8172 1668
rect 8228 1612 8240 1668
rect 8160 1348 8240 1612
rect 8160 1292 8172 1348
rect 8228 1292 8240 1348
rect 8160 1028 8240 1292
rect 8160 972 8172 1028
rect 8228 972 8240 1028
rect 8160 960 8240 972
rect 320 332 400 360
rect 320 268 328 332
rect 392 268 400 332
rect 320 252 400 268
rect 320 188 328 252
rect 392 188 400 252
rect 320 160 400 188
rect 8000 332 8080 360
rect 8000 268 8008 332
rect 8072 268 8080 332
rect 8000 252 8080 268
rect 8000 188 8008 252
rect 8072 188 8080 252
rect 8000 160 8080 188
<< via3 >>
rect 4168 5628 4232 5632
rect 4168 5572 4172 5628
rect 4172 5572 4228 5628
rect 4228 5572 4232 5628
rect 4168 5568 4232 5572
rect 4168 5548 4232 5552
rect 4168 5492 4172 5548
rect 4172 5492 4228 5548
rect 4228 5492 4232 5548
rect 4168 5488 4232 5492
rect 4168 5468 4232 5472
rect 4168 5412 4172 5468
rect 4172 5412 4228 5468
rect 4228 5412 4232 5468
rect 4168 5408 4232 5412
rect 4168 5388 4232 5392
rect 4168 5332 4172 5388
rect 4172 5332 4228 5388
rect 4228 5332 4232 5388
rect 4168 5328 4232 5332
rect 8 3988 72 3992
rect 8 3932 12 3988
rect 12 3932 68 3988
rect 68 3932 72 3988
rect 8 3928 72 3932
rect 8 3668 72 3672
rect 8 3612 12 3668
rect 12 3612 68 3668
rect 68 3612 72 3668
rect 8 3608 72 3612
rect 168 3988 232 3992
rect 168 3932 172 3988
rect 172 3932 228 3988
rect 228 3932 232 3988
rect 168 3928 232 3932
rect 168 3668 232 3672
rect 168 3612 172 3668
rect 172 3612 228 3668
rect 228 3612 232 3668
rect 168 3608 232 3612
rect 328 3988 392 3992
rect 328 3932 332 3988
rect 332 3932 388 3988
rect 388 3932 392 3988
rect 328 3928 392 3932
rect 328 3668 392 3672
rect 328 3612 332 3668
rect 332 3612 388 3668
rect 388 3612 392 3668
rect 328 3608 392 3612
rect 488 3988 552 3992
rect 488 3932 492 3988
rect 492 3932 548 3988
rect 548 3932 552 3988
rect 488 3928 552 3932
rect 488 3668 552 3672
rect 488 3612 492 3668
rect 492 3612 548 3668
rect 548 3612 552 3668
rect 488 3608 552 3612
rect 648 3988 712 3992
rect 648 3932 652 3988
rect 652 3932 708 3988
rect 708 3932 712 3988
rect 648 3928 712 3932
rect 648 3668 712 3672
rect 648 3612 652 3668
rect 652 3612 708 3668
rect 708 3612 712 3668
rect 648 3608 712 3612
rect 808 3988 872 3992
rect 808 3932 812 3988
rect 812 3932 868 3988
rect 868 3932 872 3988
rect 808 3928 872 3932
rect 808 3668 872 3672
rect 808 3612 812 3668
rect 812 3612 868 3668
rect 868 3612 872 3668
rect 808 3608 872 3612
rect 968 3988 1032 3992
rect 968 3932 972 3988
rect 972 3932 1028 3988
rect 1028 3932 1032 3988
rect 968 3928 1032 3932
rect 968 3668 1032 3672
rect 968 3612 972 3668
rect 972 3612 1028 3668
rect 1028 3612 1032 3668
rect 968 3608 1032 3612
rect 1128 3988 1192 3992
rect 1128 3932 1132 3988
rect 1132 3932 1188 3988
rect 1188 3932 1192 3988
rect 1128 3928 1192 3932
rect 1128 3668 1192 3672
rect 1128 3612 1132 3668
rect 1132 3612 1188 3668
rect 1188 3612 1192 3668
rect 1128 3608 1192 3612
rect 1448 3988 1512 3992
rect 1448 3932 1452 3988
rect 1452 3932 1508 3988
rect 1508 3932 1512 3988
rect 1448 3928 1512 3932
rect 1448 3668 1512 3672
rect 1448 3612 1452 3668
rect 1452 3612 1508 3668
rect 1508 3612 1512 3668
rect 1448 3608 1512 3612
rect 1608 3988 1672 3992
rect 1608 3932 1612 3988
rect 1612 3932 1668 3988
rect 1668 3932 1672 3988
rect 1608 3928 1672 3932
rect 1608 3668 1672 3672
rect 1608 3612 1612 3668
rect 1612 3612 1668 3668
rect 1668 3612 1672 3668
rect 1608 3608 1672 3612
rect 1768 3988 1832 3992
rect 1768 3932 1772 3988
rect 1772 3932 1828 3988
rect 1828 3932 1832 3988
rect 1768 3928 1832 3932
rect 1768 3668 1832 3672
rect 1768 3612 1772 3668
rect 1772 3612 1828 3668
rect 1828 3612 1832 3668
rect 1768 3608 1832 3612
rect 1928 3988 1992 3992
rect 1928 3932 1932 3988
rect 1932 3932 1988 3988
rect 1988 3932 1992 3988
rect 1928 3928 1992 3932
rect 1928 3668 1992 3672
rect 1928 3612 1932 3668
rect 1932 3612 1988 3668
rect 1988 3612 1992 3668
rect 1928 3608 1992 3612
rect 2088 3988 2152 3992
rect 2088 3932 2092 3988
rect 2092 3932 2148 3988
rect 2148 3932 2152 3988
rect 2088 3928 2152 3932
rect 2088 3668 2152 3672
rect 2088 3612 2092 3668
rect 2092 3612 2148 3668
rect 2148 3612 2152 3668
rect 2088 3608 2152 3612
rect 2248 3988 2312 3992
rect 2248 3932 2252 3988
rect 2252 3932 2308 3988
rect 2308 3932 2312 3988
rect 2248 3928 2312 3932
rect 2248 3668 2312 3672
rect 2248 3612 2252 3668
rect 2252 3612 2308 3668
rect 2308 3612 2312 3668
rect 2248 3608 2312 3612
rect 2408 3988 2472 3992
rect 2408 3932 2412 3988
rect 2412 3932 2468 3988
rect 2468 3932 2472 3988
rect 2408 3928 2472 3932
rect 2408 3668 2472 3672
rect 2408 3612 2412 3668
rect 2412 3612 2468 3668
rect 2468 3612 2472 3668
rect 2408 3608 2472 3612
rect 2568 3988 2632 3992
rect 2568 3932 2572 3988
rect 2572 3932 2628 3988
rect 2628 3932 2632 3988
rect 2568 3928 2632 3932
rect 2568 3668 2632 3672
rect 2568 3612 2572 3668
rect 2572 3612 2628 3668
rect 2628 3612 2632 3668
rect 2568 3608 2632 3612
rect 2728 3988 2792 3992
rect 2728 3932 2732 3988
rect 2732 3932 2788 3988
rect 2788 3932 2792 3988
rect 2728 3928 2792 3932
rect 2728 3668 2792 3672
rect 2728 3612 2732 3668
rect 2732 3612 2788 3668
rect 2788 3612 2792 3668
rect 2728 3608 2792 3612
rect 2888 3988 2952 3992
rect 2888 3932 2892 3988
rect 2892 3932 2948 3988
rect 2948 3932 2952 3988
rect 2888 3928 2952 3932
rect 2888 3668 2952 3672
rect 2888 3612 2892 3668
rect 2892 3612 2948 3668
rect 2948 3612 2952 3668
rect 2888 3608 2952 3612
rect 3048 3988 3112 3992
rect 3048 3932 3052 3988
rect 3052 3932 3108 3988
rect 3108 3932 3112 3988
rect 3048 3928 3112 3932
rect 3048 3668 3112 3672
rect 3048 3612 3052 3668
rect 3052 3612 3108 3668
rect 3108 3612 3112 3668
rect 3048 3608 3112 3612
rect 3368 3988 3432 3992
rect 3368 3932 3372 3988
rect 3372 3932 3428 3988
rect 3428 3932 3432 3988
rect 3368 3928 3432 3932
rect 3368 3668 3432 3672
rect 3368 3612 3372 3668
rect 3372 3612 3428 3668
rect 3428 3612 3432 3668
rect 3368 3608 3432 3612
rect 3528 3988 3592 3992
rect 3528 3932 3532 3988
rect 3532 3932 3588 3988
rect 3588 3932 3592 3988
rect 3528 3928 3592 3932
rect 3528 3668 3592 3672
rect 3528 3612 3532 3668
rect 3532 3612 3588 3668
rect 3588 3612 3592 3668
rect 3528 3608 3592 3612
rect 3688 3988 3752 3992
rect 3688 3932 3692 3988
rect 3692 3932 3748 3988
rect 3748 3932 3752 3988
rect 3688 3928 3752 3932
rect 3688 3668 3752 3672
rect 3688 3612 3692 3668
rect 3692 3612 3748 3668
rect 3748 3612 3752 3668
rect 3688 3608 3752 3612
rect 3848 3988 3912 3992
rect 3848 3932 3852 3988
rect 3852 3932 3908 3988
rect 3908 3932 3912 3988
rect 3848 3928 3912 3932
rect 3848 3668 3912 3672
rect 3848 3612 3852 3668
rect 3852 3612 3908 3668
rect 3908 3612 3912 3668
rect 3848 3608 3912 3612
rect 4008 3988 4072 3992
rect 4008 3932 4012 3988
rect 4012 3932 4068 3988
rect 4068 3932 4072 3988
rect 4008 3928 4072 3932
rect 4008 3668 4072 3672
rect 4008 3612 4012 3668
rect 4012 3612 4068 3668
rect 4068 3612 4072 3668
rect 4008 3608 4072 3612
rect 4168 3988 4232 3992
rect 4168 3932 4172 3988
rect 4172 3932 4228 3988
rect 4228 3932 4232 3988
rect 4168 3928 4232 3932
rect 4168 3668 4232 3672
rect 4168 3612 4172 3668
rect 4172 3612 4228 3668
rect 4228 3612 4232 3668
rect 4168 3608 4232 3612
rect 4328 3988 4392 3992
rect 4328 3932 4332 3988
rect 4332 3932 4388 3988
rect 4388 3932 4392 3988
rect 4328 3928 4392 3932
rect 4328 3668 4392 3672
rect 4328 3612 4332 3668
rect 4332 3612 4388 3668
rect 4388 3612 4392 3668
rect 4328 3608 4392 3612
rect 4488 3988 4552 3992
rect 4488 3932 4492 3988
rect 4492 3932 4548 3988
rect 4548 3932 4552 3988
rect 4488 3928 4552 3932
rect 4488 3668 4552 3672
rect 4488 3612 4492 3668
rect 4492 3612 4548 3668
rect 4548 3612 4552 3668
rect 4488 3608 4552 3612
rect 4648 3988 4712 3992
rect 4648 3932 4652 3988
rect 4652 3932 4708 3988
rect 4708 3932 4712 3988
rect 4648 3928 4712 3932
rect 4648 3668 4712 3672
rect 4648 3612 4652 3668
rect 4652 3612 4708 3668
rect 4708 3612 4712 3668
rect 4648 3608 4712 3612
rect 4808 3988 4872 3992
rect 4808 3932 4812 3988
rect 4812 3932 4868 3988
rect 4868 3932 4872 3988
rect 4808 3928 4872 3932
rect 4808 3668 4872 3672
rect 4808 3612 4812 3668
rect 4812 3612 4868 3668
rect 4868 3612 4872 3668
rect 4808 3608 4872 3612
rect 4968 3988 5032 3992
rect 4968 3932 4972 3988
rect 4972 3932 5028 3988
rect 5028 3932 5032 3988
rect 4968 3928 5032 3932
rect 4968 3668 5032 3672
rect 4968 3612 4972 3668
rect 4972 3612 5028 3668
rect 5028 3612 5032 3668
rect 4968 3608 5032 3612
rect 5288 3988 5352 3992
rect 5288 3932 5292 3988
rect 5292 3932 5348 3988
rect 5348 3932 5352 3988
rect 5288 3928 5352 3932
rect 5288 3668 5352 3672
rect 5288 3612 5292 3668
rect 5292 3612 5348 3668
rect 5348 3612 5352 3668
rect 5288 3608 5352 3612
rect 5448 3988 5512 3992
rect 5448 3932 5452 3988
rect 5452 3932 5508 3988
rect 5508 3932 5512 3988
rect 5448 3928 5512 3932
rect 5448 3668 5512 3672
rect 5448 3612 5452 3668
rect 5452 3612 5508 3668
rect 5508 3612 5512 3668
rect 5448 3608 5512 3612
rect 5608 3988 5672 3992
rect 5608 3932 5612 3988
rect 5612 3932 5668 3988
rect 5668 3932 5672 3988
rect 5608 3928 5672 3932
rect 5608 3668 5672 3672
rect 5608 3612 5612 3668
rect 5612 3612 5668 3668
rect 5668 3612 5672 3668
rect 5608 3608 5672 3612
rect 5768 3988 5832 3992
rect 5768 3932 5772 3988
rect 5772 3932 5828 3988
rect 5828 3932 5832 3988
rect 5768 3928 5832 3932
rect 5768 3668 5832 3672
rect 5768 3612 5772 3668
rect 5772 3612 5828 3668
rect 5828 3612 5832 3668
rect 5768 3608 5832 3612
rect 5928 3988 5992 3992
rect 5928 3932 5932 3988
rect 5932 3932 5988 3988
rect 5988 3932 5992 3988
rect 5928 3928 5992 3932
rect 5928 3668 5992 3672
rect 5928 3612 5932 3668
rect 5932 3612 5988 3668
rect 5988 3612 5992 3668
rect 5928 3608 5992 3612
rect 6088 3988 6152 3992
rect 6088 3932 6092 3988
rect 6092 3932 6148 3988
rect 6148 3932 6152 3988
rect 6088 3928 6152 3932
rect 6088 3668 6152 3672
rect 6088 3612 6092 3668
rect 6092 3612 6148 3668
rect 6148 3612 6152 3668
rect 6088 3608 6152 3612
rect 6248 3988 6312 3992
rect 6248 3932 6252 3988
rect 6252 3932 6308 3988
rect 6308 3932 6312 3988
rect 6248 3928 6312 3932
rect 6248 3668 6312 3672
rect 6248 3612 6252 3668
rect 6252 3612 6308 3668
rect 6308 3612 6312 3668
rect 6248 3608 6312 3612
rect 6408 3988 6472 3992
rect 6408 3932 6412 3988
rect 6412 3932 6468 3988
rect 6468 3932 6472 3988
rect 6408 3928 6472 3932
rect 6408 3668 6472 3672
rect 6408 3612 6412 3668
rect 6412 3612 6468 3668
rect 6468 3612 6472 3668
rect 6408 3608 6472 3612
rect 6568 3988 6632 3992
rect 6568 3932 6572 3988
rect 6572 3932 6628 3988
rect 6628 3932 6632 3988
rect 6568 3928 6632 3932
rect 6568 3668 6632 3672
rect 6568 3612 6572 3668
rect 6572 3612 6628 3668
rect 6628 3612 6632 3668
rect 6568 3608 6632 3612
rect 6728 3988 6792 3992
rect 6728 3932 6732 3988
rect 6732 3932 6788 3988
rect 6788 3932 6792 3988
rect 6728 3928 6792 3932
rect 6728 3668 6792 3672
rect 6728 3612 6732 3668
rect 6732 3612 6788 3668
rect 6788 3612 6792 3668
rect 6728 3608 6792 3612
rect 6888 3988 6952 3992
rect 6888 3932 6892 3988
rect 6892 3932 6948 3988
rect 6948 3932 6952 3988
rect 6888 3928 6952 3932
rect 6888 3668 6952 3672
rect 6888 3612 6892 3668
rect 6892 3612 6948 3668
rect 6948 3612 6952 3668
rect 6888 3608 6952 3612
rect 7208 3988 7272 3992
rect 7208 3932 7212 3988
rect 7212 3932 7268 3988
rect 7268 3932 7272 3988
rect 7208 3928 7272 3932
rect 7208 3668 7272 3672
rect 7208 3612 7212 3668
rect 7212 3612 7268 3668
rect 7268 3612 7272 3668
rect 7208 3608 7272 3612
rect 7368 3988 7432 3992
rect 7368 3932 7372 3988
rect 7372 3932 7428 3988
rect 7428 3932 7432 3988
rect 7368 3928 7432 3932
rect 7368 3668 7432 3672
rect 7368 3612 7372 3668
rect 7372 3612 7428 3668
rect 7428 3612 7432 3668
rect 7368 3608 7432 3612
rect 7528 3988 7592 3992
rect 7528 3932 7532 3988
rect 7532 3932 7588 3988
rect 7588 3932 7592 3988
rect 7528 3928 7592 3932
rect 7528 3668 7592 3672
rect 7528 3612 7532 3668
rect 7532 3612 7588 3668
rect 7588 3612 7592 3668
rect 7528 3608 7592 3612
rect 7688 3988 7752 3992
rect 7688 3932 7692 3988
rect 7692 3932 7748 3988
rect 7748 3932 7752 3988
rect 7688 3928 7752 3932
rect 7688 3668 7752 3672
rect 7688 3612 7692 3668
rect 7692 3612 7748 3668
rect 7748 3612 7752 3668
rect 7688 3608 7752 3612
rect 7848 3988 7912 3992
rect 7848 3932 7852 3988
rect 7852 3932 7908 3988
rect 7908 3932 7912 3988
rect 7848 3928 7912 3932
rect 7848 3668 7912 3672
rect 7848 3612 7852 3668
rect 7852 3612 7908 3668
rect 7908 3612 7912 3668
rect 7848 3608 7912 3612
rect 8008 3988 8072 3992
rect 8008 3932 8012 3988
rect 8012 3932 8068 3988
rect 8068 3932 8072 3988
rect 8008 3928 8072 3932
rect 8008 3668 8072 3672
rect 8008 3612 8012 3668
rect 8012 3612 8068 3668
rect 8068 3612 8072 3668
rect 8008 3608 8072 3612
rect 8168 3988 8232 3992
rect 8168 3932 8172 3988
rect 8172 3932 8228 3988
rect 8228 3932 8232 3988
rect 8168 3928 8232 3932
rect 8168 3668 8232 3672
rect 8168 3612 8172 3668
rect 8172 3612 8228 3668
rect 8228 3612 8232 3668
rect 8168 3608 8232 3612
rect 8328 3988 8392 3992
rect 8328 3932 8332 3988
rect 8332 3932 8388 3988
rect 8388 3932 8392 3988
rect 8328 3928 8392 3932
rect 8328 3668 8392 3672
rect 8328 3612 8332 3668
rect 8332 3612 8388 3668
rect 8388 3612 8392 3668
rect 8328 3608 8392 3612
rect 168 1348 232 1352
rect 168 1292 172 1348
rect 172 1292 228 1348
rect 228 1292 232 1348
rect 168 1288 232 1292
rect 328 328 392 332
rect 328 272 332 328
rect 332 272 388 328
rect 388 272 392 328
rect 328 268 392 272
rect 328 248 392 252
rect 328 192 332 248
rect 332 192 388 248
rect 388 192 392 248
rect 328 188 392 192
rect 8008 328 8072 332
rect 8008 272 8012 328
rect 8012 272 8068 328
rect 8068 272 8072 328
rect 8008 268 8072 272
rect 8008 248 8072 252
rect 8008 192 8012 248
rect 8012 192 8068 248
rect 8068 192 8072 248
rect 8008 188 8072 192
<< metal4 >>
rect 0 5632 8400 5680
rect 0 5598 4168 5632
rect 0 5362 242 5598
rect 478 5568 4168 5598
rect 4232 5598 8400 5632
rect 4232 5568 7922 5598
rect 478 5552 7922 5568
rect 478 5488 4168 5552
rect 4232 5488 7922 5552
rect 478 5472 7922 5488
rect 478 5408 4168 5472
rect 4232 5408 7922 5472
rect 478 5392 7922 5408
rect 478 5362 4168 5392
rect 0 5328 4168 5362
rect 4232 5362 7922 5392
rect 8158 5362 8400 5598
rect 4232 5328 8400 5362
rect 0 5280 8400 5328
rect 0 3992 8400 4000
rect 0 3928 8 3992
rect 72 3928 168 3992
rect 232 3928 328 3992
rect 392 3928 488 3992
rect 552 3928 648 3992
rect 712 3928 808 3992
rect 872 3928 968 3992
rect 1032 3928 1128 3992
rect 1192 3928 1448 3992
rect 1512 3928 1608 3992
rect 1672 3928 1768 3992
rect 1832 3928 1928 3992
rect 1992 3928 2088 3992
rect 2152 3928 2248 3992
rect 2312 3928 2408 3992
rect 2472 3928 2568 3992
rect 2632 3928 2728 3992
rect 2792 3928 2888 3992
rect 2952 3928 3048 3992
rect 3112 3928 3368 3992
rect 3432 3928 3528 3992
rect 3592 3928 3688 3992
rect 3752 3928 3848 3992
rect 3912 3928 4008 3992
rect 4072 3928 4168 3992
rect 4232 3928 4328 3992
rect 4392 3928 4488 3992
rect 4552 3928 4648 3992
rect 4712 3928 4808 3992
rect 4872 3928 4968 3992
rect 5032 3928 5288 3992
rect 5352 3928 5448 3992
rect 5512 3928 5608 3992
rect 5672 3928 5768 3992
rect 5832 3928 5928 3992
rect 5992 3928 6088 3992
rect 6152 3928 6248 3992
rect 6312 3928 6408 3992
rect 6472 3928 6568 3992
rect 6632 3928 6728 3992
rect 6792 3928 6888 3992
rect 6952 3928 7208 3992
rect 7272 3928 7368 3992
rect 7432 3928 7528 3992
rect 7592 3928 7688 3992
rect 7752 3928 7848 3992
rect 7912 3928 8008 3992
rect 8072 3928 8168 3992
rect 8232 3928 8328 3992
rect 8392 3928 8400 3992
rect 0 3918 8400 3928
rect 0 3682 1202 3918
rect 1438 3682 6962 3918
rect 7198 3682 8400 3918
rect 0 3672 8400 3682
rect 0 3608 8 3672
rect 72 3608 168 3672
rect 232 3608 328 3672
rect 392 3608 488 3672
rect 552 3608 648 3672
rect 712 3608 808 3672
rect 872 3608 968 3672
rect 1032 3608 1128 3672
rect 1192 3608 1448 3672
rect 1512 3608 1608 3672
rect 1672 3608 1768 3672
rect 1832 3608 1928 3672
rect 1992 3608 2088 3672
rect 2152 3608 2248 3672
rect 2312 3608 2408 3672
rect 2472 3608 2568 3672
rect 2632 3608 2728 3672
rect 2792 3608 2888 3672
rect 2952 3608 3048 3672
rect 3112 3608 3368 3672
rect 3432 3608 3528 3672
rect 3592 3608 3688 3672
rect 3752 3608 3848 3672
rect 3912 3608 4008 3672
rect 4072 3608 4168 3672
rect 4232 3608 4328 3672
rect 4392 3608 4488 3672
rect 4552 3608 4648 3672
rect 4712 3608 4808 3672
rect 4872 3608 4968 3672
rect 5032 3608 5288 3672
rect 5352 3608 5448 3672
rect 5512 3608 5608 3672
rect 5672 3608 5768 3672
rect 5832 3608 5928 3672
rect 5992 3608 6088 3672
rect 6152 3608 6248 3672
rect 6312 3608 6408 3672
rect 6472 3608 6568 3672
rect 6632 3608 6728 3672
rect 6792 3608 6888 3672
rect 6952 3608 7208 3672
rect 7272 3608 7368 3672
rect 7432 3608 7528 3672
rect 7592 3608 7688 3672
rect 7752 3608 7848 3672
rect 7912 3608 8008 3672
rect 8072 3608 8168 3672
rect 8232 3608 8328 3672
rect 8392 3608 8400 3672
rect 0 3600 8400 3608
rect 0 1520 80 1680
rect 8320 1520 8400 1680
rect 0 1438 8400 1520
rect 0 1352 2162 1438
rect 0 1288 168 1352
rect 232 1288 2162 1352
rect 0 1202 2162 1288
rect 2398 1202 4082 1438
rect 4318 1202 6002 1438
rect 6238 1202 8400 1438
rect 0 1120 8400 1202
rect 0 332 8400 400
rect 0 268 328 332
rect 392 318 8008 332
rect 392 268 3122 318
rect 0 252 3122 268
rect 0 188 328 252
rect 392 188 3122 252
rect 0 82 3122 188
rect 3358 82 5042 318
rect 5278 268 8008 318
rect 8072 268 8400 332
rect 5278 252 8400 268
rect 5278 188 8008 252
rect 8072 188 8400 252
rect 5278 82 8400 188
rect 0 0 8400 82
<< via4 >>
rect 242 5362 478 5598
rect 7922 5362 8158 5598
rect 1202 3682 1438 3918
rect 6962 3682 7198 3918
rect 2162 1202 2398 1438
rect 4082 1202 4318 1438
rect 6002 1202 6238 1438
rect 3122 82 3358 318
rect 5042 82 5278 318
<< metal5 >>
rect 120 5598 560 6000
rect 120 5362 242 5598
rect 478 5362 560 5598
rect 120 3080 560 5362
rect 160 0 560 3080
rect 1120 3918 1520 6000
rect 1120 3682 1202 3918
rect 1438 3682 1520 3918
rect 1120 0 1520 3682
rect 2080 1438 2480 6000
rect 2080 1202 2162 1438
rect 2398 1202 2480 1438
rect 2080 0 2480 1202
rect 3040 318 3440 6000
rect 3040 82 3122 318
rect 3358 82 3440 318
rect 3040 0 3440 82
rect 4000 1438 4400 6000
rect 4000 1202 4082 1438
rect 4318 1202 4400 1438
rect 4000 0 4400 1202
rect 4960 318 5360 6000
rect 4960 82 5042 318
rect 5278 82 5360 318
rect 4960 0 5360 82
rect 5920 1438 6320 6000
rect 5920 1202 6002 1438
rect 6238 1202 6320 1438
rect 5920 0 6320 1202
rect 6880 3918 7280 6000
rect 6880 3682 6962 3918
rect 7198 3682 7280 3918
rect 6880 0 7280 3682
rect 7840 5598 8240 6000
rect 7840 5362 7922 5598
rect 8158 5362 8240 5598
rect 7840 0 8240 5362
<< labels >>
rlabel locali s 4160 4960 4240 5040 4 xpa
rlabel metal1 s 2240 160 2320 360 4 n1
rlabel metal1 s 6080 160 6160 360 4 n2
rlabel metal1 s 6080 2840 6160 3440 4 pb2
rlabel metal1 s 2240 2840 2320 3440 4 pb1
rlabel metal1 s 6080 5080 6160 5680 4 pa2
rlabel metal1 s 2240 5080 2320 5680 4 pa1
rlabel metal2 s 0 1440 8400 1520 4 in
port 1 nsew
rlabel metal2 s 0 1120 8400 1200 4 out
port 2 nsew
rlabel metal2 s 0 2720 8400 2800 4 xpb
port 3 nsew
rlabel metal2 s 0 480 8400 560 4 xn
port 4 nsew
rlabel metal5 s 160 0 560 4000 4 vdda
port 5 nsew
rlabel metal5 s 1120 0 1520 4000 4 vddx
port 6 nsew
rlabel metal2 s 0 3760 8400 3840 4 bp
port 7 nsew
rlabel metal5 s 2080 0 2480 4000 4 gnda
port 8 nsew
rlabel metal5 s 3040 0 3440 4000 4 vssa
port 9 nsew
<< end >>
