magic
tech sky130A
timestamp 1633737718
<< metal4 >>
rect 7860 8700 13380 8720
rect 7860 8580 7880 8700
rect 8000 8580 8520 8700
rect 8640 8580 9160 8700
rect 9280 8580 11960 8700
rect 12080 8580 12600 8700
rect 12720 8580 13240 8700
rect 13360 8580 13380 8700
rect 7860 8560 13380 8580
rect 7860 8380 13380 8400
rect 7860 8260 10560 8380
rect 10680 8260 13380 8380
rect 7860 8240 13380 8260
rect 7860 8060 13380 8080
rect 7860 7940 7880 8060
rect 8000 7940 8520 8060
rect 8640 7940 9160 8060
rect 9280 7940 11960 8060
rect 12080 7940 12600 8060
rect 12720 7940 13240 8060
rect 13360 7940 13380 8060
rect 7860 7920 13380 7940
rect 9460 7740 11780 7760
rect 9460 7600 10560 7740
rect 10680 7600 11780 7740
rect 9460 7580 11780 7600
rect 8820 7400 10500 7420
rect 8820 6400 8840 7400
rect 8960 6400 10500 7400
rect 8820 6380 10500 6400
rect 10540 7400 10700 7420
rect 10540 6400 10560 7400
rect 10680 6400 10700 7400
rect 10540 6380 10700 6400
rect 10740 7400 12420 7420
rect 10740 6400 12280 7400
rect 12400 6400 12420 7400
rect 10740 6380 12420 6400
rect 8820 6200 10500 6220
rect 8820 5200 8840 6200
rect 8960 5200 10500 6200
rect 8820 5180 10500 5200
rect 10540 6200 10700 6220
rect 10540 5200 10560 6200
rect 10680 5200 10700 6200
rect 10540 5180 10700 5200
rect 10740 6200 12420 6220
rect 10740 5200 12280 6200
rect 12400 5200 12420 6200
rect 10740 5180 12420 5200
rect 8820 5000 10500 5020
rect 8820 4000 8840 5000
rect 8960 4000 10500 5000
rect 8820 3980 10500 4000
rect 10540 5000 10700 5020
rect 10540 4000 10560 5000
rect 10680 4000 10700 5000
rect 10540 3980 10700 4000
rect 10740 5000 12420 5020
rect 10740 4000 12280 5000
rect 12400 4000 12420 5000
rect 10740 3980 12420 4000
rect 8820 3800 10500 3820
rect 8820 2800 8840 3800
rect 8960 2800 10500 3800
rect 8820 2780 10500 2800
rect 10540 3800 10700 3820
rect 10540 2800 10560 3800
rect 10680 2800 10700 3800
rect 10540 2780 10700 2800
rect 10740 3800 12420 3820
rect 10740 2800 12280 3800
rect 12400 2800 12420 3800
rect 10740 2780 12420 2800
rect 8820 2600 10500 2620
rect 8820 1600 8840 2600
rect 8960 1600 10500 2600
rect 8820 1580 10500 1600
rect 10540 2600 10700 2620
rect 10540 1600 10560 2600
rect 10680 1600 10700 2600
rect 10540 1580 10700 1600
rect 10740 2600 12420 2620
rect 10740 1600 12280 2600
rect 12400 1600 12420 2600
rect 10740 1580 12420 1600
rect 8180 1400 10500 1420
rect 8180 400 8200 1400
rect 8320 400 10500 1400
rect 8180 380 10500 400
rect 10540 1400 10700 1420
rect 10540 400 10560 1400
rect 10680 400 10700 1400
rect 10540 380 10700 400
rect 10740 1400 13060 1420
rect 10740 400 12920 1400
rect 13040 400 13060 1400
rect 10740 380 13060 400
rect 8820 200 10500 220
rect 8820 -800 8840 200
rect 8960 -800 10500 200
rect 8820 -820 10500 -800
rect 10540 200 10700 220
rect 10540 -800 10560 200
rect 10680 -800 10700 200
rect 10540 -820 10700 -800
rect 10740 200 12420 220
rect 10740 -800 12280 200
rect 12400 -800 12420 200
rect 10740 -820 12420 -800
rect 8820 -1000 10500 -980
rect 8820 -2000 8840 -1000
rect 8960 -2000 10500 -1000
rect 8820 -2020 10500 -2000
rect 10540 -1000 10700 -980
rect 10540 -2000 10560 -1000
rect 10680 -2000 10700 -1000
rect 10540 -2020 10700 -2000
rect 10740 -1000 12420 -980
rect 10740 -2000 12280 -1000
rect 12400 -2000 12420 -1000
rect 10740 -2020 12420 -2000
rect 8820 -2200 10500 -2180
rect 8820 -3200 8840 -2200
rect 8960 -3200 10500 -2200
rect 8820 -3220 10500 -3200
rect 10540 -2200 10700 -2180
rect 10540 -3200 10560 -2200
rect 10680 -3200 10700 -2200
rect 10540 -3220 10700 -3200
rect 10740 -2200 12420 -2180
rect 10740 -3200 12280 -2200
rect 12400 -3200 12420 -2200
rect 10740 -3220 12420 -3200
rect 8820 -3400 10500 -3380
rect 8820 -4400 8840 -3400
rect 8960 -4400 10500 -3400
rect 8820 -4420 10500 -4400
rect 10540 -3400 10700 -3380
rect 10540 -4400 10560 -3400
rect 10680 -4400 10700 -3400
rect 10540 -4420 10700 -4400
rect 10740 -3400 12420 -3380
rect 10740 -4400 12280 -3400
rect 12400 -4400 12420 -3400
rect 10740 -4420 12420 -4400
rect 8820 -4600 10500 -4580
rect 8820 -5600 8840 -4600
rect 8960 -5600 10500 -4600
rect 8820 -5620 10500 -5600
rect 10540 -4600 10700 -4580
rect 10540 -5600 10560 -4600
rect 10680 -5600 10700 -4600
rect 10540 -5620 10700 -5600
rect 10740 -4600 12420 -4580
rect 10740 -5600 12280 -4600
rect 12400 -5600 12420 -4600
rect 10740 -5620 12420 -5600
rect 9460 -5800 11780 -5780
rect 9460 -5940 10560 -5800
rect 10680 -5940 11780 -5800
rect 9460 -5960 11780 -5940
rect 7860 -6140 13380 -6120
rect 7860 -6260 7880 -6140
rect 8000 -6260 8520 -6140
rect 8640 -6260 9160 -6140
rect 9280 -6260 11960 -6140
rect 12080 -6260 12600 -6140
rect 12720 -6260 13240 -6140
rect 13360 -6260 13380 -6140
rect 7860 -6280 13380 -6260
rect 7860 -6460 13380 -6440
rect 7860 -6580 8840 -6460
rect 8960 -6580 12280 -6460
rect 12400 -6580 13380 -6460
rect 7860 -6600 13380 -6580
rect 7860 -6780 13380 -6760
rect 7860 -6900 7880 -6780
rect 8000 -6900 8520 -6780
rect 8640 -6900 9160 -6780
rect 9280 -6900 11960 -6780
rect 12080 -6900 12600 -6780
rect 12720 -6900 13240 -6780
rect 13360 -6900 13380 -6780
rect 7860 -6920 13380 -6900
rect 7860 -7100 13380 -7080
rect 7860 -7220 8200 -7100
rect 8320 -7220 12920 -7100
rect 13040 -7220 13380 -7100
rect 7860 -7240 13380 -7220
rect 7860 -7420 13380 -7400
rect 7860 -7540 7880 -7420
rect 8000 -7540 8520 -7420
rect 8640 -7540 9160 -7420
rect 9280 -7540 11960 -7420
rect 12080 -7540 12600 -7420
rect 12720 -7540 13240 -7420
rect 13360 -7540 13380 -7420
rect 7860 -7560 13380 -7540
<< via4 >>
rect 7880 8580 8000 8700
rect 8520 8580 8640 8700
rect 9160 8580 9280 8700
rect 11960 8580 12080 8700
rect 12600 8580 12720 8700
rect 13240 8580 13360 8700
rect 10560 8260 10680 8380
rect 7880 7940 8000 8060
rect 8520 7940 8640 8060
rect 9160 7940 9280 8060
rect 11960 7940 12080 8060
rect 12600 7940 12720 8060
rect 13240 7940 13360 8060
rect 10560 7600 10680 7740
rect 8840 6400 8960 7400
rect 10560 6400 10680 7400
rect 12280 6400 12400 7400
rect 8840 5200 8960 6200
rect 10560 5200 10680 6200
rect 12280 5200 12400 6200
rect 8840 4000 8960 5000
rect 10560 4000 10680 5000
rect 12280 4000 12400 5000
rect 8840 2800 8960 3800
rect 10560 2800 10680 3800
rect 12280 2800 12400 3800
rect 8840 1600 8960 2600
rect 10560 1600 10680 2600
rect 12280 1600 12400 2600
rect 8200 400 8320 1400
rect 10560 400 10680 1400
rect 12920 400 13040 1400
rect 8840 -800 8960 200
rect 10560 -800 10680 200
rect 12280 -800 12400 200
rect 8840 -2000 8960 -1000
rect 10560 -2000 10680 -1000
rect 12280 -2000 12400 -1000
rect 8840 -3200 8960 -2200
rect 10560 -3200 10680 -2200
rect 12280 -3200 12400 -2200
rect 8840 -4400 8960 -3400
rect 10560 -4400 10680 -3400
rect 12280 -4400 12400 -3400
rect 8840 -5600 8960 -4600
rect 10560 -5600 10680 -4600
rect 12280 -5600 12400 -4600
rect 10560 -5940 10680 -5800
rect 7880 -6260 8000 -6140
rect 8520 -6260 8640 -6140
rect 9160 -6260 9280 -6140
rect 11960 -6260 12080 -6140
rect 12600 -6260 12720 -6140
rect 13240 -6260 13360 -6140
rect 8840 -6580 8960 -6460
rect 12280 -6580 12400 -6460
rect 7880 -6900 8000 -6780
rect 8520 -6900 8640 -6780
rect 9160 -6900 9280 -6780
rect 11960 -6900 12080 -6780
rect 12600 -6900 12720 -6780
rect 13240 -6900 13360 -6780
rect 8200 -7220 8320 -7100
rect 12920 -7220 13040 -7100
rect 7880 -7540 8000 -7420
rect 8520 -7540 8640 -7420
rect 9160 -7540 9280 -7420
rect 11960 -7540 12080 -7420
rect 12600 -7540 12720 -7420
rect 13240 -7540 13360 -7420
<< mimcap2 >>
rect 9480 7730 10480 7740
rect 9480 7610 9490 7730
rect 10470 7610 10480 7730
rect 9480 7600 10480 7610
rect 10760 7730 11760 7740
rect 10760 7610 10770 7730
rect 11750 7610 11760 7730
rect 10760 7600 11760 7610
rect 9480 7390 10480 7400
rect 9480 6410 9490 7390
rect 10470 6410 10480 7390
rect 9480 6400 10480 6410
rect 10760 7390 11760 7400
rect 10760 6410 10770 7390
rect 11750 6410 11760 7390
rect 10760 6400 11760 6410
rect 9480 6190 10480 6200
rect 9480 5210 9490 6190
rect 10470 5210 10480 6190
rect 9480 5200 10480 5210
rect 10760 6190 11760 6200
rect 10760 5210 10770 6190
rect 11750 5210 11760 6190
rect 10760 5200 11760 5210
rect 9480 4990 10480 5000
rect 9480 4010 9490 4990
rect 10470 4010 10480 4990
rect 9480 4000 10480 4010
rect 10760 4990 11760 5000
rect 10760 4010 10770 4990
rect 11750 4010 11760 4990
rect 10760 4000 11760 4010
rect 9480 3790 10480 3800
rect 9480 2810 9490 3790
rect 10470 2810 10480 3790
rect 9480 2800 10480 2810
rect 10760 3790 11760 3800
rect 10760 2810 10770 3790
rect 11750 2810 11760 3790
rect 10760 2800 11760 2810
rect 9480 2590 10480 2600
rect 9480 1610 9490 2590
rect 10470 1610 10480 2590
rect 9480 1600 10480 1610
rect 10760 2590 11760 2600
rect 10760 1610 10770 2590
rect 11750 1610 11760 2590
rect 10760 1600 11760 1610
rect 9480 1390 10480 1400
rect 9480 410 9490 1390
rect 10470 410 10480 1390
rect 9480 400 10480 410
rect 10760 1390 11760 1400
rect 10760 410 10770 1390
rect 11750 410 11760 1390
rect 10760 400 11760 410
rect 9480 190 10480 200
rect 9480 -790 9490 190
rect 10470 -790 10480 190
rect 9480 -800 10480 -790
rect 10760 190 11760 200
rect 10760 -790 10770 190
rect 11750 -790 11760 190
rect 10760 -800 11760 -790
rect 9480 -1010 10480 -1000
rect 9480 -1990 9490 -1010
rect 10470 -1990 10480 -1010
rect 9480 -2000 10480 -1990
rect 10760 -1010 11760 -1000
rect 10760 -1990 10770 -1010
rect 11750 -1990 11760 -1010
rect 10760 -2000 11760 -1990
rect 9480 -2210 10480 -2200
rect 9480 -3190 9490 -2210
rect 10470 -3190 10480 -2210
rect 9480 -3200 10480 -3190
rect 10760 -2210 11760 -2200
rect 10760 -3190 10770 -2210
rect 11750 -3190 11760 -2210
rect 10760 -3200 11760 -3190
rect 9480 -3410 10480 -3400
rect 9480 -4390 9490 -3410
rect 10470 -4390 10480 -3410
rect 9480 -4400 10480 -4390
rect 10760 -3410 11760 -3400
rect 10760 -4390 10770 -3410
rect 11750 -4390 11760 -3410
rect 10760 -4400 11760 -4390
rect 9480 -4610 10480 -4600
rect 9480 -5590 9490 -4610
rect 10470 -5590 10480 -4610
rect 9480 -5600 10480 -5590
rect 10760 -4610 11760 -4600
rect 10760 -5590 10770 -4610
rect 11750 -5590 11760 -4610
rect 10760 -5600 11760 -5590
rect 9480 -5810 10480 -5800
rect 9480 -5930 9490 -5810
rect 10470 -5930 10480 -5810
rect 9480 -5940 10480 -5930
rect 10760 -5810 11760 -5800
rect 10760 -5930 10770 -5810
rect 11750 -5930 11760 -5810
rect 10760 -5940 11760 -5930
<< mimcap2contact >>
rect 9490 7610 10470 7730
rect 10770 7610 11750 7730
rect 9490 6410 10470 7390
rect 10770 6410 11750 7390
rect 9490 5210 10470 6190
rect 10770 5210 11750 6190
rect 9490 4010 10470 4990
rect 10770 4010 11750 4990
rect 9490 2810 10470 3790
rect 10770 2810 11750 3790
rect 9490 1610 10470 2590
rect 10770 1610 11750 2590
rect 9490 410 10470 1390
rect 10770 410 11750 1390
rect 9490 -790 10470 190
rect 10770 -790 11750 190
rect 9490 -1990 10470 -1010
rect 10770 -1990 11750 -1010
rect 9490 -3190 10470 -2210
rect 10770 -3190 11750 -2210
rect 9490 -4390 10470 -3410
rect 10770 -4390 11750 -3410
rect 9490 -5590 10470 -4610
rect 10770 -5590 11750 -4610
rect 9490 -5930 10470 -5810
rect 10770 -5930 11750 -5810
<< metal5 >>
rect 7860 8700 8020 8720
rect 7860 8580 7880 8700
rect 8000 8580 8020 8700
rect 7860 8060 8020 8580
rect 7860 7940 7880 8060
rect 8000 7940 8020 8060
rect 7860 -6140 8020 7940
rect 8500 8700 8660 8720
rect 8500 8580 8520 8700
rect 8640 8580 8660 8700
rect 8500 8060 8660 8580
rect 8500 7940 8520 8060
rect 8640 7940 8660 8060
rect 7860 -6260 7880 -6140
rect 8000 -6260 8020 -6140
rect 7860 -6780 8020 -6260
rect 7860 -6900 7880 -6780
rect 8000 -6900 8020 -6780
rect 7860 -7420 8020 -6900
rect 7860 -7540 7880 -7420
rect 8000 -7540 8020 -7420
rect 7860 -7560 8020 -7540
rect 8180 1400 8340 7920
rect 8180 400 8200 1400
rect 8320 400 8340 1400
rect 8180 -7100 8340 400
rect 8180 -7220 8200 -7100
rect 8320 -7220 8340 -7100
rect 8180 -7560 8340 -7220
rect 8500 -6140 8660 7940
rect 9140 8700 9300 8720
rect 9140 8580 9160 8700
rect 9280 8580 9300 8700
rect 9140 8060 9300 8580
rect 9140 7940 9160 8060
rect 9280 7940 9300 8060
rect 8500 -6260 8520 -6140
rect 8640 -6260 8660 -6140
rect 8500 -6780 8660 -6260
rect 8500 -6900 8520 -6780
rect 8640 -6900 8660 -6780
rect 8500 -7420 8660 -6900
rect 8500 -7540 8520 -7420
rect 8640 -7540 8660 -7420
rect 8500 -7560 8660 -7540
rect 8820 7400 8980 7920
rect 8820 6400 8840 7400
rect 8960 6400 8980 7400
rect 8820 6200 8980 6400
rect 8820 5200 8840 6200
rect 8960 5200 8980 6200
rect 8820 5000 8980 5200
rect 8820 4000 8840 5000
rect 8960 4000 8980 5000
rect 8820 3800 8980 4000
rect 8820 2800 8840 3800
rect 8960 2800 8980 3800
rect 8820 2600 8980 2800
rect 8820 1600 8840 2600
rect 8960 1600 8980 2600
rect 8820 200 8980 1600
rect 8820 -800 8840 200
rect 8960 -800 8980 200
rect 8820 -1000 8980 -800
rect 8820 -2000 8840 -1000
rect 8960 -2000 8980 -1000
rect 8820 -2200 8980 -2000
rect 8820 -3200 8840 -2200
rect 8960 -3200 8980 -2200
rect 8820 -3400 8980 -3200
rect 8820 -4400 8840 -3400
rect 8960 -4400 8980 -3400
rect 8820 -4600 8980 -4400
rect 8820 -5600 8840 -4600
rect 8960 -5600 8980 -4600
rect 8820 -6460 8980 -5600
rect 8820 -6580 8840 -6460
rect 8960 -6580 8980 -6460
rect 8820 -7560 8980 -6580
rect 9140 -6140 9300 7940
rect 10540 8380 10700 8720
rect 10540 8260 10560 8380
rect 10680 8260 10700 8380
rect 10540 7760 10700 8260
rect 11940 8700 12100 8720
rect 11940 8580 11960 8700
rect 12080 8580 12100 8700
rect 11940 8060 12100 8580
rect 11940 7940 11960 8060
rect 12080 7940 12100 8060
rect 9460 7740 11780 7760
rect 9460 7730 10560 7740
rect 9460 7610 9490 7730
rect 10470 7610 10560 7730
rect 9460 7600 10560 7610
rect 10680 7730 11780 7740
rect 10680 7610 10770 7730
rect 11750 7610 11780 7730
rect 10680 7600 11780 7610
rect 9460 7580 11780 7600
rect 10540 7420 10700 7580
rect 9460 7400 11780 7420
rect 9460 7390 10560 7400
rect 9460 6410 9490 7390
rect 10470 6410 10560 7390
rect 9460 6400 10560 6410
rect 10680 7390 11780 7400
rect 10680 6410 10770 7390
rect 11750 6410 11780 7390
rect 10680 6400 11780 6410
rect 9460 6380 11780 6400
rect 10540 6220 10700 6380
rect 9460 6200 11780 6220
rect 9460 6190 10560 6200
rect 9460 5210 9490 6190
rect 10470 5210 10560 6190
rect 9460 5200 10560 5210
rect 10680 6190 11780 6200
rect 10680 5210 10770 6190
rect 11750 5210 11780 6190
rect 10680 5200 11780 5210
rect 9460 5180 11780 5200
rect 10540 5020 10700 5180
rect 9460 5000 11780 5020
rect 9460 4990 10560 5000
rect 9460 4010 9490 4990
rect 10470 4010 10560 4990
rect 9460 4000 10560 4010
rect 10680 4990 11780 5000
rect 10680 4010 10770 4990
rect 11750 4010 11780 4990
rect 10680 4000 11780 4010
rect 9460 3980 11780 4000
rect 10540 3820 10700 3980
rect 9460 3800 11780 3820
rect 9460 3790 10560 3800
rect 9460 2810 9490 3790
rect 10470 2810 10560 3790
rect 9460 2800 10560 2810
rect 10680 3790 11780 3800
rect 10680 2810 10770 3790
rect 11750 2810 11780 3790
rect 10680 2800 11780 2810
rect 9460 2780 11780 2800
rect 10540 2620 10700 2780
rect 9460 2600 11780 2620
rect 9460 2590 10560 2600
rect 9460 1610 9490 2590
rect 10470 1610 10560 2590
rect 9460 1600 10560 1610
rect 10680 2590 11780 2600
rect 10680 1610 10770 2590
rect 11750 1610 11780 2590
rect 10680 1600 11780 1610
rect 9460 1580 11780 1600
rect 10540 1420 10700 1580
rect 9460 1400 11780 1420
rect 9460 1390 10560 1400
rect 9460 410 9490 1390
rect 10470 410 10560 1390
rect 9460 400 10560 410
rect 10680 1390 11780 1400
rect 10680 410 10770 1390
rect 11750 410 11780 1390
rect 10680 400 11780 410
rect 9460 380 11780 400
rect 10540 220 10700 380
rect 9460 200 11780 220
rect 9460 190 10560 200
rect 9460 -790 9490 190
rect 10470 -790 10560 190
rect 9460 -800 10560 -790
rect 10680 190 11780 200
rect 10680 -790 10770 190
rect 11750 -790 11780 190
rect 10680 -800 11780 -790
rect 9460 -820 11780 -800
rect 10540 -980 10700 -820
rect 9460 -1000 11780 -980
rect 9460 -1010 10560 -1000
rect 9460 -1990 9490 -1010
rect 10470 -1990 10560 -1010
rect 9460 -2000 10560 -1990
rect 10680 -1010 11780 -1000
rect 10680 -1990 10770 -1010
rect 11750 -1990 11780 -1010
rect 10680 -2000 11780 -1990
rect 9460 -2020 11780 -2000
rect 10540 -2180 10700 -2020
rect 9460 -2200 11780 -2180
rect 9460 -2210 10560 -2200
rect 9460 -3190 9490 -2210
rect 10470 -3190 10560 -2210
rect 9460 -3200 10560 -3190
rect 10680 -2210 11780 -2200
rect 10680 -3190 10770 -2210
rect 11750 -3190 11780 -2210
rect 10680 -3200 11780 -3190
rect 9460 -3220 11780 -3200
rect 10540 -3380 10700 -3220
rect 9460 -3400 11780 -3380
rect 9460 -3410 10560 -3400
rect 9460 -4390 9490 -3410
rect 10470 -4390 10560 -3410
rect 9460 -4400 10560 -4390
rect 10680 -3410 11780 -3400
rect 10680 -4390 10770 -3410
rect 11750 -4390 11780 -3410
rect 10680 -4400 11780 -4390
rect 9460 -4420 11780 -4400
rect 10540 -4580 10700 -4420
rect 9460 -4600 11780 -4580
rect 9460 -4610 10560 -4600
rect 9460 -5590 9490 -4610
rect 10470 -5590 10560 -4610
rect 9460 -5600 10560 -5590
rect 10680 -4610 11780 -4600
rect 10680 -5590 10770 -4610
rect 11750 -5590 11780 -4610
rect 10680 -5600 11780 -5590
rect 9460 -5620 11780 -5600
rect 10540 -5780 10700 -5620
rect 9460 -5800 11780 -5780
rect 9460 -5810 10560 -5800
rect 9460 -5930 9490 -5810
rect 10470 -5930 10560 -5810
rect 9460 -5940 10560 -5930
rect 10680 -5810 11780 -5800
rect 10680 -5930 10770 -5810
rect 11750 -5930 11780 -5810
rect 10680 -5940 11780 -5930
rect 9460 -5960 11780 -5940
rect 9140 -6260 9160 -6140
rect 9280 -6260 9300 -6140
rect 9140 -6780 9300 -6260
rect 9140 -6900 9160 -6780
rect 9280 -6900 9300 -6780
rect 9140 -7420 9300 -6900
rect 9140 -7540 9160 -7420
rect 9280 -7540 9300 -7420
rect 9140 -7560 9300 -7540
rect 10540 -7560 10700 -5960
rect 11940 -6140 12100 7940
rect 12580 8700 12740 8720
rect 12580 8580 12600 8700
rect 12720 8580 12740 8700
rect 12580 8060 12740 8580
rect 12580 7940 12600 8060
rect 12720 7940 12740 8060
rect 11940 -6260 11960 -6140
rect 12080 -6260 12100 -6140
rect 11940 -6780 12100 -6260
rect 11940 -6900 11960 -6780
rect 12080 -6900 12100 -6780
rect 11940 -7420 12100 -6900
rect 11940 -7540 11960 -7420
rect 12080 -7540 12100 -7420
rect 11940 -7560 12100 -7540
rect 12260 7400 12420 7920
rect 12260 6400 12280 7400
rect 12400 6400 12420 7400
rect 12260 6200 12420 6400
rect 12260 5200 12280 6200
rect 12400 5200 12420 6200
rect 12260 5000 12420 5200
rect 12260 4000 12280 5000
rect 12400 4000 12420 5000
rect 12260 3800 12420 4000
rect 12260 2800 12280 3800
rect 12400 2800 12420 3800
rect 12260 2600 12420 2800
rect 12260 1600 12280 2600
rect 12400 1600 12420 2600
rect 12260 200 12420 1600
rect 12260 -800 12280 200
rect 12400 -800 12420 200
rect 12260 -1000 12420 -800
rect 12260 -2000 12280 -1000
rect 12400 -2000 12420 -1000
rect 12260 -2200 12420 -2000
rect 12260 -3200 12280 -2200
rect 12400 -3200 12420 -2200
rect 12260 -3400 12420 -3200
rect 12260 -4400 12280 -3400
rect 12400 -4400 12420 -3400
rect 12260 -4600 12420 -4400
rect 12260 -5600 12280 -4600
rect 12400 -5600 12420 -4600
rect 12260 -6460 12420 -5600
rect 12260 -6580 12280 -6460
rect 12400 -6580 12420 -6460
rect 12260 -7560 12420 -6580
rect 12580 -6140 12740 7940
rect 13220 8700 13380 8720
rect 13220 8580 13240 8700
rect 13360 8580 13380 8700
rect 13220 8060 13380 8580
rect 13220 7940 13240 8060
rect 13360 7940 13380 8060
rect 12580 -6260 12600 -6140
rect 12720 -6260 12740 -6140
rect 12580 -6780 12740 -6260
rect 12580 -6900 12600 -6780
rect 12720 -6900 12740 -6780
rect 12580 -7420 12740 -6900
rect 12580 -7540 12600 -7420
rect 12720 -7540 12740 -7420
rect 12580 -7560 12740 -7540
rect 12900 1400 13060 7920
rect 12900 400 12920 1400
rect 13040 400 13060 1400
rect 12900 -7100 13060 400
rect 12900 -7220 12920 -7100
rect 13040 -7220 13060 -7100
rect 12900 -7560 13060 -7220
rect 13220 -6140 13380 7940
rect 13220 -6260 13240 -6140
rect 13360 -6260 13380 -6140
rect 13220 -6780 13380 -6260
rect 13220 -6900 13240 -6780
rect 13360 -6900 13380 -6780
rect 13220 -7420 13380 -6900
rect 13220 -7540 13240 -7420
rect 13360 -7540 13380 -7420
rect 13220 -7560 13380 -7540
<< labels >>
rlabel metal5 12260 -7560 12420 -7400 1 B
port 2 n
rlabel metal5 12900 -7560 13060 -7400 1 C
port 3 n
rlabel metal5 13220 -7560 13380 -7400 1 gnd
port 4 n
rlabel metal5 10540 8560 10700 8720 1 A
port 1 n
<< end >>
