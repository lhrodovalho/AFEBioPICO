* NGSPICE file created from vga_ota.ext - technology: sky130A

.subckt p1_8 D G S B SUB
X0 x4 G x3 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X1 S G x1 B sky130_fd_pr__pfet_01v8_lvt ad=1.5e+12p pd=7e+06u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X2 x6 G x5 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X3 x2 G x1 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=0p ps=0u w=3e+06u l=8e+06u
X4 x6 G x7 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X5 x2 G x3 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X6 x4 G x5 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X7 D G x7 B sky130_fd_pr__pfet_01v8_lvt ad=1.5e+12p pd=7e+06u as=0p ps=0u w=3e+06u l=8e+06u
.ends

.subckt n1_8 D G S B
X0 a_6000_6800# G S B sky130_fd_pr__nfet_01v8_lvt ad=1e+12p pd=6e+06u as=5e+11p ps=3e+06u w=1e+06u l=8e+06u
X1 a_6000_7320# G a_5150_7190# B sky130_fd_pr__nfet_01v8_lvt ad=1e+12p pd=6e+06u as=1e+12p ps=6e+06u w=1e+06u l=8e+06u
X2 a_6000_7060# G a_5150_6930# B sky130_fd_pr__nfet_01v8_lvt ad=1e+12p pd=6e+06u as=1e+12p ps=6e+06u w=1e+06u l=8e+06u
X3 a_6000_6800# G a_5150_6930# B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X4 a_6000_7580# G D B sky130_fd_pr__nfet_01v8_lvt ad=1e+12p pd=6e+06u as=5e+11p ps=3e+06u w=1e+06u l=8e+06u
X5 a_6000_7320# G a_5150_7450# B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1e+12p ps=6e+06u w=1e+06u l=8e+06u
X6 a_6000_7060# G a_5150_7190# B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X7 a_6000_7580# G a_5150_7450# B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
.ends

.subckt vga_ota inm inp out ibias vdda gnd
Xp1_8_53 vdda ibias vdda vdda gnd p1_8
Xp1_8_42 ibias ibias a vdda gnd p1_8
Xp1_8_64 out z vdda vdda gnd p1_8
Xp1_8_31 ym inp x vdda gnd p1_8
Xp1_8_20 ibias ibias a vdda gnd p1_8
Xp1_8_5 ym inp x vdda gnd p1_8
Xp1_8_43 vdda ibias a vdda gnd p1_8
Xp1_8_21 vdda ibias a vdda gnd p1_8
Xp1_8_54 vdda z vdda vdda gnd p1_8
Xp1_8_65 out z vdda vdda gnd p1_8
Xp1_8_32 x ibias vdda vdda gnd p1_8
Xp1_8_10 vdda ibias a vdda gnd p1_8
Xn1_8_30 z yp gnd gnd n1_8
Xp1_8_22 vdda ibias a vdda gnd p1_8
Xp1_8_6 ym inp x vdda gnd p1_8
Xp1_8_33 x ibias vdda vdda gnd p1_8
Xp1_8_11 ibias ibias a vdda gnd p1_8
Xp1_8_44 vdda ibias a vdda gnd p1_8
Xp1_8_55 z z vdda vdda gnd p1_8
Xp1_8_66 z z vdda vdda gnd p1_8
Xn1_8_20 out ym gnd gnd n1_8
Xn1_8_31 out ym gnd gnd n1_8
Xp1_8_7 yp inm x vdda gnd p1_8
Xp1_8_45 ibias ibias a vdda gnd p1_8
Xp1_8_23 ibias ibias a vdda gnd p1_8
Xp1_8_56 out z vdda vdda gnd p1_8
Xp1_8_67 out z vdda vdda gnd p1_8
Xp1_8_12 yp inm x vdda gnd p1_8
Xp1_8_34 x ibias vdda vdda gnd p1_8
Xn1_8_32 z yp gnd gnd n1_8
Xn1_8_10 ym ym gnd gnd n1_8
Xn1_8_21 z yp gnd gnd n1_8
Xp1_8_8 x ibias vdda vdda gnd p1_8
Xp1_8_46 ibias ibias a vdda gnd p1_8
Xp1_8_68 z z vdda vdda gnd p1_8
Xp1_8_57 z z vdda vdda gnd p1_8
Xp1_8_13 ym inp x vdda gnd p1_8
Xp1_8_24 yp inm x vdda gnd p1_8
Xp1_8_35 x ibias vdda vdda gnd p1_8
Xn1_8_33 z yp gnd gnd n1_8
Xn1_8_11 yp yp gnd gnd n1_8
Xn1_8_22 out ym gnd gnd n1_8
Xp1_8_9 x ibias vdda vdda gnd p1_8
Xp1_8_47 ibias ibias a vdda gnd p1_8
Xp1_8_69 z z vdda vdda gnd p1_8
Xp1_8_58 out z vdda vdda gnd p1_8
Xp1_8_14 yp inm x vdda gnd p1_8
Xp1_8_25 yp inm x vdda gnd p1_8
Xp1_8_36 x ibias vdda vdda gnd p1_8
Xn1_8_34 out ym gnd gnd n1_8
Xn1_8_12 yp yp gnd gnd n1_8
Xn1_8_23 out ym gnd gnd n1_8
Xp1_8_59 out z vdda vdda gnd p1_8
Xp1_8_48 vdda ibias vdda vdda gnd p1_8
Xp1_8_15 ym inp x vdda gnd p1_8
Xp1_8_26 ym inp x vdda gnd p1_8
Xp1_8_37 x ibias vdda vdda gnd p1_8
Xn1_8_35 out ym gnd gnd n1_8
Xn1_8_13 ym ym gnd gnd n1_8
Xn1_8_24 z yp gnd gnd n1_8
Xp1_8_27 yp inm x vdda gnd p1_8
Xp1_8_49 vdda ibias vdda vdda gnd p1_8
Xp1_8_16 x ibias vdda vdda gnd p1_8
Xp1_8_38 x ibias vdda vdda gnd p1_8
Xn1_8_14 ym ym gnd gnd n1_8
Xn1_8_25 gnd ym gnd gnd n1_8
Xp1_8_28 yp inm x vdda gnd p1_8
Xp1_8_17 x ibias vdda vdda gnd p1_8
Xp1_8_39 x ibias vdda vdda gnd p1_8
Xn1_8_26 z yp gnd gnd n1_8
Xn1_8_15 ym ym gnd gnd n1_8
Xp1_8_29 ym inp x vdda gnd p1_8
Xp1_8_18 x ibias vdda vdda gnd p1_8
Xn1_8_16 gnd yp gnd gnd n1_8
Xn1_8_27 z yp gnd gnd n1_8
Xp1_8_19 x ibias vdda vdda gnd p1_8
Xn1_8_28 out ym gnd gnd n1_8
Xn1_8_17 gnd ym gnd gnd n1_8
Xn1_8_18 gnd yp gnd gnd n1_8
Xn1_8_29 out ym gnd gnd n1_8
Xn1_8_19 z yp gnd gnd n1_8
Xn1_8_0 ym yp gnd gnd n1_8
Xn1_8_1 yp yp gnd gnd n1_8
Xn1_8_2 ym ym gnd gnd n1_8
Xn1_8_3 yp yp gnd gnd n1_8
Xn1_8_4 yp yp gnd gnd n1_8
Xn1_8_5 ym ym gnd gnd n1_8
Xn1_8_6 yp yp gnd gnd n1_8
Xn1_8_7 ym ym gnd gnd n1_8
Xn1_8_8 yp yp gnd gnd n1_8
Xn1_8_9 yp yp gnd gnd n1_8
Xp1_8_70 out z vdda vdda gnd p1_8
Xp1_8_0 ibias ibias a vdda gnd p1_8
Xp1_8_71 out z vdda vdda gnd p1_8
Xp1_8_60 z z vdda vdda gnd p1_8
Xp1_8_1 vdda ibias a vdda gnd p1_8
Xp1_8_61 vdda vdda vdda vdda gnd p1_8
Xp1_8_50 vdda ibias vdda vdda gnd p1_8
Xp1_8_2 x ibias vdda vdda gnd p1_8
Xp1_8_40 vdda ibias a vdda gnd p1_8
Xp1_8_62 z z vdda vdda gnd p1_8
Xp1_8_51 vdda ibias vdda vdda gnd p1_8
Xp1_8_3 x ibias vdda vdda gnd p1_8
Xp1_8_41 vdda ibias a vdda gnd p1_8
Xp1_8_63 z z vdda vdda gnd p1_8
Xp1_8_30 ym inp x vdda gnd p1_8
Xp1_8_52 vdda ibias vdda vdda gnd p1_8
Xp1_8_4 yp inm x vdda gnd p1_8
.ends

