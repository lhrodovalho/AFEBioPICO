* symmetrical single-ended OTA open-loop testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "sym.spice"

vdda vdda 0 1.8
vssa vssa 0 0.0
egnda gnda vssa vdda vssa 0.5

vin in gnda dc 0 ac 1 SINE(0 0.4 0.5k 0 0 0)

* DUT
Xdut gnda in out ib vdda vssa sym 
IB ib vss 5n
CL out gnda 1p

.save v(in) v(out) v(ib) i(vdd)
.nodeset v(ib) 1.4
*.option gmin=1e-12
.option scale=1e-6
.control

	op
	print ib i(vdda)

	dc vin -10m 10m 100u
	wrdata sym_open_dc.txt v(in) v(out)
	plot v(in) v(out)

    
.endc

.end
