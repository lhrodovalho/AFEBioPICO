* NGSPICE file created from cap1_10.ext - technology: sky130A

.subckt cap1_10_core a b1 b2 c1 c2 gnda vssa
X0 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X5 a b2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X6 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X7 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X8 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1.2e+06u
X9 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X10 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X11 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X12 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X13 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X14 a b1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X15 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1.2e+06u
X16 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X17 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X18 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X19 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X20 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X21 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X22 a c1 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X23 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1.2e+06u
X24 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1.2e+06u
X25 a c2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt cap1_10_dummy gnda vssa
X0 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X1 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X2 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X3 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X4 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X5 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1.2e+06u
X6 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X7 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X8 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X9 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X10 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
X11 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1.2e+06u
X12 gnda gnda sky130_fd_pr__cap_mim_m3_1 l=1.2e+06u w=1e+07u
.ends

.subckt cap1_10 ip xp om im xm op gnda vssa
Xp1 xp om om ip ip gnda vssa cap1_10_core
Xp2 xp om om ip ip gnda vssa cap1_10_core
Xm1 xm op op im im gnda vssa cap1_10_core
Xm2 xm op op im im gnda vssa cap1_10_core
Xdummy1 gnda vssa cap1_10_dummy
Xdummy2 gnda vssa cap1_10_dummy
.ends

