magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< error_s >>
rect 8 31440 8392 31512
rect 8 31360 80 31440
rect 94 31400 8306 31426
rect 94 30280 120 31400
rect 160 31334 8240 31360
rect 160 30392 232 31334
rect 8214 30392 8240 31334
rect 160 30320 8240 30392
rect 8280 30280 8306 31400
rect 8320 30320 8392 31440
rect 12488 31440 20872 31512
rect 12488 31360 12560 31440
rect 12574 31400 20786 31426
rect 94 30254 8306 30280
rect 12574 30280 12600 31400
rect 12640 31334 20720 31360
rect 12640 30392 12712 31334
rect 20694 30392 20720 31334
rect 12640 30320 20720 30392
rect 20760 30280 20786 31400
rect 20800 30320 20872 31440
rect 12574 30254 20786 30280
rect 8 30000 8392 30072
rect 8 29920 80 30000
rect 94 29960 8306 29986
rect 94 28840 120 29960
rect 160 29894 8240 29920
rect 160 28952 232 29894
rect 8214 28952 8240 29894
rect 160 28880 8240 28952
rect 8280 28840 8306 29960
rect 8320 28880 8392 30000
rect 12488 30000 20872 30072
rect 12488 29920 12560 30000
rect 12574 29960 20786 29986
rect 94 28814 8306 28840
rect 12574 28840 12600 29960
rect 12640 29894 20720 29920
rect 12640 28952 12712 29894
rect 20694 28952 20720 29894
rect 12640 28880 20720 28952
rect 20760 28840 20786 29960
rect 20800 28880 20872 30000
rect 12574 28814 20786 28840
rect 8 26160 8392 26232
rect 8 26080 80 26160
rect 94 26120 8306 26146
rect 94 25000 120 26120
rect 160 26054 8240 26080
rect 160 25112 232 26054
rect 8214 25112 8240 26054
rect 160 25040 8240 25112
rect 8280 25000 8306 26120
rect 8320 25040 8392 26160
rect 12488 26160 20872 26232
rect 12488 26080 12560 26160
rect 12574 26120 20786 26146
rect 94 24974 8306 25000
rect 12574 25000 12600 26120
rect 12640 26054 20720 26080
rect 12640 25112 12712 26054
rect 20694 25112 20720 26054
rect 12640 25040 20720 25112
rect 20760 25000 20786 26120
rect 20800 25040 20872 26160
rect 12574 24974 20786 25000
rect 8 24720 8392 24792
rect 8 24640 80 24720
rect 94 24680 8306 24706
rect 94 23560 120 24680
rect 160 24614 8240 24640
rect 160 23672 232 24614
rect 8214 23672 8240 24614
rect 160 23600 8240 23672
rect 8280 23560 8306 24680
rect 8320 23600 8392 24720
rect 12488 24720 20872 24792
rect 12488 24640 12560 24720
rect 12574 24680 20786 24706
rect 94 23534 8306 23560
rect 12574 23560 12600 24680
rect 12640 24614 20720 24640
rect 12640 23672 12712 24614
rect 20694 23672 20720 24614
rect 12640 23600 20720 23672
rect 20760 23560 20786 24680
rect 20800 23600 20872 24720
rect 12574 23534 20786 23560
rect 8 23280 8392 23352
rect 8 23200 80 23280
rect 94 23240 8306 23266
rect 94 22120 120 23240
rect 160 23174 8240 23200
rect 160 22232 232 23174
rect 8214 22232 8240 23174
rect 160 22160 8240 22232
rect 8280 22120 8306 23240
rect 8320 22160 8392 23280
rect 12488 23280 20872 23352
rect 12488 23200 12560 23280
rect 12574 23240 20786 23266
rect 94 22094 8306 22120
rect 12574 22120 12600 23240
rect 12640 23174 20720 23200
rect 12640 22232 12712 23174
rect 20694 22232 20720 23174
rect 12640 22160 20720 22232
rect 20760 22120 20786 23240
rect 20800 22160 20872 23280
rect 12574 22094 20786 22120
rect 8 21840 8392 21912
rect 8 21760 80 21840
rect 94 21800 8306 21826
rect 94 20680 120 21800
rect 160 21734 8240 21760
rect 160 20792 232 21734
rect 8214 20792 8240 21734
rect 160 20720 8240 20792
rect 8280 20680 8306 21800
rect 8320 20720 8392 21840
rect 12488 21840 20872 21912
rect 12488 21760 12560 21840
rect 12574 21800 20786 21826
rect 94 20654 8306 20680
rect 12574 20680 12600 21800
rect 12640 21734 20720 21760
rect 12640 20792 12712 21734
rect 20694 20792 20720 21734
rect 12640 20720 20720 20792
rect 20760 20680 20786 21800
rect 20800 20720 20872 21840
rect 12574 20654 20786 20680
rect 8 18000 8392 18072
rect 8 17920 80 18000
rect 94 17960 8306 17986
rect 94 16840 120 17960
rect 160 17894 8240 17920
rect 160 16952 232 17894
rect 8214 16952 8240 17894
rect 160 16880 8240 16952
rect 8280 16840 8306 17960
rect 8320 16880 8392 18000
rect 12488 18000 20872 18072
rect 12488 17920 12560 18000
rect 12574 17960 20786 17986
rect 94 16814 8306 16840
rect 12574 16840 12600 17960
rect 12640 17894 20720 17920
rect 12640 16952 12712 17894
rect 20694 16952 20720 17894
rect 12640 16880 20720 16952
rect 20760 16840 20786 17960
rect 20800 16880 20872 18000
rect 12574 16814 20786 16840
rect 8 16560 8392 16632
rect 8 16480 80 16560
rect 94 16520 8306 16546
rect 94 15400 120 16520
rect 160 16454 8240 16480
rect 160 15512 232 16454
rect 8214 15512 8240 16454
rect 160 15440 8240 15512
rect 8280 15400 8306 16520
rect 8320 15440 8392 16560
rect 12488 16560 20872 16632
rect 12488 16480 12560 16560
rect 12574 16520 20786 16546
rect 94 15374 8306 15400
rect 12574 15400 12600 16520
rect 12640 16454 20720 16480
rect 12640 15512 12712 16454
rect 20694 15512 20720 16454
rect 12640 15440 20720 15512
rect 20760 15400 20786 16520
rect 20800 15440 20872 16560
rect 12574 15374 20786 15400
rect 8 15120 8392 15192
rect 8 15040 80 15120
rect 94 15080 8306 15106
rect 94 13960 120 15080
rect 160 15014 8240 15040
rect 160 14072 232 15014
rect 8214 14072 8240 15014
rect 160 14000 8240 14072
rect 8280 13960 8306 15080
rect 8320 14000 8392 15120
rect 12488 15120 20872 15192
rect 12488 15040 12560 15120
rect 12574 15080 20786 15106
rect 94 13934 8306 13960
rect 12574 13960 12600 15080
rect 12640 15014 20720 15040
rect 12640 14072 12712 15014
rect 20694 14072 20720 15014
rect 12640 14000 20720 14072
rect 20760 13960 20786 15080
rect 20800 14000 20872 15120
rect 12574 13934 20786 13960
rect 8 13680 8392 13752
rect 8 13600 80 13680
rect 94 13640 8306 13666
rect 94 12520 120 13640
rect 160 13574 8240 13600
rect 160 12632 232 13574
rect 8214 12632 8240 13574
rect 160 12560 8240 12632
rect 8280 12520 8306 13640
rect 8320 12560 8392 13680
rect 12488 13680 20872 13752
rect 12488 13600 12560 13680
rect 12574 13640 20786 13666
rect 94 12494 8306 12520
rect 12574 12520 12600 13640
rect 12640 13574 20720 13600
rect 12640 12632 12712 13574
rect 20694 12632 20720 13574
rect 12640 12560 20720 12632
rect 20760 12520 20786 13640
rect 20800 12560 20872 13680
rect 12574 12494 20786 12520
rect 8 11040 8392 11112
rect 8 10960 80 11040
rect 94 11000 8306 11026
rect 94 9880 120 11000
rect 160 10934 8240 10960
rect 160 9992 232 10934
rect 8214 9992 8240 10934
rect 160 9920 8240 9992
rect 8280 9880 8306 11000
rect 8320 9920 8392 11040
rect 12488 11040 20872 11112
rect 12488 10960 12560 11040
rect 12574 11000 20786 11026
rect 94 9854 8306 9880
rect 12574 9880 12600 11000
rect 12640 10934 20720 10960
rect 12640 9992 12712 10934
rect 20694 9992 20720 10934
rect 12640 9920 20720 9992
rect 20760 9880 20786 11000
rect 20800 9920 20872 11040
rect 12574 9854 20786 9880
rect 8 6400 8392 6472
rect 8 6320 80 6400
rect 94 6360 8306 6386
rect 94 5240 120 6360
rect 160 6294 8240 6320
rect 160 5352 232 6294
rect 8214 5352 8240 6294
rect 160 5280 8240 5352
rect 8280 5240 8306 6360
rect 8320 5280 8392 6400
rect 12488 6400 20872 6472
rect 12488 6320 12560 6400
rect 12574 6360 20786 6386
rect 94 5214 8306 5240
rect 12574 5240 12600 6360
rect 12640 6294 20720 6320
rect 12640 5352 12712 6294
rect 20694 5352 20720 6294
rect 12640 5280 20720 5352
rect 20760 5240 20786 6360
rect 20800 5280 20872 6400
rect 12574 5214 20786 5240
rect 8 4960 8392 5032
rect 8 4880 80 4960
rect 94 4920 8306 4946
rect 94 3800 120 4920
rect 160 4854 8240 4880
rect 160 3912 232 4854
rect 8214 3912 8240 4854
rect 160 3840 8240 3912
rect 8280 3800 8306 4920
rect 8320 3840 8392 4960
rect 12488 4960 20872 5032
rect 12488 4880 12560 4960
rect 12574 4920 20786 4946
rect 94 3774 8306 3800
rect 12574 3800 12600 4920
rect 12640 4854 20720 4880
rect 12640 3912 12712 4854
rect 20694 3912 20720 4854
rect 12640 3840 20720 3912
rect 20760 3800 20786 4920
rect 20800 3840 20872 4960
rect 12574 3774 20786 3800
rect 8 3520 8392 3592
rect 8 3440 80 3520
rect 94 3480 8306 3506
rect 94 2360 120 3480
rect 160 3414 8240 3440
rect 160 2472 232 3414
rect 8214 2472 8240 3414
rect 160 2400 8240 2472
rect 8280 2360 8306 3480
rect 8320 2400 8392 3520
rect 12488 3520 20872 3592
rect 12488 3440 12560 3520
rect 12574 3480 20786 3506
rect 94 2334 8306 2360
rect 12574 2360 12600 3480
rect 12640 3414 20720 3440
rect 12640 2472 12712 3414
rect 20694 2472 20720 3414
rect 12640 2400 20720 2472
rect 20760 2360 20786 3480
rect 20800 2400 20872 3520
rect 12574 2334 20786 2360
<< locali >>
rect 8480 31417 8880 31440
rect 8480 31383 8503 31417
rect 8537 31383 8663 31417
rect 8697 31383 8823 31417
rect 8857 31383 8880 31417
rect 8480 31360 8880 31383
rect 8960 31417 9360 31440
rect 8960 31383 8983 31417
rect 9017 31383 9143 31417
rect 9177 31383 9303 31417
rect 9337 31383 9360 31417
rect 8960 31360 9360 31383
rect 9440 31417 11440 31440
rect 9440 31383 9463 31417
rect 9497 31383 9623 31417
rect 9657 31383 9783 31417
rect 9817 31383 9943 31417
rect 9977 31383 10103 31417
rect 10137 31383 10263 31417
rect 10297 31383 10423 31417
rect 10457 31383 10583 31417
rect 10617 31383 10743 31417
rect 10777 31383 10903 31417
rect 10937 31383 11063 31417
rect 11097 31383 11223 31417
rect 11257 31383 11383 31417
rect 11417 31383 11440 31417
rect 9440 31360 11440 31383
rect 11520 31417 11920 31440
rect 11520 31383 11543 31417
rect 11577 31383 11703 31417
rect 11737 31383 11863 31417
rect 11897 31383 11920 31417
rect 11520 31360 11920 31383
rect 12000 31417 12400 31440
rect 12000 31383 12023 31417
rect 12057 31383 12183 31417
rect 12217 31383 12343 31417
rect 12377 31383 12400 31417
rect 12000 31360 12400 31383
rect 8480 31257 8880 31280
rect 8480 31223 8503 31257
rect 8537 31223 8663 31257
rect 8697 31223 8823 31257
rect 8857 31223 8880 31257
rect 8480 31200 8880 31223
rect 8960 31257 9360 31280
rect 8960 31223 8983 31257
rect 9017 31223 9143 31257
rect 9177 31223 9303 31257
rect 9337 31223 9360 31257
rect 8960 31200 9360 31223
rect 9440 31257 11440 31280
rect 9440 31223 9463 31257
rect 9497 31223 9623 31257
rect 9657 31223 9783 31257
rect 9817 31223 9943 31257
rect 9977 31223 10103 31257
rect 10137 31223 10263 31257
rect 10297 31223 10423 31257
rect 10457 31223 10583 31257
rect 10617 31223 10743 31257
rect 10777 31223 10903 31257
rect 10937 31223 11063 31257
rect 11097 31223 11223 31257
rect 11257 31223 11383 31257
rect 11417 31223 11440 31257
rect 9440 31200 11440 31223
rect 11520 31257 11920 31280
rect 11520 31223 11543 31257
rect 11577 31223 11703 31257
rect 11737 31223 11863 31257
rect 11897 31223 11920 31257
rect 11520 31200 11920 31223
rect 12000 31257 12400 31280
rect 12000 31223 12023 31257
rect 12057 31223 12183 31257
rect 12217 31223 12343 31257
rect 12377 31223 12400 31257
rect 12000 31200 12400 31223
rect 8480 31097 8880 31120
rect 8480 31063 8503 31097
rect 8537 31063 8663 31097
rect 8697 31063 8823 31097
rect 8857 31063 8880 31097
rect 8480 31040 8880 31063
rect 8960 31097 9360 31120
rect 8960 31063 8983 31097
rect 9017 31063 9143 31097
rect 9177 31063 9303 31097
rect 9337 31063 9360 31097
rect 8960 31040 9360 31063
rect 9440 31097 11440 31120
rect 9440 31063 9463 31097
rect 9497 31063 9623 31097
rect 9657 31063 9783 31097
rect 9817 31063 9943 31097
rect 9977 31063 10103 31097
rect 10137 31063 10263 31097
rect 10297 31063 10423 31097
rect 10457 31063 10583 31097
rect 10617 31063 10743 31097
rect 10777 31063 10903 31097
rect 10937 31063 11063 31097
rect 11097 31063 11223 31097
rect 11257 31063 11383 31097
rect 11417 31063 11440 31097
rect 9440 31040 11440 31063
rect 11520 31097 11920 31120
rect 11520 31063 11543 31097
rect 11577 31063 11703 31097
rect 11737 31063 11863 31097
rect 11897 31063 11920 31097
rect 11520 31040 11920 31063
rect 12000 31097 12400 31120
rect 12000 31063 12023 31097
rect 12057 31063 12183 31097
rect 12217 31063 12343 31097
rect 12377 31063 12400 31097
rect 12000 31040 12400 31063
rect 8480 30937 8880 30960
rect 8480 30903 8503 30937
rect 8537 30903 8663 30937
rect 8697 30903 8823 30937
rect 8857 30903 8880 30937
rect 8480 30880 8880 30903
rect 8960 30937 9360 30960
rect 8960 30903 8983 30937
rect 9017 30903 9143 30937
rect 9177 30903 9303 30937
rect 9337 30903 9360 30937
rect 8960 30880 9360 30903
rect 9440 30937 11440 30960
rect 9440 30903 9463 30937
rect 9497 30903 9623 30937
rect 9657 30903 9783 30937
rect 9817 30903 9943 30937
rect 9977 30903 10103 30937
rect 10137 30903 10263 30937
rect 10297 30903 10423 30937
rect 10457 30903 10583 30937
rect 10617 30903 10743 30937
rect 10777 30903 10903 30937
rect 10937 30903 11063 30937
rect 11097 30903 11223 30937
rect 11257 30903 11383 30937
rect 11417 30903 11440 30937
rect 9440 30880 11440 30903
rect 11520 30937 11920 30960
rect 11520 30903 11543 30937
rect 11577 30903 11703 30937
rect 11737 30903 11863 30937
rect 11897 30903 11920 30937
rect 11520 30880 11920 30903
rect 12000 30937 12400 30960
rect 12000 30903 12023 30937
rect 12057 30903 12183 30937
rect 12217 30903 12343 30937
rect 12377 30903 12400 30937
rect 12000 30880 12400 30903
rect 8480 30777 8880 30800
rect 8480 30743 8503 30777
rect 8537 30743 8663 30777
rect 8697 30743 8823 30777
rect 8857 30743 8880 30777
rect 8480 30720 8880 30743
rect 8960 30777 9360 30800
rect 8960 30743 8983 30777
rect 9017 30743 9143 30777
rect 9177 30743 9303 30777
rect 9337 30743 9360 30777
rect 8960 30720 9360 30743
rect 9440 30777 11440 30800
rect 9440 30743 9463 30777
rect 9497 30743 9623 30777
rect 9657 30743 9783 30777
rect 9817 30743 9943 30777
rect 9977 30743 10103 30777
rect 10137 30743 10263 30777
rect 10297 30743 10423 30777
rect 10457 30743 10583 30777
rect 10617 30743 10743 30777
rect 10777 30743 10903 30777
rect 10937 30743 11063 30777
rect 11097 30743 11223 30777
rect 11257 30743 11383 30777
rect 11417 30743 11440 30777
rect 9440 30720 11440 30743
rect 11520 30777 11920 30800
rect 11520 30743 11543 30777
rect 11577 30743 11703 30777
rect 11737 30743 11863 30777
rect 11897 30743 11920 30777
rect 11520 30720 11920 30743
rect 12000 30777 12400 30800
rect 12000 30743 12023 30777
rect 12057 30743 12183 30777
rect 12217 30743 12343 30777
rect 12377 30743 12400 30777
rect 12000 30720 12400 30743
rect 8480 30617 8880 30640
rect 8480 30583 8503 30617
rect 8537 30583 8663 30617
rect 8697 30583 8823 30617
rect 8857 30583 8880 30617
rect 8480 30560 8880 30583
rect 8960 30617 9360 30640
rect 8960 30583 8983 30617
rect 9017 30583 9143 30617
rect 9177 30583 9303 30617
rect 9337 30583 9360 30617
rect 8960 30560 9360 30583
rect 9440 30617 11440 30640
rect 9440 30583 9463 30617
rect 9497 30583 9623 30617
rect 9657 30583 9783 30617
rect 9817 30583 9943 30617
rect 9977 30583 10103 30617
rect 10137 30583 10263 30617
rect 10297 30583 10423 30617
rect 10457 30583 10583 30617
rect 10617 30583 10743 30617
rect 10777 30583 10903 30617
rect 10937 30583 11063 30617
rect 11097 30583 11223 30617
rect 11257 30583 11383 30617
rect 11417 30583 11440 30617
rect 9440 30560 11440 30583
rect 11520 30617 11920 30640
rect 11520 30583 11543 30617
rect 11577 30583 11703 30617
rect 11737 30583 11863 30617
rect 11897 30583 11920 30617
rect 11520 30560 11920 30583
rect 12000 30617 12400 30640
rect 12000 30583 12023 30617
rect 12057 30583 12183 30617
rect 12217 30583 12343 30617
rect 12377 30583 12400 30617
rect 12000 30560 12400 30583
rect 8480 30457 8880 30480
rect 8480 30423 8503 30457
rect 8537 30423 8663 30457
rect 8697 30423 8823 30457
rect 8857 30423 8880 30457
rect 8480 30400 8880 30423
rect 8960 30457 9360 30480
rect 8960 30423 8983 30457
rect 9017 30423 9143 30457
rect 9177 30423 9303 30457
rect 9337 30423 9360 30457
rect 8960 30400 9360 30423
rect 9440 30457 11440 30480
rect 9440 30423 9463 30457
rect 9497 30423 9623 30457
rect 9657 30423 9783 30457
rect 9817 30423 9943 30457
rect 9977 30423 10103 30457
rect 10137 30423 10263 30457
rect 10297 30423 10423 30457
rect 10457 30423 10583 30457
rect 10617 30423 10743 30457
rect 10777 30423 10903 30457
rect 10937 30423 11063 30457
rect 11097 30423 11223 30457
rect 11257 30423 11383 30457
rect 11417 30423 11440 30457
rect 9440 30400 11440 30423
rect 11520 30457 11920 30480
rect 11520 30423 11543 30457
rect 11577 30423 11703 30457
rect 11737 30423 11863 30457
rect 11897 30423 11920 30457
rect 11520 30400 11920 30423
rect 12000 30457 12400 30480
rect 12000 30423 12023 30457
rect 12057 30423 12183 30457
rect 12217 30423 12343 30457
rect 12377 30423 12400 30457
rect 12000 30400 12400 30423
rect 8480 30297 8880 30320
rect 8480 30263 8503 30297
rect 8537 30263 8663 30297
rect 8697 30263 8823 30297
rect 8857 30263 8880 30297
rect 8480 30240 8880 30263
rect 8960 30297 9360 30320
rect 8960 30263 8983 30297
rect 9017 30263 9143 30297
rect 9177 30263 9303 30297
rect 9337 30263 9360 30297
rect 8960 30240 9360 30263
rect 9440 30297 11440 30320
rect 9440 30263 9463 30297
rect 9497 30263 9623 30297
rect 9657 30263 9783 30297
rect 9817 30263 9943 30297
rect 9977 30263 10103 30297
rect 10137 30263 10263 30297
rect 10297 30263 10423 30297
rect 10457 30263 10583 30297
rect 10617 30263 10743 30297
rect 10777 30263 10903 30297
rect 10937 30263 11063 30297
rect 11097 30263 11223 30297
rect 11257 30263 11383 30297
rect 11417 30263 11440 30297
rect 9440 30240 11440 30263
rect 11520 30297 11920 30320
rect 11520 30263 11543 30297
rect 11577 30263 11703 30297
rect 11737 30263 11863 30297
rect 11897 30263 11920 30297
rect 11520 30240 11920 30263
rect 12000 30297 12400 30320
rect 12000 30263 12023 30297
rect 12057 30263 12183 30297
rect 12217 30263 12343 30297
rect 12377 30263 12400 30297
rect 12000 30240 12400 30263
rect 8480 30137 8880 30160
rect 8480 30103 8503 30137
rect 8537 30103 8663 30137
rect 8697 30103 8823 30137
rect 8857 30103 8880 30137
rect 8480 30080 8880 30103
rect 8960 30137 9360 30160
rect 8960 30103 8983 30137
rect 9017 30103 9143 30137
rect 9177 30103 9303 30137
rect 9337 30103 9360 30137
rect 8960 30080 9360 30103
rect 9440 30137 11440 30160
rect 9440 30103 9463 30137
rect 9497 30103 9623 30137
rect 9657 30103 9783 30137
rect 9817 30103 9943 30137
rect 9977 30103 10103 30137
rect 10137 30103 10263 30137
rect 10297 30103 10423 30137
rect 10457 30103 10583 30137
rect 10617 30103 10743 30137
rect 10777 30103 10903 30137
rect 10937 30103 11063 30137
rect 11097 30103 11223 30137
rect 11257 30103 11383 30137
rect 11417 30103 11440 30137
rect 9440 30080 11440 30103
rect 11520 30137 11920 30160
rect 11520 30103 11543 30137
rect 11577 30103 11703 30137
rect 11737 30103 11863 30137
rect 11897 30103 11920 30137
rect 11520 30080 11920 30103
rect 12000 30137 12400 30160
rect 12000 30103 12023 30137
rect 12057 30103 12183 30137
rect 12217 30103 12343 30137
rect 12377 30103 12400 30137
rect 12000 30080 12400 30103
rect 8480 29977 8880 30000
rect 8480 29943 8503 29977
rect 8537 29943 8663 29977
rect 8697 29943 8823 29977
rect 8857 29943 8880 29977
rect 8480 29920 8880 29943
rect 8960 29977 9360 30000
rect 8960 29943 8983 29977
rect 9017 29943 9143 29977
rect 9177 29943 9303 29977
rect 9337 29943 9360 29977
rect 8960 29920 9360 29943
rect 9440 29977 11440 30000
rect 9440 29943 9463 29977
rect 9497 29943 9623 29977
rect 9657 29943 9783 29977
rect 9817 29943 9943 29977
rect 9977 29943 10103 29977
rect 10137 29943 10263 29977
rect 10297 29943 10423 29977
rect 10457 29943 10583 29977
rect 10617 29943 10743 29977
rect 10777 29943 10903 29977
rect 10937 29943 11063 29977
rect 11097 29943 11223 29977
rect 11257 29943 11383 29977
rect 11417 29943 11440 29977
rect 9440 29920 11440 29943
rect 11520 29977 11920 30000
rect 11520 29943 11543 29977
rect 11577 29943 11703 29977
rect 11737 29943 11863 29977
rect 11897 29943 11920 29977
rect 11520 29920 11920 29943
rect 12000 29977 12400 30000
rect 12000 29943 12023 29977
rect 12057 29943 12183 29977
rect 12217 29943 12343 29977
rect 12377 29943 12400 29977
rect 12000 29920 12400 29943
rect 8480 29817 8880 29840
rect 8480 29783 8503 29817
rect 8537 29783 8663 29817
rect 8697 29783 8823 29817
rect 8857 29783 8880 29817
rect 8480 29760 8880 29783
rect 8960 29817 9360 29840
rect 8960 29783 8983 29817
rect 9017 29783 9143 29817
rect 9177 29783 9303 29817
rect 9337 29783 9360 29817
rect 8960 29760 9360 29783
rect 9440 29817 11440 29840
rect 9440 29783 9463 29817
rect 9497 29783 9623 29817
rect 9657 29783 9783 29817
rect 9817 29783 9943 29817
rect 9977 29783 10103 29817
rect 10137 29783 10263 29817
rect 10297 29783 10423 29817
rect 10457 29783 10583 29817
rect 10617 29783 10743 29817
rect 10777 29783 10903 29817
rect 10937 29783 11063 29817
rect 11097 29783 11223 29817
rect 11257 29783 11383 29817
rect 11417 29783 11440 29817
rect 9440 29760 11440 29783
rect 11520 29817 11920 29840
rect 11520 29783 11543 29817
rect 11577 29783 11703 29817
rect 11737 29783 11863 29817
rect 11897 29783 11920 29817
rect 11520 29760 11920 29783
rect 12000 29817 12400 29840
rect 12000 29783 12023 29817
rect 12057 29783 12183 29817
rect 12217 29783 12343 29817
rect 12377 29783 12400 29817
rect 12000 29760 12400 29783
rect 8480 29657 8880 29680
rect 8480 29623 8503 29657
rect 8537 29623 8663 29657
rect 8697 29623 8823 29657
rect 8857 29623 8880 29657
rect 8480 29600 8880 29623
rect 8960 29657 9360 29680
rect 8960 29623 8983 29657
rect 9017 29623 9143 29657
rect 9177 29623 9303 29657
rect 9337 29623 9360 29657
rect 8960 29600 9360 29623
rect 9440 29657 11440 29680
rect 9440 29623 9463 29657
rect 9497 29623 9623 29657
rect 9657 29623 9783 29657
rect 9817 29623 9943 29657
rect 9977 29623 10103 29657
rect 10137 29623 10263 29657
rect 10297 29623 10423 29657
rect 10457 29623 10583 29657
rect 10617 29623 10743 29657
rect 10777 29623 10903 29657
rect 10937 29623 11063 29657
rect 11097 29623 11223 29657
rect 11257 29623 11383 29657
rect 11417 29623 11440 29657
rect 9440 29600 11440 29623
rect 11520 29657 11920 29680
rect 11520 29623 11543 29657
rect 11577 29623 11703 29657
rect 11737 29623 11863 29657
rect 11897 29623 11920 29657
rect 11520 29600 11920 29623
rect 12000 29657 12400 29680
rect 12000 29623 12023 29657
rect 12057 29623 12183 29657
rect 12217 29623 12343 29657
rect 12377 29623 12400 29657
rect 12000 29600 12400 29623
rect 8480 29497 8880 29520
rect 8480 29463 8503 29497
rect 8537 29463 8663 29497
rect 8697 29463 8823 29497
rect 8857 29463 8880 29497
rect 8480 29440 8880 29463
rect 8960 29497 9360 29520
rect 8960 29463 8983 29497
rect 9017 29463 9143 29497
rect 9177 29463 9303 29497
rect 9337 29463 9360 29497
rect 8960 29440 9360 29463
rect 9440 29497 11440 29520
rect 9440 29463 9463 29497
rect 9497 29463 9623 29497
rect 9657 29463 9783 29497
rect 9817 29463 9943 29497
rect 9977 29463 10103 29497
rect 10137 29463 10263 29497
rect 10297 29463 10423 29497
rect 10457 29463 10583 29497
rect 10617 29463 10743 29497
rect 10777 29463 10903 29497
rect 10937 29463 11063 29497
rect 11097 29463 11223 29497
rect 11257 29463 11383 29497
rect 11417 29463 11440 29497
rect 9440 29440 11440 29463
rect 11520 29497 11920 29520
rect 11520 29463 11543 29497
rect 11577 29463 11703 29497
rect 11737 29463 11863 29497
rect 11897 29463 11920 29497
rect 11520 29440 11920 29463
rect 12000 29497 12400 29520
rect 12000 29463 12023 29497
rect 12057 29463 12183 29497
rect 12217 29463 12343 29497
rect 12377 29463 12400 29497
rect 12000 29440 12400 29463
rect 8480 29337 8880 29360
rect 8480 29303 8503 29337
rect 8537 29303 8663 29337
rect 8697 29303 8823 29337
rect 8857 29303 8880 29337
rect 8480 29280 8880 29303
rect 8960 29337 9360 29360
rect 8960 29303 8983 29337
rect 9017 29303 9143 29337
rect 9177 29303 9303 29337
rect 9337 29303 9360 29337
rect 8960 29280 9360 29303
rect 9440 29337 11440 29360
rect 9440 29303 9463 29337
rect 9497 29303 9623 29337
rect 9657 29303 9783 29337
rect 9817 29303 9943 29337
rect 9977 29303 10103 29337
rect 10137 29303 10263 29337
rect 10297 29303 10423 29337
rect 10457 29303 10583 29337
rect 10617 29303 10743 29337
rect 10777 29303 10903 29337
rect 10937 29303 11063 29337
rect 11097 29303 11223 29337
rect 11257 29303 11383 29337
rect 11417 29303 11440 29337
rect 9440 29280 11440 29303
rect 11520 29337 11920 29360
rect 11520 29303 11543 29337
rect 11577 29303 11703 29337
rect 11737 29303 11863 29337
rect 11897 29303 11920 29337
rect 11520 29280 11920 29303
rect 12000 29337 12400 29360
rect 12000 29303 12023 29337
rect 12057 29303 12183 29337
rect 12217 29303 12343 29337
rect 12377 29303 12400 29337
rect 12000 29280 12400 29303
rect 8480 29177 8880 29200
rect 8480 29143 8503 29177
rect 8537 29143 8663 29177
rect 8697 29143 8823 29177
rect 8857 29143 8880 29177
rect 8480 29120 8880 29143
rect 8960 29177 9360 29200
rect 8960 29143 8983 29177
rect 9017 29143 9143 29177
rect 9177 29143 9303 29177
rect 9337 29143 9360 29177
rect 8960 29120 9360 29143
rect 9440 29177 11440 29200
rect 9440 29143 9463 29177
rect 9497 29143 9623 29177
rect 9657 29143 9783 29177
rect 9817 29143 9943 29177
rect 9977 29143 10103 29177
rect 10137 29143 10263 29177
rect 10297 29143 10423 29177
rect 10457 29143 10583 29177
rect 10617 29143 10743 29177
rect 10777 29143 10903 29177
rect 10937 29143 11063 29177
rect 11097 29143 11223 29177
rect 11257 29143 11383 29177
rect 11417 29143 11440 29177
rect 9440 29120 11440 29143
rect 11520 29177 11920 29200
rect 11520 29143 11543 29177
rect 11577 29143 11703 29177
rect 11737 29143 11863 29177
rect 11897 29143 11920 29177
rect 11520 29120 11920 29143
rect 12000 29177 12400 29200
rect 12000 29143 12023 29177
rect 12057 29143 12183 29177
rect 12217 29143 12343 29177
rect 12377 29143 12400 29177
rect 12000 29120 12400 29143
rect 8480 29017 8880 29040
rect 8480 28983 8503 29017
rect 8537 28983 8663 29017
rect 8697 28983 8823 29017
rect 8857 28983 8880 29017
rect 8480 28960 8880 28983
rect 8960 29017 9360 29040
rect 8960 28983 8983 29017
rect 9017 28983 9143 29017
rect 9177 28983 9303 29017
rect 9337 28983 9360 29017
rect 8960 28960 9360 28983
rect 9440 29017 11440 29040
rect 9440 28983 9463 29017
rect 9497 28983 9623 29017
rect 9657 28983 9783 29017
rect 9817 28983 9943 29017
rect 9977 28983 10103 29017
rect 10137 28983 10263 29017
rect 10297 28983 10423 29017
rect 10457 28983 10583 29017
rect 10617 28983 10743 29017
rect 10777 28983 10903 29017
rect 10937 28983 11063 29017
rect 11097 28983 11223 29017
rect 11257 28983 11383 29017
rect 11417 28983 11440 29017
rect 9440 28960 11440 28983
rect 11520 29017 11920 29040
rect 11520 28983 11543 29017
rect 11577 28983 11703 29017
rect 11737 28983 11863 29017
rect 11897 28983 11920 29017
rect 11520 28960 11920 28983
rect 12000 29017 12400 29040
rect 12000 28983 12023 29017
rect 12057 28983 12183 29017
rect 12217 28983 12343 29017
rect 12377 28983 12400 29017
rect 12000 28960 12400 28983
rect 8480 28857 8880 28880
rect 8480 28823 8503 28857
rect 8537 28823 8663 28857
rect 8697 28823 8823 28857
rect 8857 28823 8880 28857
rect 8480 28800 8880 28823
rect 8960 28857 9360 28880
rect 8960 28823 8983 28857
rect 9017 28823 9143 28857
rect 9177 28823 9303 28857
rect 9337 28823 9360 28857
rect 8960 28800 9360 28823
rect 9440 28857 11440 28880
rect 9440 28823 9463 28857
rect 9497 28823 9623 28857
rect 9657 28823 9783 28857
rect 9817 28823 9943 28857
rect 9977 28823 10103 28857
rect 10137 28823 10263 28857
rect 10297 28823 10423 28857
rect 10457 28823 10583 28857
rect 10617 28823 10743 28857
rect 10777 28823 10903 28857
rect 10937 28823 11063 28857
rect 11097 28823 11223 28857
rect 11257 28823 11383 28857
rect 11417 28823 11440 28857
rect 9440 28800 11440 28823
rect 11520 28857 11920 28880
rect 11520 28823 11543 28857
rect 11577 28823 11703 28857
rect 11737 28823 11863 28857
rect 11897 28823 11920 28857
rect 11520 28800 11920 28823
rect 12000 28857 12400 28880
rect 12000 28823 12023 28857
rect 12057 28823 12183 28857
rect 12217 28823 12343 28857
rect 12377 28823 12400 28857
rect 12000 28800 12400 28823
rect 8480 28697 8880 28720
rect 8480 28663 8503 28697
rect 8537 28663 8663 28697
rect 8697 28663 8823 28697
rect 8857 28663 8880 28697
rect 8480 28640 8880 28663
rect 8960 28697 9360 28720
rect 8960 28663 8983 28697
rect 9017 28663 9143 28697
rect 9177 28663 9303 28697
rect 9337 28663 9360 28697
rect 8960 28640 9360 28663
rect 9440 28697 11440 28720
rect 9440 28663 9463 28697
rect 9497 28663 9623 28697
rect 9657 28663 9783 28697
rect 9817 28663 9943 28697
rect 9977 28663 10103 28697
rect 10137 28663 10263 28697
rect 10297 28663 10423 28697
rect 10457 28663 10583 28697
rect 10617 28663 10743 28697
rect 10777 28663 10903 28697
rect 10937 28663 11063 28697
rect 11097 28663 11223 28697
rect 11257 28663 11383 28697
rect 11417 28663 11440 28697
rect 9440 28640 11440 28663
rect 11520 28697 11920 28720
rect 11520 28663 11543 28697
rect 11577 28663 11703 28697
rect 11737 28663 11863 28697
rect 11897 28663 11920 28697
rect 11520 28640 11920 28663
rect 12000 28697 12400 28720
rect 12000 28663 12023 28697
rect 12057 28663 12183 28697
rect 12217 28663 12343 28697
rect 12377 28663 12400 28697
rect 12000 28640 12400 28663
rect 8480 28537 8880 28560
rect 8480 28503 8503 28537
rect 8537 28503 8663 28537
rect 8697 28503 8823 28537
rect 8857 28503 8880 28537
rect 8480 28480 8880 28503
rect 8960 28537 9360 28560
rect 8960 28503 8983 28537
rect 9017 28503 9143 28537
rect 9177 28503 9303 28537
rect 9337 28503 9360 28537
rect 8960 28480 9360 28503
rect 9440 28537 11440 28560
rect 9440 28503 9463 28537
rect 9497 28503 9623 28537
rect 9657 28503 9783 28537
rect 9817 28503 9943 28537
rect 9977 28503 10103 28537
rect 10137 28503 10263 28537
rect 10297 28503 10423 28537
rect 10457 28503 10583 28537
rect 10617 28503 10743 28537
rect 10777 28503 10903 28537
rect 10937 28503 11063 28537
rect 11097 28503 11223 28537
rect 11257 28503 11383 28537
rect 11417 28503 11440 28537
rect 9440 28480 11440 28503
rect 11520 28537 11920 28560
rect 11520 28503 11543 28537
rect 11577 28503 11703 28537
rect 11737 28503 11863 28537
rect 11897 28503 11920 28537
rect 11520 28480 11920 28503
rect 12000 28537 12400 28560
rect 12000 28503 12023 28537
rect 12057 28503 12183 28537
rect 12217 28503 12343 28537
rect 12377 28503 12400 28537
rect 12000 28480 12400 28503
rect 8480 28377 8880 28400
rect 8480 28343 8503 28377
rect 8537 28343 8663 28377
rect 8697 28343 8823 28377
rect 8857 28343 8880 28377
rect 8480 28320 8880 28343
rect 8960 28377 9360 28400
rect 8960 28343 8983 28377
rect 9017 28343 9143 28377
rect 9177 28343 9303 28377
rect 9337 28343 9360 28377
rect 8960 28320 9360 28343
rect 9440 28377 11440 28400
rect 9440 28343 9463 28377
rect 9497 28343 9623 28377
rect 9657 28343 9783 28377
rect 9817 28343 9943 28377
rect 9977 28343 10103 28377
rect 10137 28343 10263 28377
rect 10297 28343 10423 28377
rect 10457 28343 10583 28377
rect 10617 28343 10743 28377
rect 10777 28343 10903 28377
rect 10937 28343 11063 28377
rect 11097 28343 11223 28377
rect 11257 28343 11383 28377
rect 11417 28343 11440 28377
rect 9440 28320 11440 28343
rect 11520 28377 11920 28400
rect 11520 28343 11543 28377
rect 11577 28343 11703 28377
rect 11737 28343 11863 28377
rect 11897 28343 11920 28377
rect 11520 28320 11920 28343
rect 12000 28377 12400 28400
rect 12000 28343 12023 28377
rect 12057 28343 12183 28377
rect 12217 28343 12343 28377
rect 12377 28343 12400 28377
rect 12000 28320 12400 28343
rect 8480 28217 8880 28240
rect 8480 28183 8503 28217
rect 8537 28183 8663 28217
rect 8697 28183 8823 28217
rect 8857 28183 8880 28217
rect 8480 28160 8880 28183
rect 8960 28217 9360 28240
rect 8960 28183 8983 28217
rect 9017 28183 9143 28217
rect 9177 28183 9303 28217
rect 9337 28183 9360 28217
rect 8960 28160 9360 28183
rect 9440 28217 11440 28240
rect 9440 28183 9463 28217
rect 9497 28183 9623 28217
rect 9657 28183 9783 28217
rect 9817 28183 9943 28217
rect 9977 28183 10103 28217
rect 10137 28183 10263 28217
rect 10297 28183 10423 28217
rect 10457 28183 10583 28217
rect 10617 28183 10743 28217
rect 10777 28183 10903 28217
rect 10937 28183 11063 28217
rect 11097 28183 11223 28217
rect 11257 28183 11383 28217
rect 11417 28183 11440 28217
rect 9440 28160 11440 28183
rect 11520 28217 11920 28240
rect 11520 28183 11543 28217
rect 11577 28183 11703 28217
rect 11737 28183 11863 28217
rect 11897 28183 11920 28217
rect 11520 28160 11920 28183
rect 12000 28217 12400 28240
rect 12000 28183 12023 28217
rect 12057 28183 12183 28217
rect 12217 28183 12343 28217
rect 12377 28183 12400 28217
rect 12000 28160 12400 28183
rect 8480 28057 8880 28080
rect 8480 28023 8503 28057
rect 8537 28023 8663 28057
rect 8697 28023 8823 28057
rect 8857 28023 8880 28057
rect 8480 28000 8880 28023
rect 8960 28057 9360 28080
rect 8960 28023 8983 28057
rect 9017 28023 9143 28057
rect 9177 28023 9303 28057
rect 9337 28023 9360 28057
rect 8960 28000 9360 28023
rect 9440 28057 11440 28080
rect 9440 28023 9463 28057
rect 9497 28023 9623 28057
rect 9657 28023 9783 28057
rect 9817 28023 9943 28057
rect 9977 28023 10103 28057
rect 10137 28023 10263 28057
rect 10297 28023 10423 28057
rect 10457 28023 10583 28057
rect 10617 28023 10743 28057
rect 10777 28023 10903 28057
rect 10937 28023 11063 28057
rect 11097 28023 11223 28057
rect 11257 28023 11383 28057
rect 11417 28023 11440 28057
rect 9440 28000 11440 28023
rect 11520 28057 11920 28080
rect 11520 28023 11543 28057
rect 11577 28023 11703 28057
rect 11737 28023 11863 28057
rect 11897 28023 11920 28057
rect 11520 28000 11920 28023
rect 12000 28057 12400 28080
rect 12000 28023 12023 28057
rect 12057 28023 12183 28057
rect 12217 28023 12343 28057
rect 12377 28023 12400 28057
rect 12000 28000 12400 28023
rect 8480 27897 8880 27920
rect 8480 27863 8503 27897
rect 8537 27863 8663 27897
rect 8697 27863 8823 27897
rect 8857 27863 8880 27897
rect 8480 27840 8880 27863
rect 8960 27897 9360 27920
rect 8960 27863 8983 27897
rect 9017 27863 9143 27897
rect 9177 27863 9303 27897
rect 9337 27863 9360 27897
rect 8960 27840 9360 27863
rect 9440 27897 11440 27920
rect 9440 27863 9463 27897
rect 9497 27863 9623 27897
rect 9657 27863 9783 27897
rect 9817 27863 9943 27897
rect 9977 27863 10103 27897
rect 10137 27863 10263 27897
rect 10297 27863 10423 27897
rect 10457 27863 10583 27897
rect 10617 27863 10743 27897
rect 10777 27863 10903 27897
rect 10937 27863 11063 27897
rect 11097 27863 11223 27897
rect 11257 27863 11383 27897
rect 11417 27863 11440 27897
rect 9440 27840 11440 27863
rect 11520 27897 11920 27920
rect 11520 27863 11543 27897
rect 11577 27863 11703 27897
rect 11737 27863 11863 27897
rect 11897 27863 11920 27897
rect 11520 27840 11920 27863
rect 12000 27897 12400 27920
rect 12000 27863 12023 27897
rect 12057 27863 12183 27897
rect 12217 27863 12343 27897
rect 12377 27863 12400 27897
rect 12000 27840 12400 27863
rect 8480 27737 8880 27760
rect 8480 27703 8503 27737
rect 8537 27703 8663 27737
rect 8697 27703 8823 27737
rect 8857 27703 8880 27737
rect 8480 27680 8880 27703
rect 8960 27737 9360 27760
rect 8960 27703 8983 27737
rect 9017 27703 9143 27737
rect 9177 27703 9303 27737
rect 9337 27703 9360 27737
rect 8960 27680 9360 27703
rect 9440 27737 11440 27760
rect 9440 27703 9463 27737
rect 9497 27703 9623 27737
rect 9657 27703 9783 27737
rect 9817 27703 9943 27737
rect 9977 27703 10103 27737
rect 10137 27703 10263 27737
rect 10297 27703 10423 27737
rect 10457 27703 10583 27737
rect 10617 27703 10743 27737
rect 10777 27703 10903 27737
rect 10937 27703 11063 27737
rect 11097 27703 11223 27737
rect 11257 27703 11383 27737
rect 11417 27703 11440 27737
rect 9440 27680 11440 27703
rect 11520 27737 11920 27760
rect 11520 27703 11543 27737
rect 11577 27703 11703 27737
rect 11737 27703 11863 27737
rect 11897 27703 11920 27737
rect 11520 27680 11920 27703
rect 12000 27737 12400 27760
rect 12000 27703 12023 27737
rect 12057 27703 12183 27737
rect 12217 27703 12343 27737
rect 12377 27703 12400 27737
rect 12000 27680 12400 27703
rect 8480 27577 8880 27600
rect 8480 27543 8503 27577
rect 8537 27543 8663 27577
rect 8697 27543 8823 27577
rect 8857 27543 8880 27577
rect 8480 27520 8880 27543
rect 8960 27577 9360 27600
rect 8960 27543 8983 27577
rect 9017 27543 9143 27577
rect 9177 27543 9303 27577
rect 9337 27543 9360 27577
rect 8960 27520 9360 27543
rect 9440 27577 11440 27600
rect 9440 27543 9463 27577
rect 9497 27543 9623 27577
rect 9657 27543 9783 27577
rect 9817 27543 9943 27577
rect 9977 27543 10103 27577
rect 10137 27543 10263 27577
rect 10297 27543 10423 27577
rect 10457 27543 10583 27577
rect 10617 27543 10743 27577
rect 10777 27543 10903 27577
rect 10937 27543 11063 27577
rect 11097 27543 11223 27577
rect 11257 27543 11383 27577
rect 11417 27543 11440 27577
rect 9440 27520 11440 27543
rect 11520 27577 11920 27600
rect 11520 27543 11543 27577
rect 11577 27543 11703 27577
rect 11737 27543 11863 27577
rect 11897 27543 11920 27577
rect 11520 27520 11920 27543
rect 12000 27577 12400 27600
rect 12000 27543 12023 27577
rect 12057 27543 12183 27577
rect 12217 27543 12343 27577
rect 12377 27543 12400 27577
rect 12000 27520 12400 27543
rect 8480 27417 8880 27440
rect 8480 27383 8503 27417
rect 8537 27383 8663 27417
rect 8697 27383 8823 27417
rect 8857 27383 8880 27417
rect 8480 27360 8880 27383
rect 8960 27417 9360 27440
rect 8960 27383 8983 27417
rect 9017 27383 9143 27417
rect 9177 27383 9303 27417
rect 9337 27383 9360 27417
rect 8960 27360 9360 27383
rect 9440 27417 11440 27440
rect 9440 27383 9463 27417
rect 9497 27383 9623 27417
rect 9657 27383 9783 27417
rect 9817 27383 9943 27417
rect 9977 27383 10103 27417
rect 10137 27383 10263 27417
rect 10297 27383 10423 27417
rect 10457 27383 10583 27417
rect 10617 27383 10743 27417
rect 10777 27383 10903 27417
rect 10937 27383 11063 27417
rect 11097 27383 11223 27417
rect 11257 27383 11383 27417
rect 11417 27383 11440 27417
rect 9440 27360 11440 27383
rect 11520 27417 11920 27440
rect 11520 27383 11543 27417
rect 11577 27383 11703 27417
rect 11737 27383 11863 27417
rect 11897 27383 11920 27417
rect 11520 27360 11920 27383
rect 12000 27417 12400 27440
rect 12000 27383 12023 27417
rect 12057 27383 12183 27417
rect 12217 27383 12343 27417
rect 12377 27383 12400 27417
rect 12000 27360 12400 27383
rect 8480 27257 8880 27280
rect 8480 27223 8503 27257
rect 8537 27223 8663 27257
rect 8697 27223 8823 27257
rect 8857 27223 8880 27257
rect 8480 27200 8880 27223
rect 8960 27257 9360 27280
rect 8960 27223 8983 27257
rect 9017 27223 9143 27257
rect 9177 27223 9303 27257
rect 9337 27223 9360 27257
rect 8960 27200 9360 27223
rect 9440 27257 11440 27280
rect 9440 27223 9463 27257
rect 9497 27223 9623 27257
rect 9657 27223 9783 27257
rect 9817 27223 9943 27257
rect 9977 27223 10103 27257
rect 10137 27223 10263 27257
rect 10297 27223 10423 27257
rect 10457 27223 10583 27257
rect 10617 27223 10743 27257
rect 10777 27223 10903 27257
rect 10937 27223 11063 27257
rect 11097 27223 11223 27257
rect 11257 27223 11383 27257
rect 11417 27223 11440 27257
rect 9440 27200 11440 27223
rect 11520 27257 11920 27280
rect 11520 27223 11543 27257
rect 11577 27223 11703 27257
rect 11737 27223 11863 27257
rect 11897 27223 11920 27257
rect 11520 27200 11920 27223
rect 12000 27257 12400 27280
rect 12000 27223 12023 27257
rect 12057 27223 12183 27257
rect 12217 27223 12343 27257
rect 12377 27223 12400 27257
rect 12000 27200 12400 27223
rect 8480 27097 8880 27120
rect 8480 27063 8503 27097
rect 8537 27063 8663 27097
rect 8697 27063 8823 27097
rect 8857 27063 8880 27097
rect 8480 27040 8880 27063
rect 8960 27097 9360 27120
rect 8960 27063 8983 27097
rect 9017 27063 9143 27097
rect 9177 27063 9303 27097
rect 9337 27063 9360 27097
rect 8960 27040 9360 27063
rect 9440 27097 11440 27120
rect 9440 27063 9463 27097
rect 9497 27063 9623 27097
rect 9657 27063 9783 27097
rect 9817 27063 9943 27097
rect 9977 27063 10103 27097
rect 10137 27063 10263 27097
rect 10297 27063 10423 27097
rect 10457 27063 10583 27097
rect 10617 27063 10743 27097
rect 10777 27063 10903 27097
rect 10937 27063 11063 27097
rect 11097 27063 11223 27097
rect 11257 27063 11383 27097
rect 11417 27063 11440 27097
rect 9440 27040 11440 27063
rect 11520 27097 11920 27120
rect 11520 27063 11543 27097
rect 11577 27063 11703 27097
rect 11737 27063 11863 27097
rect 11897 27063 11920 27097
rect 11520 27040 11920 27063
rect 12000 27097 12400 27120
rect 12000 27063 12023 27097
rect 12057 27063 12183 27097
rect 12217 27063 12343 27097
rect 12377 27063 12400 27097
rect 12000 27040 12400 27063
rect 8480 26937 8880 26960
rect 8480 26903 8503 26937
rect 8537 26903 8663 26937
rect 8697 26903 8823 26937
rect 8857 26903 8880 26937
rect 8480 26880 8880 26903
rect 8960 26937 9360 26960
rect 8960 26903 8983 26937
rect 9017 26903 9143 26937
rect 9177 26903 9303 26937
rect 9337 26903 9360 26937
rect 8960 26880 9360 26903
rect 9440 26937 11440 26960
rect 9440 26903 9463 26937
rect 9497 26903 9623 26937
rect 9657 26903 9783 26937
rect 9817 26903 9943 26937
rect 9977 26903 10103 26937
rect 10137 26903 10263 26937
rect 10297 26903 10423 26937
rect 10457 26903 10583 26937
rect 10617 26903 10743 26937
rect 10777 26903 10903 26937
rect 10937 26903 11063 26937
rect 11097 26903 11223 26937
rect 11257 26903 11383 26937
rect 11417 26903 11440 26937
rect 9440 26880 11440 26903
rect 11520 26937 11920 26960
rect 11520 26903 11543 26937
rect 11577 26903 11703 26937
rect 11737 26903 11863 26937
rect 11897 26903 11920 26937
rect 11520 26880 11920 26903
rect 12000 26937 12400 26960
rect 12000 26903 12023 26937
rect 12057 26903 12183 26937
rect 12217 26903 12343 26937
rect 12377 26903 12400 26937
rect 12000 26880 12400 26903
rect 8480 26777 8880 26800
rect 8480 26743 8503 26777
rect 8537 26743 8663 26777
rect 8697 26743 8823 26777
rect 8857 26743 8880 26777
rect 8480 26720 8880 26743
rect 8960 26777 9360 26800
rect 8960 26743 8983 26777
rect 9017 26743 9143 26777
rect 9177 26743 9303 26777
rect 9337 26743 9360 26777
rect 8960 26720 9360 26743
rect 9440 26777 11440 26800
rect 9440 26743 9463 26777
rect 9497 26743 9623 26777
rect 9657 26743 9783 26777
rect 9817 26743 9943 26777
rect 9977 26743 10103 26777
rect 10137 26743 10263 26777
rect 10297 26743 10423 26777
rect 10457 26743 10583 26777
rect 10617 26743 10743 26777
rect 10777 26743 10903 26777
rect 10937 26743 11063 26777
rect 11097 26743 11223 26777
rect 11257 26743 11383 26777
rect 11417 26743 11440 26777
rect 9440 26720 11440 26743
rect 11520 26777 11920 26800
rect 11520 26743 11543 26777
rect 11577 26743 11703 26777
rect 11737 26743 11863 26777
rect 11897 26743 11920 26777
rect 11520 26720 11920 26743
rect 12000 26777 12400 26800
rect 12000 26743 12023 26777
rect 12057 26743 12183 26777
rect 12217 26743 12343 26777
rect 12377 26743 12400 26777
rect 12000 26720 12400 26743
rect 8480 26617 8880 26640
rect 8480 26583 8503 26617
rect 8537 26583 8663 26617
rect 8697 26583 8823 26617
rect 8857 26583 8880 26617
rect 8480 26560 8880 26583
rect 8960 26617 9360 26640
rect 8960 26583 8983 26617
rect 9017 26583 9143 26617
rect 9177 26583 9303 26617
rect 9337 26583 9360 26617
rect 8960 26560 9360 26583
rect 9440 26617 11440 26640
rect 9440 26583 9463 26617
rect 9497 26583 9623 26617
rect 9657 26583 9783 26617
rect 9817 26583 9943 26617
rect 9977 26583 10103 26617
rect 10137 26583 10263 26617
rect 10297 26583 10423 26617
rect 10457 26583 10583 26617
rect 10617 26583 10743 26617
rect 10777 26583 10903 26617
rect 10937 26583 11063 26617
rect 11097 26583 11223 26617
rect 11257 26583 11383 26617
rect 11417 26583 11440 26617
rect 9440 26560 11440 26583
rect 11520 26617 11920 26640
rect 11520 26583 11543 26617
rect 11577 26583 11703 26617
rect 11737 26583 11863 26617
rect 11897 26583 11920 26617
rect 11520 26560 11920 26583
rect 12000 26617 12400 26640
rect 12000 26583 12023 26617
rect 12057 26583 12183 26617
rect 12217 26583 12343 26617
rect 12377 26583 12400 26617
rect 12000 26560 12400 26583
rect 8480 26457 8880 26480
rect 8480 26423 8503 26457
rect 8537 26423 8663 26457
rect 8697 26423 8823 26457
rect 8857 26423 8880 26457
rect 8480 26400 8880 26423
rect 8960 26457 9360 26480
rect 8960 26423 8983 26457
rect 9017 26423 9143 26457
rect 9177 26423 9303 26457
rect 9337 26423 9360 26457
rect 8960 26400 9360 26423
rect 9440 26457 11440 26480
rect 9440 26423 9463 26457
rect 9497 26423 9623 26457
rect 9657 26423 9783 26457
rect 9817 26423 9943 26457
rect 9977 26423 10103 26457
rect 10137 26423 10263 26457
rect 10297 26423 10423 26457
rect 10457 26423 10583 26457
rect 10617 26423 10743 26457
rect 10777 26423 10903 26457
rect 10937 26423 11063 26457
rect 11097 26423 11223 26457
rect 11257 26423 11383 26457
rect 11417 26423 11440 26457
rect 9440 26400 11440 26423
rect 11520 26457 11920 26480
rect 11520 26423 11543 26457
rect 11577 26423 11703 26457
rect 11737 26423 11863 26457
rect 11897 26423 11920 26457
rect 11520 26400 11920 26423
rect 12000 26457 12400 26480
rect 12000 26423 12023 26457
rect 12057 26423 12183 26457
rect 12217 26423 12343 26457
rect 12377 26423 12400 26457
rect 12000 26400 12400 26423
rect 8480 26297 8880 26320
rect 8480 26263 8503 26297
rect 8537 26263 8663 26297
rect 8697 26263 8823 26297
rect 8857 26263 8880 26297
rect 8480 26240 8880 26263
rect 8960 26297 9360 26320
rect 8960 26263 8983 26297
rect 9017 26263 9143 26297
rect 9177 26263 9303 26297
rect 9337 26263 9360 26297
rect 8960 26240 9360 26263
rect 9440 26297 11440 26320
rect 9440 26263 9463 26297
rect 9497 26263 9623 26297
rect 9657 26263 9783 26297
rect 9817 26263 9943 26297
rect 9977 26263 10103 26297
rect 10137 26263 10263 26297
rect 10297 26263 10423 26297
rect 10457 26263 10583 26297
rect 10617 26263 10743 26297
rect 10777 26263 10903 26297
rect 10937 26263 11063 26297
rect 11097 26263 11223 26297
rect 11257 26263 11383 26297
rect 11417 26263 11440 26297
rect 9440 26240 11440 26263
rect 11520 26297 11920 26320
rect 11520 26263 11543 26297
rect 11577 26263 11703 26297
rect 11737 26263 11863 26297
rect 11897 26263 11920 26297
rect 11520 26240 11920 26263
rect 12000 26297 12400 26320
rect 12000 26263 12023 26297
rect 12057 26263 12183 26297
rect 12217 26263 12343 26297
rect 12377 26263 12400 26297
rect 12000 26240 12400 26263
rect 8480 26137 8880 26160
rect 8480 26103 8503 26137
rect 8537 26103 8663 26137
rect 8697 26103 8823 26137
rect 8857 26103 8880 26137
rect 8480 26080 8880 26103
rect 8960 26137 9360 26160
rect 8960 26103 8983 26137
rect 9017 26103 9143 26137
rect 9177 26103 9303 26137
rect 9337 26103 9360 26137
rect 8960 26080 9360 26103
rect 9440 26137 11440 26160
rect 9440 26103 9463 26137
rect 9497 26103 9623 26137
rect 9657 26103 9783 26137
rect 9817 26103 9943 26137
rect 9977 26103 10103 26137
rect 10137 26103 10263 26137
rect 10297 26103 10423 26137
rect 10457 26103 10583 26137
rect 10617 26103 10743 26137
rect 10777 26103 10903 26137
rect 10937 26103 11063 26137
rect 11097 26103 11223 26137
rect 11257 26103 11383 26137
rect 11417 26103 11440 26137
rect 9440 26080 11440 26103
rect 11520 26137 11920 26160
rect 11520 26103 11543 26137
rect 11577 26103 11703 26137
rect 11737 26103 11863 26137
rect 11897 26103 11920 26137
rect 11520 26080 11920 26103
rect 12000 26137 12400 26160
rect 12000 26103 12023 26137
rect 12057 26103 12183 26137
rect 12217 26103 12343 26137
rect 12377 26103 12400 26137
rect 12000 26080 12400 26103
rect 8480 25977 8880 26000
rect 8480 25943 8503 25977
rect 8537 25943 8663 25977
rect 8697 25943 8823 25977
rect 8857 25943 8880 25977
rect 8480 25920 8880 25943
rect 8960 25977 9360 26000
rect 8960 25943 8983 25977
rect 9017 25943 9143 25977
rect 9177 25943 9303 25977
rect 9337 25943 9360 25977
rect 8960 25920 9360 25943
rect 9440 25977 11440 26000
rect 9440 25943 9463 25977
rect 9497 25943 9623 25977
rect 9657 25943 9783 25977
rect 9817 25943 9943 25977
rect 9977 25943 10103 25977
rect 10137 25943 10263 25977
rect 10297 25943 10423 25977
rect 10457 25943 10583 25977
rect 10617 25943 10743 25977
rect 10777 25943 10903 25977
rect 10937 25943 11063 25977
rect 11097 25943 11223 25977
rect 11257 25943 11383 25977
rect 11417 25943 11440 25977
rect 9440 25920 11440 25943
rect 11520 25977 11920 26000
rect 11520 25943 11543 25977
rect 11577 25943 11703 25977
rect 11737 25943 11863 25977
rect 11897 25943 11920 25977
rect 11520 25920 11920 25943
rect 12000 25977 12400 26000
rect 12000 25943 12023 25977
rect 12057 25943 12183 25977
rect 12217 25943 12343 25977
rect 12377 25943 12400 25977
rect 12000 25920 12400 25943
rect 8480 25817 8880 25840
rect 8480 25783 8503 25817
rect 8537 25783 8663 25817
rect 8697 25783 8823 25817
rect 8857 25783 8880 25817
rect 8480 25760 8880 25783
rect 8960 25817 9360 25840
rect 8960 25783 8983 25817
rect 9017 25783 9143 25817
rect 9177 25783 9303 25817
rect 9337 25783 9360 25817
rect 8960 25760 9360 25783
rect 9440 25817 11440 25840
rect 9440 25783 9463 25817
rect 9497 25783 9623 25817
rect 9657 25783 9783 25817
rect 9817 25783 9943 25817
rect 9977 25783 10103 25817
rect 10137 25783 10263 25817
rect 10297 25783 10423 25817
rect 10457 25783 10583 25817
rect 10617 25783 10743 25817
rect 10777 25783 10903 25817
rect 10937 25783 11063 25817
rect 11097 25783 11223 25817
rect 11257 25783 11383 25817
rect 11417 25783 11440 25817
rect 9440 25760 11440 25783
rect 11520 25817 11920 25840
rect 11520 25783 11543 25817
rect 11577 25783 11703 25817
rect 11737 25783 11863 25817
rect 11897 25783 11920 25817
rect 11520 25760 11920 25783
rect 12000 25817 12400 25840
rect 12000 25783 12023 25817
rect 12057 25783 12183 25817
rect 12217 25783 12343 25817
rect 12377 25783 12400 25817
rect 12000 25760 12400 25783
rect 8480 25657 8880 25680
rect 8480 25623 8503 25657
rect 8537 25623 8663 25657
rect 8697 25623 8823 25657
rect 8857 25623 8880 25657
rect 8480 25600 8880 25623
rect 8960 25657 9360 25680
rect 8960 25623 8983 25657
rect 9017 25623 9143 25657
rect 9177 25623 9303 25657
rect 9337 25623 9360 25657
rect 8960 25600 9360 25623
rect 9440 25657 11440 25680
rect 9440 25623 9463 25657
rect 9497 25623 9623 25657
rect 9657 25623 9783 25657
rect 9817 25623 9943 25657
rect 9977 25623 10103 25657
rect 10137 25623 10263 25657
rect 10297 25623 10423 25657
rect 10457 25623 10583 25657
rect 10617 25623 10743 25657
rect 10777 25623 10903 25657
rect 10937 25623 11063 25657
rect 11097 25623 11223 25657
rect 11257 25623 11383 25657
rect 11417 25623 11440 25657
rect 9440 25600 11440 25623
rect 11520 25657 11920 25680
rect 11520 25623 11543 25657
rect 11577 25623 11703 25657
rect 11737 25623 11863 25657
rect 11897 25623 11920 25657
rect 11520 25600 11920 25623
rect 12000 25657 12400 25680
rect 12000 25623 12023 25657
rect 12057 25623 12183 25657
rect 12217 25623 12343 25657
rect 12377 25623 12400 25657
rect 12000 25600 12400 25623
rect 8480 25497 8880 25520
rect 8480 25463 8503 25497
rect 8537 25463 8663 25497
rect 8697 25463 8823 25497
rect 8857 25463 8880 25497
rect 8480 25440 8880 25463
rect 8960 25497 9360 25520
rect 8960 25463 8983 25497
rect 9017 25463 9143 25497
rect 9177 25463 9303 25497
rect 9337 25463 9360 25497
rect 8960 25440 9360 25463
rect 9440 25497 11440 25520
rect 9440 25463 9463 25497
rect 9497 25463 9623 25497
rect 9657 25463 9783 25497
rect 9817 25463 9943 25497
rect 9977 25463 10103 25497
rect 10137 25463 10263 25497
rect 10297 25463 10423 25497
rect 10457 25463 10583 25497
rect 10617 25463 10743 25497
rect 10777 25463 10903 25497
rect 10937 25463 11063 25497
rect 11097 25463 11223 25497
rect 11257 25463 11383 25497
rect 11417 25463 11440 25497
rect 9440 25440 11440 25463
rect 11520 25497 11920 25520
rect 11520 25463 11543 25497
rect 11577 25463 11703 25497
rect 11737 25463 11863 25497
rect 11897 25463 11920 25497
rect 11520 25440 11920 25463
rect 12000 25497 12400 25520
rect 12000 25463 12023 25497
rect 12057 25463 12183 25497
rect 12217 25463 12343 25497
rect 12377 25463 12400 25497
rect 12000 25440 12400 25463
rect 8480 25337 8880 25360
rect 8480 25303 8503 25337
rect 8537 25303 8663 25337
rect 8697 25303 8823 25337
rect 8857 25303 8880 25337
rect 8480 25280 8880 25303
rect 8960 25337 9360 25360
rect 8960 25303 8983 25337
rect 9017 25303 9143 25337
rect 9177 25303 9303 25337
rect 9337 25303 9360 25337
rect 8960 25280 9360 25303
rect 9440 25337 11440 25360
rect 9440 25303 9463 25337
rect 9497 25303 9623 25337
rect 9657 25303 9783 25337
rect 9817 25303 9943 25337
rect 9977 25303 10103 25337
rect 10137 25303 10263 25337
rect 10297 25303 10423 25337
rect 10457 25303 10583 25337
rect 10617 25303 10743 25337
rect 10777 25303 10903 25337
rect 10937 25303 11063 25337
rect 11097 25303 11223 25337
rect 11257 25303 11383 25337
rect 11417 25303 11440 25337
rect 9440 25280 11440 25303
rect 11520 25337 11920 25360
rect 11520 25303 11543 25337
rect 11577 25303 11703 25337
rect 11737 25303 11863 25337
rect 11897 25303 11920 25337
rect 11520 25280 11920 25303
rect 12000 25337 12400 25360
rect 12000 25303 12023 25337
rect 12057 25303 12183 25337
rect 12217 25303 12343 25337
rect 12377 25303 12400 25337
rect 12000 25280 12400 25303
rect 8480 25177 8880 25200
rect 8480 25143 8503 25177
rect 8537 25143 8663 25177
rect 8697 25143 8823 25177
rect 8857 25143 8880 25177
rect 8480 25120 8880 25143
rect 8960 25177 9360 25200
rect 8960 25143 8983 25177
rect 9017 25143 9143 25177
rect 9177 25143 9303 25177
rect 9337 25143 9360 25177
rect 8960 25120 9360 25143
rect 9440 25177 11440 25200
rect 9440 25143 9463 25177
rect 9497 25143 9623 25177
rect 9657 25143 9783 25177
rect 9817 25143 9943 25177
rect 9977 25143 10103 25177
rect 10137 25143 10263 25177
rect 10297 25143 10423 25177
rect 10457 25143 10583 25177
rect 10617 25143 10743 25177
rect 10777 25143 10903 25177
rect 10937 25143 11063 25177
rect 11097 25143 11223 25177
rect 11257 25143 11383 25177
rect 11417 25143 11440 25177
rect 9440 25120 11440 25143
rect 11520 25177 11920 25200
rect 11520 25143 11543 25177
rect 11577 25143 11703 25177
rect 11737 25143 11863 25177
rect 11897 25143 11920 25177
rect 11520 25120 11920 25143
rect 12000 25177 12400 25200
rect 12000 25143 12023 25177
rect 12057 25143 12183 25177
rect 12217 25143 12343 25177
rect 12377 25143 12400 25177
rect 12000 25120 12400 25143
rect 8480 25017 8880 25040
rect 8480 24983 8503 25017
rect 8537 24983 8663 25017
rect 8697 24983 8823 25017
rect 8857 24983 8880 25017
rect 8480 24960 8880 24983
rect 8960 25017 9360 25040
rect 8960 24983 8983 25017
rect 9017 24983 9143 25017
rect 9177 24983 9303 25017
rect 9337 24983 9360 25017
rect 8960 24960 9360 24983
rect 9440 25017 11440 25040
rect 9440 24983 9463 25017
rect 9497 24983 9623 25017
rect 9657 24983 9783 25017
rect 9817 24983 9943 25017
rect 9977 24983 10103 25017
rect 10137 24983 10263 25017
rect 10297 24983 10423 25017
rect 10457 24983 10583 25017
rect 10617 24983 10743 25017
rect 10777 24983 10903 25017
rect 10937 24983 11063 25017
rect 11097 24983 11223 25017
rect 11257 24983 11383 25017
rect 11417 24983 11440 25017
rect 9440 24960 11440 24983
rect 11520 25017 11920 25040
rect 11520 24983 11543 25017
rect 11577 24983 11703 25017
rect 11737 24983 11863 25017
rect 11897 24983 11920 25017
rect 11520 24960 11920 24983
rect 12000 25017 12400 25040
rect 12000 24983 12023 25017
rect 12057 24983 12183 25017
rect 12217 24983 12343 25017
rect 12377 24983 12400 25017
rect 12000 24960 12400 24983
rect 8480 24857 8880 24880
rect 8480 24823 8503 24857
rect 8537 24823 8663 24857
rect 8697 24823 8823 24857
rect 8857 24823 8880 24857
rect 8480 24800 8880 24823
rect 8960 24857 9360 24880
rect 8960 24823 8983 24857
rect 9017 24823 9143 24857
rect 9177 24823 9303 24857
rect 9337 24823 9360 24857
rect 8960 24800 9360 24823
rect 9440 24857 11440 24880
rect 9440 24823 9463 24857
rect 9497 24823 9623 24857
rect 9657 24823 9783 24857
rect 9817 24823 9943 24857
rect 9977 24823 10103 24857
rect 10137 24823 10263 24857
rect 10297 24823 10423 24857
rect 10457 24823 10583 24857
rect 10617 24823 10743 24857
rect 10777 24823 10903 24857
rect 10937 24823 11063 24857
rect 11097 24823 11223 24857
rect 11257 24823 11383 24857
rect 11417 24823 11440 24857
rect 9440 24800 11440 24823
rect 11520 24857 11920 24880
rect 11520 24823 11543 24857
rect 11577 24823 11703 24857
rect 11737 24823 11863 24857
rect 11897 24823 11920 24857
rect 11520 24800 11920 24823
rect 12000 24857 12400 24880
rect 12000 24823 12023 24857
rect 12057 24823 12183 24857
rect 12217 24823 12343 24857
rect 12377 24823 12400 24857
rect 12000 24800 12400 24823
rect 8480 24697 8880 24720
rect 8480 24663 8503 24697
rect 8537 24663 8663 24697
rect 8697 24663 8823 24697
rect 8857 24663 8880 24697
rect 8480 24640 8880 24663
rect 8960 24697 9360 24720
rect 8960 24663 8983 24697
rect 9017 24663 9143 24697
rect 9177 24663 9303 24697
rect 9337 24663 9360 24697
rect 8960 24640 9360 24663
rect 9440 24697 11440 24720
rect 9440 24663 9463 24697
rect 9497 24663 9623 24697
rect 9657 24663 9783 24697
rect 9817 24663 9943 24697
rect 9977 24663 10103 24697
rect 10137 24663 10263 24697
rect 10297 24663 10423 24697
rect 10457 24663 10583 24697
rect 10617 24663 10743 24697
rect 10777 24663 10903 24697
rect 10937 24663 11063 24697
rect 11097 24663 11223 24697
rect 11257 24663 11383 24697
rect 11417 24663 11440 24697
rect 9440 24640 11440 24663
rect 11520 24697 11920 24720
rect 11520 24663 11543 24697
rect 11577 24663 11703 24697
rect 11737 24663 11863 24697
rect 11897 24663 11920 24697
rect 11520 24640 11920 24663
rect 12000 24697 12400 24720
rect 12000 24663 12023 24697
rect 12057 24663 12183 24697
rect 12217 24663 12343 24697
rect 12377 24663 12400 24697
rect 12000 24640 12400 24663
rect 8480 24537 8880 24560
rect 8480 24503 8503 24537
rect 8537 24503 8663 24537
rect 8697 24503 8823 24537
rect 8857 24503 8880 24537
rect 8480 24480 8880 24503
rect 8960 24537 9360 24560
rect 8960 24503 8983 24537
rect 9017 24503 9143 24537
rect 9177 24503 9303 24537
rect 9337 24503 9360 24537
rect 8960 24480 9360 24503
rect 9440 24537 11440 24560
rect 9440 24503 9463 24537
rect 9497 24503 9623 24537
rect 9657 24503 9783 24537
rect 9817 24503 9943 24537
rect 9977 24503 10103 24537
rect 10137 24503 10263 24537
rect 10297 24503 10423 24537
rect 10457 24503 10583 24537
rect 10617 24503 10743 24537
rect 10777 24503 10903 24537
rect 10937 24503 11063 24537
rect 11097 24503 11223 24537
rect 11257 24503 11383 24537
rect 11417 24503 11440 24537
rect 9440 24480 11440 24503
rect 11520 24537 11920 24560
rect 11520 24503 11543 24537
rect 11577 24503 11703 24537
rect 11737 24503 11863 24537
rect 11897 24503 11920 24537
rect 11520 24480 11920 24503
rect 12000 24537 12400 24560
rect 12000 24503 12023 24537
rect 12057 24503 12183 24537
rect 12217 24503 12343 24537
rect 12377 24503 12400 24537
rect 12000 24480 12400 24503
rect 8480 24377 8880 24400
rect 8480 24343 8503 24377
rect 8537 24343 8663 24377
rect 8697 24343 8823 24377
rect 8857 24343 8880 24377
rect 8480 24320 8880 24343
rect 8960 24377 9360 24400
rect 8960 24343 8983 24377
rect 9017 24343 9143 24377
rect 9177 24343 9303 24377
rect 9337 24343 9360 24377
rect 8960 24320 9360 24343
rect 9440 24377 11440 24400
rect 9440 24343 9463 24377
rect 9497 24343 9623 24377
rect 9657 24343 9783 24377
rect 9817 24343 9943 24377
rect 9977 24343 10103 24377
rect 10137 24343 10263 24377
rect 10297 24343 10423 24377
rect 10457 24343 10583 24377
rect 10617 24343 10743 24377
rect 10777 24343 10903 24377
rect 10937 24343 11063 24377
rect 11097 24343 11223 24377
rect 11257 24343 11383 24377
rect 11417 24343 11440 24377
rect 9440 24320 11440 24343
rect 11520 24377 11920 24400
rect 11520 24343 11543 24377
rect 11577 24343 11703 24377
rect 11737 24343 11863 24377
rect 11897 24343 11920 24377
rect 11520 24320 11920 24343
rect 12000 24377 12400 24400
rect 12000 24343 12023 24377
rect 12057 24343 12183 24377
rect 12217 24343 12343 24377
rect 12377 24343 12400 24377
rect 12000 24320 12400 24343
rect 8480 24217 8880 24240
rect 8480 24183 8503 24217
rect 8537 24183 8663 24217
rect 8697 24183 8823 24217
rect 8857 24183 8880 24217
rect 8480 24160 8880 24183
rect 8960 24217 9360 24240
rect 8960 24183 8983 24217
rect 9017 24183 9143 24217
rect 9177 24183 9303 24217
rect 9337 24183 9360 24217
rect 8960 24160 9360 24183
rect 9440 24217 11440 24240
rect 9440 24183 9463 24217
rect 9497 24183 9623 24217
rect 9657 24183 9783 24217
rect 9817 24183 9943 24217
rect 9977 24183 10103 24217
rect 10137 24183 10263 24217
rect 10297 24183 10423 24217
rect 10457 24183 10583 24217
rect 10617 24183 10743 24217
rect 10777 24183 10903 24217
rect 10937 24183 11063 24217
rect 11097 24183 11223 24217
rect 11257 24183 11383 24217
rect 11417 24183 11440 24217
rect 9440 24160 11440 24183
rect 11520 24217 11920 24240
rect 11520 24183 11543 24217
rect 11577 24183 11703 24217
rect 11737 24183 11863 24217
rect 11897 24183 11920 24217
rect 11520 24160 11920 24183
rect 12000 24217 12400 24240
rect 12000 24183 12023 24217
rect 12057 24183 12183 24217
rect 12217 24183 12343 24217
rect 12377 24183 12400 24217
rect 12000 24160 12400 24183
rect 8480 24057 8880 24080
rect 8480 24023 8503 24057
rect 8537 24023 8663 24057
rect 8697 24023 8823 24057
rect 8857 24023 8880 24057
rect 8480 24000 8880 24023
rect 8960 24057 9360 24080
rect 8960 24023 8983 24057
rect 9017 24023 9143 24057
rect 9177 24023 9303 24057
rect 9337 24023 9360 24057
rect 8960 24000 9360 24023
rect 9440 24057 11440 24080
rect 9440 24023 9463 24057
rect 9497 24023 9623 24057
rect 9657 24023 9783 24057
rect 9817 24023 9943 24057
rect 9977 24023 10103 24057
rect 10137 24023 10263 24057
rect 10297 24023 10423 24057
rect 10457 24023 10583 24057
rect 10617 24023 10743 24057
rect 10777 24023 10903 24057
rect 10937 24023 11063 24057
rect 11097 24023 11223 24057
rect 11257 24023 11383 24057
rect 11417 24023 11440 24057
rect 9440 24000 11440 24023
rect 11520 24057 11920 24080
rect 11520 24023 11543 24057
rect 11577 24023 11703 24057
rect 11737 24023 11863 24057
rect 11897 24023 11920 24057
rect 11520 24000 11920 24023
rect 12000 24057 12400 24080
rect 12000 24023 12023 24057
rect 12057 24023 12183 24057
rect 12217 24023 12343 24057
rect 12377 24023 12400 24057
rect 12000 24000 12400 24023
rect 8480 23897 8880 23920
rect 8480 23863 8503 23897
rect 8537 23863 8663 23897
rect 8697 23863 8823 23897
rect 8857 23863 8880 23897
rect 8480 23840 8880 23863
rect 8960 23897 9360 23920
rect 8960 23863 8983 23897
rect 9017 23863 9143 23897
rect 9177 23863 9303 23897
rect 9337 23863 9360 23897
rect 8960 23840 9360 23863
rect 9440 23897 11440 23920
rect 9440 23863 9463 23897
rect 9497 23863 9623 23897
rect 9657 23863 9783 23897
rect 9817 23863 9943 23897
rect 9977 23863 10103 23897
rect 10137 23863 10263 23897
rect 10297 23863 10423 23897
rect 10457 23863 10583 23897
rect 10617 23863 10743 23897
rect 10777 23863 10903 23897
rect 10937 23863 11063 23897
rect 11097 23863 11223 23897
rect 11257 23863 11383 23897
rect 11417 23863 11440 23897
rect 9440 23840 11440 23863
rect 11520 23897 11920 23920
rect 11520 23863 11543 23897
rect 11577 23863 11703 23897
rect 11737 23863 11863 23897
rect 11897 23863 11920 23897
rect 11520 23840 11920 23863
rect 12000 23897 12400 23920
rect 12000 23863 12023 23897
rect 12057 23863 12183 23897
rect 12217 23863 12343 23897
rect 12377 23863 12400 23897
rect 12000 23840 12400 23863
rect 8480 23737 8880 23760
rect 8480 23703 8503 23737
rect 8537 23703 8663 23737
rect 8697 23703 8823 23737
rect 8857 23703 8880 23737
rect 8480 23680 8880 23703
rect 8960 23737 9360 23760
rect 8960 23703 8983 23737
rect 9017 23703 9143 23737
rect 9177 23703 9303 23737
rect 9337 23703 9360 23737
rect 8960 23680 9360 23703
rect 9440 23737 11440 23760
rect 9440 23703 9463 23737
rect 9497 23703 9623 23737
rect 9657 23703 9783 23737
rect 9817 23703 9943 23737
rect 9977 23703 10103 23737
rect 10137 23703 10263 23737
rect 10297 23703 10423 23737
rect 10457 23703 10583 23737
rect 10617 23703 10743 23737
rect 10777 23703 10903 23737
rect 10937 23703 11063 23737
rect 11097 23703 11223 23737
rect 11257 23703 11383 23737
rect 11417 23703 11440 23737
rect 9440 23680 11440 23703
rect 11520 23737 11920 23760
rect 11520 23703 11543 23737
rect 11577 23703 11703 23737
rect 11737 23703 11863 23737
rect 11897 23703 11920 23737
rect 11520 23680 11920 23703
rect 12000 23737 12400 23760
rect 12000 23703 12023 23737
rect 12057 23703 12183 23737
rect 12217 23703 12343 23737
rect 12377 23703 12400 23737
rect 12000 23680 12400 23703
rect 8480 23577 8880 23600
rect 8480 23543 8503 23577
rect 8537 23543 8663 23577
rect 8697 23543 8823 23577
rect 8857 23543 8880 23577
rect 8480 23520 8880 23543
rect 8960 23577 9360 23600
rect 8960 23543 8983 23577
rect 9017 23543 9143 23577
rect 9177 23543 9303 23577
rect 9337 23543 9360 23577
rect 8960 23520 9360 23543
rect 9440 23577 11440 23600
rect 9440 23543 9463 23577
rect 9497 23543 9623 23577
rect 9657 23543 9783 23577
rect 9817 23543 9943 23577
rect 9977 23543 10103 23577
rect 10137 23543 10263 23577
rect 10297 23543 10423 23577
rect 10457 23543 10583 23577
rect 10617 23543 10743 23577
rect 10777 23543 10903 23577
rect 10937 23543 11063 23577
rect 11097 23543 11223 23577
rect 11257 23543 11383 23577
rect 11417 23543 11440 23577
rect 9440 23520 11440 23543
rect 11520 23577 11920 23600
rect 11520 23543 11543 23577
rect 11577 23543 11703 23577
rect 11737 23543 11863 23577
rect 11897 23543 11920 23577
rect 11520 23520 11920 23543
rect 12000 23577 12400 23600
rect 12000 23543 12023 23577
rect 12057 23543 12183 23577
rect 12217 23543 12343 23577
rect 12377 23543 12400 23577
rect 12000 23520 12400 23543
rect 8480 23417 8880 23440
rect 8480 23383 8503 23417
rect 8537 23383 8663 23417
rect 8697 23383 8823 23417
rect 8857 23383 8880 23417
rect 8480 23360 8880 23383
rect 8960 23417 9360 23440
rect 8960 23383 8983 23417
rect 9017 23383 9143 23417
rect 9177 23383 9303 23417
rect 9337 23383 9360 23417
rect 8960 23360 9360 23383
rect 9440 23417 11440 23440
rect 9440 23383 9463 23417
rect 9497 23383 9623 23417
rect 9657 23383 9783 23417
rect 9817 23383 9943 23417
rect 9977 23383 10103 23417
rect 10137 23383 10263 23417
rect 10297 23383 10423 23417
rect 10457 23383 10583 23417
rect 10617 23383 10743 23417
rect 10777 23383 10903 23417
rect 10937 23383 11063 23417
rect 11097 23383 11223 23417
rect 11257 23383 11383 23417
rect 11417 23383 11440 23417
rect 9440 23360 11440 23383
rect 11520 23417 11920 23440
rect 11520 23383 11543 23417
rect 11577 23383 11703 23417
rect 11737 23383 11863 23417
rect 11897 23383 11920 23417
rect 11520 23360 11920 23383
rect 12000 23417 12400 23440
rect 12000 23383 12023 23417
rect 12057 23383 12183 23417
rect 12217 23383 12343 23417
rect 12377 23383 12400 23417
rect 12000 23360 12400 23383
rect 8480 23257 8880 23280
rect 8480 23223 8503 23257
rect 8537 23223 8663 23257
rect 8697 23223 8823 23257
rect 8857 23223 8880 23257
rect 8480 23200 8880 23223
rect 8960 23257 9360 23280
rect 8960 23223 8983 23257
rect 9017 23223 9143 23257
rect 9177 23223 9303 23257
rect 9337 23223 9360 23257
rect 8960 23200 9360 23223
rect 9440 23257 11440 23280
rect 9440 23223 9463 23257
rect 9497 23223 9623 23257
rect 9657 23223 9783 23257
rect 9817 23223 9943 23257
rect 9977 23223 10103 23257
rect 10137 23223 10263 23257
rect 10297 23223 10423 23257
rect 10457 23223 10583 23257
rect 10617 23223 10743 23257
rect 10777 23223 10903 23257
rect 10937 23223 11063 23257
rect 11097 23223 11223 23257
rect 11257 23223 11383 23257
rect 11417 23223 11440 23257
rect 9440 23200 11440 23223
rect 11520 23257 11920 23280
rect 11520 23223 11543 23257
rect 11577 23223 11703 23257
rect 11737 23223 11863 23257
rect 11897 23223 11920 23257
rect 11520 23200 11920 23223
rect 12000 23257 12400 23280
rect 12000 23223 12023 23257
rect 12057 23223 12183 23257
rect 12217 23223 12343 23257
rect 12377 23223 12400 23257
rect 12000 23200 12400 23223
rect 8480 23097 8880 23120
rect 8480 23063 8503 23097
rect 8537 23063 8663 23097
rect 8697 23063 8823 23097
rect 8857 23063 8880 23097
rect 8480 23040 8880 23063
rect 8960 23097 9360 23120
rect 8960 23063 8983 23097
rect 9017 23063 9143 23097
rect 9177 23063 9303 23097
rect 9337 23063 9360 23097
rect 8960 23040 9360 23063
rect 9440 23097 11440 23120
rect 9440 23063 9463 23097
rect 9497 23063 9623 23097
rect 9657 23063 9783 23097
rect 9817 23063 9943 23097
rect 9977 23063 10103 23097
rect 10137 23063 10263 23097
rect 10297 23063 10423 23097
rect 10457 23063 10583 23097
rect 10617 23063 10743 23097
rect 10777 23063 10903 23097
rect 10937 23063 11063 23097
rect 11097 23063 11223 23097
rect 11257 23063 11383 23097
rect 11417 23063 11440 23097
rect 9440 23040 11440 23063
rect 11520 23097 11920 23120
rect 11520 23063 11543 23097
rect 11577 23063 11703 23097
rect 11737 23063 11863 23097
rect 11897 23063 11920 23097
rect 11520 23040 11920 23063
rect 12000 23097 12400 23120
rect 12000 23063 12023 23097
rect 12057 23063 12183 23097
rect 12217 23063 12343 23097
rect 12377 23063 12400 23097
rect 12000 23040 12400 23063
rect 8480 22937 8880 22960
rect 8480 22903 8503 22937
rect 8537 22903 8663 22937
rect 8697 22903 8823 22937
rect 8857 22903 8880 22937
rect 8480 22880 8880 22903
rect 8960 22937 9360 22960
rect 8960 22903 8983 22937
rect 9017 22903 9143 22937
rect 9177 22903 9303 22937
rect 9337 22903 9360 22937
rect 8960 22880 9360 22903
rect 9440 22937 11440 22960
rect 9440 22903 9463 22937
rect 9497 22903 9623 22937
rect 9657 22903 9783 22937
rect 9817 22903 9943 22937
rect 9977 22903 10103 22937
rect 10137 22903 10263 22937
rect 10297 22903 10423 22937
rect 10457 22903 10583 22937
rect 10617 22903 10743 22937
rect 10777 22903 10903 22937
rect 10937 22903 11063 22937
rect 11097 22903 11223 22937
rect 11257 22903 11383 22937
rect 11417 22903 11440 22937
rect 9440 22880 11440 22903
rect 11520 22937 11920 22960
rect 11520 22903 11543 22937
rect 11577 22903 11703 22937
rect 11737 22903 11863 22937
rect 11897 22903 11920 22937
rect 11520 22880 11920 22903
rect 12000 22937 12400 22960
rect 12000 22903 12023 22937
rect 12057 22903 12183 22937
rect 12217 22903 12343 22937
rect 12377 22903 12400 22937
rect 12000 22880 12400 22903
rect 8480 22777 8880 22800
rect 8480 22743 8503 22777
rect 8537 22743 8663 22777
rect 8697 22743 8823 22777
rect 8857 22743 8880 22777
rect 8480 22720 8880 22743
rect 8960 22777 9360 22800
rect 8960 22743 8983 22777
rect 9017 22743 9143 22777
rect 9177 22743 9303 22777
rect 9337 22743 9360 22777
rect 8960 22720 9360 22743
rect 9440 22777 11440 22800
rect 9440 22743 9463 22777
rect 9497 22743 9623 22777
rect 9657 22743 9783 22777
rect 9817 22743 9943 22777
rect 9977 22743 10103 22777
rect 10137 22743 10263 22777
rect 10297 22743 10423 22777
rect 10457 22743 10583 22777
rect 10617 22743 10743 22777
rect 10777 22743 10903 22777
rect 10937 22743 11063 22777
rect 11097 22743 11223 22777
rect 11257 22743 11383 22777
rect 11417 22743 11440 22777
rect 9440 22720 11440 22743
rect 11520 22777 11920 22800
rect 11520 22743 11543 22777
rect 11577 22743 11703 22777
rect 11737 22743 11863 22777
rect 11897 22743 11920 22777
rect 11520 22720 11920 22743
rect 12000 22777 12400 22800
rect 12000 22743 12023 22777
rect 12057 22743 12183 22777
rect 12217 22743 12343 22777
rect 12377 22743 12400 22777
rect 12000 22720 12400 22743
rect 8480 22617 8880 22640
rect 8480 22583 8503 22617
rect 8537 22583 8663 22617
rect 8697 22583 8823 22617
rect 8857 22583 8880 22617
rect 8480 22560 8880 22583
rect 8960 22617 9360 22640
rect 8960 22583 8983 22617
rect 9017 22583 9143 22617
rect 9177 22583 9303 22617
rect 9337 22583 9360 22617
rect 8960 22560 9360 22583
rect 9440 22617 11440 22640
rect 9440 22583 9463 22617
rect 9497 22583 9623 22617
rect 9657 22583 9783 22617
rect 9817 22583 9943 22617
rect 9977 22583 10103 22617
rect 10137 22583 10263 22617
rect 10297 22583 10423 22617
rect 10457 22583 10583 22617
rect 10617 22583 10743 22617
rect 10777 22583 10903 22617
rect 10937 22583 11063 22617
rect 11097 22583 11223 22617
rect 11257 22583 11383 22617
rect 11417 22583 11440 22617
rect 9440 22560 11440 22583
rect 11520 22617 11920 22640
rect 11520 22583 11543 22617
rect 11577 22583 11703 22617
rect 11737 22583 11863 22617
rect 11897 22583 11920 22617
rect 11520 22560 11920 22583
rect 12000 22617 12400 22640
rect 12000 22583 12023 22617
rect 12057 22583 12183 22617
rect 12217 22583 12343 22617
rect 12377 22583 12400 22617
rect 12000 22560 12400 22583
rect 8480 22457 8880 22480
rect 8480 22423 8503 22457
rect 8537 22423 8663 22457
rect 8697 22423 8823 22457
rect 8857 22423 8880 22457
rect 8480 22400 8880 22423
rect 8960 22457 9360 22480
rect 8960 22423 8983 22457
rect 9017 22423 9143 22457
rect 9177 22423 9303 22457
rect 9337 22423 9360 22457
rect 8960 22400 9360 22423
rect 9440 22457 11440 22480
rect 9440 22423 9463 22457
rect 9497 22423 9623 22457
rect 9657 22423 9783 22457
rect 9817 22423 9943 22457
rect 9977 22423 10103 22457
rect 10137 22423 10263 22457
rect 10297 22423 10423 22457
rect 10457 22423 10583 22457
rect 10617 22423 10743 22457
rect 10777 22423 10903 22457
rect 10937 22423 11063 22457
rect 11097 22423 11223 22457
rect 11257 22423 11383 22457
rect 11417 22423 11440 22457
rect 9440 22400 11440 22423
rect 11520 22457 11920 22480
rect 11520 22423 11543 22457
rect 11577 22423 11703 22457
rect 11737 22423 11863 22457
rect 11897 22423 11920 22457
rect 11520 22400 11920 22423
rect 12000 22457 12400 22480
rect 12000 22423 12023 22457
rect 12057 22423 12183 22457
rect 12217 22423 12343 22457
rect 12377 22423 12400 22457
rect 12000 22400 12400 22423
rect 8480 22297 8880 22320
rect 8480 22263 8503 22297
rect 8537 22263 8663 22297
rect 8697 22263 8823 22297
rect 8857 22263 8880 22297
rect 8480 22240 8880 22263
rect 8960 22297 9360 22320
rect 8960 22263 8983 22297
rect 9017 22263 9143 22297
rect 9177 22263 9303 22297
rect 9337 22263 9360 22297
rect 8960 22240 9360 22263
rect 9440 22297 11440 22320
rect 9440 22263 9463 22297
rect 9497 22263 9623 22297
rect 9657 22263 9783 22297
rect 9817 22263 9943 22297
rect 9977 22263 10103 22297
rect 10137 22263 10263 22297
rect 10297 22263 10423 22297
rect 10457 22263 10583 22297
rect 10617 22263 10743 22297
rect 10777 22263 10903 22297
rect 10937 22263 11063 22297
rect 11097 22263 11223 22297
rect 11257 22263 11383 22297
rect 11417 22263 11440 22297
rect 9440 22240 11440 22263
rect 11520 22297 11920 22320
rect 11520 22263 11543 22297
rect 11577 22263 11703 22297
rect 11737 22263 11863 22297
rect 11897 22263 11920 22297
rect 11520 22240 11920 22263
rect 12000 22297 12400 22320
rect 12000 22263 12023 22297
rect 12057 22263 12183 22297
rect 12217 22263 12343 22297
rect 12377 22263 12400 22297
rect 12000 22240 12400 22263
rect 8480 22137 8880 22160
rect 8480 22103 8503 22137
rect 8537 22103 8663 22137
rect 8697 22103 8823 22137
rect 8857 22103 8880 22137
rect 8480 22080 8880 22103
rect 8960 22137 9360 22160
rect 8960 22103 8983 22137
rect 9017 22103 9143 22137
rect 9177 22103 9303 22137
rect 9337 22103 9360 22137
rect 8960 22080 9360 22103
rect 9440 22137 11440 22160
rect 9440 22103 9463 22137
rect 9497 22103 9623 22137
rect 9657 22103 9783 22137
rect 9817 22103 9943 22137
rect 9977 22103 10103 22137
rect 10137 22103 10263 22137
rect 10297 22103 10423 22137
rect 10457 22103 10583 22137
rect 10617 22103 10743 22137
rect 10777 22103 10903 22137
rect 10937 22103 11063 22137
rect 11097 22103 11223 22137
rect 11257 22103 11383 22137
rect 11417 22103 11440 22137
rect 9440 22080 11440 22103
rect 11520 22137 11920 22160
rect 11520 22103 11543 22137
rect 11577 22103 11703 22137
rect 11737 22103 11863 22137
rect 11897 22103 11920 22137
rect 11520 22080 11920 22103
rect 12000 22137 12400 22160
rect 12000 22103 12023 22137
rect 12057 22103 12183 22137
rect 12217 22103 12343 22137
rect 12377 22103 12400 22137
rect 12000 22080 12400 22103
rect 8480 21977 8880 22000
rect 8480 21943 8503 21977
rect 8537 21943 8663 21977
rect 8697 21943 8823 21977
rect 8857 21943 8880 21977
rect 8480 21920 8880 21943
rect 8960 21977 9360 22000
rect 8960 21943 8983 21977
rect 9017 21943 9143 21977
rect 9177 21943 9303 21977
rect 9337 21943 9360 21977
rect 8960 21920 9360 21943
rect 9440 21977 11440 22000
rect 9440 21943 9463 21977
rect 9497 21943 9623 21977
rect 9657 21943 9783 21977
rect 9817 21943 9943 21977
rect 9977 21943 10103 21977
rect 10137 21943 10263 21977
rect 10297 21943 10423 21977
rect 10457 21943 10583 21977
rect 10617 21943 10743 21977
rect 10777 21943 10903 21977
rect 10937 21943 11063 21977
rect 11097 21943 11223 21977
rect 11257 21943 11383 21977
rect 11417 21943 11440 21977
rect 9440 21920 11440 21943
rect 11520 21977 11920 22000
rect 11520 21943 11543 21977
rect 11577 21943 11703 21977
rect 11737 21943 11863 21977
rect 11897 21943 11920 21977
rect 11520 21920 11920 21943
rect 12000 21977 12400 22000
rect 12000 21943 12023 21977
rect 12057 21943 12183 21977
rect 12217 21943 12343 21977
rect 12377 21943 12400 21977
rect 12000 21920 12400 21943
rect 8480 21817 8880 21840
rect 8480 21783 8503 21817
rect 8537 21783 8663 21817
rect 8697 21783 8823 21817
rect 8857 21783 8880 21817
rect 8480 21760 8880 21783
rect 8960 21817 9360 21840
rect 8960 21783 8983 21817
rect 9017 21783 9143 21817
rect 9177 21783 9303 21817
rect 9337 21783 9360 21817
rect 8960 21760 9360 21783
rect 9440 21817 11440 21840
rect 9440 21783 9463 21817
rect 9497 21783 9623 21817
rect 9657 21783 9783 21817
rect 9817 21783 9943 21817
rect 9977 21783 10103 21817
rect 10137 21783 10263 21817
rect 10297 21783 10423 21817
rect 10457 21783 10583 21817
rect 10617 21783 10743 21817
rect 10777 21783 10903 21817
rect 10937 21783 11063 21817
rect 11097 21783 11223 21817
rect 11257 21783 11383 21817
rect 11417 21783 11440 21817
rect 9440 21760 11440 21783
rect 11520 21817 11920 21840
rect 11520 21783 11543 21817
rect 11577 21783 11703 21817
rect 11737 21783 11863 21817
rect 11897 21783 11920 21817
rect 11520 21760 11920 21783
rect 12000 21817 12400 21840
rect 12000 21783 12023 21817
rect 12057 21783 12183 21817
rect 12217 21783 12343 21817
rect 12377 21783 12400 21817
rect 12000 21760 12400 21783
rect 8480 21657 8880 21680
rect 8480 21623 8503 21657
rect 8537 21623 8663 21657
rect 8697 21623 8823 21657
rect 8857 21623 8880 21657
rect 8480 21600 8880 21623
rect 8960 21657 9360 21680
rect 8960 21623 8983 21657
rect 9017 21623 9143 21657
rect 9177 21623 9303 21657
rect 9337 21623 9360 21657
rect 8960 21600 9360 21623
rect 9440 21657 11440 21680
rect 9440 21623 9463 21657
rect 9497 21623 9623 21657
rect 9657 21623 9783 21657
rect 9817 21623 9943 21657
rect 9977 21623 10103 21657
rect 10137 21623 10263 21657
rect 10297 21623 10423 21657
rect 10457 21623 10583 21657
rect 10617 21623 10743 21657
rect 10777 21623 10903 21657
rect 10937 21623 11063 21657
rect 11097 21623 11223 21657
rect 11257 21623 11383 21657
rect 11417 21623 11440 21657
rect 9440 21600 11440 21623
rect 11520 21657 11920 21680
rect 11520 21623 11543 21657
rect 11577 21623 11703 21657
rect 11737 21623 11863 21657
rect 11897 21623 11920 21657
rect 11520 21600 11920 21623
rect 12000 21657 12400 21680
rect 12000 21623 12023 21657
rect 12057 21623 12183 21657
rect 12217 21623 12343 21657
rect 12377 21623 12400 21657
rect 12000 21600 12400 21623
rect 8480 21497 8880 21520
rect 8480 21463 8503 21497
rect 8537 21463 8663 21497
rect 8697 21463 8823 21497
rect 8857 21463 8880 21497
rect 8480 21440 8880 21463
rect 8960 21497 9360 21520
rect 8960 21463 8983 21497
rect 9017 21463 9143 21497
rect 9177 21463 9303 21497
rect 9337 21463 9360 21497
rect 8960 21440 9360 21463
rect 9440 21497 11440 21520
rect 9440 21463 9463 21497
rect 9497 21463 9623 21497
rect 9657 21463 9783 21497
rect 9817 21463 9943 21497
rect 9977 21463 10103 21497
rect 10137 21463 10263 21497
rect 10297 21463 10423 21497
rect 10457 21463 10583 21497
rect 10617 21463 10743 21497
rect 10777 21463 10903 21497
rect 10937 21463 11063 21497
rect 11097 21463 11223 21497
rect 11257 21463 11383 21497
rect 11417 21463 11440 21497
rect 9440 21440 11440 21463
rect 11520 21497 11920 21520
rect 11520 21463 11543 21497
rect 11577 21463 11703 21497
rect 11737 21463 11863 21497
rect 11897 21463 11920 21497
rect 11520 21440 11920 21463
rect 12000 21497 12400 21520
rect 12000 21463 12023 21497
rect 12057 21463 12183 21497
rect 12217 21463 12343 21497
rect 12377 21463 12400 21497
rect 12000 21440 12400 21463
rect 8480 21337 8880 21360
rect 8480 21303 8503 21337
rect 8537 21303 8663 21337
rect 8697 21303 8823 21337
rect 8857 21303 8880 21337
rect 8480 21280 8880 21303
rect 8960 21337 9360 21360
rect 8960 21303 8983 21337
rect 9017 21303 9143 21337
rect 9177 21303 9303 21337
rect 9337 21303 9360 21337
rect 8960 21280 9360 21303
rect 9440 21337 11440 21360
rect 9440 21303 9463 21337
rect 9497 21303 9623 21337
rect 9657 21303 9783 21337
rect 9817 21303 9943 21337
rect 9977 21303 10103 21337
rect 10137 21303 10263 21337
rect 10297 21303 10423 21337
rect 10457 21303 10583 21337
rect 10617 21303 10743 21337
rect 10777 21303 10903 21337
rect 10937 21303 11063 21337
rect 11097 21303 11223 21337
rect 11257 21303 11383 21337
rect 11417 21303 11440 21337
rect 9440 21280 11440 21303
rect 11520 21337 11920 21360
rect 11520 21303 11543 21337
rect 11577 21303 11703 21337
rect 11737 21303 11863 21337
rect 11897 21303 11920 21337
rect 11520 21280 11920 21303
rect 12000 21337 12400 21360
rect 12000 21303 12023 21337
rect 12057 21303 12183 21337
rect 12217 21303 12343 21337
rect 12377 21303 12400 21337
rect 12000 21280 12400 21303
rect 8480 21177 8880 21200
rect 8480 21143 8503 21177
rect 8537 21143 8663 21177
rect 8697 21143 8823 21177
rect 8857 21143 8880 21177
rect 8480 21120 8880 21143
rect 8960 21177 9360 21200
rect 8960 21143 8983 21177
rect 9017 21143 9143 21177
rect 9177 21143 9303 21177
rect 9337 21143 9360 21177
rect 8960 21120 9360 21143
rect 9440 21177 11440 21200
rect 9440 21143 9463 21177
rect 9497 21143 9623 21177
rect 9657 21143 9783 21177
rect 9817 21143 9943 21177
rect 9977 21143 10103 21177
rect 10137 21143 10263 21177
rect 10297 21143 10423 21177
rect 10457 21143 10583 21177
rect 10617 21143 10743 21177
rect 10777 21143 10903 21177
rect 10937 21143 11063 21177
rect 11097 21143 11223 21177
rect 11257 21143 11383 21177
rect 11417 21143 11440 21177
rect 9440 21120 11440 21143
rect 11520 21177 11920 21200
rect 11520 21143 11543 21177
rect 11577 21143 11703 21177
rect 11737 21143 11863 21177
rect 11897 21143 11920 21177
rect 11520 21120 11920 21143
rect 12000 21177 12400 21200
rect 12000 21143 12023 21177
rect 12057 21143 12183 21177
rect 12217 21143 12343 21177
rect 12377 21143 12400 21177
rect 12000 21120 12400 21143
rect 8480 21017 8880 21040
rect 8480 20983 8503 21017
rect 8537 20983 8663 21017
rect 8697 20983 8823 21017
rect 8857 20983 8880 21017
rect 8480 20960 8880 20983
rect 8960 21017 9360 21040
rect 8960 20983 8983 21017
rect 9017 20983 9143 21017
rect 9177 20983 9303 21017
rect 9337 20983 9360 21017
rect 8960 20960 9360 20983
rect 9440 21017 11440 21040
rect 9440 20983 9463 21017
rect 9497 20983 9623 21017
rect 9657 20983 9783 21017
rect 9817 20983 9943 21017
rect 9977 20983 10103 21017
rect 10137 20983 10263 21017
rect 10297 20983 10423 21017
rect 10457 20983 10583 21017
rect 10617 20983 10743 21017
rect 10777 20983 10903 21017
rect 10937 20983 11063 21017
rect 11097 20983 11223 21017
rect 11257 20983 11383 21017
rect 11417 20983 11440 21017
rect 9440 20960 11440 20983
rect 11520 21017 11920 21040
rect 11520 20983 11543 21017
rect 11577 20983 11703 21017
rect 11737 20983 11863 21017
rect 11897 20983 11920 21017
rect 11520 20960 11920 20983
rect 12000 21017 12400 21040
rect 12000 20983 12023 21017
rect 12057 20983 12183 21017
rect 12217 20983 12343 21017
rect 12377 20983 12400 21017
rect 12000 20960 12400 20983
rect 8480 20857 8880 20880
rect 8480 20823 8503 20857
rect 8537 20823 8663 20857
rect 8697 20823 8823 20857
rect 8857 20823 8880 20857
rect 8480 20800 8880 20823
rect 8960 20857 9360 20880
rect 8960 20823 8983 20857
rect 9017 20823 9143 20857
rect 9177 20823 9303 20857
rect 9337 20823 9360 20857
rect 8960 20800 9360 20823
rect 9440 20857 11440 20880
rect 9440 20823 9463 20857
rect 9497 20823 9623 20857
rect 9657 20823 9783 20857
rect 9817 20823 9943 20857
rect 9977 20823 10103 20857
rect 10137 20823 10263 20857
rect 10297 20823 10423 20857
rect 10457 20823 10583 20857
rect 10617 20823 10743 20857
rect 10777 20823 10903 20857
rect 10937 20823 11063 20857
rect 11097 20823 11223 20857
rect 11257 20823 11383 20857
rect 11417 20823 11440 20857
rect 9440 20800 11440 20823
rect 11520 20857 11920 20880
rect 11520 20823 11543 20857
rect 11577 20823 11703 20857
rect 11737 20823 11863 20857
rect 11897 20823 11920 20857
rect 11520 20800 11920 20823
rect 12000 20857 12400 20880
rect 12000 20823 12023 20857
rect 12057 20823 12183 20857
rect 12217 20823 12343 20857
rect 12377 20823 12400 20857
rect 12000 20800 12400 20823
rect 8480 20697 8880 20720
rect 8480 20663 8503 20697
rect 8537 20663 8663 20697
rect 8697 20663 8823 20697
rect 8857 20663 8880 20697
rect 8480 20640 8880 20663
rect 8960 20697 9360 20720
rect 8960 20663 8983 20697
rect 9017 20663 9143 20697
rect 9177 20663 9303 20697
rect 9337 20663 9360 20697
rect 8960 20640 9360 20663
rect 9440 20697 11440 20720
rect 9440 20663 9463 20697
rect 9497 20663 9623 20697
rect 9657 20663 9783 20697
rect 9817 20663 9943 20697
rect 9977 20663 10103 20697
rect 10137 20663 10263 20697
rect 10297 20663 10423 20697
rect 10457 20663 10583 20697
rect 10617 20663 10743 20697
rect 10777 20663 10903 20697
rect 10937 20663 11063 20697
rect 11097 20663 11223 20697
rect 11257 20663 11383 20697
rect 11417 20663 11440 20697
rect 9440 20640 11440 20663
rect 11520 20697 11920 20720
rect 11520 20663 11543 20697
rect 11577 20663 11703 20697
rect 11737 20663 11863 20697
rect 11897 20663 11920 20697
rect 11520 20640 11920 20663
rect 12000 20697 12400 20720
rect 12000 20663 12023 20697
rect 12057 20663 12183 20697
rect 12217 20663 12343 20697
rect 12377 20663 12400 20697
rect 12000 20640 12400 20663
rect 8480 20537 8880 20560
rect 8480 20503 8503 20537
rect 8537 20503 8663 20537
rect 8697 20503 8823 20537
rect 8857 20503 8880 20537
rect 8480 20480 8880 20503
rect 8960 20537 9360 20560
rect 8960 20503 8983 20537
rect 9017 20503 9143 20537
rect 9177 20503 9303 20537
rect 9337 20503 9360 20537
rect 8960 20480 9360 20503
rect 9440 20537 11440 20560
rect 9440 20503 9463 20537
rect 9497 20503 9623 20537
rect 9657 20503 9783 20537
rect 9817 20503 9943 20537
rect 9977 20503 10103 20537
rect 10137 20503 10263 20537
rect 10297 20503 10423 20537
rect 10457 20503 10583 20537
rect 10617 20503 10743 20537
rect 10777 20503 10903 20537
rect 10937 20503 11063 20537
rect 11097 20503 11223 20537
rect 11257 20503 11383 20537
rect 11417 20503 11440 20537
rect 9440 20480 11440 20503
rect 11520 20537 11920 20560
rect 11520 20503 11543 20537
rect 11577 20503 11703 20537
rect 11737 20503 11863 20537
rect 11897 20503 11920 20537
rect 11520 20480 11920 20503
rect 12000 20537 12400 20560
rect 12000 20503 12023 20537
rect 12057 20503 12183 20537
rect 12217 20503 12343 20537
rect 12377 20503 12400 20537
rect 12000 20480 12400 20503
rect 8480 20377 8880 20400
rect 8480 20343 8503 20377
rect 8537 20343 8663 20377
rect 8697 20343 8823 20377
rect 8857 20343 8880 20377
rect 8480 20320 8880 20343
rect 8960 20377 9360 20400
rect 8960 20343 8983 20377
rect 9017 20343 9143 20377
rect 9177 20343 9303 20377
rect 9337 20343 9360 20377
rect 8960 20320 9360 20343
rect 9440 20377 11440 20400
rect 9440 20343 9463 20377
rect 9497 20343 9623 20377
rect 9657 20343 9783 20377
rect 9817 20343 9943 20377
rect 9977 20343 10103 20377
rect 10137 20343 10263 20377
rect 10297 20343 10423 20377
rect 10457 20343 10583 20377
rect 10617 20343 10743 20377
rect 10777 20343 10903 20377
rect 10937 20343 11063 20377
rect 11097 20343 11223 20377
rect 11257 20343 11383 20377
rect 11417 20343 11440 20377
rect 9440 20320 11440 20343
rect 11520 20377 11920 20400
rect 11520 20343 11543 20377
rect 11577 20343 11703 20377
rect 11737 20343 11863 20377
rect 11897 20343 11920 20377
rect 11520 20320 11920 20343
rect 12000 20377 12400 20400
rect 12000 20343 12023 20377
rect 12057 20343 12183 20377
rect 12217 20343 12343 20377
rect 12377 20343 12400 20377
rect 12000 20320 12400 20343
rect 8480 20217 8880 20240
rect 8480 20183 8503 20217
rect 8537 20183 8663 20217
rect 8697 20183 8823 20217
rect 8857 20183 8880 20217
rect 8480 20160 8880 20183
rect 8960 20217 9360 20240
rect 8960 20183 8983 20217
rect 9017 20183 9143 20217
rect 9177 20183 9303 20217
rect 9337 20183 9360 20217
rect 8960 20160 9360 20183
rect 9440 20217 11440 20240
rect 9440 20183 9463 20217
rect 9497 20183 9623 20217
rect 9657 20183 9783 20217
rect 9817 20183 9943 20217
rect 9977 20183 10103 20217
rect 10137 20183 10263 20217
rect 10297 20183 10423 20217
rect 10457 20183 10583 20217
rect 10617 20183 10743 20217
rect 10777 20183 10903 20217
rect 10937 20183 11063 20217
rect 11097 20183 11223 20217
rect 11257 20183 11383 20217
rect 11417 20183 11440 20217
rect 9440 20160 11440 20183
rect 11520 20217 11920 20240
rect 11520 20183 11543 20217
rect 11577 20183 11703 20217
rect 11737 20183 11863 20217
rect 11897 20183 11920 20217
rect 11520 20160 11920 20183
rect 12000 20217 12400 20240
rect 12000 20183 12023 20217
rect 12057 20183 12183 20217
rect 12217 20183 12343 20217
rect 12377 20183 12400 20217
rect 12000 20160 12400 20183
rect 8480 20057 8880 20080
rect 8480 20023 8503 20057
rect 8537 20023 8663 20057
rect 8697 20023 8823 20057
rect 8857 20023 8880 20057
rect 8480 20000 8880 20023
rect 8960 20057 9360 20080
rect 8960 20023 8983 20057
rect 9017 20023 9143 20057
rect 9177 20023 9303 20057
rect 9337 20023 9360 20057
rect 8960 20000 9360 20023
rect 9440 20057 11440 20080
rect 9440 20023 9463 20057
rect 9497 20023 9623 20057
rect 9657 20023 9783 20057
rect 9817 20023 9943 20057
rect 9977 20023 10103 20057
rect 10137 20023 10263 20057
rect 10297 20023 10423 20057
rect 10457 20023 10583 20057
rect 10617 20023 10743 20057
rect 10777 20023 10903 20057
rect 10937 20023 11063 20057
rect 11097 20023 11223 20057
rect 11257 20023 11383 20057
rect 11417 20023 11440 20057
rect 9440 20000 11440 20023
rect 11520 20057 11920 20080
rect 11520 20023 11543 20057
rect 11577 20023 11703 20057
rect 11737 20023 11863 20057
rect 11897 20023 11920 20057
rect 11520 20000 11920 20023
rect 12000 20057 12400 20080
rect 12000 20023 12023 20057
rect 12057 20023 12183 20057
rect 12217 20023 12343 20057
rect 12377 20023 12400 20057
rect 12000 20000 12400 20023
rect 8480 19897 8880 19920
rect 8480 19863 8503 19897
rect 8537 19863 8663 19897
rect 8697 19863 8823 19897
rect 8857 19863 8880 19897
rect 8480 19840 8880 19863
rect 8960 19897 9360 19920
rect 8960 19863 8983 19897
rect 9017 19863 9143 19897
rect 9177 19863 9303 19897
rect 9337 19863 9360 19897
rect 8960 19840 9360 19863
rect 9440 19897 11440 19920
rect 9440 19863 9463 19897
rect 9497 19863 9623 19897
rect 9657 19863 9783 19897
rect 9817 19863 9943 19897
rect 9977 19863 10103 19897
rect 10137 19863 10263 19897
rect 10297 19863 10423 19897
rect 10457 19863 10583 19897
rect 10617 19863 10743 19897
rect 10777 19863 10903 19897
rect 10937 19863 11063 19897
rect 11097 19863 11223 19897
rect 11257 19863 11383 19897
rect 11417 19863 11440 19897
rect 9440 19840 11440 19863
rect 11520 19897 11920 19920
rect 11520 19863 11543 19897
rect 11577 19863 11703 19897
rect 11737 19863 11863 19897
rect 11897 19863 11920 19897
rect 11520 19840 11920 19863
rect 12000 19897 12400 19920
rect 12000 19863 12023 19897
rect 12057 19863 12183 19897
rect 12217 19863 12343 19897
rect 12377 19863 12400 19897
rect 12000 19840 12400 19863
rect 8480 19737 8880 19760
rect 8480 19703 8503 19737
rect 8537 19703 8663 19737
rect 8697 19703 8823 19737
rect 8857 19703 8880 19737
rect 8480 19680 8880 19703
rect 8960 19737 9360 19760
rect 8960 19703 8983 19737
rect 9017 19703 9143 19737
rect 9177 19703 9303 19737
rect 9337 19703 9360 19737
rect 8960 19680 9360 19703
rect 9440 19737 11440 19760
rect 9440 19703 9463 19737
rect 9497 19703 9623 19737
rect 9657 19703 9783 19737
rect 9817 19703 9943 19737
rect 9977 19703 10103 19737
rect 10137 19703 10263 19737
rect 10297 19703 10423 19737
rect 10457 19703 10583 19737
rect 10617 19703 10743 19737
rect 10777 19703 10903 19737
rect 10937 19703 11063 19737
rect 11097 19703 11223 19737
rect 11257 19703 11383 19737
rect 11417 19703 11440 19737
rect 9440 19680 11440 19703
rect 11520 19737 11920 19760
rect 11520 19703 11543 19737
rect 11577 19703 11703 19737
rect 11737 19703 11863 19737
rect 11897 19703 11920 19737
rect 11520 19680 11920 19703
rect 12000 19737 12400 19760
rect 12000 19703 12023 19737
rect 12057 19703 12183 19737
rect 12217 19703 12343 19737
rect 12377 19703 12400 19737
rect 12000 19680 12400 19703
rect 8480 19577 8880 19600
rect 8480 19543 8503 19577
rect 8537 19543 8663 19577
rect 8697 19543 8823 19577
rect 8857 19543 8880 19577
rect 8480 19520 8880 19543
rect 8960 19577 9360 19600
rect 8960 19543 8983 19577
rect 9017 19543 9143 19577
rect 9177 19543 9303 19577
rect 9337 19543 9360 19577
rect 8960 19520 9360 19543
rect 9440 19577 11440 19600
rect 9440 19543 9463 19577
rect 9497 19543 9623 19577
rect 9657 19543 9783 19577
rect 9817 19543 9943 19577
rect 9977 19543 10103 19577
rect 10137 19543 10263 19577
rect 10297 19543 10423 19577
rect 10457 19543 10583 19577
rect 10617 19543 10743 19577
rect 10777 19543 10903 19577
rect 10937 19543 11063 19577
rect 11097 19543 11223 19577
rect 11257 19543 11383 19577
rect 11417 19543 11440 19577
rect 9440 19520 11440 19543
rect 11520 19577 11920 19600
rect 11520 19543 11543 19577
rect 11577 19543 11703 19577
rect 11737 19543 11863 19577
rect 11897 19543 11920 19577
rect 11520 19520 11920 19543
rect 12000 19577 12400 19600
rect 12000 19543 12023 19577
rect 12057 19543 12183 19577
rect 12217 19543 12343 19577
rect 12377 19543 12400 19577
rect 12000 19520 12400 19543
rect 8480 19417 8880 19440
rect 8480 19383 8503 19417
rect 8537 19383 8663 19417
rect 8697 19383 8823 19417
rect 8857 19383 8880 19417
rect 8480 19360 8880 19383
rect 8960 19417 9360 19440
rect 8960 19383 8983 19417
rect 9017 19383 9143 19417
rect 9177 19383 9303 19417
rect 9337 19383 9360 19417
rect 8960 19360 9360 19383
rect 9440 19417 11440 19440
rect 9440 19383 9463 19417
rect 9497 19383 9623 19417
rect 9657 19383 9783 19417
rect 9817 19383 9943 19417
rect 9977 19383 10103 19417
rect 10137 19383 10263 19417
rect 10297 19383 10423 19417
rect 10457 19383 10583 19417
rect 10617 19383 10743 19417
rect 10777 19383 10903 19417
rect 10937 19383 11063 19417
rect 11097 19383 11223 19417
rect 11257 19383 11383 19417
rect 11417 19383 11440 19417
rect 9440 19360 11440 19383
rect 11520 19417 11920 19440
rect 11520 19383 11543 19417
rect 11577 19383 11703 19417
rect 11737 19383 11863 19417
rect 11897 19383 11920 19417
rect 11520 19360 11920 19383
rect 12000 19417 12400 19440
rect 12000 19383 12023 19417
rect 12057 19383 12183 19417
rect 12217 19383 12343 19417
rect 12377 19383 12400 19417
rect 12000 19360 12400 19383
rect 8480 19257 8880 19280
rect 8480 19223 8503 19257
rect 8537 19223 8663 19257
rect 8697 19223 8823 19257
rect 8857 19223 8880 19257
rect 8480 19200 8880 19223
rect 8960 19257 9360 19280
rect 8960 19223 8983 19257
rect 9017 19223 9143 19257
rect 9177 19223 9303 19257
rect 9337 19223 9360 19257
rect 8960 19200 9360 19223
rect 9440 19257 11440 19280
rect 9440 19223 9463 19257
rect 9497 19223 9623 19257
rect 9657 19223 9783 19257
rect 9817 19223 9943 19257
rect 9977 19223 10103 19257
rect 10137 19223 10263 19257
rect 10297 19223 10423 19257
rect 10457 19223 10583 19257
rect 10617 19223 10743 19257
rect 10777 19223 10903 19257
rect 10937 19223 11063 19257
rect 11097 19223 11223 19257
rect 11257 19223 11383 19257
rect 11417 19223 11440 19257
rect 9440 19200 11440 19223
rect 11520 19257 11920 19280
rect 11520 19223 11543 19257
rect 11577 19223 11703 19257
rect 11737 19223 11863 19257
rect 11897 19223 11920 19257
rect 11520 19200 11920 19223
rect 12000 19257 12400 19280
rect 12000 19223 12023 19257
rect 12057 19223 12183 19257
rect 12217 19223 12343 19257
rect 12377 19223 12400 19257
rect 12000 19200 12400 19223
rect 8480 19097 8880 19120
rect 8480 19063 8503 19097
rect 8537 19063 8663 19097
rect 8697 19063 8823 19097
rect 8857 19063 8880 19097
rect 8480 19040 8880 19063
rect 8960 19097 9360 19120
rect 8960 19063 8983 19097
rect 9017 19063 9143 19097
rect 9177 19063 9303 19097
rect 9337 19063 9360 19097
rect 8960 19040 9360 19063
rect 9440 19097 11440 19120
rect 9440 19063 9463 19097
rect 9497 19063 9623 19097
rect 9657 19063 9783 19097
rect 9817 19063 9943 19097
rect 9977 19063 10103 19097
rect 10137 19063 10263 19097
rect 10297 19063 10423 19097
rect 10457 19063 10583 19097
rect 10617 19063 10743 19097
rect 10777 19063 10903 19097
rect 10937 19063 11063 19097
rect 11097 19063 11223 19097
rect 11257 19063 11383 19097
rect 11417 19063 11440 19097
rect 9440 19040 11440 19063
rect 11520 19097 11920 19120
rect 11520 19063 11543 19097
rect 11577 19063 11703 19097
rect 11737 19063 11863 19097
rect 11897 19063 11920 19097
rect 11520 19040 11920 19063
rect 12000 19097 12400 19120
rect 12000 19063 12023 19097
rect 12057 19063 12183 19097
rect 12217 19063 12343 19097
rect 12377 19063 12400 19097
rect 12000 19040 12400 19063
rect 8480 18937 8880 18960
rect 8480 18903 8503 18937
rect 8537 18903 8663 18937
rect 8697 18903 8823 18937
rect 8857 18903 8880 18937
rect 8480 18880 8880 18903
rect 8960 18937 9360 18960
rect 8960 18903 8983 18937
rect 9017 18903 9143 18937
rect 9177 18903 9303 18937
rect 9337 18903 9360 18937
rect 8960 18880 9360 18903
rect 9440 18937 11440 18960
rect 9440 18903 9463 18937
rect 9497 18903 9623 18937
rect 9657 18903 9783 18937
rect 9817 18903 9943 18937
rect 9977 18903 10103 18937
rect 10137 18903 10263 18937
rect 10297 18903 10423 18937
rect 10457 18903 10583 18937
rect 10617 18903 10743 18937
rect 10777 18903 10903 18937
rect 10937 18903 11063 18937
rect 11097 18903 11223 18937
rect 11257 18903 11383 18937
rect 11417 18903 11440 18937
rect 9440 18880 11440 18903
rect 11520 18937 11920 18960
rect 11520 18903 11543 18937
rect 11577 18903 11703 18937
rect 11737 18903 11863 18937
rect 11897 18903 11920 18937
rect 11520 18880 11920 18903
rect 12000 18937 12400 18960
rect 12000 18903 12023 18937
rect 12057 18903 12183 18937
rect 12217 18903 12343 18937
rect 12377 18903 12400 18937
rect 12000 18880 12400 18903
rect 8480 18777 8880 18800
rect 8480 18743 8503 18777
rect 8537 18743 8663 18777
rect 8697 18743 8823 18777
rect 8857 18743 8880 18777
rect 8480 18720 8880 18743
rect 8960 18777 9360 18800
rect 8960 18743 8983 18777
rect 9017 18743 9143 18777
rect 9177 18743 9303 18777
rect 9337 18743 9360 18777
rect 8960 18720 9360 18743
rect 9440 18777 11440 18800
rect 9440 18743 9463 18777
rect 9497 18743 9623 18777
rect 9657 18743 9783 18777
rect 9817 18743 9943 18777
rect 9977 18743 10103 18777
rect 10137 18743 10263 18777
rect 10297 18743 10423 18777
rect 10457 18743 10583 18777
rect 10617 18743 10743 18777
rect 10777 18743 10903 18777
rect 10937 18743 11063 18777
rect 11097 18743 11223 18777
rect 11257 18743 11383 18777
rect 11417 18743 11440 18777
rect 9440 18720 11440 18743
rect 11520 18777 11920 18800
rect 11520 18743 11543 18777
rect 11577 18743 11703 18777
rect 11737 18743 11863 18777
rect 11897 18743 11920 18777
rect 11520 18720 11920 18743
rect 12000 18777 12400 18800
rect 12000 18743 12023 18777
rect 12057 18743 12183 18777
rect 12217 18743 12343 18777
rect 12377 18743 12400 18777
rect 12000 18720 12400 18743
rect 8480 18617 8880 18640
rect 8480 18583 8503 18617
rect 8537 18583 8663 18617
rect 8697 18583 8823 18617
rect 8857 18583 8880 18617
rect 8480 18560 8880 18583
rect 8960 18617 9360 18640
rect 8960 18583 8983 18617
rect 9017 18583 9143 18617
rect 9177 18583 9303 18617
rect 9337 18583 9360 18617
rect 8960 18560 9360 18583
rect 9440 18617 11440 18640
rect 9440 18583 9463 18617
rect 9497 18583 9623 18617
rect 9657 18583 9783 18617
rect 9817 18583 9943 18617
rect 9977 18583 10103 18617
rect 10137 18583 10263 18617
rect 10297 18583 10423 18617
rect 10457 18583 10583 18617
rect 10617 18583 10743 18617
rect 10777 18583 10903 18617
rect 10937 18583 11063 18617
rect 11097 18583 11223 18617
rect 11257 18583 11383 18617
rect 11417 18583 11440 18617
rect 9440 18560 11440 18583
rect 11520 18617 11920 18640
rect 11520 18583 11543 18617
rect 11577 18583 11703 18617
rect 11737 18583 11863 18617
rect 11897 18583 11920 18617
rect 11520 18560 11920 18583
rect 12000 18617 12400 18640
rect 12000 18583 12023 18617
rect 12057 18583 12183 18617
rect 12217 18583 12343 18617
rect 12377 18583 12400 18617
rect 12000 18560 12400 18583
rect 8480 18457 8880 18480
rect 8480 18423 8503 18457
rect 8537 18423 8663 18457
rect 8697 18423 8823 18457
rect 8857 18423 8880 18457
rect 8480 18400 8880 18423
rect 8960 18457 9360 18480
rect 8960 18423 8983 18457
rect 9017 18423 9143 18457
rect 9177 18423 9303 18457
rect 9337 18423 9360 18457
rect 8960 18400 9360 18423
rect 9440 18457 11440 18480
rect 9440 18423 9463 18457
rect 9497 18423 9623 18457
rect 9657 18423 9783 18457
rect 9817 18423 9943 18457
rect 9977 18423 10103 18457
rect 10137 18423 10263 18457
rect 10297 18423 10423 18457
rect 10457 18423 10583 18457
rect 10617 18423 10743 18457
rect 10777 18423 10903 18457
rect 10937 18423 11063 18457
rect 11097 18423 11223 18457
rect 11257 18423 11383 18457
rect 11417 18423 11440 18457
rect 9440 18400 11440 18423
rect 11520 18457 11920 18480
rect 11520 18423 11543 18457
rect 11577 18423 11703 18457
rect 11737 18423 11863 18457
rect 11897 18423 11920 18457
rect 11520 18400 11920 18423
rect 12000 18457 12400 18480
rect 12000 18423 12023 18457
rect 12057 18423 12183 18457
rect 12217 18423 12343 18457
rect 12377 18423 12400 18457
rect 12000 18400 12400 18423
rect 8480 18297 8880 18320
rect 8480 18263 8503 18297
rect 8537 18263 8663 18297
rect 8697 18263 8823 18297
rect 8857 18263 8880 18297
rect 8480 18240 8880 18263
rect 8960 18297 9360 18320
rect 8960 18263 8983 18297
rect 9017 18263 9143 18297
rect 9177 18263 9303 18297
rect 9337 18263 9360 18297
rect 8960 18240 9360 18263
rect 9440 18297 11440 18320
rect 9440 18263 9463 18297
rect 9497 18263 9623 18297
rect 9657 18263 9783 18297
rect 9817 18263 9943 18297
rect 9977 18263 10103 18297
rect 10137 18263 10263 18297
rect 10297 18263 10423 18297
rect 10457 18263 10583 18297
rect 10617 18263 10743 18297
rect 10777 18263 10903 18297
rect 10937 18263 11063 18297
rect 11097 18263 11223 18297
rect 11257 18263 11383 18297
rect 11417 18263 11440 18297
rect 9440 18240 11440 18263
rect 11520 18297 11920 18320
rect 11520 18263 11543 18297
rect 11577 18263 11703 18297
rect 11737 18263 11863 18297
rect 11897 18263 11920 18297
rect 11520 18240 11920 18263
rect 12000 18297 12400 18320
rect 12000 18263 12023 18297
rect 12057 18263 12183 18297
rect 12217 18263 12343 18297
rect 12377 18263 12400 18297
rect 12000 18240 12400 18263
rect 8480 18137 8880 18160
rect 8480 18103 8503 18137
rect 8537 18103 8663 18137
rect 8697 18103 8823 18137
rect 8857 18103 8880 18137
rect 8480 18080 8880 18103
rect 8960 18137 9360 18160
rect 8960 18103 8983 18137
rect 9017 18103 9143 18137
rect 9177 18103 9303 18137
rect 9337 18103 9360 18137
rect 8960 18080 9360 18103
rect 9440 18137 11440 18160
rect 9440 18103 9463 18137
rect 9497 18103 9623 18137
rect 9657 18103 9783 18137
rect 9817 18103 9943 18137
rect 9977 18103 10103 18137
rect 10137 18103 10263 18137
rect 10297 18103 10423 18137
rect 10457 18103 10583 18137
rect 10617 18103 10743 18137
rect 10777 18103 10903 18137
rect 10937 18103 11063 18137
rect 11097 18103 11223 18137
rect 11257 18103 11383 18137
rect 11417 18103 11440 18137
rect 9440 18080 11440 18103
rect 11520 18137 11920 18160
rect 11520 18103 11543 18137
rect 11577 18103 11703 18137
rect 11737 18103 11863 18137
rect 11897 18103 11920 18137
rect 11520 18080 11920 18103
rect 12000 18137 12400 18160
rect 12000 18103 12023 18137
rect 12057 18103 12183 18137
rect 12217 18103 12343 18137
rect 12377 18103 12400 18137
rect 12000 18080 12400 18103
rect 8480 17977 8880 18000
rect 8480 17943 8503 17977
rect 8537 17943 8663 17977
rect 8697 17943 8823 17977
rect 8857 17943 8880 17977
rect 8480 17920 8880 17943
rect 8960 17977 9360 18000
rect 8960 17943 8983 17977
rect 9017 17943 9143 17977
rect 9177 17943 9303 17977
rect 9337 17943 9360 17977
rect 8960 17920 9360 17943
rect 9440 17977 11440 18000
rect 9440 17943 9463 17977
rect 9497 17943 9623 17977
rect 9657 17943 9783 17977
rect 9817 17943 9943 17977
rect 9977 17943 10103 17977
rect 10137 17943 10263 17977
rect 10297 17943 10423 17977
rect 10457 17943 10583 17977
rect 10617 17943 10743 17977
rect 10777 17943 10903 17977
rect 10937 17943 11063 17977
rect 11097 17943 11223 17977
rect 11257 17943 11383 17977
rect 11417 17943 11440 17977
rect 9440 17920 11440 17943
rect 11520 17977 11920 18000
rect 11520 17943 11543 17977
rect 11577 17943 11703 17977
rect 11737 17943 11863 17977
rect 11897 17943 11920 17977
rect 11520 17920 11920 17943
rect 12000 17977 12400 18000
rect 12000 17943 12023 17977
rect 12057 17943 12183 17977
rect 12217 17943 12343 17977
rect 12377 17943 12400 17977
rect 12000 17920 12400 17943
rect 8480 17817 8880 17840
rect 8480 17783 8503 17817
rect 8537 17783 8663 17817
rect 8697 17783 8823 17817
rect 8857 17783 8880 17817
rect 8480 17760 8880 17783
rect 8960 17817 9360 17840
rect 8960 17783 8983 17817
rect 9017 17783 9143 17817
rect 9177 17783 9303 17817
rect 9337 17783 9360 17817
rect 8960 17760 9360 17783
rect 9440 17817 11440 17840
rect 9440 17783 9463 17817
rect 9497 17783 9623 17817
rect 9657 17783 9783 17817
rect 9817 17783 9943 17817
rect 9977 17783 10103 17817
rect 10137 17783 10263 17817
rect 10297 17783 10423 17817
rect 10457 17783 10583 17817
rect 10617 17783 10743 17817
rect 10777 17783 10903 17817
rect 10937 17783 11063 17817
rect 11097 17783 11223 17817
rect 11257 17783 11383 17817
rect 11417 17783 11440 17817
rect 9440 17760 11440 17783
rect 11520 17817 11920 17840
rect 11520 17783 11543 17817
rect 11577 17783 11703 17817
rect 11737 17783 11863 17817
rect 11897 17783 11920 17817
rect 11520 17760 11920 17783
rect 12000 17817 12400 17840
rect 12000 17783 12023 17817
rect 12057 17783 12183 17817
rect 12217 17783 12343 17817
rect 12377 17783 12400 17817
rect 12000 17760 12400 17783
rect 8480 17657 8880 17680
rect 8480 17623 8503 17657
rect 8537 17623 8663 17657
rect 8697 17623 8823 17657
rect 8857 17623 8880 17657
rect 8480 17600 8880 17623
rect 8960 17657 9360 17680
rect 8960 17623 8983 17657
rect 9017 17623 9143 17657
rect 9177 17623 9303 17657
rect 9337 17623 9360 17657
rect 8960 17600 9360 17623
rect 9440 17657 11440 17680
rect 9440 17623 9463 17657
rect 9497 17623 9623 17657
rect 9657 17623 9783 17657
rect 9817 17623 9943 17657
rect 9977 17623 10103 17657
rect 10137 17623 10263 17657
rect 10297 17623 10423 17657
rect 10457 17623 10583 17657
rect 10617 17623 10743 17657
rect 10777 17623 10903 17657
rect 10937 17623 11063 17657
rect 11097 17623 11223 17657
rect 11257 17623 11383 17657
rect 11417 17623 11440 17657
rect 9440 17600 11440 17623
rect 11520 17657 11920 17680
rect 11520 17623 11543 17657
rect 11577 17623 11703 17657
rect 11737 17623 11863 17657
rect 11897 17623 11920 17657
rect 11520 17600 11920 17623
rect 12000 17657 12400 17680
rect 12000 17623 12023 17657
rect 12057 17623 12183 17657
rect 12217 17623 12343 17657
rect 12377 17623 12400 17657
rect 12000 17600 12400 17623
rect 8480 17497 8880 17520
rect 8480 17463 8503 17497
rect 8537 17463 8663 17497
rect 8697 17463 8823 17497
rect 8857 17463 8880 17497
rect 8480 17440 8880 17463
rect 8960 17497 9360 17520
rect 8960 17463 8983 17497
rect 9017 17463 9143 17497
rect 9177 17463 9303 17497
rect 9337 17463 9360 17497
rect 8960 17440 9360 17463
rect 9440 17497 11440 17520
rect 9440 17463 9463 17497
rect 9497 17463 9623 17497
rect 9657 17463 9783 17497
rect 9817 17463 9943 17497
rect 9977 17463 10103 17497
rect 10137 17463 10263 17497
rect 10297 17463 10423 17497
rect 10457 17463 10583 17497
rect 10617 17463 10743 17497
rect 10777 17463 10903 17497
rect 10937 17463 11063 17497
rect 11097 17463 11223 17497
rect 11257 17463 11383 17497
rect 11417 17463 11440 17497
rect 9440 17440 11440 17463
rect 11520 17497 11920 17520
rect 11520 17463 11543 17497
rect 11577 17463 11703 17497
rect 11737 17463 11863 17497
rect 11897 17463 11920 17497
rect 11520 17440 11920 17463
rect 12000 17497 12400 17520
rect 12000 17463 12023 17497
rect 12057 17463 12183 17497
rect 12217 17463 12343 17497
rect 12377 17463 12400 17497
rect 12000 17440 12400 17463
rect 8480 17337 8880 17360
rect 8480 17303 8503 17337
rect 8537 17303 8663 17337
rect 8697 17303 8823 17337
rect 8857 17303 8880 17337
rect 8480 17280 8880 17303
rect 8960 17337 9360 17360
rect 8960 17303 8983 17337
rect 9017 17303 9143 17337
rect 9177 17303 9303 17337
rect 9337 17303 9360 17337
rect 8960 17280 9360 17303
rect 9440 17337 11440 17360
rect 9440 17303 9463 17337
rect 9497 17303 9623 17337
rect 9657 17303 9783 17337
rect 9817 17303 9943 17337
rect 9977 17303 10103 17337
rect 10137 17303 10263 17337
rect 10297 17303 10423 17337
rect 10457 17303 10583 17337
rect 10617 17303 10743 17337
rect 10777 17303 10903 17337
rect 10937 17303 11063 17337
rect 11097 17303 11223 17337
rect 11257 17303 11383 17337
rect 11417 17303 11440 17337
rect 9440 17280 11440 17303
rect 11520 17337 11920 17360
rect 11520 17303 11543 17337
rect 11577 17303 11703 17337
rect 11737 17303 11863 17337
rect 11897 17303 11920 17337
rect 11520 17280 11920 17303
rect 12000 17337 12400 17360
rect 12000 17303 12023 17337
rect 12057 17303 12183 17337
rect 12217 17303 12343 17337
rect 12377 17303 12400 17337
rect 12000 17280 12400 17303
rect 8480 17177 8880 17200
rect 8480 17143 8503 17177
rect 8537 17143 8663 17177
rect 8697 17143 8823 17177
rect 8857 17143 8880 17177
rect 8480 17120 8880 17143
rect 8960 17177 9360 17200
rect 8960 17143 8983 17177
rect 9017 17143 9143 17177
rect 9177 17143 9303 17177
rect 9337 17143 9360 17177
rect 8960 17120 9360 17143
rect 9440 17177 11440 17200
rect 9440 17143 9463 17177
rect 9497 17143 9623 17177
rect 9657 17143 9783 17177
rect 9817 17143 9943 17177
rect 9977 17143 10103 17177
rect 10137 17143 10263 17177
rect 10297 17143 10423 17177
rect 10457 17143 10583 17177
rect 10617 17143 10743 17177
rect 10777 17143 10903 17177
rect 10937 17143 11063 17177
rect 11097 17143 11223 17177
rect 11257 17143 11383 17177
rect 11417 17143 11440 17177
rect 9440 17120 11440 17143
rect 11520 17177 11920 17200
rect 11520 17143 11543 17177
rect 11577 17143 11703 17177
rect 11737 17143 11863 17177
rect 11897 17143 11920 17177
rect 11520 17120 11920 17143
rect 12000 17177 12400 17200
rect 12000 17143 12023 17177
rect 12057 17143 12183 17177
rect 12217 17143 12343 17177
rect 12377 17143 12400 17177
rect 12000 17120 12400 17143
rect 8480 17017 8880 17040
rect 8480 16983 8503 17017
rect 8537 16983 8663 17017
rect 8697 16983 8823 17017
rect 8857 16983 8880 17017
rect 8480 16960 8880 16983
rect 8960 17017 9360 17040
rect 8960 16983 8983 17017
rect 9017 16983 9143 17017
rect 9177 16983 9303 17017
rect 9337 16983 9360 17017
rect 8960 16960 9360 16983
rect 9440 17017 11440 17040
rect 9440 16983 9463 17017
rect 9497 16983 9623 17017
rect 9657 16983 9783 17017
rect 9817 16983 9943 17017
rect 9977 16983 10103 17017
rect 10137 16983 10263 17017
rect 10297 16983 10423 17017
rect 10457 16983 10583 17017
rect 10617 16983 10743 17017
rect 10777 16983 10903 17017
rect 10937 16983 11063 17017
rect 11097 16983 11223 17017
rect 11257 16983 11383 17017
rect 11417 16983 11440 17017
rect 9440 16960 11440 16983
rect 11520 17017 11920 17040
rect 11520 16983 11543 17017
rect 11577 16983 11703 17017
rect 11737 16983 11863 17017
rect 11897 16983 11920 17017
rect 11520 16960 11920 16983
rect 12000 17017 12400 17040
rect 12000 16983 12023 17017
rect 12057 16983 12183 17017
rect 12217 16983 12343 17017
rect 12377 16983 12400 17017
rect 12000 16960 12400 16983
rect 8480 16857 8880 16880
rect 8480 16823 8503 16857
rect 8537 16823 8663 16857
rect 8697 16823 8823 16857
rect 8857 16823 8880 16857
rect 8480 16800 8880 16823
rect 8960 16857 9360 16880
rect 8960 16823 8983 16857
rect 9017 16823 9143 16857
rect 9177 16823 9303 16857
rect 9337 16823 9360 16857
rect 8960 16800 9360 16823
rect 9440 16857 11440 16880
rect 9440 16823 9463 16857
rect 9497 16823 9623 16857
rect 9657 16823 9783 16857
rect 9817 16823 9943 16857
rect 9977 16823 10103 16857
rect 10137 16823 10263 16857
rect 10297 16823 10423 16857
rect 10457 16823 10583 16857
rect 10617 16823 10743 16857
rect 10777 16823 10903 16857
rect 10937 16823 11063 16857
rect 11097 16823 11223 16857
rect 11257 16823 11383 16857
rect 11417 16823 11440 16857
rect 9440 16800 11440 16823
rect 11520 16857 11920 16880
rect 11520 16823 11543 16857
rect 11577 16823 11703 16857
rect 11737 16823 11863 16857
rect 11897 16823 11920 16857
rect 11520 16800 11920 16823
rect 12000 16857 12400 16880
rect 12000 16823 12023 16857
rect 12057 16823 12183 16857
rect 12217 16823 12343 16857
rect 12377 16823 12400 16857
rect 12000 16800 12400 16823
rect 8480 16697 8880 16720
rect 8480 16663 8503 16697
rect 8537 16663 8663 16697
rect 8697 16663 8823 16697
rect 8857 16663 8880 16697
rect 8480 16640 8880 16663
rect 8960 16697 9360 16720
rect 8960 16663 8983 16697
rect 9017 16663 9143 16697
rect 9177 16663 9303 16697
rect 9337 16663 9360 16697
rect 8960 16640 9360 16663
rect 9440 16697 11440 16720
rect 9440 16663 9463 16697
rect 9497 16663 9623 16697
rect 9657 16663 9783 16697
rect 9817 16663 9943 16697
rect 9977 16663 10103 16697
rect 10137 16663 10263 16697
rect 10297 16663 10423 16697
rect 10457 16663 10583 16697
rect 10617 16663 10743 16697
rect 10777 16663 10903 16697
rect 10937 16663 11063 16697
rect 11097 16663 11223 16697
rect 11257 16663 11383 16697
rect 11417 16663 11440 16697
rect 9440 16640 11440 16663
rect 11520 16697 11920 16720
rect 11520 16663 11543 16697
rect 11577 16663 11703 16697
rect 11737 16663 11863 16697
rect 11897 16663 11920 16697
rect 11520 16640 11920 16663
rect 12000 16697 12400 16720
rect 12000 16663 12023 16697
rect 12057 16663 12183 16697
rect 12217 16663 12343 16697
rect 12377 16663 12400 16697
rect 12000 16640 12400 16663
rect 8480 16537 8880 16560
rect 8480 16503 8503 16537
rect 8537 16503 8663 16537
rect 8697 16503 8823 16537
rect 8857 16503 8880 16537
rect 8480 16480 8880 16503
rect 8960 16537 9360 16560
rect 8960 16503 8983 16537
rect 9017 16503 9143 16537
rect 9177 16503 9303 16537
rect 9337 16503 9360 16537
rect 8960 16480 9360 16503
rect 9440 16537 11440 16560
rect 9440 16503 9463 16537
rect 9497 16503 9623 16537
rect 9657 16503 9783 16537
rect 9817 16503 9943 16537
rect 9977 16503 10103 16537
rect 10137 16503 10263 16537
rect 10297 16503 10423 16537
rect 10457 16503 10583 16537
rect 10617 16503 10743 16537
rect 10777 16503 10903 16537
rect 10937 16503 11063 16537
rect 11097 16503 11223 16537
rect 11257 16503 11383 16537
rect 11417 16503 11440 16537
rect 9440 16480 11440 16503
rect 11520 16537 11920 16560
rect 11520 16503 11543 16537
rect 11577 16503 11703 16537
rect 11737 16503 11863 16537
rect 11897 16503 11920 16537
rect 11520 16480 11920 16503
rect 12000 16537 12400 16560
rect 12000 16503 12023 16537
rect 12057 16503 12183 16537
rect 12217 16503 12343 16537
rect 12377 16503 12400 16537
rect 12000 16480 12400 16503
rect 8480 16377 8880 16400
rect 8480 16343 8503 16377
rect 8537 16343 8663 16377
rect 8697 16343 8823 16377
rect 8857 16343 8880 16377
rect 8480 16320 8880 16343
rect 8960 16377 9360 16400
rect 8960 16343 8983 16377
rect 9017 16343 9143 16377
rect 9177 16343 9303 16377
rect 9337 16343 9360 16377
rect 8960 16320 9360 16343
rect 9440 16377 11440 16400
rect 9440 16343 9463 16377
rect 9497 16343 9623 16377
rect 9657 16343 9783 16377
rect 9817 16343 9943 16377
rect 9977 16343 10103 16377
rect 10137 16343 10263 16377
rect 10297 16343 10423 16377
rect 10457 16343 10583 16377
rect 10617 16343 10743 16377
rect 10777 16343 10903 16377
rect 10937 16343 11063 16377
rect 11097 16343 11223 16377
rect 11257 16343 11383 16377
rect 11417 16343 11440 16377
rect 9440 16320 11440 16343
rect 11520 16377 11920 16400
rect 11520 16343 11543 16377
rect 11577 16343 11703 16377
rect 11737 16343 11863 16377
rect 11897 16343 11920 16377
rect 11520 16320 11920 16343
rect 12000 16377 12400 16400
rect 12000 16343 12023 16377
rect 12057 16343 12183 16377
rect 12217 16343 12343 16377
rect 12377 16343 12400 16377
rect 12000 16320 12400 16343
rect 8480 16217 8880 16240
rect 8480 16183 8503 16217
rect 8537 16183 8663 16217
rect 8697 16183 8823 16217
rect 8857 16183 8880 16217
rect 8480 16160 8880 16183
rect 8960 16217 9360 16240
rect 8960 16183 8983 16217
rect 9017 16183 9143 16217
rect 9177 16183 9303 16217
rect 9337 16183 9360 16217
rect 8960 16160 9360 16183
rect 9440 16217 11440 16240
rect 9440 16183 9463 16217
rect 9497 16183 9623 16217
rect 9657 16183 9783 16217
rect 9817 16183 9943 16217
rect 9977 16183 10103 16217
rect 10137 16183 10263 16217
rect 10297 16183 10423 16217
rect 10457 16183 10583 16217
rect 10617 16183 10743 16217
rect 10777 16183 10903 16217
rect 10937 16183 11063 16217
rect 11097 16183 11223 16217
rect 11257 16183 11383 16217
rect 11417 16183 11440 16217
rect 9440 16160 11440 16183
rect 11520 16217 11920 16240
rect 11520 16183 11543 16217
rect 11577 16183 11703 16217
rect 11737 16183 11863 16217
rect 11897 16183 11920 16217
rect 11520 16160 11920 16183
rect 12000 16217 12400 16240
rect 12000 16183 12023 16217
rect 12057 16183 12183 16217
rect 12217 16183 12343 16217
rect 12377 16183 12400 16217
rect 12000 16160 12400 16183
rect 8480 16057 8880 16080
rect 8480 16023 8503 16057
rect 8537 16023 8663 16057
rect 8697 16023 8823 16057
rect 8857 16023 8880 16057
rect 8480 16000 8880 16023
rect 8960 16057 9360 16080
rect 8960 16023 8983 16057
rect 9017 16023 9143 16057
rect 9177 16023 9303 16057
rect 9337 16023 9360 16057
rect 8960 16000 9360 16023
rect 9440 16057 11440 16080
rect 9440 16023 9463 16057
rect 9497 16023 9623 16057
rect 9657 16023 9783 16057
rect 9817 16023 9943 16057
rect 9977 16023 10103 16057
rect 10137 16023 10263 16057
rect 10297 16023 10423 16057
rect 10457 16023 10583 16057
rect 10617 16023 10743 16057
rect 10777 16023 10903 16057
rect 10937 16023 11063 16057
rect 11097 16023 11223 16057
rect 11257 16023 11383 16057
rect 11417 16023 11440 16057
rect 9440 16000 11440 16023
rect 11520 16057 11920 16080
rect 11520 16023 11543 16057
rect 11577 16023 11703 16057
rect 11737 16023 11863 16057
rect 11897 16023 11920 16057
rect 11520 16000 11920 16023
rect 12000 16057 12400 16080
rect 12000 16023 12023 16057
rect 12057 16023 12183 16057
rect 12217 16023 12343 16057
rect 12377 16023 12400 16057
rect 12000 16000 12400 16023
rect 8480 15897 8880 15920
rect 8480 15863 8503 15897
rect 8537 15863 8663 15897
rect 8697 15863 8823 15897
rect 8857 15863 8880 15897
rect 8480 15840 8880 15863
rect 8960 15897 9360 15920
rect 8960 15863 8983 15897
rect 9017 15863 9143 15897
rect 9177 15863 9303 15897
rect 9337 15863 9360 15897
rect 8960 15840 9360 15863
rect 9440 15897 11440 15920
rect 9440 15863 9463 15897
rect 9497 15863 9623 15897
rect 9657 15863 9783 15897
rect 9817 15863 9943 15897
rect 9977 15863 10103 15897
rect 10137 15863 10263 15897
rect 10297 15863 10423 15897
rect 10457 15863 10583 15897
rect 10617 15863 10743 15897
rect 10777 15863 10903 15897
rect 10937 15863 11063 15897
rect 11097 15863 11223 15897
rect 11257 15863 11383 15897
rect 11417 15863 11440 15897
rect 9440 15840 11440 15863
rect 11520 15897 11920 15920
rect 11520 15863 11543 15897
rect 11577 15863 11703 15897
rect 11737 15863 11863 15897
rect 11897 15863 11920 15897
rect 11520 15840 11920 15863
rect 12000 15897 12400 15920
rect 12000 15863 12023 15897
rect 12057 15863 12183 15897
rect 12217 15863 12343 15897
rect 12377 15863 12400 15897
rect 12000 15840 12400 15863
rect 8480 15737 8880 15760
rect 8480 15703 8503 15737
rect 8537 15703 8663 15737
rect 8697 15703 8823 15737
rect 8857 15703 8880 15737
rect 8480 15680 8880 15703
rect 8960 15737 9360 15760
rect 8960 15703 8983 15737
rect 9017 15703 9143 15737
rect 9177 15703 9303 15737
rect 9337 15703 9360 15737
rect 8960 15680 9360 15703
rect 9440 15737 11440 15760
rect 9440 15703 9463 15737
rect 9497 15703 9623 15737
rect 9657 15703 9783 15737
rect 9817 15703 9943 15737
rect 9977 15703 10103 15737
rect 10137 15703 10263 15737
rect 10297 15703 10423 15737
rect 10457 15703 10583 15737
rect 10617 15703 10743 15737
rect 10777 15703 10903 15737
rect 10937 15703 11063 15737
rect 11097 15703 11223 15737
rect 11257 15703 11383 15737
rect 11417 15703 11440 15737
rect 9440 15680 11440 15703
rect 11520 15737 11920 15760
rect 11520 15703 11543 15737
rect 11577 15703 11703 15737
rect 11737 15703 11863 15737
rect 11897 15703 11920 15737
rect 11520 15680 11920 15703
rect 12000 15737 12400 15760
rect 12000 15703 12023 15737
rect 12057 15703 12183 15737
rect 12217 15703 12343 15737
rect 12377 15703 12400 15737
rect 12000 15680 12400 15703
rect 8480 15577 8880 15600
rect 8480 15543 8503 15577
rect 8537 15543 8663 15577
rect 8697 15543 8823 15577
rect 8857 15543 8880 15577
rect 8480 15520 8880 15543
rect 8960 15577 9360 15600
rect 8960 15543 8983 15577
rect 9017 15543 9143 15577
rect 9177 15543 9303 15577
rect 9337 15543 9360 15577
rect 8960 15520 9360 15543
rect 9440 15577 11440 15600
rect 9440 15543 9463 15577
rect 9497 15543 9623 15577
rect 9657 15543 9783 15577
rect 9817 15543 9943 15577
rect 9977 15543 10103 15577
rect 10137 15543 10263 15577
rect 10297 15543 10423 15577
rect 10457 15543 10583 15577
rect 10617 15543 10743 15577
rect 10777 15543 10903 15577
rect 10937 15543 11063 15577
rect 11097 15543 11223 15577
rect 11257 15543 11383 15577
rect 11417 15543 11440 15577
rect 9440 15520 11440 15543
rect 11520 15577 11920 15600
rect 11520 15543 11543 15577
rect 11577 15543 11703 15577
rect 11737 15543 11863 15577
rect 11897 15543 11920 15577
rect 11520 15520 11920 15543
rect 12000 15577 12400 15600
rect 12000 15543 12023 15577
rect 12057 15543 12183 15577
rect 12217 15543 12343 15577
rect 12377 15543 12400 15577
rect 12000 15520 12400 15543
rect 8480 15417 8880 15440
rect 8480 15383 8503 15417
rect 8537 15383 8663 15417
rect 8697 15383 8823 15417
rect 8857 15383 8880 15417
rect 8480 15360 8880 15383
rect 8960 15417 9360 15440
rect 8960 15383 8983 15417
rect 9017 15383 9143 15417
rect 9177 15383 9303 15417
rect 9337 15383 9360 15417
rect 8960 15360 9360 15383
rect 9440 15417 11440 15440
rect 9440 15383 9463 15417
rect 9497 15383 9623 15417
rect 9657 15383 9783 15417
rect 9817 15383 9943 15417
rect 9977 15383 10103 15417
rect 10137 15383 10263 15417
rect 10297 15383 10423 15417
rect 10457 15383 10583 15417
rect 10617 15383 10743 15417
rect 10777 15383 10903 15417
rect 10937 15383 11063 15417
rect 11097 15383 11223 15417
rect 11257 15383 11383 15417
rect 11417 15383 11440 15417
rect 9440 15360 11440 15383
rect 11520 15417 11920 15440
rect 11520 15383 11543 15417
rect 11577 15383 11703 15417
rect 11737 15383 11863 15417
rect 11897 15383 11920 15417
rect 11520 15360 11920 15383
rect 12000 15417 12400 15440
rect 12000 15383 12023 15417
rect 12057 15383 12183 15417
rect 12217 15383 12343 15417
rect 12377 15383 12400 15417
rect 12000 15360 12400 15383
rect 8480 15257 8880 15280
rect 8480 15223 8503 15257
rect 8537 15223 8663 15257
rect 8697 15223 8823 15257
rect 8857 15223 8880 15257
rect 8480 15200 8880 15223
rect 8960 15257 9360 15280
rect 8960 15223 8983 15257
rect 9017 15223 9143 15257
rect 9177 15223 9303 15257
rect 9337 15223 9360 15257
rect 8960 15200 9360 15223
rect 9440 15257 11440 15280
rect 9440 15223 9463 15257
rect 9497 15223 9623 15257
rect 9657 15223 9783 15257
rect 9817 15223 9943 15257
rect 9977 15223 10103 15257
rect 10137 15223 10263 15257
rect 10297 15223 10423 15257
rect 10457 15223 10583 15257
rect 10617 15223 10743 15257
rect 10777 15223 10903 15257
rect 10937 15223 11063 15257
rect 11097 15223 11223 15257
rect 11257 15223 11383 15257
rect 11417 15223 11440 15257
rect 9440 15200 11440 15223
rect 11520 15257 11920 15280
rect 11520 15223 11543 15257
rect 11577 15223 11703 15257
rect 11737 15223 11863 15257
rect 11897 15223 11920 15257
rect 11520 15200 11920 15223
rect 12000 15257 12400 15280
rect 12000 15223 12023 15257
rect 12057 15223 12183 15257
rect 12217 15223 12343 15257
rect 12377 15223 12400 15257
rect 12000 15200 12400 15223
rect 8480 15097 8880 15120
rect 8480 15063 8503 15097
rect 8537 15063 8663 15097
rect 8697 15063 8823 15097
rect 8857 15063 8880 15097
rect 8480 15040 8880 15063
rect 8960 15097 9360 15120
rect 8960 15063 8983 15097
rect 9017 15063 9143 15097
rect 9177 15063 9303 15097
rect 9337 15063 9360 15097
rect 8960 15040 9360 15063
rect 9440 15097 11440 15120
rect 9440 15063 9463 15097
rect 9497 15063 9623 15097
rect 9657 15063 9783 15097
rect 9817 15063 9943 15097
rect 9977 15063 10103 15097
rect 10137 15063 10263 15097
rect 10297 15063 10423 15097
rect 10457 15063 10583 15097
rect 10617 15063 10743 15097
rect 10777 15063 10903 15097
rect 10937 15063 11063 15097
rect 11097 15063 11223 15097
rect 11257 15063 11383 15097
rect 11417 15063 11440 15097
rect 9440 15040 11440 15063
rect 11520 15097 11920 15120
rect 11520 15063 11543 15097
rect 11577 15063 11703 15097
rect 11737 15063 11863 15097
rect 11897 15063 11920 15097
rect 11520 15040 11920 15063
rect 12000 15097 12400 15120
rect 12000 15063 12023 15097
rect 12057 15063 12183 15097
rect 12217 15063 12343 15097
rect 12377 15063 12400 15097
rect 12000 15040 12400 15063
rect 8480 14937 8880 14960
rect 8480 14903 8503 14937
rect 8537 14903 8663 14937
rect 8697 14903 8823 14937
rect 8857 14903 8880 14937
rect 8480 14880 8880 14903
rect 8960 14937 9360 14960
rect 8960 14903 8983 14937
rect 9017 14903 9143 14937
rect 9177 14903 9303 14937
rect 9337 14903 9360 14937
rect 8960 14880 9360 14903
rect 9440 14937 11440 14960
rect 9440 14903 9463 14937
rect 9497 14903 9623 14937
rect 9657 14903 9783 14937
rect 9817 14903 9943 14937
rect 9977 14903 10103 14937
rect 10137 14903 10263 14937
rect 10297 14903 10423 14937
rect 10457 14903 10583 14937
rect 10617 14903 10743 14937
rect 10777 14903 10903 14937
rect 10937 14903 11063 14937
rect 11097 14903 11223 14937
rect 11257 14903 11383 14937
rect 11417 14903 11440 14937
rect 9440 14880 11440 14903
rect 11520 14937 11920 14960
rect 11520 14903 11543 14937
rect 11577 14903 11703 14937
rect 11737 14903 11863 14937
rect 11897 14903 11920 14937
rect 11520 14880 11920 14903
rect 12000 14937 12400 14960
rect 12000 14903 12023 14937
rect 12057 14903 12183 14937
rect 12217 14903 12343 14937
rect 12377 14903 12400 14937
rect 12000 14880 12400 14903
rect 8480 14777 8880 14800
rect 8480 14743 8503 14777
rect 8537 14743 8663 14777
rect 8697 14743 8823 14777
rect 8857 14743 8880 14777
rect 8480 14720 8880 14743
rect 8960 14777 9360 14800
rect 8960 14743 8983 14777
rect 9017 14743 9143 14777
rect 9177 14743 9303 14777
rect 9337 14743 9360 14777
rect 8960 14720 9360 14743
rect 9440 14777 11440 14800
rect 9440 14743 9463 14777
rect 9497 14743 9623 14777
rect 9657 14743 9783 14777
rect 9817 14743 9943 14777
rect 9977 14743 10103 14777
rect 10137 14743 10263 14777
rect 10297 14743 10423 14777
rect 10457 14743 10583 14777
rect 10617 14743 10743 14777
rect 10777 14743 10903 14777
rect 10937 14743 11063 14777
rect 11097 14743 11223 14777
rect 11257 14743 11383 14777
rect 11417 14743 11440 14777
rect 9440 14720 11440 14743
rect 11520 14777 11920 14800
rect 11520 14743 11543 14777
rect 11577 14743 11703 14777
rect 11737 14743 11863 14777
rect 11897 14743 11920 14777
rect 11520 14720 11920 14743
rect 12000 14777 12400 14800
rect 12000 14743 12023 14777
rect 12057 14743 12183 14777
rect 12217 14743 12343 14777
rect 12377 14743 12400 14777
rect 12000 14720 12400 14743
rect 8480 14617 8880 14640
rect 8480 14583 8503 14617
rect 8537 14583 8663 14617
rect 8697 14583 8823 14617
rect 8857 14583 8880 14617
rect 8480 14560 8880 14583
rect 8960 14617 9360 14640
rect 8960 14583 8983 14617
rect 9017 14583 9143 14617
rect 9177 14583 9303 14617
rect 9337 14583 9360 14617
rect 8960 14560 9360 14583
rect 9440 14617 11440 14640
rect 9440 14583 9463 14617
rect 9497 14583 9623 14617
rect 9657 14583 9783 14617
rect 9817 14583 9943 14617
rect 9977 14583 10103 14617
rect 10137 14583 10263 14617
rect 10297 14583 10423 14617
rect 10457 14583 10583 14617
rect 10617 14583 10743 14617
rect 10777 14583 10903 14617
rect 10937 14583 11063 14617
rect 11097 14583 11223 14617
rect 11257 14583 11383 14617
rect 11417 14583 11440 14617
rect 9440 14560 11440 14583
rect 11520 14617 11920 14640
rect 11520 14583 11543 14617
rect 11577 14583 11703 14617
rect 11737 14583 11863 14617
rect 11897 14583 11920 14617
rect 11520 14560 11920 14583
rect 12000 14617 12400 14640
rect 12000 14583 12023 14617
rect 12057 14583 12183 14617
rect 12217 14583 12343 14617
rect 12377 14583 12400 14617
rect 12000 14560 12400 14583
rect 8480 14457 8880 14480
rect 8480 14423 8503 14457
rect 8537 14423 8663 14457
rect 8697 14423 8823 14457
rect 8857 14423 8880 14457
rect 8480 14400 8880 14423
rect 8960 14457 9360 14480
rect 8960 14423 8983 14457
rect 9017 14423 9143 14457
rect 9177 14423 9303 14457
rect 9337 14423 9360 14457
rect 8960 14400 9360 14423
rect 9440 14457 11440 14480
rect 9440 14423 9463 14457
rect 9497 14423 9623 14457
rect 9657 14423 9783 14457
rect 9817 14423 9943 14457
rect 9977 14423 10103 14457
rect 10137 14423 10263 14457
rect 10297 14423 10423 14457
rect 10457 14423 10583 14457
rect 10617 14423 10743 14457
rect 10777 14423 10903 14457
rect 10937 14423 11063 14457
rect 11097 14423 11223 14457
rect 11257 14423 11383 14457
rect 11417 14423 11440 14457
rect 9440 14400 11440 14423
rect 11520 14457 11920 14480
rect 11520 14423 11543 14457
rect 11577 14423 11703 14457
rect 11737 14423 11863 14457
rect 11897 14423 11920 14457
rect 11520 14400 11920 14423
rect 12000 14457 12400 14480
rect 12000 14423 12023 14457
rect 12057 14423 12183 14457
rect 12217 14423 12343 14457
rect 12377 14423 12400 14457
rect 12000 14400 12400 14423
rect 8480 14297 8880 14320
rect 8480 14263 8503 14297
rect 8537 14263 8663 14297
rect 8697 14263 8823 14297
rect 8857 14263 8880 14297
rect 8480 14240 8880 14263
rect 8960 14297 9360 14320
rect 8960 14263 8983 14297
rect 9017 14263 9143 14297
rect 9177 14263 9303 14297
rect 9337 14263 9360 14297
rect 8960 14240 9360 14263
rect 9440 14297 11440 14320
rect 9440 14263 9463 14297
rect 9497 14263 9623 14297
rect 9657 14263 9783 14297
rect 9817 14263 9943 14297
rect 9977 14263 10103 14297
rect 10137 14263 10263 14297
rect 10297 14263 10423 14297
rect 10457 14263 10583 14297
rect 10617 14263 10743 14297
rect 10777 14263 10903 14297
rect 10937 14263 11063 14297
rect 11097 14263 11223 14297
rect 11257 14263 11383 14297
rect 11417 14263 11440 14297
rect 9440 14240 11440 14263
rect 11520 14297 11920 14320
rect 11520 14263 11543 14297
rect 11577 14263 11703 14297
rect 11737 14263 11863 14297
rect 11897 14263 11920 14297
rect 11520 14240 11920 14263
rect 12000 14297 12400 14320
rect 12000 14263 12023 14297
rect 12057 14263 12183 14297
rect 12217 14263 12343 14297
rect 12377 14263 12400 14297
rect 12000 14240 12400 14263
rect 8480 14137 8880 14160
rect 8480 14103 8503 14137
rect 8537 14103 8663 14137
rect 8697 14103 8823 14137
rect 8857 14103 8880 14137
rect 8480 14080 8880 14103
rect 8960 14137 9360 14160
rect 8960 14103 8983 14137
rect 9017 14103 9143 14137
rect 9177 14103 9303 14137
rect 9337 14103 9360 14137
rect 8960 14080 9360 14103
rect 9440 14137 11440 14160
rect 9440 14103 9463 14137
rect 9497 14103 9623 14137
rect 9657 14103 9783 14137
rect 9817 14103 9943 14137
rect 9977 14103 10103 14137
rect 10137 14103 10263 14137
rect 10297 14103 10423 14137
rect 10457 14103 10583 14137
rect 10617 14103 10743 14137
rect 10777 14103 10903 14137
rect 10937 14103 11063 14137
rect 11097 14103 11223 14137
rect 11257 14103 11383 14137
rect 11417 14103 11440 14137
rect 9440 14080 11440 14103
rect 11520 14137 11920 14160
rect 11520 14103 11543 14137
rect 11577 14103 11703 14137
rect 11737 14103 11863 14137
rect 11897 14103 11920 14137
rect 11520 14080 11920 14103
rect 12000 14137 12400 14160
rect 12000 14103 12023 14137
rect 12057 14103 12183 14137
rect 12217 14103 12343 14137
rect 12377 14103 12400 14137
rect 12000 14080 12400 14103
rect 8480 13977 8880 14000
rect 8480 13943 8503 13977
rect 8537 13943 8663 13977
rect 8697 13943 8823 13977
rect 8857 13943 8880 13977
rect 8480 13920 8880 13943
rect 8960 13977 9360 14000
rect 8960 13943 8983 13977
rect 9017 13943 9143 13977
rect 9177 13943 9303 13977
rect 9337 13943 9360 13977
rect 8960 13920 9360 13943
rect 9440 13977 11440 14000
rect 9440 13943 9463 13977
rect 9497 13943 9623 13977
rect 9657 13943 9783 13977
rect 9817 13943 9943 13977
rect 9977 13943 10103 13977
rect 10137 13943 10263 13977
rect 10297 13943 10423 13977
rect 10457 13943 10583 13977
rect 10617 13943 10743 13977
rect 10777 13943 10903 13977
rect 10937 13943 11063 13977
rect 11097 13943 11223 13977
rect 11257 13943 11383 13977
rect 11417 13943 11440 13977
rect 9440 13920 11440 13943
rect 11520 13977 11920 14000
rect 11520 13943 11543 13977
rect 11577 13943 11703 13977
rect 11737 13943 11863 13977
rect 11897 13943 11920 13977
rect 11520 13920 11920 13943
rect 12000 13977 12400 14000
rect 12000 13943 12023 13977
rect 12057 13943 12183 13977
rect 12217 13943 12343 13977
rect 12377 13943 12400 13977
rect 12000 13920 12400 13943
rect 8480 13817 8880 13840
rect 8480 13783 8503 13817
rect 8537 13783 8663 13817
rect 8697 13783 8823 13817
rect 8857 13783 8880 13817
rect 8480 13760 8880 13783
rect 8960 13817 9360 13840
rect 8960 13783 8983 13817
rect 9017 13783 9143 13817
rect 9177 13783 9303 13817
rect 9337 13783 9360 13817
rect 8960 13760 9360 13783
rect 9440 13817 11440 13840
rect 9440 13783 9463 13817
rect 9497 13783 9623 13817
rect 9657 13783 9783 13817
rect 9817 13783 9943 13817
rect 9977 13783 10103 13817
rect 10137 13783 10263 13817
rect 10297 13783 10423 13817
rect 10457 13783 10583 13817
rect 10617 13783 10743 13817
rect 10777 13783 10903 13817
rect 10937 13783 11063 13817
rect 11097 13783 11223 13817
rect 11257 13783 11383 13817
rect 11417 13783 11440 13817
rect 9440 13760 11440 13783
rect 11520 13817 11920 13840
rect 11520 13783 11543 13817
rect 11577 13783 11703 13817
rect 11737 13783 11863 13817
rect 11897 13783 11920 13817
rect 11520 13760 11920 13783
rect 12000 13817 12400 13840
rect 12000 13783 12023 13817
rect 12057 13783 12183 13817
rect 12217 13783 12343 13817
rect 12377 13783 12400 13817
rect 12000 13760 12400 13783
rect 8480 13657 8880 13680
rect 8480 13623 8503 13657
rect 8537 13623 8663 13657
rect 8697 13623 8823 13657
rect 8857 13623 8880 13657
rect 8480 13600 8880 13623
rect 8960 13657 9360 13680
rect 8960 13623 8983 13657
rect 9017 13623 9143 13657
rect 9177 13623 9303 13657
rect 9337 13623 9360 13657
rect 8960 13600 9360 13623
rect 9440 13657 11440 13680
rect 9440 13623 9463 13657
rect 9497 13623 9623 13657
rect 9657 13623 9783 13657
rect 9817 13623 9943 13657
rect 9977 13623 10103 13657
rect 10137 13623 10263 13657
rect 10297 13623 10423 13657
rect 10457 13623 10583 13657
rect 10617 13623 10743 13657
rect 10777 13623 10903 13657
rect 10937 13623 11063 13657
rect 11097 13623 11223 13657
rect 11257 13623 11383 13657
rect 11417 13623 11440 13657
rect 9440 13600 11440 13623
rect 11520 13657 11920 13680
rect 11520 13623 11543 13657
rect 11577 13623 11703 13657
rect 11737 13623 11863 13657
rect 11897 13623 11920 13657
rect 11520 13600 11920 13623
rect 12000 13657 12400 13680
rect 12000 13623 12023 13657
rect 12057 13623 12183 13657
rect 12217 13623 12343 13657
rect 12377 13623 12400 13657
rect 12000 13600 12400 13623
rect 8480 13497 8880 13520
rect 8480 13463 8503 13497
rect 8537 13463 8663 13497
rect 8697 13463 8823 13497
rect 8857 13463 8880 13497
rect 8480 13440 8880 13463
rect 8960 13497 9360 13520
rect 8960 13463 8983 13497
rect 9017 13463 9143 13497
rect 9177 13463 9303 13497
rect 9337 13463 9360 13497
rect 8960 13440 9360 13463
rect 9440 13497 11440 13520
rect 9440 13463 9463 13497
rect 9497 13463 9623 13497
rect 9657 13463 9783 13497
rect 9817 13463 9943 13497
rect 9977 13463 10103 13497
rect 10137 13463 10263 13497
rect 10297 13463 10423 13497
rect 10457 13463 10583 13497
rect 10617 13463 10743 13497
rect 10777 13463 10903 13497
rect 10937 13463 11063 13497
rect 11097 13463 11223 13497
rect 11257 13463 11383 13497
rect 11417 13463 11440 13497
rect 9440 13440 11440 13463
rect 11520 13497 11920 13520
rect 11520 13463 11543 13497
rect 11577 13463 11703 13497
rect 11737 13463 11863 13497
rect 11897 13463 11920 13497
rect 11520 13440 11920 13463
rect 12000 13497 12400 13520
rect 12000 13463 12023 13497
rect 12057 13463 12183 13497
rect 12217 13463 12343 13497
rect 12377 13463 12400 13497
rect 12000 13440 12400 13463
rect 8480 13337 8880 13360
rect 8480 13303 8503 13337
rect 8537 13303 8663 13337
rect 8697 13303 8823 13337
rect 8857 13303 8880 13337
rect 8480 13280 8880 13303
rect 8960 13337 9360 13360
rect 8960 13303 8983 13337
rect 9017 13303 9143 13337
rect 9177 13303 9303 13337
rect 9337 13303 9360 13337
rect 8960 13280 9360 13303
rect 9440 13337 11440 13360
rect 9440 13303 9463 13337
rect 9497 13303 9623 13337
rect 9657 13303 9783 13337
rect 9817 13303 9943 13337
rect 9977 13303 10103 13337
rect 10137 13303 10263 13337
rect 10297 13303 10423 13337
rect 10457 13303 10583 13337
rect 10617 13303 10743 13337
rect 10777 13303 10903 13337
rect 10937 13303 11063 13337
rect 11097 13303 11223 13337
rect 11257 13303 11383 13337
rect 11417 13303 11440 13337
rect 9440 13280 11440 13303
rect 11520 13337 11920 13360
rect 11520 13303 11543 13337
rect 11577 13303 11703 13337
rect 11737 13303 11863 13337
rect 11897 13303 11920 13337
rect 11520 13280 11920 13303
rect 12000 13337 12400 13360
rect 12000 13303 12023 13337
rect 12057 13303 12183 13337
rect 12217 13303 12343 13337
rect 12377 13303 12400 13337
rect 12000 13280 12400 13303
rect 8480 13177 8880 13200
rect 8480 13143 8503 13177
rect 8537 13143 8663 13177
rect 8697 13143 8823 13177
rect 8857 13143 8880 13177
rect 8480 13120 8880 13143
rect 8960 13177 9360 13200
rect 8960 13143 8983 13177
rect 9017 13143 9143 13177
rect 9177 13143 9303 13177
rect 9337 13143 9360 13177
rect 8960 13120 9360 13143
rect 9440 13177 11440 13200
rect 9440 13143 9463 13177
rect 9497 13143 9623 13177
rect 9657 13143 9783 13177
rect 9817 13143 9943 13177
rect 9977 13143 10103 13177
rect 10137 13143 10263 13177
rect 10297 13143 10423 13177
rect 10457 13143 10583 13177
rect 10617 13143 10743 13177
rect 10777 13143 10903 13177
rect 10937 13143 11063 13177
rect 11097 13143 11223 13177
rect 11257 13143 11383 13177
rect 11417 13143 11440 13177
rect 9440 13120 11440 13143
rect 11520 13177 11920 13200
rect 11520 13143 11543 13177
rect 11577 13143 11703 13177
rect 11737 13143 11863 13177
rect 11897 13143 11920 13177
rect 11520 13120 11920 13143
rect 12000 13177 12400 13200
rect 12000 13143 12023 13177
rect 12057 13143 12183 13177
rect 12217 13143 12343 13177
rect 12377 13143 12400 13177
rect 12000 13120 12400 13143
rect 8480 13017 8880 13040
rect 8480 12983 8503 13017
rect 8537 12983 8663 13017
rect 8697 12983 8823 13017
rect 8857 12983 8880 13017
rect 8480 12960 8880 12983
rect 8960 13017 9360 13040
rect 8960 12983 8983 13017
rect 9017 12983 9143 13017
rect 9177 12983 9303 13017
rect 9337 12983 9360 13017
rect 8960 12960 9360 12983
rect 9440 13017 11440 13040
rect 9440 12983 9463 13017
rect 9497 12983 9623 13017
rect 9657 12983 9783 13017
rect 9817 12983 9943 13017
rect 9977 12983 10103 13017
rect 10137 12983 10263 13017
rect 10297 12983 10423 13017
rect 10457 12983 10583 13017
rect 10617 12983 10743 13017
rect 10777 12983 10903 13017
rect 10937 12983 11063 13017
rect 11097 12983 11223 13017
rect 11257 12983 11383 13017
rect 11417 12983 11440 13017
rect 9440 12960 11440 12983
rect 11520 13017 11920 13040
rect 11520 12983 11543 13017
rect 11577 12983 11703 13017
rect 11737 12983 11863 13017
rect 11897 12983 11920 13017
rect 11520 12960 11920 12983
rect 12000 13017 12400 13040
rect 12000 12983 12023 13017
rect 12057 12983 12183 13017
rect 12217 12983 12343 13017
rect 12377 12983 12400 13017
rect 12000 12960 12400 12983
rect 8480 12857 8880 12880
rect 8480 12823 8503 12857
rect 8537 12823 8663 12857
rect 8697 12823 8823 12857
rect 8857 12823 8880 12857
rect 8480 12800 8880 12823
rect 8960 12857 9360 12880
rect 8960 12823 8983 12857
rect 9017 12823 9143 12857
rect 9177 12823 9303 12857
rect 9337 12823 9360 12857
rect 8960 12800 9360 12823
rect 9440 12857 11440 12880
rect 9440 12823 9463 12857
rect 9497 12823 9623 12857
rect 9657 12823 9783 12857
rect 9817 12823 9943 12857
rect 9977 12823 10103 12857
rect 10137 12823 10263 12857
rect 10297 12823 10423 12857
rect 10457 12823 10583 12857
rect 10617 12823 10743 12857
rect 10777 12823 10903 12857
rect 10937 12823 11063 12857
rect 11097 12823 11223 12857
rect 11257 12823 11383 12857
rect 11417 12823 11440 12857
rect 9440 12800 11440 12823
rect 11520 12857 11920 12880
rect 11520 12823 11543 12857
rect 11577 12823 11703 12857
rect 11737 12823 11863 12857
rect 11897 12823 11920 12857
rect 11520 12800 11920 12823
rect 12000 12857 12400 12880
rect 12000 12823 12023 12857
rect 12057 12823 12183 12857
rect 12217 12823 12343 12857
rect 12377 12823 12400 12857
rect 12000 12800 12400 12823
rect 8480 12697 8880 12720
rect 8480 12663 8503 12697
rect 8537 12663 8663 12697
rect 8697 12663 8823 12697
rect 8857 12663 8880 12697
rect 8480 12640 8880 12663
rect 8960 12697 9360 12720
rect 8960 12663 8983 12697
rect 9017 12663 9143 12697
rect 9177 12663 9303 12697
rect 9337 12663 9360 12697
rect 8960 12640 9360 12663
rect 9440 12697 11440 12720
rect 9440 12663 9463 12697
rect 9497 12663 9623 12697
rect 9657 12663 9783 12697
rect 9817 12663 9943 12697
rect 9977 12663 10103 12697
rect 10137 12663 10263 12697
rect 10297 12663 10423 12697
rect 10457 12663 10583 12697
rect 10617 12663 10743 12697
rect 10777 12663 10903 12697
rect 10937 12663 11063 12697
rect 11097 12663 11223 12697
rect 11257 12663 11383 12697
rect 11417 12663 11440 12697
rect 9440 12640 11440 12663
rect 11520 12697 11920 12720
rect 11520 12663 11543 12697
rect 11577 12663 11703 12697
rect 11737 12663 11863 12697
rect 11897 12663 11920 12697
rect 11520 12640 11920 12663
rect 12000 12697 12400 12720
rect 12000 12663 12023 12697
rect 12057 12663 12183 12697
rect 12217 12663 12343 12697
rect 12377 12663 12400 12697
rect 12000 12640 12400 12663
rect 8480 12537 8880 12560
rect 8480 12503 8503 12537
rect 8537 12503 8663 12537
rect 8697 12503 8823 12537
rect 8857 12503 8880 12537
rect 8480 12480 8880 12503
rect 8960 12537 9360 12560
rect 8960 12503 8983 12537
rect 9017 12503 9143 12537
rect 9177 12503 9303 12537
rect 9337 12503 9360 12537
rect 8960 12480 9360 12503
rect 9440 12537 11440 12560
rect 9440 12503 9463 12537
rect 9497 12503 9623 12537
rect 9657 12503 9783 12537
rect 9817 12503 9943 12537
rect 9977 12503 10103 12537
rect 10137 12503 10263 12537
rect 10297 12503 10423 12537
rect 10457 12503 10583 12537
rect 10617 12503 10743 12537
rect 10777 12503 10903 12537
rect 10937 12503 11063 12537
rect 11097 12503 11223 12537
rect 11257 12503 11383 12537
rect 11417 12503 11440 12537
rect 9440 12480 11440 12503
rect 11520 12537 11920 12560
rect 11520 12503 11543 12537
rect 11577 12503 11703 12537
rect 11737 12503 11863 12537
rect 11897 12503 11920 12537
rect 11520 12480 11920 12503
rect 12000 12537 12400 12560
rect 12000 12503 12023 12537
rect 12057 12503 12183 12537
rect 12217 12503 12343 12537
rect 12377 12503 12400 12537
rect 12000 12480 12400 12503
rect 8480 12377 8880 12400
rect 8480 12343 8503 12377
rect 8537 12343 8663 12377
rect 8697 12343 8823 12377
rect 8857 12343 8880 12377
rect 8480 12320 8880 12343
rect 8960 12377 9360 12400
rect 8960 12343 8983 12377
rect 9017 12343 9143 12377
rect 9177 12343 9303 12377
rect 9337 12343 9360 12377
rect 8960 12320 9360 12343
rect 9440 12377 11440 12400
rect 9440 12343 9463 12377
rect 9497 12343 9623 12377
rect 9657 12343 9783 12377
rect 9817 12343 9943 12377
rect 9977 12343 10103 12377
rect 10137 12343 10263 12377
rect 10297 12343 10423 12377
rect 10457 12343 10583 12377
rect 10617 12343 10743 12377
rect 10777 12343 10903 12377
rect 10937 12343 11063 12377
rect 11097 12343 11223 12377
rect 11257 12343 11383 12377
rect 11417 12343 11440 12377
rect 9440 12320 11440 12343
rect 11520 12377 11920 12400
rect 11520 12343 11543 12377
rect 11577 12343 11703 12377
rect 11737 12343 11863 12377
rect 11897 12343 11920 12377
rect 11520 12320 11920 12343
rect 12000 12377 12400 12400
rect 12000 12343 12023 12377
rect 12057 12343 12183 12377
rect 12217 12343 12343 12377
rect 12377 12343 12400 12377
rect 12000 12320 12400 12343
rect 8480 12217 8880 12240
rect 8480 12183 8503 12217
rect 8537 12183 8663 12217
rect 8697 12183 8823 12217
rect 8857 12183 8880 12217
rect 8480 12160 8880 12183
rect 8960 12217 9360 12240
rect 8960 12183 8983 12217
rect 9017 12183 9143 12217
rect 9177 12183 9303 12217
rect 9337 12183 9360 12217
rect 8960 12160 9360 12183
rect 9440 12217 11440 12240
rect 9440 12183 9463 12217
rect 9497 12183 9623 12217
rect 9657 12183 9783 12217
rect 9817 12183 9943 12217
rect 9977 12183 10103 12217
rect 10137 12183 10263 12217
rect 10297 12183 10423 12217
rect 10457 12183 10583 12217
rect 10617 12183 10743 12217
rect 10777 12183 10903 12217
rect 10937 12183 11063 12217
rect 11097 12183 11223 12217
rect 11257 12183 11383 12217
rect 11417 12183 11440 12217
rect 9440 12160 11440 12183
rect 11520 12217 11920 12240
rect 11520 12183 11543 12217
rect 11577 12183 11703 12217
rect 11737 12183 11863 12217
rect 11897 12183 11920 12217
rect 11520 12160 11920 12183
rect 12000 12217 12400 12240
rect 12000 12183 12023 12217
rect 12057 12183 12183 12217
rect 12217 12183 12343 12217
rect 12377 12183 12400 12217
rect 12000 12160 12400 12183
rect 8480 12057 8880 12080
rect 8480 12023 8503 12057
rect 8537 12023 8663 12057
rect 8697 12023 8823 12057
rect 8857 12023 8880 12057
rect 8480 12000 8880 12023
rect 8960 12057 9360 12080
rect 8960 12023 8983 12057
rect 9017 12023 9143 12057
rect 9177 12023 9303 12057
rect 9337 12023 9360 12057
rect 8960 12000 9360 12023
rect 9440 12057 11440 12080
rect 9440 12023 9463 12057
rect 9497 12023 9623 12057
rect 9657 12023 9783 12057
rect 9817 12023 9943 12057
rect 9977 12023 10103 12057
rect 10137 12023 10263 12057
rect 10297 12023 10423 12057
rect 10457 12023 10583 12057
rect 10617 12023 10743 12057
rect 10777 12023 10903 12057
rect 10937 12023 11063 12057
rect 11097 12023 11223 12057
rect 11257 12023 11383 12057
rect 11417 12023 11440 12057
rect 9440 12000 11440 12023
rect 11520 12057 11920 12080
rect 11520 12023 11543 12057
rect 11577 12023 11703 12057
rect 11737 12023 11863 12057
rect 11897 12023 11920 12057
rect 11520 12000 11920 12023
rect 12000 12057 12400 12080
rect 12000 12023 12023 12057
rect 12057 12023 12183 12057
rect 12217 12023 12343 12057
rect 12377 12023 12400 12057
rect 12000 12000 12400 12023
rect 8480 11897 8880 11920
rect 8480 11863 8503 11897
rect 8537 11863 8663 11897
rect 8697 11863 8823 11897
rect 8857 11863 8880 11897
rect 8480 11840 8880 11863
rect 8960 11897 9360 11920
rect 8960 11863 8983 11897
rect 9017 11863 9143 11897
rect 9177 11863 9303 11897
rect 9337 11863 9360 11897
rect 8960 11840 9360 11863
rect 9440 11897 11440 11920
rect 9440 11863 9463 11897
rect 9497 11863 9623 11897
rect 9657 11863 9783 11897
rect 9817 11863 9943 11897
rect 9977 11863 10103 11897
rect 10137 11863 10263 11897
rect 10297 11863 10423 11897
rect 10457 11863 10583 11897
rect 10617 11863 10743 11897
rect 10777 11863 10903 11897
rect 10937 11863 11063 11897
rect 11097 11863 11223 11897
rect 11257 11863 11383 11897
rect 11417 11863 11440 11897
rect 9440 11840 11440 11863
rect 11520 11897 11920 11920
rect 11520 11863 11543 11897
rect 11577 11863 11703 11897
rect 11737 11863 11863 11897
rect 11897 11863 11920 11897
rect 11520 11840 11920 11863
rect 12000 11897 12400 11920
rect 12000 11863 12023 11897
rect 12057 11863 12183 11897
rect 12217 11863 12343 11897
rect 12377 11863 12400 11897
rect 12000 11840 12400 11863
rect 8480 11737 8880 11760
rect 8480 11703 8503 11737
rect 8537 11703 8663 11737
rect 8697 11703 8823 11737
rect 8857 11703 8880 11737
rect 8480 11680 8880 11703
rect 8960 11737 9360 11760
rect 8960 11703 8983 11737
rect 9017 11703 9143 11737
rect 9177 11703 9303 11737
rect 9337 11703 9360 11737
rect 8960 11680 9360 11703
rect 9440 11737 11440 11760
rect 9440 11703 9463 11737
rect 9497 11703 9623 11737
rect 9657 11703 9783 11737
rect 9817 11703 9943 11737
rect 9977 11703 10103 11737
rect 10137 11703 10263 11737
rect 10297 11703 10423 11737
rect 10457 11703 10583 11737
rect 10617 11703 10743 11737
rect 10777 11703 10903 11737
rect 10937 11703 11063 11737
rect 11097 11703 11223 11737
rect 11257 11703 11383 11737
rect 11417 11703 11440 11737
rect 9440 11680 11440 11703
rect 11520 11737 11920 11760
rect 11520 11703 11543 11737
rect 11577 11703 11703 11737
rect 11737 11703 11863 11737
rect 11897 11703 11920 11737
rect 11520 11680 11920 11703
rect 12000 11737 12400 11760
rect 12000 11703 12023 11737
rect 12057 11703 12183 11737
rect 12217 11703 12343 11737
rect 12377 11703 12400 11737
rect 12000 11680 12400 11703
rect 8480 11577 8880 11600
rect 8480 11543 8503 11577
rect 8537 11543 8663 11577
rect 8697 11543 8823 11577
rect 8857 11543 8880 11577
rect 8480 11520 8880 11543
rect 8960 11577 9360 11600
rect 8960 11543 8983 11577
rect 9017 11543 9143 11577
rect 9177 11543 9303 11577
rect 9337 11543 9360 11577
rect 8960 11520 9360 11543
rect 9440 11577 11440 11600
rect 9440 11543 9463 11577
rect 9497 11543 9623 11577
rect 9657 11543 9783 11577
rect 9817 11543 9943 11577
rect 9977 11543 10103 11577
rect 10137 11543 10263 11577
rect 10297 11543 10423 11577
rect 10457 11543 10583 11577
rect 10617 11543 10743 11577
rect 10777 11543 10903 11577
rect 10937 11543 11063 11577
rect 11097 11543 11223 11577
rect 11257 11543 11383 11577
rect 11417 11543 11440 11577
rect 9440 11520 11440 11543
rect 11520 11577 11920 11600
rect 11520 11543 11543 11577
rect 11577 11543 11703 11577
rect 11737 11543 11863 11577
rect 11897 11543 11920 11577
rect 11520 11520 11920 11543
rect 12000 11577 12400 11600
rect 12000 11543 12023 11577
rect 12057 11543 12183 11577
rect 12217 11543 12343 11577
rect 12377 11543 12400 11577
rect 12000 11520 12400 11543
rect 8480 11417 8880 11440
rect 8480 11383 8503 11417
rect 8537 11383 8663 11417
rect 8697 11383 8823 11417
rect 8857 11383 8880 11417
rect 8480 11360 8880 11383
rect 8960 11417 9360 11440
rect 8960 11383 8983 11417
rect 9017 11383 9143 11417
rect 9177 11383 9303 11417
rect 9337 11383 9360 11417
rect 8960 11360 9360 11383
rect 9440 11417 11440 11440
rect 9440 11383 9463 11417
rect 9497 11383 9623 11417
rect 9657 11383 9783 11417
rect 9817 11383 9943 11417
rect 9977 11383 10103 11417
rect 10137 11383 10263 11417
rect 10297 11383 10423 11417
rect 10457 11383 10583 11417
rect 10617 11383 10743 11417
rect 10777 11383 10903 11417
rect 10937 11383 11063 11417
rect 11097 11383 11223 11417
rect 11257 11383 11383 11417
rect 11417 11383 11440 11417
rect 9440 11360 11440 11383
rect 11520 11417 11920 11440
rect 11520 11383 11543 11417
rect 11577 11383 11703 11417
rect 11737 11383 11863 11417
rect 11897 11383 11920 11417
rect 11520 11360 11920 11383
rect 12000 11417 12400 11440
rect 12000 11383 12023 11417
rect 12057 11383 12183 11417
rect 12217 11383 12343 11417
rect 12377 11383 12400 11417
rect 12000 11360 12400 11383
rect 8480 11257 8880 11280
rect 8480 11223 8503 11257
rect 8537 11223 8663 11257
rect 8697 11223 8823 11257
rect 8857 11223 8880 11257
rect 8480 11200 8880 11223
rect 8960 11257 9360 11280
rect 8960 11223 8983 11257
rect 9017 11223 9143 11257
rect 9177 11223 9303 11257
rect 9337 11223 9360 11257
rect 8960 11200 9360 11223
rect 9440 11257 11440 11280
rect 9440 11223 9463 11257
rect 9497 11223 9623 11257
rect 9657 11223 9783 11257
rect 9817 11223 9943 11257
rect 9977 11223 10103 11257
rect 10137 11223 10263 11257
rect 10297 11223 10423 11257
rect 10457 11223 10583 11257
rect 10617 11223 10743 11257
rect 10777 11223 10903 11257
rect 10937 11223 11063 11257
rect 11097 11223 11223 11257
rect 11257 11223 11383 11257
rect 11417 11223 11440 11257
rect 9440 11200 11440 11223
rect 11520 11257 11920 11280
rect 11520 11223 11543 11257
rect 11577 11223 11703 11257
rect 11737 11223 11863 11257
rect 11897 11223 11920 11257
rect 11520 11200 11920 11223
rect 12000 11257 12400 11280
rect 12000 11223 12023 11257
rect 12057 11223 12183 11257
rect 12217 11223 12343 11257
rect 12377 11223 12400 11257
rect 12000 11200 12400 11223
rect 8480 11097 8880 11120
rect 8480 11063 8503 11097
rect 8537 11063 8663 11097
rect 8697 11063 8823 11097
rect 8857 11063 8880 11097
rect 8480 11040 8880 11063
rect 8960 11097 9360 11120
rect 8960 11063 8983 11097
rect 9017 11063 9143 11097
rect 9177 11063 9303 11097
rect 9337 11063 9360 11097
rect 8960 11040 9360 11063
rect 9440 11097 11440 11120
rect 9440 11063 9463 11097
rect 9497 11063 9623 11097
rect 9657 11063 9783 11097
rect 9817 11063 9943 11097
rect 9977 11063 10103 11097
rect 10137 11063 10263 11097
rect 10297 11063 10423 11097
rect 10457 11063 10583 11097
rect 10617 11063 10743 11097
rect 10777 11063 10903 11097
rect 10937 11063 11063 11097
rect 11097 11063 11223 11097
rect 11257 11063 11383 11097
rect 11417 11063 11440 11097
rect 9440 11040 11440 11063
rect 11520 11097 11920 11120
rect 11520 11063 11543 11097
rect 11577 11063 11703 11097
rect 11737 11063 11863 11097
rect 11897 11063 11920 11097
rect 11520 11040 11920 11063
rect 12000 11097 12400 11120
rect 12000 11063 12023 11097
rect 12057 11063 12183 11097
rect 12217 11063 12343 11097
rect 12377 11063 12400 11097
rect 12000 11040 12400 11063
rect 8480 10937 8880 10960
rect 8480 10903 8503 10937
rect 8537 10903 8663 10937
rect 8697 10903 8823 10937
rect 8857 10903 8880 10937
rect 8480 10880 8880 10903
rect 8960 10937 9360 10960
rect 8960 10903 8983 10937
rect 9017 10903 9143 10937
rect 9177 10903 9303 10937
rect 9337 10903 9360 10937
rect 8960 10880 9360 10903
rect 9440 10937 11440 10960
rect 9440 10903 9463 10937
rect 9497 10903 9623 10937
rect 9657 10903 9783 10937
rect 9817 10903 9943 10937
rect 9977 10903 10103 10937
rect 10137 10903 10263 10937
rect 10297 10903 10423 10937
rect 10457 10903 10583 10937
rect 10617 10903 10743 10937
rect 10777 10903 10903 10937
rect 10937 10903 11063 10937
rect 11097 10903 11223 10937
rect 11257 10903 11383 10937
rect 11417 10903 11440 10937
rect 9440 10880 11440 10903
rect 11520 10937 11920 10960
rect 11520 10903 11543 10937
rect 11577 10903 11703 10937
rect 11737 10903 11863 10937
rect 11897 10903 11920 10937
rect 11520 10880 11920 10903
rect 12000 10937 12400 10960
rect 12000 10903 12023 10937
rect 12057 10903 12183 10937
rect 12217 10903 12343 10937
rect 12377 10903 12400 10937
rect 12000 10880 12400 10903
rect 8480 10777 8880 10800
rect 8480 10743 8503 10777
rect 8537 10743 8663 10777
rect 8697 10743 8823 10777
rect 8857 10743 8880 10777
rect 8480 10720 8880 10743
rect 8960 10777 9360 10800
rect 8960 10743 8983 10777
rect 9017 10743 9143 10777
rect 9177 10743 9303 10777
rect 9337 10743 9360 10777
rect 8960 10720 9360 10743
rect 9440 10777 11440 10800
rect 9440 10743 9463 10777
rect 9497 10743 9623 10777
rect 9657 10743 9783 10777
rect 9817 10743 9943 10777
rect 9977 10743 10103 10777
rect 10137 10743 10263 10777
rect 10297 10743 10423 10777
rect 10457 10743 10583 10777
rect 10617 10743 10743 10777
rect 10777 10743 10903 10777
rect 10937 10743 11063 10777
rect 11097 10743 11223 10777
rect 11257 10743 11383 10777
rect 11417 10743 11440 10777
rect 9440 10720 11440 10743
rect 11520 10777 11920 10800
rect 11520 10743 11543 10777
rect 11577 10743 11703 10777
rect 11737 10743 11863 10777
rect 11897 10743 11920 10777
rect 11520 10720 11920 10743
rect 12000 10777 12400 10800
rect 12000 10743 12023 10777
rect 12057 10743 12183 10777
rect 12217 10743 12343 10777
rect 12377 10743 12400 10777
rect 12000 10720 12400 10743
rect 8480 10617 8880 10640
rect 8480 10583 8503 10617
rect 8537 10583 8663 10617
rect 8697 10583 8823 10617
rect 8857 10583 8880 10617
rect 8480 10560 8880 10583
rect 8960 10617 9360 10640
rect 8960 10583 8983 10617
rect 9017 10583 9143 10617
rect 9177 10583 9303 10617
rect 9337 10583 9360 10617
rect 8960 10560 9360 10583
rect 9440 10617 11440 10640
rect 9440 10583 9463 10617
rect 9497 10583 9623 10617
rect 9657 10583 9783 10617
rect 9817 10583 9943 10617
rect 9977 10583 10103 10617
rect 10137 10583 10263 10617
rect 10297 10583 10423 10617
rect 10457 10583 10583 10617
rect 10617 10583 10743 10617
rect 10777 10583 10903 10617
rect 10937 10583 11063 10617
rect 11097 10583 11223 10617
rect 11257 10583 11383 10617
rect 11417 10583 11440 10617
rect 9440 10560 11440 10583
rect 11520 10617 11920 10640
rect 11520 10583 11543 10617
rect 11577 10583 11703 10617
rect 11737 10583 11863 10617
rect 11897 10583 11920 10617
rect 11520 10560 11920 10583
rect 12000 10617 12400 10640
rect 12000 10583 12023 10617
rect 12057 10583 12183 10617
rect 12217 10583 12343 10617
rect 12377 10583 12400 10617
rect 12000 10560 12400 10583
rect 8480 10457 8880 10480
rect 8480 10423 8503 10457
rect 8537 10423 8663 10457
rect 8697 10423 8823 10457
rect 8857 10423 8880 10457
rect 8480 10400 8880 10423
rect 8960 10457 9360 10480
rect 8960 10423 8983 10457
rect 9017 10423 9143 10457
rect 9177 10423 9303 10457
rect 9337 10423 9360 10457
rect 8960 10400 9360 10423
rect 9440 10457 11440 10480
rect 9440 10423 9463 10457
rect 9497 10423 9623 10457
rect 9657 10423 9783 10457
rect 9817 10423 9943 10457
rect 9977 10423 10103 10457
rect 10137 10423 10263 10457
rect 10297 10423 10423 10457
rect 10457 10423 10583 10457
rect 10617 10423 10743 10457
rect 10777 10423 10903 10457
rect 10937 10423 11063 10457
rect 11097 10423 11223 10457
rect 11257 10423 11383 10457
rect 11417 10423 11440 10457
rect 9440 10400 11440 10423
rect 11520 10457 11920 10480
rect 11520 10423 11543 10457
rect 11577 10423 11703 10457
rect 11737 10423 11863 10457
rect 11897 10423 11920 10457
rect 11520 10400 11920 10423
rect 12000 10457 12400 10480
rect 12000 10423 12023 10457
rect 12057 10423 12183 10457
rect 12217 10423 12343 10457
rect 12377 10423 12400 10457
rect 12000 10400 12400 10423
rect 8480 10297 8880 10320
rect 8480 10263 8503 10297
rect 8537 10263 8663 10297
rect 8697 10263 8823 10297
rect 8857 10263 8880 10297
rect 8480 10240 8880 10263
rect 8960 10297 9360 10320
rect 8960 10263 8983 10297
rect 9017 10263 9143 10297
rect 9177 10263 9303 10297
rect 9337 10263 9360 10297
rect 8960 10240 9360 10263
rect 9440 10297 11440 10320
rect 9440 10263 9463 10297
rect 9497 10263 9623 10297
rect 9657 10263 9783 10297
rect 9817 10263 9943 10297
rect 9977 10263 10103 10297
rect 10137 10263 10263 10297
rect 10297 10263 10423 10297
rect 10457 10263 10583 10297
rect 10617 10263 10743 10297
rect 10777 10263 10903 10297
rect 10937 10263 11063 10297
rect 11097 10263 11223 10297
rect 11257 10263 11383 10297
rect 11417 10263 11440 10297
rect 9440 10240 11440 10263
rect 11520 10297 11920 10320
rect 11520 10263 11543 10297
rect 11577 10263 11703 10297
rect 11737 10263 11863 10297
rect 11897 10263 11920 10297
rect 11520 10240 11920 10263
rect 12000 10297 12400 10320
rect 12000 10263 12023 10297
rect 12057 10263 12183 10297
rect 12217 10263 12343 10297
rect 12377 10263 12400 10297
rect 12000 10240 12400 10263
rect 8480 10137 8880 10160
rect 8480 10103 8503 10137
rect 8537 10103 8663 10137
rect 8697 10103 8823 10137
rect 8857 10103 8880 10137
rect 8480 10080 8880 10103
rect 8960 10137 9360 10160
rect 8960 10103 8983 10137
rect 9017 10103 9143 10137
rect 9177 10103 9303 10137
rect 9337 10103 9360 10137
rect 8960 10080 9360 10103
rect 9440 10137 11440 10160
rect 9440 10103 9463 10137
rect 9497 10103 9623 10137
rect 9657 10103 9783 10137
rect 9817 10103 9943 10137
rect 9977 10103 10103 10137
rect 10137 10103 10263 10137
rect 10297 10103 10423 10137
rect 10457 10103 10583 10137
rect 10617 10103 10743 10137
rect 10777 10103 10903 10137
rect 10937 10103 11063 10137
rect 11097 10103 11223 10137
rect 11257 10103 11383 10137
rect 11417 10103 11440 10137
rect 9440 10080 11440 10103
rect 11520 10137 11920 10160
rect 11520 10103 11543 10137
rect 11577 10103 11703 10137
rect 11737 10103 11863 10137
rect 11897 10103 11920 10137
rect 11520 10080 11920 10103
rect 12000 10137 12400 10160
rect 12000 10103 12023 10137
rect 12057 10103 12183 10137
rect 12217 10103 12343 10137
rect 12377 10103 12400 10137
rect 12000 10080 12400 10103
rect 8480 9977 8880 10000
rect 8480 9943 8503 9977
rect 8537 9943 8663 9977
rect 8697 9943 8823 9977
rect 8857 9943 8880 9977
rect 8480 9920 8880 9943
rect 8960 9977 9360 10000
rect 8960 9943 8983 9977
rect 9017 9943 9143 9977
rect 9177 9943 9303 9977
rect 9337 9943 9360 9977
rect 8960 9920 9360 9943
rect 9440 9977 11440 10000
rect 9440 9943 9463 9977
rect 9497 9943 9623 9977
rect 9657 9943 9783 9977
rect 9817 9943 9943 9977
rect 9977 9943 10103 9977
rect 10137 9943 10263 9977
rect 10297 9943 10423 9977
rect 10457 9943 10583 9977
rect 10617 9943 10743 9977
rect 10777 9943 10903 9977
rect 10937 9943 11063 9977
rect 11097 9943 11223 9977
rect 11257 9943 11383 9977
rect 11417 9943 11440 9977
rect 9440 9920 11440 9943
rect 11520 9977 11920 10000
rect 11520 9943 11543 9977
rect 11577 9943 11703 9977
rect 11737 9943 11863 9977
rect 11897 9943 11920 9977
rect 11520 9920 11920 9943
rect 12000 9977 12400 10000
rect 12000 9943 12023 9977
rect 12057 9943 12183 9977
rect 12217 9943 12343 9977
rect 12377 9943 12400 9977
rect 12000 9920 12400 9943
rect 8480 9817 8880 9840
rect 8480 9783 8503 9817
rect 8537 9783 8663 9817
rect 8697 9783 8823 9817
rect 8857 9783 8880 9817
rect 8480 9760 8880 9783
rect 8960 9817 9360 9840
rect 8960 9783 8983 9817
rect 9017 9783 9143 9817
rect 9177 9783 9303 9817
rect 9337 9783 9360 9817
rect 8960 9760 9360 9783
rect 9440 9817 11440 9840
rect 9440 9783 9463 9817
rect 9497 9783 9623 9817
rect 9657 9783 9783 9817
rect 9817 9783 9943 9817
rect 9977 9783 10103 9817
rect 10137 9783 10263 9817
rect 10297 9783 10423 9817
rect 10457 9783 10583 9817
rect 10617 9783 10743 9817
rect 10777 9783 10903 9817
rect 10937 9783 11063 9817
rect 11097 9783 11223 9817
rect 11257 9783 11383 9817
rect 11417 9783 11440 9817
rect 9440 9760 11440 9783
rect 11520 9817 11920 9840
rect 11520 9783 11543 9817
rect 11577 9783 11703 9817
rect 11737 9783 11863 9817
rect 11897 9783 11920 9817
rect 11520 9760 11920 9783
rect 12000 9817 12400 9840
rect 12000 9783 12023 9817
rect 12057 9783 12183 9817
rect 12217 9783 12343 9817
rect 12377 9783 12400 9817
rect 12000 9760 12400 9783
rect 8480 9657 8880 9680
rect 8480 9623 8503 9657
rect 8537 9623 8663 9657
rect 8697 9623 8823 9657
rect 8857 9623 8880 9657
rect 8480 9600 8880 9623
rect 8960 9657 9360 9680
rect 8960 9623 8983 9657
rect 9017 9623 9143 9657
rect 9177 9623 9303 9657
rect 9337 9623 9360 9657
rect 8960 9600 9360 9623
rect 9440 9657 11440 9680
rect 9440 9623 9463 9657
rect 9497 9623 9623 9657
rect 9657 9623 9783 9657
rect 9817 9623 9943 9657
rect 9977 9623 10103 9657
rect 10137 9623 10263 9657
rect 10297 9623 10423 9657
rect 10457 9623 10583 9657
rect 10617 9623 10743 9657
rect 10777 9623 10903 9657
rect 10937 9623 11063 9657
rect 11097 9623 11223 9657
rect 11257 9623 11383 9657
rect 11417 9623 11440 9657
rect 9440 9600 11440 9623
rect 11520 9657 11920 9680
rect 11520 9623 11543 9657
rect 11577 9623 11703 9657
rect 11737 9623 11863 9657
rect 11897 9623 11920 9657
rect 11520 9600 11920 9623
rect 12000 9657 12400 9680
rect 12000 9623 12023 9657
rect 12057 9623 12183 9657
rect 12217 9623 12343 9657
rect 12377 9623 12400 9657
rect 12000 9600 12400 9623
rect 8480 9497 8880 9520
rect 8480 9463 8503 9497
rect 8537 9463 8663 9497
rect 8697 9463 8823 9497
rect 8857 9463 8880 9497
rect 8480 9440 8880 9463
rect 8960 9497 9360 9520
rect 8960 9463 8983 9497
rect 9017 9463 9143 9497
rect 9177 9463 9303 9497
rect 9337 9463 9360 9497
rect 8960 9440 9360 9463
rect 9440 9497 11440 9520
rect 9440 9463 9463 9497
rect 9497 9463 9623 9497
rect 9657 9463 9783 9497
rect 9817 9463 9943 9497
rect 9977 9463 10103 9497
rect 10137 9463 10263 9497
rect 10297 9463 10423 9497
rect 10457 9463 10583 9497
rect 10617 9463 10743 9497
rect 10777 9463 10903 9497
rect 10937 9463 11063 9497
rect 11097 9463 11223 9497
rect 11257 9463 11383 9497
rect 11417 9463 11440 9497
rect 9440 9440 11440 9463
rect 11520 9497 11920 9520
rect 11520 9463 11543 9497
rect 11577 9463 11703 9497
rect 11737 9463 11863 9497
rect 11897 9463 11920 9497
rect 11520 9440 11920 9463
rect 12000 9497 12400 9520
rect 12000 9463 12023 9497
rect 12057 9463 12183 9497
rect 12217 9463 12343 9497
rect 12377 9463 12400 9497
rect 12000 9440 12400 9463
rect 8480 9337 8880 9360
rect 8480 9303 8503 9337
rect 8537 9303 8663 9337
rect 8697 9303 8823 9337
rect 8857 9303 8880 9337
rect 8480 9280 8880 9303
rect 8960 9337 9360 9360
rect 8960 9303 8983 9337
rect 9017 9303 9143 9337
rect 9177 9303 9303 9337
rect 9337 9303 9360 9337
rect 8960 9280 9360 9303
rect 9440 9337 11440 9360
rect 9440 9303 9463 9337
rect 9497 9303 9623 9337
rect 9657 9303 9783 9337
rect 9817 9303 9943 9337
rect 9977 9303 10103 9337
rect 10137 9303 10263 9337
rect 10297 9303 10423 9337
rect 10457 9303 10583 9337
rect 10617 9303 10743 9337
rect 10777 9303 10903 9337
rect 10937 9303 11063 9337
rect 11097 9303 11223 9337
rect 11257 9303 11383 9337
rect 11417 9303 11440 9337
rect 9440 9280 11440 9303
rect 11520 9337 11920 9360
rect 11520 9303 11543 9337
rect 11577 9303 11703 9337
rect 11737 9303 11863 9337
rect 11897 9303 11920 9337
rect 11520 9280 11920 9303
rect 12000 9337 12400 9360
rect 12000 9303 12023 9337
rect 12057 9303 12183 9337
rect 12217 9303 12343 9337
rect 12377 9303 12400 9337
rect 12000 9280 12400 9303
rect 8480 9177 8880 9200
rect 8480 9143 8503 9177
rect 8537 9143 8663 9177
rect 8697 9143 8823 9177
rect 8857 9143 8880 9177
rect 8480 9120 8880 9143
rect 8960 9177 9360 9200
rect 8960 9143 8983 9177
rect 9017 9143 9143 9177
rect 9177 9143 9303 9177
rect 9337 9143 9360 9177
rect 8960 9120 9360 9143
rect 9440 9177 11440 9200
rect 9440 9143 9463 9177
rect 9497 9143 9623 9177
rect 9657 9143 9783 9177
rect 9817 9143 9943 9177
rect 9977 9143 10103 9177
rect 10137 9143 10263 9177
rect 10297 9143 10423 9177
rect 10457 9143 10583 9177
rect 10617 9143 10743 9177
rect 10777 9143 10903 9177
rect 10937 9143 11063 9177
rect 11097 9143 11223 9177
rect 11257 9143 11383 9177
rect 11417 9143 11440 9177
rect 9440 9120 11440 9143
rect 11520 9177 11920 9200
rect 11520 9143 11543 9177
rect 11577 9143 11703 9177
rect 11737 9143 11863 9177
rect 11897 9143 11920 9177
rect 11520 9120 11920 9143
rect 12000 9177 12400 9200
rect 12000 9143 12023 9177
rect 12057 9143 12183 9177
rect 12217 9143 12343 9177
rect 12377 9143 12400 9177
rect 12000 9120 12400 9143
rect 8480 9017 8880 9040
rect 8480 8983 8503 9017
rect 8537 8983 8663 9017
rect 8697 8983 8823 9017
rect 8857 8983 8880 9017
rect 8480 8960 8880 8983
rect 8960 9017 9360 9040
rect 8960 8983 8983 9017
rect 9017 8983 9143 9017
rect 9177 8983 9303 9017
rect 9337 8983 9360 9017
rect 8960 8960 9360 8983
rect 9440 9017 11440 9040
rect 9440 8983 9463 9017
rect 9497 8983 9623 9017
rect 9657 8983 9783 9017
rect 9817 8983 9943 9017
rect 9977 8983 10103 9017
rect 10137 8983 10263 9017
rect 10297 8983 10423 9017
rect 10457 8983 10583 9017
rect 10617 8983 10743 9017
rect 10777 8983 10903 9017
rect 10937 8983 11063 9017
rect 11097 8983 11223 9017
rect 11257 8983 11383 9017
rect 11417 8983 11440 9017
rect 9440 8960 11440 8983
rect 11520 9017 11920 9040
rect 11520 8983 11543 9017
rect 11577 8983 11703 9017
rect 11737 8983 11863 9017
rect 11897 8983 11920 9017
rect 11520 8960 11920 8983
rect 12000 9017 12400 9040
rect 12000 8983 12023 9017
rect 12057 8983 12183 9017
rect 12217 8983 12343 9017
rect 12377 8983 12400 9017
rect 12000 8960 12400 8983
rect 8480 8857 8880 8880
rect 8480 8823 8503 8857
rect 8537 8823 8663 8857
rect 8697 8823 8823 8857
rect 8857 8823 8880 8857
rect 8480 8800 8880 8823
rect 8960 8857 9360 8880
rect 8960 8823 8983 8857
rect 9017 8823 9143 8857
rect 9177 8823 9303 8857
rect 9337 8823 9360 8857
rect 8960 8800 9360 8823
rect 9440 8857 11440 8880
rect 9440 8823 9463 8857
rect 9497 8823 9623 8857
rect 9657 8823 9783 8857
rect 9817 8823 9943 8857
rect 9977 8823 10103 8857
rect 10137 8823 10263 8857
rect 10297 8823 10423 8857
rect 10457 8823 10583 8857
rect 10617 8823 10743 8857
rect 10777 8823 10903 8857
rect 10937 8823 11063 8857
rect 11097 8823 11223 8857
rect 11257 8823 11383 8857
rect 11417 8823 11440 8857
rect 9440 8800 11440 8823
rect 11520 8857 11920 8880
rect 11520 8823 11543 8857
rect 11577 8823 11703 8857
rect 11737 8823 11863 8857
rect 11897 8823 11920 8857
rect 11520 8800 11920 8823
rect 12000 8857 12400 8880
rect 12000 8823 12023 8857
rect 12057 8823 12183 8857
rect 12217 8823 12343 8857
rect 12377 8823 12400 8857
rect 12000 8800 12400 8823
rect 8480 8697 8880 8720
rect 8480 8663 8503 8697
rect 8537 8663 8663 8697
rect 8697 8663 8823 8697
rect 8857 8663 8880 8697
rect 8480 8640 8880 8663
rect 8960 8697 9360 8720
rect 8960 8663 8983 8697
rect 9017 8663 9143 8697
rect 9177 8663 9303 8697
rect 9337 8663 9360 8697
rect 8960 8640 9360 8663
rect 9440 8697 11440 8720
rect 9440 8663 9463 8697
rect 9497 8663 9623 8697
rect 9657 8663 9783 8697
rect 9817 8663 9943 8697
rect 9977 8663 10103 8697
rect 10137 8663 10263 8697
rect 10297 8663 10423 8697
rect 10457 8663 10583 8697
rect 10617 8663 10743 8697
rect 10777 8663 10903 8697
rect 10937 8663 11063 8697
rect 11097 8663 11223 8697
rect 11257 8663 11383 8697
rect 11417 8663 11440 8697
rect 9440 8640 11440 8663
rect 11520 8697 11920 8720
rect 11520 8663 11543 8697
rect 11577 8663 11703 8697
rect 11737 8663 11863 8697
rect 11897 8663 11920 8697
rect 11520 8640 11920 8663
rect 12000 8697 12400 8720
rect 12000 8663 12023 8697
rect 12057 8663 12183 8697
rect 12217 8663 12343 8697
rect 12377 8663 12400 8697
rect 12000 8640 12400 8663
rect 8480 8537 8880 8560
rect 8480 8503 8503 8537
rect 8537 8503 8663 8537
rect 8697 8503 8823 8537
rect 8857 8503 8880 8537
rect 8480 8480 8880 8503
rect 8960 8537 9360 8560
rect 8960 8503 8983 8537
rect 9017 8503 9143 8537
rect 9177 8503 9303 8537
rect 9337 8503 9360 8537
rect 8960 8480 9360 8503
rect 9440 8537 11440 8560
rect 9440 8503 9463 8537
rect 9497 8503 9623 8537
rect 9657 8503 9783 8537
rect 9817 8503 9943 8537
rect 9977 8503 10103 8537
rect 10137 8503 10263 8537
rect 10297 8503 10423 8537
rect 10457 8503 10583 8537
rect 10617 8503 10743 8537
rect 10777 8503 10903 8537
rect 10937 8503 11063 8537
rect 11097 8503 11223 8537
rect 11257 8503 11383 8537
rect 11417 8503 11440 8537
rect 9440 8480 11440 8503
rect 11520 8537 11920 8560
rect 11520 8503 11543 8537
rect 11577 8503 11703 8537
rect 11737 8503 11863 8537
rect 11897 8503 11920 8537
rect 11520 8480 11920 8503
rect 12000 8537 12400 8560
rect 12000 8503 12023 8537
rect 12057 8503 12183 8537
rect 12217 8503 12343 8537
rect 12377 8503 12400 8537
rect 12000 8480 12400 8503
rect 8480 8377 8880 8400
rect 8480 8343 8503 8377
rect 8537 8343 8663 8377
rect 8697 8343 8823 8377
rect 8857 8343 8880 8377
rect 8480 8320 8880 8343
rect 8960 8377 9360 8400
rect 8960 8343 8983 8377
rect 9017 8343 9143 8377
rect 9177 8343 9303 8377
rect 9337 8343 9360 8377
rect 8960 8320 9360 8343
rect 9440 8377 11440 8400
rect 9440 8343 9463 8377
rect 9497 8343 9623 8377
rect 9657 8343 9783 8377
rect 9817 8343 9943 8377
rect 9977 8343 10103 8377
rect 10137 8343 10263 8377
rect 10297 8343 10423 8377
rect 10457 8343 10583 8377
rect 10617 8343 10743 8377
rect 10777 8343 10903 8377
rect 10937 8343 11063 8377
rect 11097 8343 11223 8377
rect 11257 8343 11383 8377
rect 11417 8343 11440 8377
rect 9440 8320 11440 8343
rect 11520 8377 11920 8400
rect 11520 8343 11543 8377
rect 11577 8343 11703 8377
rect 11737 8343 11863 8377
rect 11897 8343 11920 8377
rect 11520 8320 11920 8343
rect 12000 8377 12400 8400
rect 12000 8343 12023 8377
rect 12057 8343 12183 8377
rect 12217 8343 12343 8377
rect 12377 8343 12400 8377
rect 12000 8320 12400 8343
rect 8480 8217 8880 8240
rect 8480 8183 8503 8217
rect 8537 8183 8663 8217
rect 8697 8183 8823 8217
rect 8857 8183 8880 8217
rect 8480 8160 8880 8183
rect 8960 8217 9360 8240
rect 8960 8183 8983 8217
rect 9017 8183 9143 8217
rect 9177 8183 9303 8217
rect 9337 8183 9360 8217
rect 8960 8160 9360 8183
rect 9440 8217 11440 8240
rect 9440 8183 9463 8217
rect 9497 8183 9623 8217
rect 9657 8183 9783 8217
rect 9817 8183 9943 8217
rect 9977 8183 10103 8217
rect 10137 8183 10263 8217
rect 10297 8183 10423 8217
rect 10457 8183 10583 8217
rect 10617 8183 10743 8217
rect 10777 8183 10903 8217
rect 10937 8183 11063 8217
rect 11097 8183 11223 8217
rect 11257 8183 11383 8217
rect 11417 8183 11440 8217
rect 9440 8160 11440 8183
rect 11520 8217 11920 8240
rect 11520 8183 11543 8217
rect 11577 8183 11703 8217
rect 11737 8183 11863 8217
rect 11897 8183 11920 8217
rect 11520 8160 11920 8183
rect 12000 8217 12400 8240
rect 12000 8183 12023 8217
rect 12057 8183 12183 8217
rect 12217 8183 12343 8217
rect 12377 8183 12400 8217
rect 12000 8160 12400 8183
rect 8480 8057 8880 8080
rect 8480 8023 8503 8057
rect 8537 8023 8663 8057
rect 8697 8023 8823 8057
rect 8857 8023 8880 8057
rect 8480 8000 8880 8023
rect 8960 8057 9360 8080
rect 8960 8023 8983 8057
rect 9017 8023 9143 8057
rect 9177 8023 9303 8057
rect 9337 8023 9360 8057
rect 8960 8000 9360 8023
rect 9440 8057 11440 8080
rect 9440 8023 9463 8057
rect 9497 8023 9623 8057
rect 9657 8023 9783 8057
rect 9817 8023 9943 8057
rect 9977 8023 10103 8057
rect 10137 8023 10263 8057
rect 10297 8023 10423 8057
rect 10457 8023 10583 8057
rect 10617 8023 10743 8057
rect 10777 8023 10903 8057
rect 10937 8023 11063 8057
rect 11097 8023 11223 8057
rect 11257 8023 11383 8057
rect 11417 8023 11440 8057
rect 9440 8000 11440 8023
rect 11520 8057 11920 8080
rect 11520 8023 11543 8057
rect 11577 8023 11703 8057
rect 11737 8023 11863 8057
rect 11897 8023 11920 8057
rect 11520 8000 11920 8023
rect 12000 8057 12400 8080
rect 12000 8023 12023 8057
rect 12057 8023 12183 8057
rect 12217 8023 12343 8057
rect 12377 8023 12400 8057
rect 12000 8000 12400 8023
rect 8480 7897 8880 7920
rect 8480 7863 8503 7897
rect 8537 7863 8663 7897
rect 8697 7863 8823 7897
rect 8857 7863 8880 7897
rect 8480 7840 8880 7863
rect 8960 7897 9360 7920
rect 8960 7863 8983 7897
rect 9017 7863 9143 7897
rect 9177 7863 9303 7897
rect 9337 7863 9360 7897
rect 8960 7840 9360 7863
rect 9440 7897 11440 7920
rect 9440 7863 9463 7897
rect 9497 7863 9623 7897
rect 9657 7863 9783 7897
rect 9817 7863 9943 7897
rect 9977 7863 10103 7897
rect 10137 7863 10263 7897
rect 10297 7863 10423 7897
rect 10457 7863 10583 7897
rect 10617 7863 10743 7897
rect 10777 7863 10903 7897
rect 10937 7863 11063 7897
rect 11097 7863 11223 7897
rect 11257 7863 11383 7897
rect 11417 7863 11440 7897
rect 9440 7840 11440 7863
rect 11520 7897 11920 7920
rect 11520 7863 11543 7897
rect 11577 7863 11703 7897
rect 11737 7863 11863 7897
rect 11897 7863 11920 7897
rect 11520 7840 11920 7863
rect 12000 7897 12400 7920
rect 12000 7863 12023 7897
rect 12057 7863 12183 7897
rect 12217 7863 12343 7897
rect 12377 7863 12400 7897
rect 12000 7840 12400 7863
rect 8480 7737 8880 7760
rect 8480 7703 8503 7737
rect 8537 7703 8663 7737
rect 8697 7703 8823 7737
rect 8857 7703 8880 7737
rect 8480 7680 8880 7703
rect 8960 7737 9360 7760
rect 8960 7703 8983 7737
rect 9017 7703 9143 7737
rect 9177 7703 9303 7737
rect 9337 7703 9360 7737
rect 8960 7680 9360 7703
rect 9440 7737 11440 7760
rect 9440 7703 9463 7737
rect 9497 7703 9623 7737
rect 9657 7703 9783 7737
rect 9817 7703 9943 7737
rect 9977 7703 10103 7737
rect 10137 7703 10263 7737
rect 10297 7703 10423 7737
rect 10457 7703 10583 7737
rect 10617 7703 10743 7737
rect 10777 7703 10903 7737
rect 10937 7703 11063 7737
rect 11097 7703 11223 7737
rect 11257 7703 11383 7737
rect 11417 7703 11440 7737
rect 9440 7680 11440 7703
rect 11520 7737 11920 7760
rect 11520 7703 11543 7737
rect 11577 7703 11703 7737
rect 11737 7703 11863 7737
rect 11897 7703 11920 7737
rect 11520 7680 11920 7703
rect 12000 7737 12400 7760
rect 12000 7703 12023 7737
rect 12057 7703 12183 7737
rect 12217 7703 12343 7737
rect 12377 7703 12400 7737
rect 12000 7680 12400 7703
rect 8480 7577 8880 7600
rect 8480 7543 8503 7577
rect 8537 7543 8663 7577
rect 8697 7543 8823 7577
rect 8857 7543 8880 7577
rect 8480 7520 8880 7543
rect 8960 7577 9360 7600
rect 8960 7543 8983 7577
rect 9017 7543 9143 7577
rect 9177 7543 9303 7577
rect 9337 7543 9360 7577
rect 8960 7520 9360 7543
rect 9440 7577 11440 7600
rect 9440 7543 9463 7577
rect 9497 7543 9623 7577
rect 9657 7543 9783 7577
rect 9817 7543 9943 7577
rect 9977 7543 10103 7577
rect 10137 7543 10263 7577
rect 10297 7543 10423 7577
rect 10457 7543 10583 7577
rect 10617 7543 10743 7577
rect 10777 7543 10903 7577
rect 10937 7543 11063 7577
rect 11097 7543 11223 7577
rect 11257 7543 11383 7577
rect 11417 7543 11440 7577
rect 9440 7520 11440 7543
rect 11520 7577 11920 7600
rect 11520 7543 11543 7577
rect 11577 7543 11703 7577
rect 11737 7543 11863 7577
rect 11897 7543 11920 7577
rect 11520 7520 11920 7543
rect 12000 7577 12400 7600
rect 12000 7543 12023 7577
rect 12057 7543 12183 7577
rect 12217 7543 12343 7577
rect 12377 7543 12400 7577
rect 12000 7520 12400 7543
rect 8480 7417 8880 7440
rect 8480 7383 8503 7417
rect 8537 7383 8663 7417
rect 8697 7383 8823 7417
rect 8857 7383 8880 7417
rect 8480 7360 8880 7383
rect 8960 7417 9360 7440
rect 8960 7383 8983 7417
rect 9017 7383 9143 7417
rect 9177 7383 9303 7417
rect 9337 7383 9360 7417
rect 8960 7360 9360 7383
rect 9440 7417 11440 7440
rect 9440 7383 9463 7417
rect 9497 7383 9623 7417
rect 9657 7383 9783 7417
rect 9817 7383 9943 7417
rect 9977 7383 10103 7417
rect 10137 7383 10263 7417
rect 10297 7383 10423 7417
rect 10457 7383 10583 7417
rect 10617 7383 10743 7417
rect 10777 7383 10903 7417
rect 10937 7383 11063 7417
rect 11097 7383 11223 7417
rect 11257 7383 11383 7417
rect 11417 7383 11440 7417
rect 9440 7360 11440 7383
rect 11520 7417 11920 7440
rect 11520 7383 11543 7417
rect 11577 7383 11703 7417
rect 11737 7383 11863 7417
rect 11897 7383 11920 7417
rect 11520 7360 11920 7383
rect 12000 7417 12400 7440
rect 12000 7383 12023 7417
rect 12057 7383 12183 7417
rect 12217 7383 12343 7417
rect 12377 7383 12400 7417
rect 12000 7360 12400 7383
rect 8480 7257 8880 7280
rect 8480 7223 8503 7257
rect 8537 7223 8663 7257
rect 8697 7223 8823 7257
rect 8857 7223 8880 7257
rect 8480 7200 8880 7223
rect 8960 7257 9360 7280
rect 8960 7223 8983 7257
rect 9017 7223 9143 7257
rect 9177 7223 9303 7257
rect 9337 7223 9360 7257
rect 8960 7200 9360 7223
rect 9440 7257 11440 7280
rect 9440 7223 9463 7257
rect 9497 7223 9623 7257
rect 9657 7223 9783 7257
rect 9817 7223 9943 7257
rect 9977 7223 10103 7257
rect 10137 7223 10263 7257
rect 10297 7223 10423 7257
rect 10457 7223 10583 7257
rect 10617 7223 10743 7257
rect 10777 7223 10903 7257
rect 10937 7223 11063 7257
rect 11097 7223 11223 7257
rect 11257 7223 11383 7257
rect 11417 7223 11440 7257
rect 9440 7200 11440 7223
rect 11520 7257 11920 7280
rect 11520 7223 11543 7257
rect 11577 7223 11703 7257
rect 11737 7223 11863 7257
rect 11897 7223 11920 7257
rect 11520 7200 11920 7223
rect 12000 7257 12400 7280
rect 12000 7223 12023 7257
rect 12057 7223 12183 7257
rect 12217 7223 12343 7257
rect 12377 7223 12400 7257
rect 12000 7200 12400 7223
rect 8480 7097 8880 7120
rect 8480 7063 8503 7097
rect 8537 7063 8663 7097
rect 8697 7063 8823 7097
rect 8857 7063 8880 7097
rect 8480 7040 8880 7063
rect 8960 7097 9360 7120
rect 8960 7063 8983 7097
rect 9017 7063 9143 7097
rect 9177 7063 9303 7097
rect 9337 7063 9360 7097
rect 8960 7040 9360 7063
rect 9440 7097 11440 7120
rect 9440 7063 9463 7097
rect 9497 7063 9623 7097
rect 9657 7063 9783 7097
rect 9817 7063 9943 7097
rect 9977 7063 10103 7097
rect 10137 7063 10263 7097
rect 10297 7063 10423 7097
rect 10457 7063 10583 7097
rect 10617 7063 10743 7097
rect 10777 7063 10903 7097
rect 10937 7063 11063 7097
rect 11097 7063 11223 7097
rect 11257 7063 11383 7097
rect 11417 7063 11440 7097
rect 9440 7040 11440 7063
rect 11520 7097 11920 7120
rect 11520 7063 11543 7097
rect 11577 7063 11703 7097
rect 11737 7063 11863 7097
rect 11897 7063 11920 7097
rect 11520 7040 11920 7063
rect 12000 7097 12400 7120
rect 12000 7063 12023 7097
rect 12057 7063 12183 7097
rect 12217 7063 12343 7097
rect 12377 7063 12400 7097
rect 12000 7040 12400 7063
rect 8480 6937 8880 6960
rect 8480 6903 8503 6937
rect 8537 6903 8663 6937
rect 8697 6903 8823 6937
rect 8857 6903 8880 6937
rect 8480 6880 8880 6903
rect 8960 6937 9360 6960
rect 8960 6903 8983 6937
rect 9017 6903 9143 6937
rect 9177 6903 9303 6937
rect 9337 6903 9360 6937
rect 8960 6880 9360 6903
rect 9440 6937 11440 6960
rect 9440 6903 9463 6937
rect 9497 6903 9623 6937
rect 9657 6903 9783 6937
rect 9817 6903 9943 6937
rect 9977 6903 10103 6937
rect 10137 6903 10263 6937
rect 10297 6903 10423 6937
rect 10457 6903 10583 6937
rect 10617 6903 10743 6937
rect 10777 6903 10903 6937
rect 10937 6903 11063 6937
rect 11097 6903 11223 6937
rect 11257 6903 11383 6937
rect 11417 6903 11440 6937
rect 9440 6880 11440 6903
rect 11520 6937 11920 6960
rect 11520 6903 11543 6937
rect 11577 6903 11703 6937
rect 11737 6903 11863 6937
rect 11897 6903 11920 6937
rect 11520 6880 11920 6903
rect 12000 6937 12400 6960
rect 12000 6903 12023 6937
rect 12057 6903 12183 6937
rect 12217 6903 12343 6937
rect 12377 6903 12400 6937
rect 12000 6880 12400 6903
rect 8480 6777 8880 6800
rect 8480 6743 8503 6777
rect 8537 6743 8663 6777
rect 8697 6743 8823 6777
rect 8857 6743 8880 6777
rect 8480 6720 8880 6743
rect 8960 6777 9360 6800
rect 8960 6743 8983 6777
rect 9017 6743 9143 6777
rect 9177 6743 9303 6777
rect 9337 6743 9360 6777
rect 8960 6720 9360 6743
rect 9440 6777 11440 6800
rect 9440 6743 9463 6777
rect 9497 6743 9623 6777
rect 9657 6743 9783 6777
rect 9817 6743 9943 6777
rect 9977 6743 10103 6777
rect 10137 6743 10263 6777
rect 10297 6743 10423 6777
rect 10457 6743 10583 6777
rect 10617 6743 10743 6777
rect 10777 6743 10903 6777
rect 10937 6743 11063 6777
rect 11097 6743 11223 6777
rect 11257 6743 11383 6777
rect 11417 6743 11440 6777
rect 9440 6720 11440 6743
rect 11520 6777 11920 6800
rect 11520 6743 11543 6777
rect 11577 6743 11703 6777
rect 11737 6743 11863 6777
rect 11897 6743 11920 6777
rect 11520 6720 11920 6743
rect 12000 6777 12400 6800
rect 12000 6743 12023 6777
rect 12057 6743 12183 6777
rect 12217 6743 12343 6777
rect 12377 6743 12400 6777
rect 12000 6720 12400 6743
rect 8480 6617 8880 6640
rect 8480 6583 8503 6617
rect 8537 6583 8663 6617
rect 8697 6583 8823 6617
rect 8857 6583 8880 6617
rect 8480 6560 8880 6583
rect 8960 6617 9360 6640
rect 8960 6583 8983 6617
rect 9017 6583 9143 6617
rect 9177 6583 9303 6617
rect 9337 6583 9360 6617
rect 8960 6560 9360 6583
rect 9440 6617 11440 6640
rect 9440 6583 9463 6617
rect 9497 6583 9623 6617
rect 9657 6583 9783 6617
rect 9817 6583 9943 6617
rect 9977 6583 10103 6617
rect 10137 6583 10263 6617
rect 10297 6583 10423 6617
rect 10457 6583 10583 6617
rect 10617 6583 10743 6617
rect 10777 6583 10903 6617
rect 10937 6583 11063 6617
rect 11097 6583 11223 6617
rect 11257 6583 11383 6617
rect 11417 6583 11440 6617
rect 9440 6560 11440 6583
rect 11520 6617 11920 6640
rect 11520 6583 11543 6617
rect 11577 6583 11703 6617
rect 11737 6583 11863 6617
rect 11897 6583 11920 6617
rect 11520 6560 11920 6583
rect 12000 6617 12400 6640
rect 12000 6583 12023 6617
rect 12057 6583 12183 6617
rect 12217 6583 12343 6617
rect 12377 6583 12400 6617
rect 12000 6560 12400 6583
rect 8480 6457 8880 6480
rect 8480 6423 8503 6457
rect 8537 6423 8663 6457
rect 8697 6423 8823 6457
rect 8857 6423 8880 6457
rect 8480 6400 8880 6423
rect 8960 6457 9360 6480
rect 8960 6423 8983 6457
rect 9017 6423 9143 6457
rect 9177 6423 9303 6457
rect 9337 6423 9360 6457
rect 8960 6400 9360 6423
rect 9440 6457 11440 6480
rect 9440 6423 9463 6457
rect 9497 6423 9623 6457
rect 9657 6423 9783 6457
rect 9817 6423 9943 6457
rect 9977 6423 10103 6457
rect 10137 6423 10263 6457
rect 10297 6423 10423 6457
rect 10457 6423 10583 6457
rect 10617 6423 10743 6457
rect 10777 6423 10903 6457
rect 10937 6423 11063 6457
rect 11097 6423 11223 6457
rect 11257 6423 11383 6457
rect 11417 6423 11440 6457
rect 9440 6400 11440 6423
rect 11520 6457 11920 6480
rect 11520 6423 11543 6457
rect 11577 6423 11703 6457
rect 11737 6423 11863 6457
rect 11897 6423 11920 6457
rect 11520 6400 11920 6423
rect 12000 6457 12400 6480
rect 12000 6423 12023 6457
rect 12057 6423 12183 6457
rect 12217 6423 12343 6457
rect 12377 6423 12400 6457
rect 12000 6400 12400 6423
rect 8480 6297 8880 6320
rect 8480 6263 8503 6297
rect 8537 6263 8663 6297
rect 8697 6263 8823 6297
rect 8857 6263 8880 6297
rect 8480 6240 8880 6263
rect 8960 6297 9360 6320
rect 8960 6263 8983 6297
rect 9017 6263 9143 6297
rect 9177 6263 9303 6297
rect 9337 6263 9360 6297
rect 8960 6240 9360 6263
rect 9440 6297 11440 6320
rect 9440 6263 9463 6297
rect 9497 6263 9623 6297
rect 9657 6263 9783 6297
rect 9817 6263 9943 6297
rect 9977 6263 10103 6297
rect 10137 6263 10263 6297
rect 10297 6263 10423 6297
rect 10457 6263 10583 6297
rect 10617 6263 10743 6297
rect 10777 6263 10903 6297
rect 10937 6263 11063 6297
rect 11097 6263 11223 6297
rect 11257 6263 11383 6297
rect 11417 6263 11440 6297
rect 9440 6240 11440 6263
rect 11520 6297 11920 6320
rect 11520 6263 11543 6297
rect 11577 6263 11703 6297
rect 11737 6263 11863 6297
rect 11897 6263 11920 6297
rect 11520 6240 11920 6263
rect 12000 6297 12400 6320
rect 12000 6263 12023 6297
rect 12057 6263 12183 6297
rect 12217 6263 12343 6297
rect 12377 6263 12400 6297
rect 12000 6240 12400 6263
rect 8480 6137 8880 6160
rect 8480 6103 8503 6137
rect 8537 6103 8663 6137
rect 8697 6103 8823 6137
rect 8857 6103 8880 6137
rect 8480 6080 8880 6103
rect 8960 6137 9360 6160
rect 8960 6103 8983 6137
rect 9017 6103 9143 6137
rect 9177 6103 9303 6137
rect 9337 6103 9360 6137
rect 8960 6080 9360 6103
rect 9440 6137 11440 6160
rect 9440 6103 9463 6137
rect 9497 6103 9623 6137
rect 9657 6103 9783 6137
rect 9817 6103 9943 6137
rect 9977 6103 10103 6137
rect 10137 6103 10263 6137
rect 10297 6103 10423 6137
rect 10457 6103 10583 6137
rect 10617 6103 10743 6137
rect 10777 6103 10903 6137
rect 10937 6103 11063 6137
rect 11097 6103 11223 6137
rect 11257 6103 11383 6137
rect 11417 6103 11440 6137
rect 9440 6080 11440 6103
rect 11520 6137 11920 6160
rect 11520 6103 11543 6137
rect 11577 6103 11703 6137
rect 11737 6103 11863 6137
rect 11897 6103 11920 6137
rect 11520 6080 11920 6103
rect 12000 6137 12400 6160
rect 12000 6103 12023 6137
rect 12057 6103 12183 6137
rect 12217 6103 12343 6137
rect 12377 6103 12400 6137
rect 12000 6080 12400 6103
rect 8480 5977 8880 6000
rect 8480 5943 8503 5977
rect 8537 5943 8663 5977
rect 8697 5943 8823 5977
rect 8857 5943 8880 5977
rect 8480 5920 8880 5943
rect 8960 5977 9360 6000
rect 8960 5943 8983 5977
rect 9017 5943 9143 5977
rect 9177 5943 9303 5977
rect 9337 5943 9360 5977
rect 8960 5920 9360 5943
rect 9440 5977 11440 6000
rect 9440 5943 9463 5977
rect 9497 5943 9623 5977
rect 9657 5943 9783 5977
rect 9817 5943 9943 5977
rect 9977 5943 10103 5977
rect 10137 5943 10263 5977
rect 10297 5943 10423 5977
rect 10457 5943 10583 5977
rect 10617 5943 10743 5977
rect 10777 5943 10903 5977
rect 10937 5943 11063 5977
rect 11097 5943 11223 5977
rect 11257 5943 11383 5977
rect 11417 5943 11440 5977
rect 9440 5920 11440 5943
rect 11520 5977 11920 6000
rect 11520 5943 11543 5977
rect 11577 5943 11703 5977
rect 11737 5943 11863 5977
rect 11897 5943 11920 5977
rect 11520 5920 11920 5943
rect 12000 5977 12400 6000
rect 12000 5943 12023 5977
rect 12057 5943 12183 5977
rect 12217 5943 12343 5977
rect 12377 5943 12400 5977
rect 12000 5920 12400 5943
rect 8480 5817 8880 5840
rect 8480 5783 8503 5817
rect 8537 5783 8663 5817
rect 8697 5783 8823 5817
rect 8857 5783 8880 5817
rect 8480 5760 8880 5783
rect 8960 5817 9360 5840
rect 8960 5783 8983 5817
rect 9017 5783 9143 5817
rect 9177 5783 9303 5817
rect 9337 5783 9360 5817
rect 8960 5760 9360 5783
rect 9440 5817 11440 5840
rect 9440 5783 9463 5817
rect 9497 5783 9623 5817
rect 9657 5783 9783 5817
rect 9817 5783 9943 5817
rect 9977 5783 10103 5817
rect 10137 5783 10263 5817
rect 10297 5783 10423 5817
rect 10457 5783 10583 5817
rect 10617 5783 10743 5817
rect 10777 5783 10903 5817
rect 10937 5783 11063 5817
rect 11097 5783 11223 5817
rect 11257 5783 11383 5817
rect 11417 5783 11440 5817
rect 9440 5760 11440 5783
rect 11520 5817 11920 5840
rect 11520 5783 11543 5817
rect 11577 5783 11703 5817
rect 11737 5783 11863 5817
rect 11897 5783 11920 5817
rect 11520 5760 11920 5783
rect 12000 5817 12400 5840
rect 12000 5783 12023 5817
rect 12057 5783 12183 5817
rect 12217 5783 12343 5817
rect 12377 5783 12400 5817
rect 12000 5760 12400 5783
rect 8480 5657 8880 5680
rect 8480 5623 8503 5657
rect 8537 5623 8663 5657
rect 8697 5623 8823 5657
rect 8857 5623 8880 5657
rect 8480 5600 8880 5623
rect 8960 5657 9360 5680
rect 8960 5623 8983 5657
rect 9017 5623 9143 5657
rect 9177 5623 9303 5657
rect 9337 5623 9360 5657
rect 8960 5600 9360 5623
rect 9440 5657 11440 5680
rect 9440 5623 9463 5657
rect 9497 5623 9623 5657
rect 9657 5623 9783 5657
rect 9817 5623 9943 5657
rect 9977 5623 10103 5657
rect 10137 5623 10263 5657
rect 10297 5623 10423 5657
rect 10457 5623 10583 5657
rect 10617 5623 10743 5657
rect 10777 5623 10903 5657
rect 10937 5623 11063 5657
rect 11097 5623 11223 5657
rect 11257 5623 11383 5657
rect 11417 5623 11440 5657
rect 9440 5600 11440 5623
rect 11520 5657 11920 5680
rect 11520 5623 11543 5657
rect 11577 5623 11703 5657
rect 11737 5623 11863 5657
rect 11897 5623 11920 5657
rect 11520 5600 11920 5623
rect 12000 5657 12400 5680
rect 12000 5623 12023 5657
rect 12057 5623 12183 5657
rect 12217 5623 12343 5657
rect 12377 5623 12400 5657
rect 12000 5600 12400 5623
rect 8480 5497 8880 5520
rect 8480 5463 8503 5497
rect 8537 5463 8663 5497
rect 8697 5463 8823 5497
rect 8857 5463 8880 5497
rect 8480 5440 8880 5463
rect 8960 5497 9360 5520
rect 8960 5463 8983 5497
rect 9017 5463 9143 5497
rect 9177 5463 9303 5497
rect 9337 5463 9360 5497
rect 8960 5440 9360 5463
rect 9440 5497 11440 5520
rect 9440 5463 9463 5497
rect 9497 5463 9623 5497
rect 9657 5463 9783 5497
rect 9817 5463 9943 5497
rect 9977 5463 10103 5497
rect 10137 5463 10263 5497
rect 10297 5463 10423 5497
rect 10457 5463 10583 5497
rect 10617 5463 10743 5497
rect 10777 5463 10903 5497
rect 10937 5463 11063 5497
rect 11097 5463 11223 5497
rect 11257 5463 11383 5497
rect 11417 5463 11440 5497
rect 9440 5440 11440 5463
rect 11520 5497 11920 5520
rect 11520 5463 11543 5497
rect 11577 5463 11703 5497
rect 11737 5463 11863 5497
rect 11897 5463 11920 5497
rect 11520 5440 11920 5463
rect 12000 5497 12400 5520
rect 12000 5463 12023 5497
rect 12057 5463 12183 5497
rect 12217 5463 12343 5497
rect 12377 5463 12400 5497
rect 12000 5440 12400 5463
rect 8480 5337 8880 5360
rect 8480 5303 8503 5337
rect 8537 5303 8663 5337
rect 8697 5303 8823 5337
rect 8857 5303 8880 5337
rect 8480 5280 8880 5303
rect 8960 5337 9360 5360
rect 8960 5303 8983 5337
rect 9017 5303 9143 5337
rect 9177 5303 9303 5337
rect 9337 5303 9360 5337
rect 8960 5280 9360 5303
rect 9440 5337 11440 5360
rect 9440 5303 9463 5337
rect 9497 5303 9623 5337
rect 9657 5303 9783 5337
rect 9817 5303 9943 5337
rect 9977 5303 10103 5337
rect 10137 5303 10263 5337
rect 10297 5303 10423 5337
rect 10457 5303 10583 5337
rect 10617 5303 10743 5337
rect 10777 5303 10903 5337
rect 10937 5303 11063 5337
rect 11097 5303 11223 5337
rect 11257 5303 11383 5337
rect 11417 5303 11440 5337
rect 9440 5280 11440 5303
rect 11520 5337 11920 5360
rect 11520 5303 11543 5337
rect 11577 5303 11703 5337
rect 11737 5303 11863 5337
rect 11897 5303 11920 5337
rect 11520 5280 11920 5303
rect 12000 5337 12400 5360
rect 12000 5303 12023 5337
rect 12057 5303 12183 5337
rect 12217 5303 12343 5337
rect 12377 5303 12400 5337
rect 12000 5280 12400 5303
rect 8480 5177 8880 5200
rect 8480 5143 8503 5177
rect 8537 5143 8663 5177
rect 8697 5143 8823 5177
rect 8857 5143 8880 5177
rect 8480 5120 8880 5143
rect 8960 5177 9360 5200
rect 8960 5143 8983 5177
rect 9017 5143 9143 5177
rect 9177 5143 9303 5177
rect 9337 5143 9360 5177
rect 8960 5120 9360 5143
rect 9440 5177 11440 5200
rect 9440 5143 9463 5177
rect 9497 5143 9623 5177
rect 9657 5143 9783 5177
rect 9817 5143 9943 5177
rect 9977 5143 10103 5177
rect 10137 5143 10263 5177
rect 10297 5143 10423 5177
rect 10457 5143 10583 5177
rect 10617 5143 10743 5177
rect 10777 5143 10903 5177
rect 10937 5143 11063 5177
rect 11097 5143 11223 5177
rect 11257 5143 11383 5177
rect 11417 5143 11440 5177
rect 9440 5120 11440 5143
rect 11520 5177 11920 5200
rect 11520 5143 11543 5177
rect 11577 5143 11703 5177
rect 11737 5143 11863 5177
rect 11897 5143 11920 5177
rect 11520 5120 11920 5143
rect 12000 5177 12400 5200
rect 12000 5143 12023 5177
rect 12057 5143 12183 5177
rect 12217 5143 12343 5177
rect 12377 5143 12400 5177
rect 12000 5120 12400 5143
rect 8480 5017 8880 5040
rect 8480 4983 8503 5017
rect 8537 4983 8663 5017
rect 8697 4983 8823 5017
rect 8857 4983 8880 5017
rect 8480 4960 8880 4983
rect 8960 5017 9360 5040
rect 8960 4983 8983 5017
rect 9017 4983 9143 5017
rect 9177 4983 9303 5017
rect 9337 4983 9360 5017
rect 8960 4960 9360 4983
rect 9440 5017 11440 5040
rect 9440 4983 9463 5017
rect 9497 4983 9623 5017
rect 9657 4983 9783 5017
rect 9817 4983 9943 5017
rect 9977 4983 10103 5017
rect 10137 4983 10263 5017
rect 10297 4983 10423 5017
rect 10457 4983 10583 5017
rect 10617 4983 10743 5017
rect 10777 4983 10903 5017
rect 10937 4983 11063 5017
rect 11097 4983 11223 5017
rect 11257 4983 11383 5017
rect 11417 4983 11440 5017
rect 9440 4960 11440 4983
rect 11520 5017 11920 5040
rect 11520 4983 11543 5017
rect 11577 4983 11703 5017
rect 11737 4983 11863 5017
rect 11897 4983 11920 5017
rect 11520 4960 11920 4983
rect 12000 5017 12400 5040
rect 12000 4983 12023 5017
rect 12057 4983 12183 5017
rect 12217 4983 12343 5017
rect 12377 4983 12400 5017
rect 12000 4960 12400 4983
rect 8480 4857 8880 4880
rect 8480 4823 8503 4857
rect 8537 4823 8663 4857
rect 8697 4823 8823 4857
rect 8857 4823 8880 4857
rect 8480 4800 8880 4823
rect 8960 4857 9360 4880
rect 8960 4823 8983 4857
rect 9017 4823 9143 4857
rect 9177 4823 9303 4857
rect 9337 4823 9360 4857
rect 8960 4800 9360 4823
rect 9440 4857 11440 4880
rect 9440 4823 9463 4857
rect 9497 4823 9623 4857
rect 9657 4823 9783 4857
rect 9817 4823 9943 4857
rect 9977 4823 10103 4857
rect 10137 4823 10263 4857
rect 10297 4823 10423 4857
rect 10457 4823 10583 4857
rect 10617 4823 10743 4857
rect 10777 4823 10903 4857
rect 10937 4823 11063 4857
rect 11097 4823 11223 4857
rect 11257 4823 11383 4857
rect 11417 4823 11440 4857
rect 9440 4800 11440 4823
rect 11520 4857 11920 4880
rect 11520 4823 11543 4857
rect 11577 4823 11703 4857
rect 11737 4823 11863 4857
rect 11897 4823 11920 4857
rect 11520 4800 11920 4823
rect 12000 4857 12400 4880
rect 12000 4823 12023 4857
rect 12057 4823 12183 4857
rect 12217 4823 12343 4857
rect 12377 4823 12400 4857
rect 12000 4800 12400 4823
rect 8480 4697 8880 4720
rect 8480 4663 8503 4697
rect 8537 4663 8663 4697
rect 8697 4663 8823 4697
rect 8857 4663 8880 4697
rect 8480 4640 8880 4663
rect 8960 4697 9360 4720
rect 8960 4663 8983 4697
rect 9017 4663 9143 4697
rect 9177 4663 9303 4697
rect 9337 4663 9360 4697
rect 8960 4640 9360 4663
rect 9440 4697 11440 4720
rect 9440 4663 9463 4697
rect 9497 4663 9623 4697
rect 9657 4663 9783 4697
rect 9817 4663 9943 4697
rect 9977 4663 10103 4697
rect 10137 4663 10263 4697
rect 10297 4663 10423 4697
rect 10457 4663 10583 4697
rect 10617 4663 10743 4697
rect 10777 4663 10903 4697
rect 10937 4663 11063 4697
rect 11097 4663 11223 4697
rect 11257 4663 11383 4697
rect 11417 4663 11440 4697
rect 9440 4640 11440 4663
rect 11520 4697 11920 4720
rect 11520 4663 11543 4697
rect 11577 4663 11703 4697
rect 11737 4663 11863 4697
rect 11897 4663 11920 4697
rect 11520 4640 11920 4663
rect 12000 4697 12400 4720
rect 12000 4663 12023 4697
rect 12057 4663 12183 4697
rect 12217 4663 12343 4697
rect 12377 4663 12400 4697
rect 12000 4640 12400 4663
rect 8480 4537 8880 4560
rect 8480 4503 8503 4537
rect 8537 4503 8663 4537
rect 8697 4503 8823 4537
rect 8857 4503 8880 4537
rect 8480 4480 8880 4503
rect 8960 4537 9360 4560
rect 8960 4503 8983 4537
rect 9017 4503 9143 4537
rect 9177 4503 9303 4537
rect 9337 4503 9360 4537
rect 8960 4480 9360 4503
rect 9440 4537 11440 4560
rect 9440 4503 9463 4537
rect 9497 4503 9623 4537
rect 9657 4503 9783 4537
rect 9817 4503 9943 4537
rect 9977 4503 10103 4537
rect 10137 4503 10263 4537
rect 10297 4503 10423 4537
rect 10457 4503 10583 4537
rect 10617 4503 10743 4537
rect 10777 4503 10903 4537
rect 10937 4503 11063 4537
rect 11097 4503 11223 4537
rect 11257 4503 11383 4537
rect 11417 4503 11440 4537
rect 9440 4480 11440 4503
rect 11520 4537 11920 4560
rect 11520 4503 11543 4537
rect 11577 4503 11703 4537
rect 11737 4503 11863 4537
rect 11897 4503 11920 4537
rect 11520 4480 11920 4503
rect 12000 4537 12400 4560
rect 12000 4503 12023 4537
rect 12057 4503 12183 4537
rect 12217 4503 12343 4537
rect 12377 4503 12400 4537
rect 12000 4480 12400 4503
rect 8480 4377 8880 4400
rect 8480 4343 8503 4377
rect 8537 4343 8663 4377
rect 8697 4343 8823 4377
rect 8857 4343 8880 4377
rect 8480 4320 8880 4343
rect 8960 4377 9360 4400
rect 8960 4343 8983 4377
rect 9017 4343 9143 4377
rect 9177 4343 9303 4377
rect 9337 4343 9360 4377
rect 8960 4320 9360 4343
rect 9440 4377 11440 4400
rect 9440 4343 9463 4377
rect 9497 4343 9623 4377
rect 9657 4343 9783 4377
rect 9817 4343 9943 4377
rect 9977 4343 10103 4377
rect 10137 4343 10263 4377
rect 10297 4343 10423 4377
rect 10457 4343 10583 4377
rect 10617 4343 10743 4377
rect 10777 4343 10903 4377
rect 10937 4343 11063 4377
rect 11097 4343 11223 4377
rect 11257 4343 11383 4377
rect 11417 4343 11440 4377
rect 9440 4320 11440 4343
rect 11520 4377 11920 4400
rect 11520 4343 11543 4377
rect 11577 4343 11703 4377
rect 11737 4343 11863 4377
rect 11897 4343 11920 4377
rect 11520 4320 11920 4343
rect 12000 4377 12400 4400
rect 12000 4343 12023 4377
rect 12057 4343 12183 4377
rect 12217 4343 12343 4377
rect 12377 4343 12400 4377
rect 12000 4320 12400 4343
rect 8480 4217 8880 4240
rect 8480 4183 8503 4217
rect 8537 4183 8663 4217
rect 8697 4183 8823 4217
rect 8857 4183 8880 4217
rect 8480 4160 8880 4183
rect 8960 4217 9360 4240
rect 8960 4183 8983 4217
rect 9017 4183 9143 4217
rect 9177 4183 9303 4217
rect 9337 4183 9360 4217
rect 8960 4160 9360 4183
rect 9440 4217 11440 4240
rect 9440 4183 9463 4217
rect 9497 4183 9623 4217
rect 9657 4183 9783 4217
rect 9817 4183 9943 4217
rect 9977 4183 10103 4217
rect 10137 4183 10263 4217
rect 10297 4183 10423 4217
rect 10457 4183 10583 4217
rect 10617 4183 10743 4217
rect 10777 4183 10903 4217
rect 10937 4183 11063 4217
rect 11097 4183 11223 4217
rect 11257 4183 11383 4217
rect 11417 4183 11440 4217
rect 9440 4160 11440 4183
rect 11520 4217 11920 4240
rect 11520 4183 11543 4217
rect 11577 4183 11703 4217
rect 11737 4183 11863 4217
rect 11897 4183 11920 4217
rect 11520 4160 11920 4183
rect 12000 4217 12400 4240
rect 12000 4183 12023 4217
rect 12057 4183 12183 4217
rect 12217 4183 12343 4217
rect 12377 4183 12400 4217
rect 12000 4160 12400 4183
rect 8480 4057 8880 4080
rect 8480 4023 8503 4057
rect 8537 4023 8663 4057
rect 8697 4023 8823 4057
rect 8857 4023 8880 4057
rect 8480 4000 8880 4023
rect 8960 4057 9360 4080
rect 8960 4023 8983 4057
rect 9017 4023 9143 4057
rect 9177 4023 9303 4057
rect 9337 4023 9360 4057
rect 8960 4000 9360 4023
rect 9440 4057 11440 4080
rect 9440 4023 9463 4057
rect 9497 4023 9623 4057
rect 9657 4023 9783 4057
rect 9817 4023 9943 4057
rect 9977 4023 10103 4057
rect 10137 4023 10263 4057
rect 10297 4023 10423 4057
rect 10457 4023 10583 4057
rect 10617 4023 10743 4057
rect 10777 4023 10903 4057
rect 10937 4023 11063 4057
rect 11097 4023 11223 4057
rect 11257 4023 11383 4057
rect 11417 4023 11440 4057
rect 9440 4000 11440 4023
rect 11520 4057 11920 4080
rect 11520 4023 11543 4057
rect 11577 4023 11703 4057
rect 11737 4023 11863 4057
rect 11897 4023 11920 4057
rect 11520 4000 11920 4023
rect 12000 4057 12400 4080
rect 12000 4023 12023 4057
rect 12057 4023 12183 4057
rect 12217 4023 12343 4057
rect 12377 4023 12400 4057
rect 12000 4000 12400 4023
rect 8480 3897 8880 3920
rect 8480 3863 8503 3897
rect 8537 3863 8663 3897
rect 8697 3863 8823 3897
rect 8857 3863 8880 3897
rect 8480 3840 8880 3863
rect 8960 3897 9360 3920
rect 8960 3863 8983 3897
rect 9017 3863 9143 3897
rect 9177 3863 9303 3897
rect 9337 3863 9360 3897
rect 8960 3840 9360 3863
rect 9440 3897 11440 3920
rect 9440 3863 9463 3897
rect 9497 3863 9623 3897
rect 9657 3863 9783 3897
rect 9817 3863 9943 3897
rect 9977 3863 10103 3897
rect 10137 3863 10263 3897
rect 10297 3863 10423 3897
rect 10457 3863 10583 3897
rect 10617 3863 10743 3897
rect 10777 3863 10903 3897
rect 10937 3863 11063 3897
rect 11097 3863 11223 3897
rect 11257 3863 11383 3897
rect 11417 3863 11440 3897
rect 9440 3840 11440 3863
rect 11520 3897 11920 3920
rect 11520 3863 11543 3897
rect 11577 3863 11703 3897
rect 11737 3863 11863 3897
rect 11897 3863 11920 3897
rect 11520 3840 11920 3863
rect 12000 3897 12400 3920
rect 12000 3863 12023 3897
rect 12057 3863 12183 3897
rect 12217 3863 12343 3897
rect 12377 3863 12400 3897
rect 12000 3840 12400 3863
rect 8480 3737 8880 3760
rect 8480 3703 8503 3737
rect 8537 3703 8663 3737
rect 8697 3703 8823 3737
rect 8857 3703 8880 3737
rect 8480 3680 8880 3703
rect 8960 3737 9360 3760
rect 8960 3703 8983 3737
rect 9017 3703 9143 3737
rect 9177 3703 9303 3737
rect 9337 3703 9360 3737
rect 8960 3680 9360 3703
rect 9440 3737 11440 3760
rect 9440 3703 9463 3737
rect 9497 3703 9623 3737
rect 9657 3703 9783 3737
rect 9817 3703 9943 3737
rect 9977 3703 10103 3737
rect 10137 3703 10263 3737
rect 10297 3703 10423 3737
rect 10457 3703 10583 3737
rect 10617 3703 10743 3737
rect 10777 3703 10903 3737
rect 10937 3703 11063 3737
rect 11097 3703 11223 3737
rect 11257 3703 11383 3737
rect 11417 3703 11440 3737
rect 9440 3680 11440 3703
rect 11520 3737 11920 3760
rect 11520 3703 11543 3737
rect 11577 3703 11703 3737
rect 11737 3703 11863 3737
rect 11897 3703 11920 3737
rect 11520 3680 11920 3703
rect 12000 3737 12400 3760
rect 12000 3703 12023 3737
rect 12057 3703 12183 3737
rect 12217 3703 12343 3737
rect 12377 3703 12400 3737
rect 12000 3680 12400 3703
rect 8480 3577 8880 3600
rect 8480 3543 8503 3577
rect 8537 3543 8663 3577
rect 8697 3543 8823 3577
rect 8857 3543 8880 3577
rect 8480 3520 8880 3543
rect 8960 3577 9360 3600
rect 8960 3543 8983 3577
rect 9017 3543 9143 3577
rect 9177 3543 9303 3577
rect 9337 3543 9360 3577
rect 8960 3520 9360 3543
rect 9440 3577 11440 3600
rect 9440 3543 9463 3577
rect 9497 3543 9623 3577
rect 9657 3543 9783 3577
rect 9817 3543 9943 3577
rect 9977 3543 10103 3577
rect 10137 3543 10263 3577
rect 10297 3543 10423 3577
rect 10457 3543 10583 3577
rect 10617 3543 10743 3577
rect 10777 3543 10903 3577
rect 10937 3543 11063 3577
rect 11097 3543 11223 3577
rect 11257 3543 11383 3577
rect 11417 3543 11440 3577
rect 9440 3520 11440 3543
rect 11520 3577 11920 3600
rect 11520 3543 11543 3577
rect 11577 3543 11703 3577
rect 11737 3543 11863 3577
rect 11897 3543 11920 3577
rect 11520 3520 11920 3543
rect 12000 3577 12400 3600
rect 12000 3543 12023 3577
rect 12057 3543 12183 3577
rect 12217 3543 12343 3577
rect 12377 3543 12400 3577
rect 12000 3520 12400 3543
rect 8480 3417 8880 3440
rect 8480 3383 8503 3417
rect 8537 3383 8663 3417
rect 8697 3383 8823 3417
rect 8857 3383 8880 3417
rect 8480 3360 8880 3383
rect 8960 3417 9360 3440
rect 8960 3383 8983 3417
rect 9017 3383 9143 3417
rect 9177 3383 9303 3417
rect 9337 3383 9360 3417
rect 8960 3360 9360 3383
rect 9440 3417 11440 3440
rect 9440 3383 9463 3417
rect 9497 3383 9623 3417
rect 9657 3383 9783 3417
rect 9817 3383 9943 3417
rect 9977 3383 10103 3417
rect 10137 3383 10263 3417
rect 10297 3383 10423 3417
rect 10457 3383 10583 3417
rect 10617 3383 10743 3417
rect 10777 3383 10903 3417
rect 10937 3383 11063 3417
rect 11097 3383 11223 3417
rect 11257 3383 11383 3417
rect 11417 3383 11440 3417
rect 9440 3360 11440 3383
rect 11520 3417 11920 3440
rect 11520 3383 11543 3417
rect 11577 3383 11703 3417
rect 11737 3383 11863 3417
rect 11897 3383 11920 3417
rect 11520 3360 11920 3383
rect 12000 3417 12400 3440
rect 12000 3383 12023 3417
rect 12057 3383 12183 3417
rect 12217 3383 12343 3417
rect 12377 3383 12400 3417
rect 12000 3360 12400 3383
rect 8480 3257 8880 3280
rect 8480 3223 8503 3257
rect 8537 3223 8663 3257
rect 8697 3223 8823 3257
rect 8857 3223 8880 3257
rect 8480 3200 8880 3223
rect 8960 3257 9360 3280
rect 8960 3223 8983 3257
rect 9017 3223 9143 3257
rect 9177 3223 9303 3257
rect 9337 3223 9360 3257
rect 8960 3200 9360 3223
rect 9440 3257 11440 3280
rect 9440 3223 9463 3257
rect 9497 3223 9623 3257
rect 9657 3223 9783 3257
rect 9817 3223 9943 3257
rect 9977 3223 10103 3257
rect 10137 3223 10263 3257
rect 10297 3223 10423 3257
rect 10457 3223 10583 3257
rect 10617 3223 10743 3257
rect 10777 3223 10903 3257
rect 10937 3223 11063 3257
rect 11097 3223 11223 3257
rect 11257 3223 11383 3257
rect 11417 3223 11440 3257
rect 9440 3200 11440 3223
rect 11520 3257 11920 3280
rect 11520 3223 11543 3257
rect 11577 3223 11703 3257
rect 11737 3223 11863 3257
rect 11897 3223 11920 3257
rect 11520 3200 11920 3223
rect 12000 3257 12400 3280
rect 12000 3223 12023 3257
rect 12057 3223 12183 3257
rect 12217 3223 12343 3257
rect 12377 3223 12400 3257
rect 12000 3200 12400 3223
rect 8480 3097 8880 3120
rect 8480 3063 8503 3097
rect 8537 3063 8663 3097
rect 8697 3063 8823 3097
rect 8857 3063 8880 3097
rect 8480 3040 8880 3063
rect 8960 3097 9360 3120
rect 8960 3063 8983 3097
rect 9017 3063 9143 3097
rect 9177 3063 9303 3097
rect 9337 3063 9360 3097
rect 8960 3040 9360 3063
rect 9440 3097 11440 3120
rect 9440 3063 9463 3097
rect 9497 3063 9623 3097
rect 9657 3063 9783 3097
rect 9817 3063 9943 3097
rect 9977 3063 10103 3097
rect 10137 3063 10263 3097
rect 10297 3063 10423 3097
rect 10457 3063 10583 3097
rect 10617 3063 10743 3097
rect 10777 3063 10903 3097
rect 10937 3063 11063 3097
rect 11097 3063 11223 3097
rect 11257 3063 11383 3097
rect 11417 3063 11440 3097
rect 9440 3040 11440 3063
rect 11520 3097 11920 3120
rect 11520 3063 11543 3097
rect 11577 3063 11703 3097
rect 11737 3063 11863 3097
rect 11897 3063 11920 3097
rect 11520 3040 11920 3063
rect 12000 3097 12400 3120
rect 12000 3063 12023 3097
rect 12057 3063 12183 3097
rect 12217 3063 12343 3097
rect 12377 3063 12400 3097
rect 12000 3040 12400 3063
rect 8480 2937 8880 2960
rect 8480 2903 8503 2937
rect 8537 2903 8663 2937
rect 8697 2903 8823 2937
rect 8857 2903 8880 2937
rect 8480 2880 8880 2903
rect 8960 2937 9360 2960
rect 8960 2903 8983 2937
rect 9017 2903 9143 2937
rect 9177 2903 9303 2937
rect 9337 2903 9360 2937
rect 8960 2880 9360 2903
rect 9440 2937 11440 2960
rect 9440 2903 9463 2937
rect 9497 2903 9623 2937
rect 9657 2903 9783 2937
rect 9817 2903 9943 2937
rect 9977 2903 10103 2937
rect 10137 2903 10263 2937
rect 10297 2903 10423 2937
rect 10457 2903 10583 2937
rect 10617 2903 10743 2937
rect 10777 2903 10903 2937
rect 10937 2903 11063 2937
rect 11097 2903 11223 2937
rect 11257 2903 11383 2937
rect 11417 2903 11440 2937
rect 9440 2880 11440 2903
rect 11520 2937 11920 2960
rect 11520 2903 11543 2937
rect 11577 2903 11703 2937
rect 11737 2903 11863 2937
rect 11897 2903 11920 2937
rect 11520 2880 11920 2903
rect 12000 2937 12400 2960
rect 12000 2903 12023 2937
rect 12057 2903 12183 2937
rect 12217 2903 12343 2937
rect 12377 2903 12400 2937
rect 12000 2880 12400 2903
rect 8480 2777 8880 2800
rect 8480 2743 8503 2777
rect 8537 2743 8663 2777
rect 8697 2743 8823 2777
rect 8857 2743 8880 2777
rect 8480 2720 8880 2743
rect 8960 2777 9360 2800
rect 8960 2743 8983 2777
rect 9017 2743 9143 2777
rect 9177 2743 9303 2777
rect 9337 2743 9360 2777
rect 8960 2720 9360 2743
rect 9440 2777 11440 2800
rect 9440 2743 9463 2777
rect 9497 2743 9623 2777
rect 9657 2743 9783 2777
rect 9817 2743 9943 2777
rect 9977 2743 10103 2777
rect 10137 2743 10263 2777
rect 10297 2743 10423 2777
rect 10457 2743 10583 2777
rect 10617 2743 10743 2777
rect 10777 2743 10903 2777
rect 10937 2743 11063 2777
rect 11097 2743 11223 2777
rect 11257 2743 11383 2777
rect 11417 2743 11440 2777
rect 9440 2720 11440 2743
rect 11520 2777 11920 2800
rect 11520 2743 11543 2777
rect 11577 2743 11703 2777
rect 11737 2743 11863 2777
rect 11897 2743 11920 2777
rect 11520 2720 11920 2743
rect 12000 2777 12400 2800
rect 12000 2743 12023 2777
rect 12057 2743 12183 2777
rect 12217 2743 12343 2777
rect 12377 2743 12400 2777
rect 12000 2720 12400 2743
rect 8480 2617 8880 2640
rect 8480 2583 8503 2617
rect 8537 2583 8663 2617
rect 8697 2583 8823 2617
rect 8857 2583 8880 2617
rect 8480 2560 8880 2583
rect 8960 2617 9360 2640
rect 8960 2583 8983 2617
rect 9017 2583 9143 2617
rect 9177 2583 9303 2617
rect 9337 2583 9360 2617
rect 8960 2560 9360 2583
rect 9440 2617 11440 2640
rect 9440 2583 9463 2617
rect 9497 2583 9623 2617
rect 9657 2583 9783 2617
rect 9817 2583 9943 2617
rect 9977 2583 10103 2617
rect 10137 2583 10263 2617
rect 10297 2583 10423 2617
rect 10457 2583 10583 2617
rect 10617 2583 10743 2617
rect 10777 2583 10903 2617
rect 10937 2583 11063 2617
rect 11097 2583 11223 2617
rect 11257 2583 11383 2617
rect 11417 2583 11440 2617
rect 9440 2560 11440 2583
rect 11520 2617 11920 2640
rect 11520 2583 11543 2617
rect 11577 2583 11703 2617
rect 11737 2583 11863 2617
rect 11897 2583 11920 2617
rect 11520 2560 11920 2583
rect 12000 2617 12400 2640
rect 12000 2583 12023 2617
rect 12057 2583 12183 2617
rect 12217 2583 12343 2617
rect 12377 2583 12400 2617
rect 12000 2560 12400 2583
rect 8480 2457 8880 2480
rect 8480 2423 8503 2457
rect 8537 2423 8663 2457
rect 8697 2423 8823 2457
rect 8857 2423 8880 2457
rect 8480 2400 8880 2423
rect 8960 2457 9360 2480
rect 8960 2423 8983 2457
rect 9017 2423 9143 2457
rect 9177 2423 9303 2457
rect 9337 2423 9360 2457
rect 8960 2400 9360 2423
rect 9440 2457 11440 2480
rect 9440 2423 9463 2457
rect 9497 2423 9623 2457
rect 9657 2423 9783 2457
rect 9817 2423 9943 2457
rect 9977 2423 10103 2457
rect 10137 2423 10263 2457
rect 10297 2423 10423 2457
rect 10457 2423 10583 2457
rect 10617 2423 10743 2457
rect 10777 2423 10903 2457
rect 10937 2423 11063 2457
rect 11097 2423 11223 2457
rect 11257 2423 11383 2457
rect 11417 2423 11440 2457
rect 9440 2400 11440 2423
rect 11520 2457 11920 2480
rect 11520 2423 11543 2457
rect 11577 2423 11703 2457
rect 11737 2423 11863 2457
rect 11897 2423 11920 2457
rect 11520 2400 11920 2423
rect 12000 2457 12400 2480
rect 12000 2423 12023 2457
rect 12057 2423 12183 2457
rect 12217 2423 12343 2457
rect 12377 2423 12400 2457
rect 12000 2400 12400 2423
rect 8480 2297 8880 2320
rect 8480 2263 8503 2297
rect 8537 2263 8663 2297
rect 8697 2263 8823 2297
rect 8857 2263 8880 2297
rect 8480 2240 8880 2263
rect 8960 2297 9360 2320
rect 8960 2263 8983 2297
rect 9017 2263 9143 2297
rect 9177 2263 9303 2297
rect 9337 2263 9360 2297
rect 8960 2240 9360 2263
rect 9440 2297 11440 2320
rect 9440 2263 9463 2297
rect 9497 2263 9623 2297
rect 9657 2263 9783 2297
rect 9817 2263 9943 2297
rect 9977 2263 10103 2297
rect 10137 2263 10263 2297
rect 10297 2263 10423 2297
rect 10457 2263 10583 2297
rect 10617 2263 10743 2297
rect 10777 2263 10903 2297
rect 10937 2263 11063 2297
rect 11097 2263 11223 2297
rect 11257 2263 11383 2297
rect 11417 2263 11440 2297
rect 9440 2240 11440 2263
rect 11520 2297 11920 2320
rect 11520 2263 11543 2297
rect 11577 2263 11703 2297
rect 11737 2263 11863 2297
rect 11897 2263 11920 2297
rect 11520 2240 11920 2263
rect 12000 2297 12400 2320
rect 12000 2263 12023 2297
rect 12057 2263 12183 2297
rect 12217 2263 12343 2297
rect 12377 2263 12400 2297
rect 12000 2240 12400 2263
rect 8480 2137 8880 2160
rect 8480 2103 8503 2137
rect 8537 2103 8663 2137
rect 8697 2103 8823 2137
rect 8857 2103 8880 2137
rect 8480 2080 8880 2103
rect 8960 2137 9360 2160
rect 8960 2103 8983 2137
rect 9017 2103 9143 2137
rect 9177 2103 9303 2137
rect 9337 2103 9360 2137
rect 8960 2080 9360 2103
rect 9440 2137 11440 2160
rect 9440 2103 9463 2137
rect 9497 2103 9623 2137
rect 9657 2103 9783 2137
rect 9817 2103 9943 2137
rect 9977 2103 10103 2137
rect 10137 2103 10263 2137
rect 10297 2103 10423 2137
rect 10457 2103 10583 2137
rect 10617 2103 10743 2137
rect 10777 2103 10903 2137
rect 10937 2103 11063 2137
rect 11097 2103 11223 2137
rect 11257 2103 11383 2137
rect 11417 2103 11440 2137
rect 9440 2080 11440 2103
rect 11520 2137 11920 2160
rect 11520 2103 11543 2137
rect 11577 2103 11703 2137
rect 11737 2103 11863 2137
rect 11897 2103 11920 2137
rect 11520 2080 11920 2103
rect 12000 2137 12400 2160
rect 12000 2103 12023 2137
rect 12057 2103 12183 2137
rect 12217 2103 12343 2137
rect 12377 2103 12400 2137
rect 12000 2080 12400 2103
rect 8480 1977 8880 2000
rect 8480 1943 8503 1977
rect 8537 1943 8663 1977
rect 8697 1943 8823 1977
rect 8857 1943 8880 1977
rect 8480 1920 8880 1943
rect 8960 1977 9360 2000
rect 8960 1943 8983 1977
rect 9017 1943 9143 1977
rect 9177 1943 9303 1977
rect 9337 1943 9360 1977
rect 8960 1920 9360 1943
rect 9440 1977 11440 2000
rect 9440 1943 9463 1977
rect 9497 1943 9623 1977
rect 9657 1943 9783 1977
rect 9817 1943 9943 1977
rect 9977 1943 10103 1977
rect 10137 1943 10263 1977
rect 10297 1943 10423 1977
rect 10457 1943 10583 1977
rect 10617 1943 10743 1977
rect 10777 1943 10903 1977
rect 10937 1943 11063 1977
rect 11097 1943 11223 1977
rect 11257 1943 11383 1977
rect 11417 1943 11440 1977
rect 9440 1920 11440 1943
rect 11520 1977 11920 2000
rect 11520 1943 11543 1977
rect 11577 1943 11703 1977
rect 11737 1943 11863 1977
rect 11897 1943 11920 1977
rect 11520 1920 11920 1943
rect 12000 1977 12400 2000
rect 12000 1943 12023 1977
rect 12057 1943 12183 1977
rect 12217 1943 12343 1977
rect 12377 1943 12400 1977
rect 12000 1920 12400 1943
rect 8480 1817 8880 1840
rect 8480 1783 8503 1817
rect 8537 1783 8663 1817
rect 8697 1783 8823 1817
rect 8857 1783 8880 1817
rect 8480 1760 8880 1783
rect 8960 1817 9360 1840
rect 8960 1783 8983 1817
rect 9017 1783 9143 1817
rect 9177 1783 9303 1817
rect 9337 1783 9360 1817
rect 8960 1760 9360 1783
rect 9440 1817 11440 1840
rect 9440 1783 9463 1817
rect 9497 1783 9623 1817
rect 9657 1783 9783 1817
rect 9817 1783 9943 1817
rect 9977 1783 10103 1817
rect 10137 1783 10263 1817
rect 10297 1783 10423 1817
rect 10457 1783 10583 1817
rect 10617 1783 10743 1817
rect 10777 1783 10903 1817
rect 10937 1783 11063 1817
rect 11097 1783 11223 1817
rect 11257 1783 11383 1817
rect 11417 1783 11440 1817
rect 9440 1760 11440 1783
rect 11520 1817 11920 1840
rect 11520 1783 11543 1817
rect 11577 1783 11703 1817
rect 11737 1783 11863 1817
rect 11897 1783 11920 1817
rect 11520 1760 11920 1783
rect 12000 1817 12400 1840
rect 12000 1783 12023 1817
rect 12057 1783 12183 1817
rect 12217 1783 12343 1817
rect 12377 1783 12400 1817
rect 12000 1760 12400 1783
rect 8480 1657 8880 1680
rect 8480 1623 8503 1657
rect 8537 1623 8663 1657
rect 8697 1623 8823 1657
rect 8857 1623 8880 1657
rect 8480 1600 8880 1623
rect 8960 1657 9360 1680
rect 8960 1623 8983 1657
rect 9017 1623 9143 1657
rect 9177 1623 9303 1657
rect 9337 1623 9360 1657
rect 8960 1600 9360 1623
rect 9440 1657 11440 1680
rect 9440 1623 9463 1657
rect 9497 1623 9623 1657
rect 9657 1623 9783 1657
rect 9817 1623 9943 1657
rect 9977 1623 10103 1657
rect 10137 1623 10263 1657
rect 10297 1623 10423 1657
rect 10457 1623 10583 1657
rect 10617 1623 10743 1657
rect 10777 1623 10903 1657
rect 10937 1623 11063 1657
rect 11097 1623 11223 1657
rect 11257 1623 11383 1657
rect 11417 1623 11440 1657
rect 9440 1600 11440 1623
rect 11520 1657 11920 1680
rect 11520 1623 11543 1657
rect 11577 1623 11703 1657
rect 11737 1623 11863 1657
rect 11897 1623 11920 1657
rect 11520 1600 11920 1623
rect 12000 1657 12400 1680
rect 12000 1623 12023 1657
rect 12057 1623 12183 1657
rect 12217 1623 12343 1657
rect 12377 1623 12400 1657
rect 12000 1600 12400 1623
rect 8480 1497 8880 1520
rect 8480 1463 8503 1497
rect 8537 1463 8663 1497
rect 8697 1463 8823 1497
rect 8857 1463 8880 1497
rect 8480 1440 8880 1463
rect 8960 1497 9360 1520
rect 8960 1463 8983 1497
rect 9017 1463 9143 1497
rect 9177 1463 9303 1497
rect 9337 1463 9360 1497
rect 8960 1440 9360 1463
rect 9440 1497 11440 1520
rect 9440 1463 9463 1497
rect 9497 1463 9623 1497
rect 9657 1463 9783 1497
rect 9817 1463 9943 1497
rect 9977 1463 10103 1497
rect 10137 1463 10263 1497
rect 10297 1463 10423 1497
rect 10457 1463 10583 1497
rect 10617 1463 10743 1497
rect 10777 1463 10903 1497
rect 10937 1463 11063 1497
rect 11097 1463 11223 1497
rect 11257 1463 11383 1497
rect 11417 1463 11440 1497
rect 9440 1440 11440 1463
rect 11520 1497 11920 1520
rect 11520 1463 11543 1497
rect 11577 1463 11703 1497
rect 11737 1463 11863 1497
rect 11897 1463 11920 1497
rect 11520 1440 11920 1463
rect 12000 1497 12400 1520
rect 12000 1463 12023 1497
rect 12057 1463 12183 1497
rect 12217 1463 12343 1497
rect 12377 1463 12400 1497
rect 12000 1440 12400 1463
rect 8480 1337 8880 1360
rect 8480 1303 8503 1337
rect 8537 1303 8663 1337
rect 8697 1303 8823 1337
rect 8857 1303 8880 1337
rect 8480 1280 8880 1303
rect 8960 1337 9360 1360
rect 8960 1303 8983 1337
rect 9017 1303 9143 1337
rect 9177 1303 9303 1337
rect 9337 1303 9360 1337
rect 8960 1280 9360 1303
rect 9440 1337 11440 1360
rect 9440 1303 9463 1337
rect 9497 1303 9623 1337
rect 9657 1303 9783 1337
rect 9817 1303 9943 1337
rect 9977 1303 10103 1337
rect 10137 1303 10263 1337
rect 10297 1303 10423 1337
rect 10457 1303 10583 1337
rect 10617 1303 10743 1337
rect 10777 1303 10903 1337
rect 10937 1303 11063 1337
rect 11097 1303 11223 1337
rect 11257 1303 11383 1337
rect 11417 1303 11440 1337
rect 9440 1280 11440 1303
rect 11520 1337 11920 1360
rect 11520 1303 11543 1337
rect 11577 1303 11703 1337
rect 11737 1303 11863 1337
rect 11897 1303 11920 1337
rect 11520 1280 11920 1303
rect 12000 1337 12400 1360
rect 12000 1303 12023 1337
rect 12057 1303 12183 1337
rect 12217 1303 12343 1337
rect 12377 1303 12400 1337
rect 12000 1280 12400 1303
rect 8480 1177 8880 1200
rect 8480 1143 8503 1177
rect 8537 1143 8663 1177
rect 8697 1143 8823 1177
rect 8857 1143 8880 1177
rect 8480 1120 8880 1143
rect 8960 1177 9360 1200
rect 8960 1143 8983 1177
rect 9017 1143 9143 1177
rect 9177 1143 9303 1177
rect 9337 1143 9360 1177
rect 8960 1120 9360 1143
rect 9440 1177 11440 1200
rect 9440 1143 9463 1177
rect 9497 1143 9623 1177
rect 9657 1143 9783 1177
rect 9817 1143 9943 1177
rect 9977 1143 10103 1177
rect 10137 1143 10263 1177
rect 10297 1143 10423 1177
rect 10457 1143 10583 1177
rect 10617 1143 10743 1177
rect 10777 1143 10903 1177
rect 10937 1143 11063 1177
rect 11097 1143 11223 1177
rect 11257 1143 11383 1177
rect 11417 1143 11440 1177
rect 9440 1120 11440 1143
rect 11520 1177 11920 1200
rect 11520 1143 11543 1177
rect 11577 1143 11703 1177
rect 11737 1143 11863 1177
rect 11897 1143 11920 1177
rect 11520 1120 11920 1143
rect 12000 1177 12400 1200
rect 12000 1143 12023 1177
rect 12057 1143 12183 1177
rect 12217 1143 12343 1177
rect 12377 1143 12400 1177
rect 12000 1120 12400 1143
rect 8480 1017 8880 1040
rect 8480 983 8503 1017
rect 8537 983 8663 1017
rect 8697 983 8823 1017
rect 8857 983 8880 1017
rect 8480 960 8880 983
rect 8960 1017 9360 1040
rect 8960 983 8983 1017
rect 9017 983 9143 1017
rect 9177 983 9303 1017
rect 9337 983 9360 1017
rect 8960 960 9360 983
rect 9440 1017 11440 1040
rect 9440 983 9463 1017
rect 9497 983 9623 1017
rect 9657 983 9783 1017
rect 9817 983 9943 1017
rect 9977 983 10103 1017
rect 10137 983 10263 1017
rect 10297 983 10423 1017
rect 10457 983 10583 1017
rect 10617 983 10743 1017
rect 10777 983 10903 1017
rect 10937 983 11063 1017
rect 11097 983 11223 1017
rect 11257 983 11383 1017
rect 11417 983 11440 1017
rect 9440 960 11440 983
rect 11520 1017 11920 1040
rect 11520 983 11543 1017
rect 11577 983 11703 1017
rect 11737 983 11863 1017
rect 11897 983 11920 1017
rect 11520 960 11920 983
rect 12000 1017 12400 1040
rect 12000 983 12023 1017
rect 12057 983 12183 1017
rect 12217 983 12343 1017
rect 12377 983 12400 1017
rect 12000 960 12400 983
rect 8480 857 8880 880
rect 8480 823 8503 857
rect 8537 823 8663 857
rect 8697 823 8823 857
rect 8857 823 8880 857
rect 8480 800 8880 823
rect 8960 857 9360 880
rect 8960 823 8983 857
rect 9017 823 9143 857
rect 9177 823 9303 857
rect 9337 823 9360 857
rect 8960 800 9360 823
rect 9440 857 11440 880
rect 9440 823 9463 857
rect 9497 823 9623 857
rect 9657 823 9783 857
rect 9817 823 9943 857
rect 9977 823 10103 857
rect 10137 823 10263 857
rect 10297 823 10423 857
rect 10457 823 10583 857
rect 10617 823 10743 857
rect 10777 823 10903 857
rect 10937 823 11063 857
rect 11097 823 11223 857
rect 11257 823 11383 857
rect 11417 823 11440 857
rect 9440 800 11440 823
rect 11520 857 11920 880
rect 11520 823 11543 857
rect 11577 823 11703 857
rect 11737 823 11863 857
rect 11897 823 11920 857
rect 11520 800 11920 823
rect 12000 857 12400 880
rect 12000 823 12023 857
rect 12057 823 12183 857
rect 12217 823 12343 857
rect 12377 823 12400 857
rect 12000 800 12400 823
rect 8480 697 8880 720
rect 8480 663 8503 697
rect 8537 663 8663 697
rect 8697 663 8823 697
rect 8857 663 8880 697
rect 8480 640 8880 663
rect 8960 697 9360 720
rect 8960 663 8983 697
rect 9017 663 9143 697
rect 9177 663 9303 697
rect 9337 663 9360 697
rect 8960 640 9360 663
rect 9440 697 11440 720
rect 9440 663 9463 697
rect 9497 663 9623 697
rect 9657 663 9783 697
rect 9817 663 9943 697
rect 9977 663 10103 697
rect 10137 663 10263 697
rect 10297 663 10423 697
rect 10457 663 10583 697
rect 10617 663 10743 697
rect 10777 663 10903 697
rect 10937 663 11063 697
rect 11097 663 11223 697
rect 11257 663 11383 697
rect 11417 663 11440 697
rect 9440 640 11440 663
rect 11520 697 11920 720
rect 11520 663 11543 697
rect 11577 663 11703 697
rect 11737 663 11863 697
rect 11897 663 11920 697
rect 11520 640 11920 663
rect 12000 697 12400 720
rect 12000 663 12023 697
rect 12057 663 12183 697
rect 12217 663 12343 697
rect 12377 663 12400 697
rect 12000 640 12400 663
rect 8480 537 8880 560
rect 8480 503 8503 537
rect 8537 503 8663 537
rect 8697 503 8823 537
rect 8857 503 8880 537
rect 8480 480 8880 503
rect 8960 537 9360 560
rect 8960 503 8983 537
rect 9017 503 9143 537
rect 9177 503 9303 537
rect 9337 503 9360 537
rect 8960 480 9360 503
rect 9440 537 11440 560
rect 9440 503 9463 537
rect 9497 503 9623 537
rect 9657 503 9783 537
rect 9817 503 9943 537
rect 9977 503 10103 537
rect 10137 503 10263 537
rect 10297 503 10423 537
rect 10457 503 10583 537
rect 10617 503 10743 537
rect 10777 503 10903 537
rect 10937 503 11063 537
rect 11097 503 11223 537
rect 11257 503 11383 537
rect 11417 503 11440 537
rect 9440 480 11440 503
rect 11520 537 11920 560
rect 11520 503 11543 537
rect 11577 503 11703 537
rect 11737 503 11863 537
rect 11897 503 11920 537
rect 11520 480 11920 503
rect 12000 537 12400 560
rect 12000 503 12023 537
rect 12057 503 12183 537
rect 12217 503 12343 537
rect 12377 503 12400 537
rect 12000 480 12400 503
rect 8480 377 8880 400
rect 8480 343 8503 377
rect 8537 343 8663 377
rect 8697 343 8823 377
rect 8857 343 8880 377
rect 8480 320 8880 343
rect 8960 377 9360 400
rect 8960 343 8983 377
rect 9017 343 9143 377
rect 9177 343 9303 377
rect 9337 343 9360 377
rect 8960 320 9360 343
rect 9440 377 11440 400
rect 9440 343 9463 377
rect 9497 343 9623 377
rect 9657 343 9783 377
rect 9817 343 9943 377
rect 9977 343 10103 377
rect 10137 343 10263 377
rect 10297 343 10423 377
rect 10457 343 10583 377
rect 10617 343 10743 377
rect 10777 343 10903 377
rect 10937 343 11063 377
rect 11097 343 11223 377
rect 11257 343 11383 377
rect 11417 343 11440 377
rect 9440 320 11440 343
rect 11520 377 11920 400
rect 11520 343 11543 377
rect 11577 343 11703 377
rect 11737 343 11863 377
rect 11897 343 11920 377
rect 11520 320 11920 343
rect 12000 377 12400 400
rect 12000 343 12023 377
rect 12057 343 12183 377
rect 12217 343 12343 377
rect 12377 343 12400 377
rect 12000 320 12400 343
rect 8480 217 8880 240
rect 8480 183 8503 217
rect 8537 183 8663 217
rect 8697 183 8823 217
rect 8857 183 8880 217
rect 8480 160 8880 183
rect 8960 217 9360 240
rect 8960 183 8983 217
rect 9017 183 9143 217
rect 9177 183 9303 217
rect 9337 183 9360 217
rect 8960 160 9360 183
rect 9440 217 11440 240
rect 9440 183 9463 217
rect 9497 183 9623 217
rect 9657 183 9783 217
rect 9817 183 9943 217
rect 9977 183 10103 217
rect 10137 183 10263 217
rect 10297 183 10423 217
rect 10457 183 10583 217
rect 10617 183 10743 217
rect 10777 183 10903 217
rect 10937 183 11063 217
rect 11097 183 11223 217
rect 11257 183 11383 217
rect 11417 183 11440 217
rect 9440 160 11440 183
rect 11520 217 11920 240
rect 11520 183 11543 217
rect 11577 183 11703 217
rect 11737 183 11863 217
rect 11897 183 11920 217
rect 11520 160 11920 183
rect 12000 217 12400 240
rect 12000 183 12023 217
rect 12057 183 12183 217
rect 12217 183 12343 217
rect 12377 183 12400 217
rect 12000 160 12400 183
rect 8480 57 8880 80
rect 8480 23 8503 57
rect 8537 23 8663 57
rect 8697 23 8823 57
rect 8857 23 8880 57
rect 8480 0 8880 23
rect 8960 57 9360 80
rect 8960 23 8983 57
rect 9017 23 9143 57
rect 9177 23 9303 57
rect 9337 23 9360 57
rect 8960 0 9360 23
rect 9440 57 11440 80
rect 9440 23 9463 57
rect 9497 23 9623 57
rect 9657 23 9783 57
rect 9817 23 9943 57
rect 9977 23 10103 57
rect 10137 23 10263 57
rect 10297 23 10423 57
rect 10457 23 10583 57
rect 10617 23 10743 57
rect 10777 23 10903 57
rect 10937 23 11063 57
rect 11097 23 11223 57
rect 11257 23 11383 57
rect 11417 23 11440 57
rect 9440 0 11440 23
rect 11520 57 11920 80
rect 11520 23 11543 57
rect 11577 23 11703 57
rect 11737 23 11863 57
rect 11897 23 11920 57
rect 11520 0 11920 23
rect 12000 57 12400 80
rect 12000 23 12023 57
rect 12057 23 12183 57
rect 12217 23 12343 57
rect 12377 23 12400 57
rect 12000 0 12400 23
<< viali >>
rect 8503 31383 8537 31417
rect 8663 31383 8697 31417
rect 8823 31383 8857 31417
rect 8983 31383 9017 31417
rect 9143 31383 9177 31417
rect 9303 31383 9337 31417
rect 9463 31383 9497 31417
rect 9623 31383 9657 31417
rect 9783 31383 9817 31417
rect 9943 31383 9977 31417
rect 10103 31383 10137 31417
rect 10263 31383 10297 31417
rect 10423 31383 10457 31417
rect 10583 31383 10617 31417
rect 10743 31383 10777 31417
rect 10903 31383 10937 31417
rect 11063 31383 11097 31417
rect 11223 31383 11257 31417
rect 11383 31383 11417 31417
rect 11543 31383 11577 31417
rect 11703 31383 11737 31417
rect 11863 31383 11897 31417
rect 12023 31383 12057 31417
rect 12183 31383 12217 31417
rect 12343 31383 12377 31417
rect 8503 31223 8537 31257
rect 8663 31223 8697 31257
rect 8823 31223 8857 31257
rect 8983 31223 9017 31257
rect 9143 31223 9177 31257
rect 9303 31223 9337 31257
rect 9463 31223 9497 31257
rect 9623 31223 9657 31257
rect 9783 31223 9817 31257
rect 9943 31223 9977 31257
rect 10103 31223 10137 31257
rect 10263 31223 10297 31257
rect 10423 31223 10457 31257
rect 10583 31223 10617 31257
rect 10743 31223 10777 31257
rect 10903 31223 10937 31257
rect 11063 31223 11097 31257
rect 11223 31223 11257 31257
rect 11383 31223 11417 31257
rect 11543 31223 11577 31257
rect 11703 31223 11737 31257
rect 11863 31223 11897 31257
rect 12023 31223 12057 31257
rect 12183 31223 12217 31257
rect 12343 31223 12377 31257
rect 8503 31063 8537 31097
rect 8663 31063 8697 31097
rect 8823 31063 8857 31097
rect 8983 31063 9017 31097
rect 9143 31063 9177 31097
rect 9303 31063 9337 31097
rect 9463 31063 9497 31097
rect 9623 31063 9657 31097
rect 9783 31063 9817 31097
rect 9943 31063 9977 31097
rect 10103 31063 10137 31097
rect 10263 31063 10297 31097
rect 10423 31063 10457 31097
rect 10583 31063 10617 31097
rect 10743 31063 10777 31097
rect 10903 31063 10937 31097
rect 11063 31063 11097 31097
rect 11223 31063 11257 31097
rect 11383 31063 11417 31097
rect 11543 31063 11577 31097
rect 11703 31063 11737 31097
rect 11863 31063 11897 31097
rect 12023 31063 12057 31097
rect 12183 31063 12217 31097
rect 12343 31063 12377 31097
rect 8503 30903 8537 30937
rect 8663 30903 8697 30937
rect 8823 30903 8857 30937
rect 8983 30903 9017 30937
rect 9143 30903 9177 30937
rect 9303 30903 9337 30937
rect 9463 30903 9497 30937
rect 9623 30903 9657 30937
rect 9783 30903 9817 30937
rect 9943 30903 9977 30937
rect 10103 30903 10137 30937
rect 10263 30903 10297 30937
rect 10423 30903 10457 30937
rect 10583 30903 10617 30937
rect 10743 30903 10777 30937
rect 10903 30903 10937 30937
rect 11063 30903 11097 30937
rect 11223 30903 11257 30937
rect 11383 30903 11417 30937
rect 11543 30903 11577 30937
rect 11703 30903 11737 30937
rect 11863 30903 11897 30937
rect 12023 30903 12057 30937
rect 12183 30903 12217 30937
rect 12343 30903 12377 30937
rect 8503 30743 8537 30777
rect 8663 30743 8697 30777
rect 8823 30743 8857 30777
rect 8983 30743 9017 30777
rect 9143 30743 9177 30777
rect 9303 30743 9337 30777
rect 9463 30743 9497 30777
rect 9623 30743 9657 30777
rect 9783 30743 9817 30777
rect 9943 30743 9977 30777
rect 10103 30743 10137 30777
rect 10263 30743 10297 30777
rect 10423 30743 10457 30777
rect 10583 30743 10617 30777
rect 10743 30743 10777 30777
rect 10903 30743 10937 30777
rect 11063 30743 11097 30777
rect 11223 30743 11257 30777
rect 11383 30743 11417 30777
rect 11543 30743 11577 30777
rect 11703 30743 11737 30777
rect 11863 30743 11897 30777
rect 12023 30743 12057 30777
rect 12183 30743 12217 30777
rect 12343 30743 12377 30777
rect 8503 30583 8537 30617
rect 8663 30583 8697 30617
rect 8823 30583 8857 30617
rect 8983 30583 9017 30617
rect 9143 30583 9177 30617
rect 9303 30583 9337 30617
rect 9463 30583 9497 30617
rect 9623 30583 9657 30617
rect 9783 30583 9817 30617
rect 9943 30583 9977 30617
rect 10103 30583 10137 30617
rect 10263 30583 10297 30617
rect 10423 30583 10457 30617
rect 10583 30583 10617 30617
rect 10743 30583 10777 30617
rect 10903 30583 10937 30617
rect 11063 30583 11097 30617
rect 11223 30583 11257 30617
rect 11383 30583 11417 30617
rect 11543 30583 11577 30617
rect 11703 30583 11737 30617
rect 11863 30583 11897 30617
rect 12023 30583 12057 30617
rect 12183 30583 12217 30617
rect 12343 30583 12377 30617
rect 8503 30423 8537 30457
rect 8663 30423 8697 30457
rect 8823 30423 8857 30457
rect 8983 30423 9017 30457
rect 9143 30423 9177 30457
rect 9303 30423 9337 30457
rect 9463 30423 9497 30457
rect 9623 30423 9657 30457
rect 9783 30423 9817 30457
rect 9943 30423 9977 30457
rect 10103 30423 10137 30457
rect 10263 30423 10297 30457
rect 10423 30423 10457 30457
rect 10583 30423 10617 30457
rect 10743 30423 10777 30457
rect 10903 30423 10937 30457
rect 11063 30423 11097 30457
rect 11223 30423 11257 30457
rect 11383 30423 11417 30457
rect 11543 30423 11577 30457
rect 11703 30423 11737 30457
rect 11863 30423 11897 30457
rect 12023 30423 12057 30457
rect 12183 30423 12217 30457
rect 12343 30423 12377 30457
rect 8503 30263 8537 30297
rect 8663 30263 8697 30297
rect 8823 30263 8857 30297
rect 8983 30263 9017 30297
rect 9143 30263 9177 30297
rect 9303 30263 9337 30297
rect 9463 30263 9497 30297
rect 9623 30263 9657 30297
rect 9783 30263 9817 30297
rect 9943 30263 9977 30297
rect 10103 30263 10137 30297
rect 10263 30263 10297 30297
rect 10423 30263 10457 30297
rect 10583 30263 10617 30297
rect 10743 30263 10777 30297
rect 10903 30263 10937 30297
rect 11063 30263 11097 30297
rect 11223 30263 11257 30297
rect 11383 30263 11417 30297
rect 11543 30263 11577 30297
rect 11703 30263 11737 30297
rect 11863 30263 11897 30297
rect 12023 30263 12057 30297
rect 12183 30263 12217 30297
rect 12343 30263 12377 30297
rect 8503 30103 8537 30137
rect 8663 30103 8697 30137
rect 8823 30103 8857 30137
rect 8983 30103 9017 30137
rect 9143 30103 9177 30137
rect 9303 30103 9337 30137
rect 9463 30103 9497 30137
rect 9623 30103 9657 30137
rect 9783 30103 9817 30137
rect 9943 30103 9977 30137
rect 10103 30103 10137 30137
rect 10263 30103 10297 30137
rect 10423 30103 10457 30137
rect 10583 30103 10617 30137
rect 10743 30103 10777 30137
rect 10903 30103 10937 30137
rect 11063 30103 11097 30137
rect 11223 30103 11257 30137
rect 11383 30103 11417 30137
rect 11543 30103 11577 30137
rect 11703 30103 11737 30137
rect 11863 30103 11897 30137
rect 12023 30103 12057 30137
rect 12183 30103 12217 30137
rect 12343 30103 12377 30137
rect 8503 29943 8537 29977
rect 8663 29943 8697 29977
rect 8823 29943 8857 29977
rect 8983 29943 9017 29977
rect 9143 29943 9177 29977
rect 9303 29943 9337 29977
rect 9463 29943 9497 29977
rect 9623 29943 9657 29977
rect 9783 29943 9817 29977
rect 9943 29943 9977 29977
rect 10103 29943 10137 29977
rect 10263 29943 10297 29977
rect 10423 29943 10457 29977
rect 10583 29943 10617 29977
rect 10743 29943 10777 29977
rect 10903 29943 10937 29977
rect 11063 29943 11097 29977
rect 11223 29943 11257 29977
rect 11383 29943 11417 29977
rect 11543 29943 11577 29977
rect 11703 29943 11737 29977
rect 11863 29943 11897 29977
rect 12023 29943 12057 29977
rect 12183 29943 12217 29977
rect 12343 29943 12377 29977
rect 8503 29783 8537 29817
rect 8663 29783 8697 29817
rect 8823 29783 8857 29817
rect 8983 29783 9017 29817
rect 9143 29783 9177 29817
rect 9303 29783 9337 29817
rect 9463 29783 9497 29817
rect 9623 29783 9657 29817
rect 9783 29783 9817 29817
rect 9943 29783 9977 29817
rect 10103 29783 10137 29817
rect 10263 29783 10297 29817
rect 10423 29783 10457 29817
rect 10583 29783 10617 29817
rect 10743 29783 10777 29817
rect 10903 29783 10937 29817
rect 11063 29783 11097 29817
rect 11223 29783 11257 29817
rect 11383 29783 11417 29817
rect 11543 29783 11577 29817
rect 11703 29783 11737 29817
rect 11863 29783 11897 29817
rect 12023 29783 12057 29817
rect 12183 29783 12217 29817
rect 12343 29783 12377 29817
rect 8503 29623 8537 29657
rect 8663 29623 8697 29657
rect 8823 29623 8857 29657
rect 8983 29623 9017 29657
rect 9143 29623 9177 29657
rect 9303 29623 9337 29657
rect 9463 29623 9497 29657
rect 9623 29623 9657 29657
rect 9783 29623 9817 29657
rect 9943 29623 9977 29657
rect 10103 29623 10137 29657
rect 10263 29623 10297 29657
rect 10423 29623 10457 29657
rect 10583 29623 10617 29657
rect 10743 29623 10777 29657
rect 10903 29623 10937 29657
rect 11063 29623 11097 29657
rect 11223 29623 11257 29657
rect 11383 29623 11417 29657
rect 11543 29623 11577 29657
rect 11703 29623 11737 29657
rect 11863 29623 11897 29657
rect 12023 29623 12057 29657
rect 12183 29623 12217 29657
rect 12343 29623 12377 29657
rect 8503 29463 8537 29497
rect 8663 29463 8697 29497
rect 8823 29463 8857 29497
rect 8983 29463 9017 29497
rect 9143 29463 9177 29497
rect 9303 29463 9337 29497
rect 9463 29463 9497 29497
rect 9623 29463 9657 29497
rect 9783 29463 9817 29497
rect 9943 29463 9977 29497
rect 10103 29463 10137 29497
rect 10263 29463 10297 29497
rect 10423 29463 10457 29497
rect 10583 29463 10617 29497
rect 10743 29463 10777 29497
rect 10903 29463 10937 29497
rect 11063 29463 11097 29497
rect 11223 29463 11257 29497
rect 11383 29463 11417 29497
rect 11543 29463 11577 29497
rect 11703 29463 11737 29497
rect 11863 29463 11897 29497
rect 12023 29463 12057 29497
rect 12183 29463 12217 29497
rect 12343 29463 12377 29497
rect 8503 29303 8537 29337
rect 8663 29303 8697 29337
rect 8823 29303 8857 29337
rect 8983 29303 9017 29337
rect 9143 29303 9177 29337
rect 9303 29303 9337 29337
rect 9463 29303 9497 29337
rect 9623 29303 9657 29337
rect 9783 29303 9817 29337
rect 9943 29303 9977 29337
rect 10103 29303 10137 29337
rect 10263 29303 10297 29337
rect 10423 29303 10457 29337
rect 10583 29303 10617 29337
rect 10743 29303 10777 29337
rect 10903 29303 10937 29337
rect 11063 29303 11097 29337
rect 11223 29303 11257 29337
rect 11383 29303 11417 29337
rect 11543 29303 11577 29337
rect 11703 29303 11737 29337
rect 11863 29303 11897 29337
rect 12023 29303 12057 29337
rect 12183 29303 12217 29337
rect 12343 29303 12377 29337
rect 8503 29143 8537 29177
rect 8663 29143 8697 29177
rect 8823 29143 8857 29177
rect 8983 29143 9017 29177
rect 9143 29143 9177 29177
rect 9303 29143 9337 29177
rect 9463 29143 9497 29177
rect 9623 29143 9657 29177
rect 9783 29143 9817 29177
rect 9943 29143 9977 29177
rect 10103 29143 10137 29177
rect 10263 29143 10297 29177
rect 10423 29143 10457 29177
rect 10583 29143 10617 29177
rect 10743 29143 10777 29177
rect 10903 29143 10937 29177
rect 11063 29143 11097 29177
rect 11223 29143 11257 29177
rect 11383 29143 11417 29177
rect 11543 29143 11577 29177
rect 11703 29143 11737 29177
rect 11863 29143 11897 29177
rect 12023 29143 12057 29177
rect 12183 29143 12217 29177
rect 12343 29143 12377 29177
rect 8503 28983 8537 29017
rect 8663 28983 8697 29017
rect 8823 28983 8857 29017
rect 8983 28983 9017 29017
rect 9143 28983 9177 29017
rect 9303 28983 9337 29017
rect 9463 28983 9497 29017
rect 9623 28983 9657 29017
rect 9783 28983 9817 29017
rect 9943 28983 9977 29017
rect 10103 28983 10137 29017
rect 10263 28983 10297 29017
rect 10423 28983 10457 29017
rect 10583 28983 10617 29017
rect 10743 28983 10777 29017
rect 10903 28983 10937 29017
rect 11063 28983 11097 29017
rect 11223 28983 11257 29017
rect 11383 28983 11417 29017
rect 11543 28983 11577 29017
rect 11703 28983 11737 29017
rect 11863 28983 11897 29017
rect 12023 28983 12057 29017
rect 12183 28983 12217 29017
rect 12343 28983 12377 29017
rect 8503 28823 8537 28857
rect 8663 28823 8697 28857
rect 8823 28823 8857 28857
rect 8983 28823 9017 28857
rect 9143 28823 9177 28857
rect 9303 28823 9337 28857
rect 9463 28823 9497 28857
rect 9623 28823 9657 28857
rect 9783 28823 9817 28857
rect 9943 28823 9977 28857
rect 10103 28823 10137 28857
rect 10263 28823 10297 28857
rect 10423 28823 10457 28857
rect 10583 28823 10617 28857
rect 10743 28823 10777 28857
rect 10903 28823 10937 28857
rect 11063 28823 11097 28857
rect 11223 28823 11257 28857
rect 11383 28823 11417 28857
rect 11543 28823 11577 28857
rect 11703 28823 11737 28857
rect 11863 28823 11897 28857
rect 12023 28823 12057 28857
rect 12183 28823 12217 28857
rect 12343 28823 12377 28857
rect 8503 28663 8537 28697
rect 8663 28663 8697 28697
rect 8823 28663 8857 28697
rect 8983 28663 9017 28697
rect 9143 28663 9177 28697
rect 9303 28663 9337 28697
rect 9463 28663 9497 28697
rect 9623 28663 9657 28697
rect 9783 28663 9817 28697
rect 9943 28663 9977 28697
rect 10103 28663 10137 28697
rect 10263 28663 10297 28697
rect 10423 28663 10457 28697
rect 10583 28663 10617 28697
rect 10743 28663 10777 28697
rect 10903 28663 10937 28697
rect 11063 28663 11097 28697
rect 11223 28663 11257 28697
rect 11383 28663 11417 28697
rect 11543 28663 11577 28697
rect 11703 28663 11737 28697
rect 11863 28663 11897 28697
rect 12023 28663 12057 28697
rect 12183 28663 12217 28697
rect 12343 28663 12377 28697
rect 8503 28503 8537 28537
rect 8663 28503 8697 28537
rect 8823 28503 8857 28537
rect 8983 28503 9017 28537
rect 9143 28503 9177 28537
rect 9303 28503 9337 28537
rect 9463 28503 9497 28537
rect 9623 28503 9657 28537
rect 9783 28503 9817 28537
rect 9943 28503 9977 28537
rect 10103 28503 10137 28537
rect 10263 28503 10297 28537
rect 10423 28503 10457 28537
rect 10583 28503 10617 28537
rect 10743 28503 10777 28537
rect 10903 28503 10937 28537
rect 11063 28503 11097 28537
rect 11223 28503 11257 28537
rect 11383 28503 11417 28537
rect 11543 28503 11577 28537
rect 11703 28503 11737 28537
rect 11863 28503 11897 28537
rect 12023 28503 12057 28537
rect 12183 28503 12217 28537
rect 12343 28503 12377 28537
rect 8503 28343 8537 28377
rect 8663 28343 8697 28377
rect 8823 28343 8857 28377
rect 8983 28343 9017 28377
rect 9143 28343 9177 28377
rect 9303 28343 9337 28377
rect 9463 28343 9497 28377
rect 9623 28343 9657 28377
rect 9783 28343 9817 28377
rect 9943 28343 9977 28377
rect 10103 28343 10137 28377
rect 10263 28343 10297 28377
rect 10423 28343 10457 28377
rect 10583 28343 10617 28377
rect 10743 28343 10777 28377
rect 10903 28343 10937 28377
rect 11063 28343 11097 28377
rect 11223 28343 11257 28377
rect 11383 28343 11417 28377
rect 11543 28343 11577 28377
rect 11703 28343 11737 28377
rect 11863 28343 11897 28377
rect 12023 28343 12057 28377
rect 12183 28343 12217 28377
rect 12343 28343 12377 28377
rect 8503 28183 8537 28217
rect 8663 28183 8697 28217
rect 8823 28183 8857 28217
rect 8983 28183 9017 28217
rect 9143 28183 9177 28217
rect 9303 28183 9337 28217
rect 9463 28183 9497 28217
rect 9623 28183 9657 28217
rect 9783 28183 9817 28217
rect 9943 28183 9977 28217
rect 10103 28183 10137 28217
rect 10263 28183 10297 28217
rect 10423 28183 10457 28217
rect 10583 28183 10617 28217
rect 10743 28183 10777 28217
rect 10903 28183 10937 28217
rect 11063 28183 11097 28217
rect 11223 28183 11257 28217
rect 11383 28183 11417 28217
rect 11543 28183 11577 28217
rect 11703 28183 11737 28217
rect 11863 28183 11897 28217
rect 12023 28183 12057 28217
rect 12183 28183 12217 28217
rect 12343 28183 12377 28217
rect 8503 28023 8537 28057
rect 8663 28023 8697 28057
rect 8823 28023 8857 28057
rect 8983 28023 9017 28057
rect 9143 28023 9177 28057
rect 9303 28023 9337 28057
rect 9463 28023 9497 28057
rect 9623 28023 9657 28057
rect 9783 28023 9817 28057
rect 9943 28023 9977 28057
rect 10103 28023 10137 28057
rect 10263 28023 10297 28057
rect 10423 28023 10457 28057
rect 10583 28023 10617 28057
rect 10743 28023 10777 28057
rect 10903 28023 10937 28057
rect 11063 28023 11097 28057
rect 11223 28023 11257 28057
rect 11383 28023 11417 28057
rect 11543 28023 11577 28057
rect 11703 28023 11737 28057
rect 11863 28023 11897 28057
rect 12023 28023 12057 28057
rect 12183 28023 12217 28057
rect 12343 28023 12377 28057
rect 8503 27863 8537 27897
rect 8663 27863 8697 27897
rect 8823 27863 8857 27897
rect 8983 27863 9017 27897
rect 9143 27863 9177 27897
rect 9303 27863 9337 27897
rect 9463 27863 9497 27897
rect 9623 27863 9657 27897
rect 9783 27863 9817 27897
rect 9943 27863 9977 27897
rect 10103 27863 10137 27897
rect 10263 27863 10297 27897
rect 10423 27863 10457 27897
rect 10583 27863 10617 27897
rect 10743 27863 10777 27897
rect 10903 27863 10937 27897
rect 11063 27863 11097 27897
rect 11223 27863 11257 27897
rect 11383 27863 11417 27897
rect 11543 27863 11577 27897
rect 11703 27863 11737 27897
rect 11863 27863 11897 27897
rect 12023 27863 12057 27897
rect 12183 27863 12217 27897
rect 12343 27863 12377 27897
rect 8503 27703 8537 27737
rect 8663 27703 8697 27737
rect 8823 27703 8857 27737
rect 8983 27703 9017 27737
rect 9143 27703 9177 27737
rect 9303 27703 9337 27737
rect 9463 27703 9497 27737
rect 9623 27703 9657 27737
rect 9783 27703 9817 27737
rect 9943 27703 9977 27737
rect 10103 27703 10137 27737
rect 10263 27703 10297 27737
rect 10423 27703 10457 27737
rect 10583 27703 10617 27737
rect 10743 27703 10777 27737
rect 10903 27703 10937 27737
rect 11063 27703 11097 27737
rect 11223 27703 11257 27737
rect 11383 27703 11417 27737
rect 11543 27703 11577 27737
rect 11703 27703 11737 27737
rect 11863 27703 11897 27737
rect 12023 27703 12057 27737
rect 12183 27703 12217 27737
rect 12343 27703 12377 27737
rect 8503 27543 8537 27577
rect 8663 27543 8697 27577
rect 8823 27543 8857 27577
rect 8983 27543 9017 27577
rect 9143 27543 9177 27577
rect 9303 27543 9337 27577
rect 9463 27543 9497 27577
rect 9623 27543 9657 27577
rect 9783 27543 9817 27577
rect 9943 27543 9977 27577
rect 10103 27543 10137 27577
rect 10263 27543 10297 27577
rect 10423 27543 10457 27577
rect 10583 27543 10617 27577
rect 10743 27543 10777 27577
rect 10903 27543 10937 27577
rect 11063 27543 11097 27577
rect 11223 27543 11257 27577
rect 11383 27543 11417 27577
rect 11543 27543 11577 27577
rect 11703 27543 11737 27577
rect 11863 27543 11897 27577
rect 12023 27543 12057 27577
rect 12183 27543 12217 27577
rect 12343 27543 12377 27577
rect 8503 27383 8537 27417
rect 8663 27383 8697 27417
rect 8823 27383 8857 27417
rect 8983 27383 9017 27417
rect 9143 27383 9177 27417
rect 9303 27383 9337 27417
rect 9463 27383 9497 27417
rect 9623 27383 9657 27417
rect 9783 27383 9817 27417
rect 9943 27383 9977 27417
rect 10103 27383 10137 27417
rect 10263 27383 10297 27417
rect 10423 27383 10457 27417
rect 10583 27383 10617 27417
rect 10743 27383 10777 27417
rect 10903 27383 10937 27417
rect 11063 27383 11097 27417
rect 11223 27383 11257 27417
rect 11383 27383 11417 27417
rect 11543 27383 11577 27417
rect 11703 27383 11737 27417
rect 11863 27383 11897 27417
rect 12023 27383 12057 27417
rect 12183 27383 12217 27417
rect 12343 27383 12377 27417
rect 8503 27223 8537 27257
rect 8663 27223 8697 27257
rect 8823 27223 8857 27257
rect 8983 27223 9017 27257
rect 9143 27223 9177 27257
rect 9303 27223 9337 27257
rect 9463 27223 9497 27257
rect 9623 27223 9657 27257
rect 9783 27223 9817 27257
rect 9943 27223 9977 27257
rect 10103 27223 10137 27257
rect 10263 27223 10297 27257
rect 10423 27223 10457 27257
rect 10583 27223 10617 27257
rect 10743 27223 10777 27257
rect 10903 27223 10937 27257
rect 11063 27223 11097 27257
rect 11223 27223 11257 27257
rect 11383 27223 11417 27257
rect 11543 27223 11577 27257
rect 11703 27223 11737 27257
rect 11863 27223 11897 27257
rect 12023 27223 12057 27257
rect 12183 27223 12217 27257
rect 12343 27223 12377 27257
rect 8503 27063 8537 27097
rect 8663 27063 8697 27097
rect 8823 27063 8857 27097
rect 8983 27063 9017 27097
rect 9143 27063 9177 27097
rect 9303 27063 9337 27097
rect 9463 27063 9497 27097
rect 9623 27063 9657 27097
rect 9783 27063 9817 27097
rect 9943 27063 9977 27097
rect 10103 27063 10137 27097
rect 10263 27063 10297 27097
rect 10423 27063 10457 27097
rect 10583 27063 10617 27097
rect 10743 27063 10777 27097
rect 10903 27063 10937 27097
rect 11063 27063 11097 27097
rect 11223 27063 11257 27097
rect 11383 27063 11417 27097
rect 11543 27063 11577 27097
rect 11703 27063 11737 27097
rect 11863 27063 11897 27097
rect 12023 27063 12057 27097
rect 12183 27063 12217 27097
rect 12343 27063 12377 27097
rect 8503 26903 8537 26937
rect 8663 26903 8697 26937
rect 8823 26903 8857 26937
rect 8983 26903 9017 26937
rect 9143 26903 9177 26937
rect 9303 26903 9337 26937
rect 9463 26903 9497 26937
rect 9623 26903 9657 26937
rect 9783 26903 9817 26937
rect 9943 26903 9977 26937
rect 10103 26903 10137 26937
rect 10263 26903 10297 26937
rect 10423 26903 10457 26937
rect 10583 26903 10617 26937
rect 10743 26903 10777 26937
rect 10903 26903 10937 26937
rect 11063 26903 11097 26937
rect 11223 26903 11257 26937
rect 11383 26903 11417 26937
rect 11543 26903 11577 26937
rect 11703 26903 11737 26937
rect 11863 26903 11897 26937
rect 12023 26903 12057 26937
rect 12183 26903 12217 26937
rect 12343 26903 12377 26937
rect 8503 26743 8537 26777
rect 8663 26743 8697 26777
rect 8823 26743 8857 26777
rect 8983 26743 9017 26777
rect 9143 26743 9177 26777
rect 9303 26743 9337 26777
rect 9463 26743 9497 26777
rect 9623 26743 9657 26777
rect 9783 26743 9817 26777
rect 9943 26743 9977 26777
rect 10103 26743 10137 26777
rect 10263 26743 10297 26777
rect 10423 26743 10457 26777
rect 10583 26743 10617 26777
rect 10743 26743 10777 26777
rect 10903 26743 10937 26777
rect 11063 26743 11097 26777
rect 11223 26743 11257 26777
rect 11383 26743 11417 26777
rect 11543 26743 11577 26777
rect 11703 26743 11737 26777
rect 11863 26743 11897 26777
rect 12023 26743 12057 26777
rect 12183 26743 12217 26777
rect 12343 26743 12377 26777
rect 8503 26583 8537 26617
rect 8663 26583 8697 26617
rect 8823 26583 8857 26617
rect 8983 26583 9017 26617
rect 9143 26583 9177 26617
rect 9303 26583 9337 26617
rect 9463 26583 9497 26617
rect 9623 26583 9657 26617
rect 9783 26583 9817 26617
rect 9943 26583 9977 26617
rect 10103 26583 10137 26617
rect 10263 26583 10297 26617
rect 10423 26583 10457 26617
rect 10583 26583 10617 26617
rect 10743 26583 10777 26617
rect 10903 26583 10937 26617
rect 11063 26583 11097 26617
rect 11223 26583 11257 26617
rect 11383 26583 11417 26617
rect 11543 26583 11577 26617
rect 11703 26583 11737 26617
rect 11863 26583 11897 26617
rect 12023 26583 12057 26617
rect 12183 26583 12217 26617
rect 12343 26583 12377 26617
rect 8503 26423 8537 26457
rect 8663 26423 8697 26457
rect 8823 26423 8857 26457
rect 8983 26423 9017 26457
rect 9143 26423 9177 26457
rect 9303 26423 9337 26457
rect 9463 26423 9497 26457
rect 9623 26423 9657 26457
rect 9783 26423 9817 26457
rect 9943 26423 9977 26457
rect 10103 26423 10137 26457
rect 10263 26423 10297 26457
rect 10423 26423 10457 26457
rect 10583 26423 10617 26457
rect 10743 26423 10777 26457
rect 10903 26423 10937 26457
rect 11063 26423 11097 26457
rect 11223 26423 11257 26457
rect 11383 26423 11417 26457
rect 11543 26423 11577 26457
rect 11703 26423 11737 26457
rect 11863 26423 11897 26457
rect 12023 26423 12057 26457
rect 12183 26423 12217 26457
rect 12343 26423 12377 26457
rect 8503 26263 8537 26297
rect 8663 26263 8697 26297
rect 8823 26263 8857 26297
rect 8983 26263 9017 26297
rect 9143 26263 9177 26297
rect 9303 26263 9337 26297
rect 9463 26263 9497 26297
rect 9623 26263 9657 26297
rect 9783 26263 9817 26297
rect 9943 26263 9977 26297
rect 10103 26263 10137 26297
rect 10263 26263 10297 26297
rect 10423 26263 10457 26297
rect 10583 26263 10617 26297
rect 10743 26263 10777 26297
rect 10903 26263 10937 26297
rect 11063 26263 11097 26297
rect 11223 26263 11257 26297
rect 11383 26263 11417 26297
rect 11543 26263 11577 26297
rect 11703 26263 11737 26297
rect 11863 26263 11897 26297
rect 12023 26263 12057 26297
rect 12183 26263 12217 26297
rect 12343 26263 12377 26297
rect 8503 26103 8537 26137
rect 8663 26103 8697 26137
rect 8823 26103 8857 26137
rect 8983 26103 9017 26137
rect 9143 26103 9177 26137
rect 9303 26103 9337 26137
rect 9463 26103 9497 26137
rect 9623 26103 9657 26137
rect 9783 26103 9817 26137
rect 9943 26103 9977 26137
rect 10103 26103 10137 26137
rect 10263 26103 10297 26137
rect 10423 26103 10457 26137
rect 10583 26103 10617 26137
rect 10743 26103 10777 26137
rect 10903 26103 10937 26137
rect 11063 26103 11097 26137
rect 11223 26103 11257 26137
rect 11383 26103 11417 26137
rect 11543 26103 11577 26137
rect 11703 26103 11737 26137
rect 11863 26103 11897 26137
rect 12023 26103 12057 26137
rect 12183 26103 12217 26137
rect 12343 26103 12377 26137
rect 8503 25943 8537 25977
rect 8663 25943 8697 25977
rect 8823 25943 8857 25977
rect 8983 25943 9017 25977
rect 9143 25943 9177 25977
rect 9303 25943 9337 25977
rect 9463 25943 9497 25977
rect 9623 25943 9657 25977
rect 9783 25943 9817 25977
rect 9943 25943 9977 25977
rect 10103 25943 10137 25977
rect 10263 25943 10297 25977
rect 10423 25943 10457 25977
rect 10583 25943 10617 25977
rect 10743 25943 10777 25977
rect 10903 25943 10937 25977
rect 11063 25943 11097 25977
rect 11223 25943 11257 25977
rect 11383 25943 11417 25977
rect 11543 25943 11577 25977
rect 11703 25943 11737 25977
rect 11863 25943 11897 25977
rect 12023 25943 12057 25977
rect 12183 25943 12217 25977
rect 12343 25943 12377 25977
rect 8503 25783 8537 25817
rect 8663 25783 8697 25817
rect 8823 25783 8857 25817
rect 8983 25783 9017 25817
rect 9143 25783 9177 25817
rect 9303 25783 9337 25817
rect 9463 25783 9497 25817
rect 9623 25783 9657 25817
rect 9783 25783 9817 25817
rect 9943 25783 9977 25817
rect 10103 25783 10137 25817
rect 10263 25783 10297 25817
rect 10423 25783 10457 25817
rect 10583 25783 10617 25817
rect 10743 25783 10777 25817
rect 10903 25783 10937 25817
rect 11063 25783 11097 25817
rect 11223 25783 11257 25817
rect 11383 25783 11417 25817
rect 11543 25783 11577 25817
rect 11703 25783 11737 25817
rect 11863 25783 11897 25817
rect 12023 25783 12057 25817
rect 12183 25783 12217 25817
rect 12343 25783 12377 25817
rect 8503 25623 8537 25657
rect 8663 25623 8697 25657
rect 8823 25623 8857 25657
rect 8983 25623 9017 25657
rect 9143 25623 9177 25657
rect 9303 25623 9337 25657
rect 9463 25623 9497 25657
rect 9623 25623 9657 25657
rect 9783 25623 9817 25657
rect 9943 25623 9977 25657
rect 10103 25623 10137 25657
rect 10263 25623 10297 25657
rect 10423 25623 10457 25657
rect 10583 25623 10617 25657
rect 10743 25623 10777 25657
rect 10903 25623 10937 25657
rect 11063 25623 11097 25657
rect 11223 25623 11257 25657
rect 11383 25623 11417 25657
rect 11543 25623 11577 25657
rect 11703 25623 11737 25657
rect 11863 25623 11897 25657
rect 12023 25623 12057 25657
rect 12183 25623 12217 25657
rect 12343 25623 12377 25657
rect 8503 25463 8537 25497
rect 8663 25463 8697 25497
rect 8823 25463 8857 25497
rect 8983 25463 9017 25497
rect 9143 25463 9177 25497
rect 9303 25463 9337 25497
rect 9463 25463 9497 25497
rect 9623 25463 9657 25497
rect 9783 25463 9817 25497
rect 9943 25463 9977 25497
rect 10103 25463 10137 25497
rect 10263 25463 10297 25497
rect 10423 25463 10457 25497
rect 10583 25463 10617 25497
rect 10743 25463 10777 25497
rect 10903 25463 10937 25497
rect 11063 25463 11097 25497
rect 11223 25463 11257 25497
rect 11383 25463 11417 25497
rect 11543 25463 11577 25497
rect 11703 25463 11737 25497
rect 11863 25463 11897 25497
rect 12023 25463 12057 25497
rect 12183 25463 12217 25497
rect 12343 25463 12377 25497
rect 8503 25303 8537 25337
rect 8663 25303 8697 25337
rect 8823 25303 8857 25337
rect 8983 25303 9017 25337
rect 9143 25303 9177 25337
rect 9303 25303 9337 25337
rect 9463 25303 9497 25337
rect 9623 25303 9657 25337
rect 9783 25303 9817 25337
rect 9943 25303 9977 25337
rect 10103 25303 10137 25337
rect 10263 25303 10297 25337
rect 10423 25303 10457 25337
rect 10583 25303 10617 25337
rect 10743 25303 10777 25337
rect 10903 25303 10937 25337
rect 11063 25303 11097 25337
rect 11223 25303 11257 25337
rect 11383 25303 11417 25337
rect 11543 25303 11577 25337
rect 11703 25303 11737 25337
rect 11863 25303 11897 25337
rect 12023 25303 12057 25337
rect 12183 25303 12217 25337
rect 12343 25303 12377 25337
rect 8503 25143 8537 25177
rect 8663 25143 8697 25177
rect 8823 25143 8857 25177
rect 8983 25143 9017 25177
rect 9143 25143 9177 25177
rect 9303 25143 9337 25177
rect 9463 25143 9497 25177
rect 9623 25143 9657 25177
rect 9783 25143 9817 25177
rect 9943 25143 9977 25177
rect 10103 25143 10137 25177
rect 10263 25143 10297 25177
rect 10423 25143 10457 25177
rect 10583 25143 10617 25177
rect 10743 25143 10777 25177
rect 10903 25143 10937 25177
rect 11063 25143 11097 25177
rect 11223 25143 11257 25177
rect 11383 25143 11417 25177
rect 11543 25143 11577 25177
rect 11703 25143 11737 25177
rect 11863 25143 11897 25177
rect 12023 25143 12057 25177
rect 12183 25143 12217 25177
rect 12343 25143 12377 25177
rect 8503 24983 8537 25017
rect 8663 24983 8697 25017
rect 8823 24983 8857 25017
rect 8983 24983 9017 25017
rect 9143 24983 9177 25017
rect 9303 24983 9337 25017
rect 9463 24983 9497 25017
rect 9623 24983 9657 25017
rect 9783 24983 9817 25017
rect 9943 24983 9977 25017
rect 10103 24983 10137 25017
rect 10263 24983 10297 25017
rect 10423 24983 10457 25017
rect 10583 24983 10617 25017
rect 10743 24983 10777 25017
rect 10903 24983 10937 25017
rect 11063 24983 11097 25017
rect 11223 24983 11257 25017
rect 11383 24983 11417 25017
rect 11543 24983 11577 25017
rect 11703 24983 11737 25017
rect 11863 24983 11897 25017
rect 12023 24983 12057 25017
rect 12183 24983 12217 25017
rect 12343 24983 12377 25017
rect 8503 24823 8537 24857
rect 8663 24823 8697 24857
rect 8823 24823 8857 24857
rect 8983 24823 9017 24857
rect 9143 24823 9177 24857
rect 9303 24823 9337 24857
rect 9463 24823 9497 24857
rect 9623 24823 9657 24857
rect 9783 24823 9817 24857
rect 9943 24823 9977 24857
rect 10103 24823 10137 24857
rect 10263 24823 10297 24857
rect 10423 24823 10457 24857
rect 10583 24823 10617 24857
rect 10743 24823 10777 24857
rect 10903 24823 10937 24857
rect 11063 24823 11097 24857
rect 11223 24823 11257 24857
rect 11383 24823 11417 24857
rect 11543 24823 11577 24857
rect 11703 24823 11737 24857
rect 11863 24823 11897 24857
rect 12023 24823 12057 24857
rect 12183 24823 12217 24857
rect 12343 24823 12377 24857
rect 8503 24663 8537 24697
rect 8663 24663 8697 24697
rect 8823 24663 8857 24697
rect 8983 24663 9017 24697
rect 9143 24663 9177 24697
rect 9303 24663 9337 24697
rect 9463 24663 9497 24697
rect 9623 24663 9657 24697
rect 9783 24663 9817 24697
rect 9943 24663 9977 24697
rect 10103 24663 10137 24697
rect 10263 24663 10297 24697
rect 10423 24663 10457 24697
rect 10583 24663 10617 24697
rect 10743 24663 10777 24697
rect 10903 24663 10937 24697
rect 11063 24663 11097 24697
rect 11223 24663 11257 24697
rect 11383 24663 11417 24697
rect 11543 24663 11577 24697
rect 11703 24663 11737 24697
rect 11863 24663 11897 24697
rect 12023 24663 12057 24697
rect 12183 24663 12217 24697
rect 12343 24663 12377 24697
rect 8503 24503 8537 24537
rect 8663 24503 8697 24537
rect 8823 24503 8857 24537
rect 8983 24503 9017 24537
rect 9143 24503 9177 24537
rect 9303 24503 9337 24537
rect 9463 24503 9497 24537
rect 9623 24503 9657 24537
rect 9783 24503 9817 24537
rect 9943 24503 9977 24537
rect 10103 24503 10137 24537
rect 10263 24503 10297 24537
rect 10423 24503 10457 24537
rect 10583 24503 10617 24537
rect 10743 24503 10777 24537
rect 10903 24503 10937 24537
rect 11063 24503 11097 24537
rect 11223 24503 11257 24537
rect 11383 24503 11417 24537
rect 11543 24503 11577 24537
rect 11703 24503 11737 24537
rect 11863 24503 11897 24537
rect 12023 24503 12057 24537
rect 12183 24503 12217 24537
rect 12343 24503 12377 24537
rect 8503 24343 8537 24377
rect 8663 24343 8697 24377
rect 8823 24343 8857 24377
rect 8983 24343 9017 24377
rect 9143 24343 9177 24377
rect 9303 24343 9337 24377
rect 9463 24343 9497 24377
rect 9623 24343 9657 24377
rect 9783 24343 9817 24377
rect 9943 24343 9977 24377
rect 10103 24343 10137 24377
rect 10263 24343 10297 24377
rect 10423 24343 10457 24377
rect 10583 24343 10617 24377
rect 10743 24343 10777 24377
rect 10903 24343 10937 24377
rect 11063 24343 11097 24377
rect 11223 24343 11257 24377
rect 11383 24343 11417 24377
rect 11543 24343 11577 24377
rect 11703 24343 11737 24377
rect 11863 24343 11897 24377
rect 12023 24343 12057 24377
rect 12183 24343 12217 24377
rect 12343 24343 12377 24377
rect 8503 24183 8537 24217
rect 8663 24183 8697 24217
rect 8823 24183 8857 24217
rect 8983 24183 9017 24217
rect 9143 24183 9177 24217
rect 9303 24183 9337 24217
rect 9463 24183 9497 24217
rect 9623 24183 9657 24217
rect 9783 24183 9817 24217
rect 9943 24183 9977 24217
rect 10103 24183 10137 24217
rect 10263 24183 10297 24217
rect 10423 24183 10457 24217
rect 10583 24183 10617 24217
rect 10743 24183 10777 24217
rect 10903 24183 10937 24217
rect 11063 24183 11097 24217
rect 11223 24183 11257 24217
rect 11383 24183 11417 24217
rect 11543 24183 11577 24217
rect 11703 24183 11737 24217
rect 11863 24183 11897 24217
rect 12023 24183 12057 24217
rect 12183 24183 12217 24217
rect 12343 24183 12377 24217
rect 8503 24023 8537 24057
rect 8663 24023 8697 24057
rect 8823 24023 8857 24057
rect 8983 24023 9017 24057
rect 9143 24023 9177 24057
rect 9303 24023 9337 24057
rect 9463 24023 9497 24057
rect 9623 24023 9657 24057
rect 9783 24023 9817 24057
rect 9943 24023 9977 24057
rect 10103 24023 10137 24057
rect 10263 24023 10297 24057
rect 10423 24023 10457 24057
rect 10583 24023 10617 24057
rect 10743 24023 10777 24057
rect 10903 24023 10937 24057
rect 11063 24023 11097 24057
rect 11223 24023 11257 24057
rect 11383 24023 11417 24057
rect 11543 24023 11577 24057
rect 11703 24023 11737 24057
rect 11863 24023 11897 24057
rect 12023 24023 12057 24057
rect 12183 24023 12217 24057
rect 12343 24023 12377 24057
rect 8503 23863 8537 23897
rect 8663 23863 8697 23897
rect 8823 23863 8857 23897
rect 8983 23863 9017 23897
rect 9143 23863 9177 23897
rect 9303 23863 9337 23897
rect 9463 23863 9497 23897
rect 9623 23863 9657 23897
rect 9783 23863 9817 23897
rect 9943 23863 9977 23897
rect 10103 23863 10137 23897
rect 10263 23863 10297 23897
rect 10423 23863 10457 23897
rect 10583 23863 10617 23897
rect 10743 23863 10777 23897
rect 10903 23863 10937 23897
rect 11063 23863 11097 23897
rect 11223 23863 11257 23897
rect 11383 23863 11417 23897
rect 11543 23863 11577 23897
rect 11703 23863 11737 23897
rect 11863 23863 11897 23897
rect 12023 23863 12057 23897
rect 12183 23863 12217 23897
rect 12343 23863 12377 23897
rect 8503 23703 8537 23737
rect 8663 23703 8697 23737
rect 8823 23703 8857 23737
rect 8983 23703 9017 23737
rect 9143 23703 9177 23737
rect 9303 23703 9337 23737
rect 9463 23703 9497 23737
rect 9623 23703 9657 23737
rect 9783 23703 9817 23737
rect 9943 23703 9977 23737
rect 10103 23703 10137 23737
rect 10263 23703 10297 23737
rect 10423 23703 10457 23737
rect 10583 23703 10617 23737
rect 10743 23703 10777 23737
rect 10903 23703 10937 23737
rect 11063 23703 11097 23737
rect 11223 23703 11257 23737
rect 11383 23703 11417 23737
rect 11543 23703 11577 23737
rect 11703 23703 11737 23737
rect 11863 23703 11897 23737
rect 12023 23703 12057 23737
rect 12183 23703 12217 23737
rect 12343 23703 12377 23737
rect 8503 23543 8537 23577
rect 8663 23543 8697 23577
rect 8823 23543 8857 23577
rect 8983 23543 9017 23577
rect 9143 23543 9177 23577
rect 9303 23543 9337 23577
rect 9463 23543 9497 23577
rect 9623 23543 9657 23577
rect 9783 23543 9817 23577
rect 9943 23543 9977 23577
rect 10103 23543 10137 23577
rect 10263 23543 10297 23577
rect 10423 23543 10457 23577
rect 10583 23543 10617 23577
rect 10743 23543 10777 23577
rect 10903 23543 10937 23577
rect 11063 23543 11097 23577
rect 11223 23543 11257 23577
rect 11383 23543 11417 23577
rect 11543 23543 11577 23577
rect 11703 23543 11737 23577
rect 11863 23543 11897 23577
rect 12023 23543 12057 23577
rect 12183 23543 12217 23577
rect 12343 23543 12377 23577
rect 8503 23383 8537 23417
rect 8663 23383 8697 23417
rect 8823 23383 8857 23417
rect 8983 23383 9017 23417
rect 9143 23383 9177 23417
rect 9303 23383 9337 23417
rect 9463 23383 9497 23417
rect 9623 23383 9657 23417
rect 9783 23383 9817 23417
rect 9943 23383 9977 23417
rect 10103 23383 10137 23417
rect 10263 23383 10297 23417
rect 10423 23383 10457 23417
rect 10583 23383 10617 23417
rect 10743 23383 10777 23417
rect 10903 23383 10937 23417
rect 11063 23383 11097 23417
rect 11223 23383 11257 23417
rect 11383 23383 11417 23417
rect 11543 23383 11577 23417
rect 11703 23383 11737 23417
rect 11863 23383 11897 23417
rect 12023 23383 12057 23417
rect 12183 23383 12217 23417
rect 12343 23383 12377 23417
rect 8503 23223 8537 23257
rect 8663 23223 8697 23257
rect 8823 23223 8857 23257
rect 8983 23223 9017 23257
rect 9143 23223 9177 23257
rect 9303 23223 9337 23257
rect 9463 23223 9497 23257
rect 9623 23223 9657 23257
rect 9783 23223 9817 23257
rect 9943 23223 9977 23257
rect 10103 23223 10137 23257
rect 10263 23223 10297 23257
rect 10423 23223 10457 23257
rect 10583 23223 10617 23257
rect 10743 23223 10777 23257
rect 10903 23223 10937 23257
rect 11063 23223 11097 23257
rect 11223 23223 11257 23257
rect 11383 23223 11417 23257
rect 11543 23223 11577 23257
rect 11703 23223 11737 23257
rect 11863 23223 11897 23257
rect 12023 23223 12057 23257
rect 12183 23223 12217 23257
rect 12343 23223 12377 23257
rect 8503 23063 8537 23097
rect 8663 23063 8697 23097
rect 8823 23063 8857 23097
rect 8983 23063 9017 23097
rect 9143 23063 9177 23097
rect 9303 23063 9337 23097
rect 9463 23063 9497 23097
rect 9623 23063 9657 23097
rect 9783 23063 9817 23097
rect 9943 23063 9977 23097
rect 10103 23063 10137 23097
rect 10263 23063 10297 23097
rect 10423 23063 10457 23097
rect 10583 23063 10617 23097
rect 10743 23063 10777 23097
rect 10903 23063 10937 23097
rect 11063 23063 11097 23097
rect 11223 23063 11257 23097
rect 11383 23063 11417 23097
rect 11543 23063 11577 23097
rect 11703 23063 11737 23097
rect 11863 23063 11897 23097
rect 12023 23063 12057 23097
rect 12183 23063 12217 23097
rect 12343 23063 12377 23097
rect 8503 22903 8537 22937
rect 8663 22903 8697 22937
rect 8823 22903 8857 22937
rect 8983 22903 9017 22937
rect 9143 22903 9177 22937
rect 9303 22903 9337 22937
rect 9463 22903 9497 22937
rect 9623 22903 9657 22937
rect 9783 22903 9817 22937
rect 9943 22903 9977 22937
rect 10103 22903 10137 22937
rect 10263 22903 10297 22937
rect 10423 22903 10457 22937
rect 10583 22903 10617 22937
rect 10743 22903 10777 22937
rect 10903 22903 10937 22937
rect 11063 22903 11097 22937
rect 11223 22903 11257 22937
rect 11383 22903 11417 22937
rect 11543 22903 11577 22937
rect 11703 22903 11737 22937
rect 11863 22903 11897 22937
rect 12023 22903 12057 22937
rect 12183 22903 12217 22937
rect 12343 22903 12377 22937
rect 8503 22743 8537 22777
rect 8663 22743 8697 22777
rect 8823 22743 8857 22777
rect 8983 22743 9017 22777
rect 9143 22743 9177 22777
rect 9303 22743 9337 22777
rect 9463 22743 9497 22777
rect 9623 22743 9657 22777
rect 9783 22743 9817 22777
rect 9943 22743 9977 22777
rect 10103 22743 10137 22777
rect 10263 22743 10297 22777
rect 10423 22743 10457 22777
rect 10583 22743 10617 22777
rect 10743 22743 10777 22777
rect 10903 22743 10937 22777
rect 11063 22743 11097 22777
rect 11223 22743 11257 22777
rect 11383 22743 11417 22777
rect 11543 22743 11577 22777
rect 11703 22743 11737 22777
rect 11863 22743 11897 22777
rect 12023 22743 12057 22777
rect 12183 22743 12217 22777
rect 12343 22743 12377 22777
rect 8503 22583 8537 22617
rect 8663 22583 8697 22617
rect 8823 22583 8857 22617
rect 8983 22583 9017 22617
rect 9143 22583 9177 22617
rect 9303 22583 9337 22617
rect 9463 22583 9497 22617
rect 9623 22583 9657 22617
rect 9783 22583 9817 22617
rect 9943 22583 9977 22617
rect 10103 22583 10137 22617
rect 10263 22583 10297 22617
rect 10423 22583 10457 22617
rect 10583 22583 10617 22617
rect 10743 22583 10777 22617
rect 10903 22583 10937 22617
rect 11063 22583 11097 22617
rect 11223 22583 11257 22617
rect 11383 22583 11417 22617
rect 11543 22583 11577 22617
rect 11703 22583 11737 22617
rect 11863 22583 11897 22617
rect 12023 22583 12057 22617
rect 12183 22583 12217 22617
rect 12343 22583 12377 22617
rect 8503 22423 8537 22457
rect 8663 22423 8697 22457
rect 8823 22423 8857 22457
rect 8983 22423 9017 22457
rect 9143 22423 9177 22457
rect 9303 22423 9337 22457
rect 9463 22423 9497 22457
rect 9623 22423 9657 22457
rect 9783 22423 9817 22457
rect 9943 22423 9977 22457
rect 10103 22423 10137 22457
rect 10263 22423 10297 22457
rect 10423 22423 10457 22457
rect 10583 22423 10617 22457
rect 10743 22423 10777 22457
rect 10903 22423 10937 22457
rect 11063 22423 11097 22457
rect 11223 22423 11257 22457
rect 11383 22423 11417 22457
rect 11543 22423 11577 22457
rect 11703 22423 11737 22457
rect 11863 22423 11897 22457
rect 12023 22423 12057 22457
rect 12183 22423 12217 22457
rect 12343 22423 12377 22457
rect 8503 22263 8537 22297
rect 8663 22263 8697 22297
rect 8823 22263 8857 22297
rect 8983 22263 9017 22297
rect 9143 22263 9177 22297
rect 9303 22263 9337 22297
rect 9463 22263 9497 22297
rect 9623 22263 9657 22297
rect 9783 22263 9817 22297
rect 9943 22263 9977 22297
rect 10103 22263 10137 22297
rect 10263 22263 10297 22297
rect 10423 22263 10457 22297
rect 10583 22263 10617 22297
rect 10743 22263 10777 22297
rect 10903 22263 10937 22297
rect 11063 22263 11097 22297
rect 11223 22263 11257 22297
rect 11383 22263 11417 22297
rect 11543 22263 11577 22297
rect 11703 22263 11737 22297
rect 11863 22263 11897 22297
rect 12023 22263 12057 22297
rect 12183 22263 12217 22297
rect 12343 22263 12377 22297
rect 8503 22103 8537 22137
rect 8663 22103 8697 22137
rect 8823 22103 8857 22137
rect 8983 22103 9017 22137
rect 9143 22103 9177 22137
rect 9303 22103 9337 22137
rect 9463 22103 9497 22137
rect 9623 22103 9657 22137
rect 9783 22103 9817 22137
rect 9943 22103 9977 22137
rect 10103 22103 10137 22137
rect 10263 22103 10297 22137
rect 10423 22103 10457 22137
rect 10583 22103 10617 22137
rect 10743 22103 10777 22137
rect 10903 22103 10937 22137
rect 11063 22103 11097 22137
rect 11223 22103 11257 22137
rect 11383 22103 11417 22137
rect 11543 22103 11577 22137
rect 11703 22103 11737 22137
rect 11863 22103 11897 22137
rect 12023 22103 12057 22137
rect 12183 22103 12217 22137
rect 12343 22103 12377 22137
rect 8503 21943 8537 21977
rect 8663 21943 8697 21977
rect 8823 21943 8857 21977
rect 8983 21943 9017 21977
rect 9143 21943 9177 21977
rect 9303 21943 9337 21977
rect 9463 21943 9497 21977
rect 9623 21943 9657 21977
rect 9783 21943 9817 21977
rect 9943 21943 9977 21977
rect 10103 21943 10137 21977
rect 10263 21943 10297 21977
rect 10423 21943 10457 21977
rect 10583 21943 10617 21977
rect 10743 21943 10777 21977
rect 10903 21943 10937 21977
rect 11063 21943 11097 21977
rect 11223 21943 11257 21977
rect 11383 21943 11417 21977
rect 11543 21943 11577 21977
rect 11703 21943 11737 21977
rect 11863 21943 11897 21977
rect 12023 21943 12057 21977
rect 12183 21943 12217 21977
rect 12343 21943 12377 21977
rect 8503 21783 8537 21817
rect 8663 21783 8697 21817
rect 8823 21783 8857 21817
rect 8983 21783 9017 21817
rect 9143 21783 9177 21817
rect 9303 21783 9337 21817
rect 9463 21783 9497 21817
rect 9623 21783 9657 21817
rect 9783 21783 9817 21817
rect 9943 21783 9977 21817
rect 10103 21783 10137 21817
rect 10263 21783 10297 21817
rect 10423 21783 10457 21817
rect 10583 21783 10617 21817
rect 10743 21783 10777 21817
rect 10903 21783 10937 21817
rect 11063 21783 11097 21817
rect 11223 21783 11257 21817
rect 11383 21783 11417 21817
rect 11543 21783 11577 21817
rect 11703 21783 11737 21817
rect 11863 21783 11897 21817
rect 12023 21783 12057 21817
rect 12183 21783 12217 21817
rect 12343 21783 12377 21817
rect 8503 21623 8537 21657
rect 8663 21623 8697 21657
rect 8823 21623 8857 21657
rect 8983 21623 9017 21657
rect 9143 21623 9177 21657
rect 9303 21623 9337 21657
rect 9463 21623 9497 21657
rect 9623 21623 9657 21657
rect 9783 21623 9817 21657
rect 9943 21623 9977 21657
rect 10103 21623 10137 21657
rect 10263 21623 10297 21657
rect 10423 21623 10457 21657
rect 10583 21623 10617 21657
rect 10743 21623 10777 21657
rect 10903 21623 10937 21657
rect 11063 21623 11097 21657
rect 11223 21623 11257 21657
rect 11383 21623 11417 21657
rect 11543 21623 11577 21657
rect 11703 21623 11737 21657
rect 11863 21623 11897 21657
rect 12023 21623 12057 21657
rect 12183 21623 12217 21657
rect 12343 21623 12377 21657
rect 8503 21463 8537 21497
rect 8663 21463 8697 21497
rect 8823 21463 8857 21497
rect 8983 21463 9017 21497
rect 9143 21463 9177 21497
rect 9303 21463 9337 21497
rect 9463 21463 9497 21497
rect 9623 21463 9657 21497
rect 9783 21463 9817 21497
rect 9943 21463 9977 21497
rect 10103 21463 10137 21497
rect 10263 21463 10297 21497
rect 10423 21463 10457 21497
rect 10583 21463 10617 21497
rect 10743 21463 10777 21497
rect 10903 21463 10937 21497
rect 11063 21463 11097 21497
rect 11223 21463 11257 21497
rect 11383 21463 11417 21497
rect 11543 21463 11577 21497
rect 11703 21463 11737 21497
rect 11863 21463 11897 21497
rect 12023 21463 12057 21497
rect 12183 21463 12217 21497
rect 12343 21463 12377 21497
rect 8503 21303 8537 21337
rect 8663 21303 8697 21337
rect 8823 21303 8857 21337
rect 8983 21303 9017 21337
rect 9143 21303 9177 21337
rect 9303 21303 9337 21337
rect 9463 21303 9497 21337
rect 9623 21303 9657 21337
rect 9783 21303 9817 21337
rect 9943 21303 9977 21337
rect 10103 21303 10137 21337
rect 10263 21303 10297 21337
rect 10423 21303 10457 21337
rect 10583 21303 10617 21337
rect 10743 21303 10777 21337
rect 10903 21303 10937 21337
rect 11063 21303 11097 21337
rect 11223 21303 11257 21337
rect 11383 21303 11417 21337
rect 11543 21303 11577 21337
rect 11703 21303 11737 21337
rect 11863 21303 11897 21337
rect 12023 21303 12057 21337
rect 12183 21303 12217 21337
rect 12343 21303 12377 21337
rect 8503 21143 8537 21177
rect 8663 21143 8697 21177
rect 8823 21143 8857 21177
rect 8983 21143 9017 21177
rect 9143 21143 9177 21177
rect 9303 21143 9337 21177
rect 9463 21143 9497 21177
rect 9623 21143 9657 21177
rect 9783 21143 9817 21177
rect 9943 21143 9977 21177
rect 10103 21143 10137 21177
rect 10263 21143 10297 21177
rect 10423 21143 10457 21177
rect 10583 21143 10617 21177
rect 10743 21143 10777 21177
rect 10903 21143 10937 21177
rect 11063 21143 11097 21177
rect 11223 21143 11257 21177
rect 11383 21143 11417 21177
rect 11543 21143 11577 21177
rect 11703 21143 11737 21177
rect 11863 21143 11897 21177
rect 12023 21143 12057 21177
rect 12183 21143 12217 21177
rect 12343 21143 12377 21177
rect 8503 20983 8537 21017
rect 8663 20983 8697 21017
rect 8823 20983 8857 21017
rect 8983 20983 9017 21017
rect 9143 20983 9177 21017
rect 9303 20983 9337 21017
rect 9463 20983 9497 21017
rect 9623 20983 9657 21017
rect 9783 20983 9817 21017
rect 9943 20983 9977 21017
rect 10103 20983 10137 21017
rect 10263 20983 10297 21017
rect 10423 20983 10457 21017
rect 10583 20983 10617 21017
rect 10743 20983 10777 21017
rect 10903 20983 10937 21017
rect 11063 20983 11097 21017
rect 11223 20983 11257 21017
rect 11383 20983 11417 21017
rect 11543 20983 11577 21017
rect 11703 20983 11737 21017
rect 11863 20983 11897 21017
rect 12023 20983 12057 21017
rect 12183 20983 12217 21017
rect 12343 20983 12377 21017
rect 8503 20823 8537 20857
rect 8663 20823 8697 20857
rect 8823 20823 8857 20857
rect 8983 20823 9017 20857
rect 9143 20823 9177 20857
rect 9303 20823 9337 20857
rect 9463 20823 9497 20857
rect 9623 20823 9657 20857
rect 9783 20823 9817 20857
rect 9943 20823 9977 20857
rect 10103 20823 10137 20857
rect 10263 20823 10297 20857
rect 10423 20823 10457 20857
rect 10583 20823 10617 20857
rect 10743 20823 10777 20857
rect 10903 20823 10937 20857
rect 11063 20823 11097 20857
rect 11223 20823 11257 20857
rect 11383 20823 11417 20857
rect 11543 20823 11577 20857
rect 11703 20823 11737 20857
rect 11863 20823 11897 20857
rect 12023 20823 12057 20857
rect 12183 20823 12217 20857
rect 12343 20823 12377 20857
rect 8503 20663 8537 20697
rect 8663 20663 8697 20697
rect 8823 20663 8857 20697
rect 8983 20663 9017 20697
rect 9143 20663 9177 20697
rect 9303 20663 9337 20697
rect 9463 20663 9497 20697
rect 9623 20663 9657 20697
rect 9783 20663 9817 20697
rect 9943 20663 9977 20697
rect 10103 20663 10137 20697
rect 10263 20663 10297 20697
rect 10423 20663 10457 20697
rect 10583 20663 10617 20697
rect 10743 20663 10777 20697
rect 10903 20663 10937 20697
rect 11063 20663 11097 20697
rect 11223 20663 11257 20697
rect 11383 20663 11417 20697
rect 11543 20663 11577 20697
rect 11703 20663 11737 20697
rect 11863 20663 11897 20697
rect 12023 20663 12057 20697
rect 12183 20663 12217 20697
rect 12343 20663 12377 20697
rect 8503 20503 8537 20537
rect 8663 20503 8697 20537
rect 8823 20503 8857 20537
rect 8983 20503 9017 20537
rect 9143 20503 9177 20537
rect 9303 20503 9337 20537
rect 9463 20503 9497 20537
rect 9623 20503 9657 20537
rect 9783 20503 9817 20537
rect 9943 20503 9977 20537
rect 10103 20503 10137 20537
rect 10263 20503 10297 20537
rect 10423 20503 10457 20537
rect 10583 20503 10617 20537
rect 10743 20503 10777 20537
rect 10903 20503 10937 20537
rect 11063 20503 11097 20537
rect 11223 20503 11257 20537
rect 11383 20503 11417 20537
rect 11543 20503 11577 20537
rect 11703 20503 11737 20537
rect 11863 20503 11897 20537
rect 12023 20503 12057 20537
rect 12183 20503 12217 20537
rect 12343 20503 12377 20537
rect 8503 20343 8537 20377
rect 8663 20343 8697 20377
rect 8823 20343 8857 20377
rect 8983 20343 9017 20377
rect 9143 20343 9177 20377
rect 9303 20343 9337 20377
rect 9463 20343 9497 20377
rect 9623 20343 9657 20377
rect 9783 20343 9817 20377
rect 9943 20343 9977 20377
rect 10103 20343 10137 20377
rect 10263 20343 10297 20377
rect 10423 20343 10457 20377
rect 10583 20343 10617 20377
rect 10743 20343 10777 20377
rect 10903 20343 10937 20377
rect 11063 20343 11097 20377
rect 11223 20343 11257 20377
rect 11383 20343 11417 20377
rect 11543 20343 11577 20377
rect 11703 20343 11737 20377
rect 11863 20343 11897 20377
rect 12023 20343 12057 20377
rect 12183 20343 12217 20377
rect 12343 20343 12377 20377
rect 8503 20183 8537 20217
rect 8663 20183 8697 20217
rect 8823 20183 8857 20217
rect 8983 20183 9017 20217
rect 9143 20183 9177 20217
rect 9303 20183 9337 20217
rect 9463 20183 9497 20217
rect 9623 20183 9657 20217
rect 9783 20183 9817 20217
rect 9943 20183 9977 20217
rect 10103 20183 10137 20217
rect 10263 20183 10297 20217
rect 10423 20183 10457 20217
rect 10583 20183 10617 20217
rect 10743 20183 10777 20217
rect 10903 20183 10937 20217
rect 11063 20183 11097 20217
rect 11223 20183 11257 20217
rect 11383 20183 11417 20217
rect 11543 20183 11577 20217
rect 11703 20183 11737 20217
rect 11863 20183 11897 20217
rect 12023 20183 12057 20217
rect 12183 20183 12217 20217
rect 12343 20183 12377 20217
rect 8503 20023 8537 20057
rect 8663 20023 8697 20057
rect 8823 20023 8857 20057
rect 8983 20023 9017 20057
rect 9143 20023 9177 20057
rect 9303 20023 9337 20057
rect 9463 20023 9497 20057
rect 9623 20023 9657 20057
rect 9783 20023 9817 20057
rect 9943 20023 9977 20057
rect 10103 20023 10137 20057
rect 10263 20023 10297 20057
rect 10423 20023 10457 20057
rect 10583 20023 10617 20057
rect 10743 20023 10777 20057
rect 10903 20023 10937 20057
rect 11063 20023 11097 20057
rect 11223 20023 11257 20057
rect 11383 20023 11417 20057
rect 11543 20023 11577 20057
rect 11703 20023 11737 20057
rect 11863 20023 11897 20057
rect 12023 20023 12057 20057
rect 12183 20023 12217 20057
rect 12343 20023 12377 20057
rect 8503 19863 8537 19897
rect 8663 19863 8697 19897
rect 8823 19863 8857 19897
rect 8983 19863 9017 19897
rect 9143 19863 9177 19897
rect 9303 19863 9337 19897
rect 9463 19863 9497 19897
rect 9623 19863 9657 19897
rect 9783 19863 9817 19897
rect 9943 19863 9977 19897
rect 10103 19863 10137 19897
rect 10263 19863 10297 19897
rect 10423 19863 10457 19897
rect 10583 19863 10617 19897
rect 10743 19863 10777 19897
rect 10903 19863 10937 19897
rect 11063 19863 11097 19897
rect 11223 19863 11257 19897
rect 11383 19863 11417 19897
rect 11543 19863 11577 19897
rect 11703 19863 11737 19897
rect 11863 19863 11897 19897
rect 12023 19863 12057 19897
rect 12183 19863 12217 19897
rect 12343 19863 12377 19897
rect 8503 19703 8537 19737
rect 8663 19703 8697 19737
rect 8823 19703 8857 19737
rect 8983 19703 9017 19737
rect 9143 19703 9177 19737
rect 9303 19703 9337 19737
rect 9463 19703 9497 19737
rect 9623 19703 9657 19737
rect 9783 19703 9817 19737
rect 9943 19703 9977 19737
rect 10103 19703 10137 19737
rect 10263 19703 10297 19737
rect 10423 19703 10457 19737
rect 10583 19703 10617 19737
rect 10743 19703 10777 19737
rect 10903 19703 10937 19737
rect 11063 19703 11097 19737
rect 11223 19703 11257 19737
rect 11383 19703 11417 19737
rect 11543 19703 11577 19737
rect 11703 19703 11737 19737
rect 11863 19703 11897 19737
rect 12023 19703 12057 19737
rect 12183 19703 12217 19737
rect 12343 19703 12377 19737
rect 8503 19543 8537 19577
rect 8663 19543 8697 19577
rect 8823 19543 8857 19577
rect 8983 19543 9017 19577
rect 9143 19543 9177 19577
rect 9303 19543 9337 19577
rect 9463 19543 9497 19577
rect 9623 19543 9657 19577
rect 9783 19543 9817 19577
rect 9943 19543 9977 19577
rect 10103 19543 10137 19577
rect 10263 19543 10297 19577
rect 10423 19543 10457 19577
rect 10583 19543 10617 19577
rect 10743 19543 10777 19577
rect 10903 19543 10937 19577
rect 11063 19543 11097 19577
rect 11223 19543 11257 19577
rect 11383 19543 11417 19577
rect 11543 19543 11577 19577
rect 11703 19543 11737 19577
rect 11863 19543 11897 19577
rect 12023 19543 12057 19577
rect 12183 19543 12217 19577
rect 12343 19543 12377 19577
rect 8503 19383 8537 19417
rect 8663 19383 8697 19417
rect 8823 19383 8857 19417
rect 8983 19383 9017 19417
rect 9143 19383 9177 19417
rect 9303 19383 9337 19417
rect 9463 19383 9497 19417
rect 9623 19383 9657 19417
rect 9783 19383 9817 19417
rect 9943 19383 9977 19417
rect 10103 19383 10137 19417
rect 10263 19383 10297 19417
rect 10423 19383 10457 19417
rect 10583 19383 10617 19417
rect 10743 19383 10777 19417
rect 10903 19383 10937 19417
rect 11063 19383 11097 19417
rect 11223 19383 11257 19417
rect 11383 19383 11417 19417
rect 11543 19383 11577 19417
rect 11703 19383 11737 19417
rect 11863 19383 11897 19417
rect 12023 19383 12057 19417
rect 12183 19383 12217 19417
rect 12343 19383 12377 19417
rect 8503 19223 8537 19257
rect 8663 19223 8697 19257
rect 8823 19223 8857 19257
rect 8983 19223 9017 19257
rect 9143 19223 9177 19257
rect 9303 19223 9337 19257
rect 9463 19223 9497 19257
rect 9623 19223 9657 19257
rect 9783 19223 9817 19257
rect 9943 19223 9977 19257
rect 10103 19223 10137 19257
rect 10263 19223 10297 19257
rect 10423 19223 10457 19257
rect 10583 19223 10617 19257
rect 10743 19223 10777 19257
rect 10903 19223 10937 19257
rect 11063 19223 11097 19257
rect 11223 19223 11257 19257
rect 11383 19223 11417 19257
rect 11543 19223 11577 19257
rect 11703 19223 11737 19257
rect 11863 19223 11897 19257
rect 12023 19223 12057 19257
rect 12183 19223 12217 19257
rect 12343 19223 12377 19257
rect 8503 19063 8537 19097
rect 8663 19063 8697 19097
rect 8823 19063 8857 19097
rect 8983 19063 9017 19097
rect 9143 19063 9177 19097
rect 9303 19063 9337 19097
rect 9463 19063 9497 19097
rect 9623 19063 9657 19097
rect 9783 19063 9817 19097
rect 9943 19063 9977 19097
rect 10103 19063 10137 19097
rect 10263 19063 10297 19097
rect 10423 19063 10457 19097
rect 10583 19063 10617 19097
rect 10743 19063 10777 19097
rect 10903 19063 10937 19097
rect 11063 19063 11097 19097
rect 11223 19063 11257 19097
rect 11383 19063 11417 19097
rect 11543 19063 11577 19097
rect 11703 19063 11737 19097
rect 11863 19063 11897 19097
rect 12023 19063 12057 19097
rect 12183 19063 12217 19097
rect 12343 19063 12377 19097
rect 8503 18903 8537 18937
rect 8663 18903 8697 18937
rect 8823 18903 8857 18937
rect 8983 18903 9017 18937
rect 9143 18903 9177 18937
rect 9303 18903 9337 18937
rect 9463 18903 9497 18937
rect 9623 18903 9657 18937
rect 9783 18903 9817 18937
rect 9943 18903 9977 18937
rect 10103 18903 10137 18937
rect 10263 18903 10297 18937
rect 10423 18903 10457 18937
rect 10583 18903 10617 18937
rect 10743 18903 10777 18937
rect 10903 18903 10937 18937
rect 11063 18903 11097 18937
rect 11223 18903 11257 18937
rect 11383 18903 11417 18937
rect 11543 18903 11577 18937
rect 11703 18903 11737 18937
rect 11863 18903 11897 18937
rect 12023 18903 12057 18937
rect 12183 18903 12217 18937
rect 12343 18903 12377 18937
rect 8503 18743 8537 18777
rect 8663 18743 8697 18777
rect 8823 18743 8857 18777
rect 8983 18743 9017 18777
rect 9143 18743 9177 18777
rect 9303 18743 9337 18777
rect 9463 18743 9497 18777
rect 9623 18743 9657 18777
rect 9783 18743 9817 18777
rect 9943 18743 9977 18777
rect 10103 18743 10137 18777
rect 10263 18743 10297 18777
rect 10423 18743 10457 18777
rect 10583 18743 10617 18777
rect 10743 18743 10777 18777
rect 10903 18743 10937 18777
rect 11063 18743 11097 18777
rect 11223 18743 11257 18777
rect 11383 18743 11417 18777
rect 11543 18743 11577 18777
rect 11703 18743 11737 18777
rect 11863 18743 11897 18777
rect 12023 18743 12057 18777
rect 12183 18743 12217 18777
rect 12343 18743 12377 18777
rect 8503 18583 8537 18617
rect 8663 18583 8697 18617
rect 8823 18583 8857 18617
rect 8983 18583 9017 18617
rect 9143 18583 9177 18617
rect 9303 18583 9337 18617
rect 9463 18583 9497 18617
rect 9623 18583 9657 18617
rect 9783 18583 9817 18617
rect 9943 18583 9977 18617
rect 10103 18583 10137 18617
rect 10263 18583 10297 18617
rect 10423 18583 10457 18617
rect 10583 18583 10617 18617
rect 10743 18583 10777 18617
rect 10903 18583 10937 18617
rect 11063 18583 11097 18617
rect 11223 18583 11257 18617
rect 11383 18583 11417 18617
rect 11543 18583 11577 18617
rect 11703 18583 11737 18617
rect 11863 18583 11897 18617
rect 12023 18583 12057 18617
rect 12183 18583 12217 18617
rect 12343 18583 12377 18617
rect 8503 18423 8537 18457
rect 8663 18423 8697 18457
rect 8823 18423 8857 18457
rect 8983 18423 9017 18457
rect 9143 18423 9177 18457
rect 9303 18423 9337 18457
rect 9463 18423 9497 18457
rect 9623 18423 9657 18457
rect 9783 18423 9817 18457
rect 9943 18423 9977 18457
rect 10103 18423 10137 18457
rect 10263 18423 10297 18457
rect 10423 18423 10457 18457
rect 10583 18423 10617 18457
rect 10743 18423 10777 18457
rect 10903 18423 10937 18457
rect 11063 18423 11097 18457
rect 11223 18423 11257 18457
rect 11383 18423 11417 18457
rect 11543 18423 11577 18457
rect 11703 18423 11737 18457
rect 11863 18423 11897 18457
rect 12023 18423 12057 18457
rect 12183 18423 12217 18457
rect 12343 18423 12377 18457
rect 8503 18263 8537 18297
rect 8663 18263 8697 18297
rect 8823 18263 8857 18297
rect 8983 18263 9017 18297
rect 9143 18263 9177 18297
rect 9303 18263 9337 18297
rect 9463 18263 9497 18297
rect 9623 18263 9657 18297
rect 9783 18263 9817 18297
rect 9943 18263 9977 18297
rect 10103 18263 10137 18297
rect 10263 18263 10297 18297
rect 10423 18263 10457 18297
rect 10583 18263 10617 18297
rect 10743 18263 10777 18297
rect 10903 18263 10937 18297
rect 11063 18263 11097 18297
rect 11223 18263 11257 18297
rect 11383 18263 11417 18297
rect 11543 18263 11577 18297
rect 11703 18263 11737 18297
rect 11863 18263 11897 18297
rect 12023 18263 12057 18297
rect 12183 18263 12217 18297
rect 12343 18263 12377 18297
rect 8503 18103 8537 18137
rect 8663 18103 8697 18137
rect 8823 18103 8857 18137
rect 8983 18103 9017 18137
rect 9143 18103 9177 18137
rect 9303 18103 9337 18137
rect 9463 18103 9497 18137
rect 9623 18103 9657 18137
rect 9783 18103 9817 18137
rect 9943 18103 9977 18137
rect 10103 18103 10137 18137
rect 10263 18103 10297 18137
rect 10423 18103 10457 18137
rect 10583 18103 10617 18137
rect 10743 18103 10777 18137
rect 10903 18103 10937 18137
rect 11063 18103 11097 18137
rect 11223 18103 11257 18137
rect 11383 18103 11417 18137
rect 11543 18103 11577 18137
rect 11703 18103 11737 18137
rect 11863 18103 11897 18137
rect 12023 18103 12057 18137
rect 12183 18103 12217 18137
rect 12343 18103 12377 18137
rect 8503 17943 8537 17977
rect 8663 17943 8697 17977
rect 8823 17943 8857 17977
rect 8983 17943 9017 17977
rect 9143 17943 9177 17977
rect 9303 17943 9337 17977
rect 9463 17943 9497 17977
rect 9623 17943 9657 17977
rect 9783 17943 9817 17977
rect 9943 17943 9977 17977
rect 10103 17943 10137 17977
rect 10263 17943 10297 17977
rect 10423 17943 10457 17977
rect 10583 17943 10617 17977
rect 10743 17943 10777 17977
rect 10903 17943 10937 17977
rect 11063 17943 11097 17977
rect 11223 17943 11257 17977
rect 11383 17943 11417 17977
rect 11543 17943 11577 17977
rect 11703 17943 11737 17977
rect 11863 17943 11897 17977
rect 12023 17943 12057 17977
rect 12183 17943 12217 17977
rect 12343 17943 12377 17977
rect 8503 17783 8537 17817
rect 8663 17783 8697 17817
rect 8823 17783 8857 17817
rect 8983 17783 9017 17817
rect 9143 17783 9177 17817
rect 9303 17783 9337 17817
rect 9463 17783 9497 17817
rect 9623 17783 9657 17817
rect 9783 17783 9817 17817
rect 9943 17783 9977 17817
rect 10103 17783 10137 17817
rect 10263 17783 10297 17817
rect 10423 17783 10457 17817
rect 10583 17783 10617 17817
rect 10743 17783 10777 17817
rect 10903 17783 10937 17817
rect 11063 17783 11097 17817
rect 11223 17783 11257 17817
rect 11383 17783 11417 17817
rect 11543 17783 11577 17817
rect 11703 17783 11737 17817
rect 11863 17783 11897 17817
rect 12023 17783 12057 17817
rect 12183 17783 12217 17817
rect 12343 17783 12377 17817
rect 8503 17623 8537 17657
rect 8663 17623 8697 17657
rect 8823 17623 8857 17657
rect 8983 17623 9017 17657
rect 9143 17623 9177 17657
rect 9303 17623 9337 17657
rect 9463 17623 9497 17657
rect 9623 17623 9657 17657
rect 9783 17623 9817 17657
rect 9943 17623 9977 17657
rect 10103 17623 10137 17657
rect 10263 17623 10297 17657
rect 10423 17623 10457 17657
rect 10583 17623 10617 17657
rect 10743 17623 10777 17657
rect 10903 17623 10937 17657
rect 11063 17623 11097 17657
rect 11223 17623 11257 17657
rect 11383 17623 11417 17657
rect 11543 17623 11577 17657
rect 11703 17623 11737 17657
rect 11863 17623 11897 17657
rect 12023 17623 12057 17657
rect 12183 17623 12217 17657
rect 12343 17623 12377 17657
rect 8503 17463 8537 17497
rect 8663 17463 8697 17497
rect 8823 17463 8857 17497
rect 8983 17463 9017 17497
rect 9143 17463 9177 17497
rect 9303 17463 9337 17497
rect 9463 17463 9497 17497
rect 9623 17463 9657 17497
rect 9783 17463 9817 17497
rect 9943 17463 9977 17497
rect 10103 17463 10137 17497
rect 10263 17463 10297 17497
rect 10423 17463 10457 17497
rect 10583 17463 10617 17497
rect 10743 17463 10777 17497
rect 10903 17463 10937 17497
rect 11063 17463 11097 17497
rect 11223 17463 11257 17497
rect 11383 17463 11417 17497
rect 11543 17463 11577 17497
rect 11703 17463 11737 17497
rect 11863 17463 11897 17497
rect 12023 17463 12057 17497
rect 12183 17463 12217 17497
rect 12343 17463 12377 17497
rect 8503 17303 8537 17337
rect 8663 17303 8697 17337
rect 8823 17303 8857 17337
rect 8983 17303 9017 17337
rect 9143 17303 9177 17337
rect 9303 17303 9337 17337
rect 9463 17303 9497 17337
rect 9623 17303 9657 17337
rect 9783 17303 9817 17337
rect 9943 17303 9977 17337
rect 10103 17303 10137 17337
rect 10263 17303 10297 17337
rect 10423 17303 10457 17337
rect 10583 17303 10617 17337
rect 10743 17303 10777 17337
rect 10903 17303 10937 17337
rect 11063 17303 11097 17337
rect 11223 17303 11257 17337
rect 11383 17303 11417 17337
rect 11543 17303 11577 17337
rect 11703 17303 11737 17337
rect 11863 17303 11897 17337
rect 12023 17303 12057 17337
rect 12183 17303 12217 17337
rect 12343 17303 12377 17337
rect 8503 17143 8537 17177
rect 8663 17143 8697 17177
rect 8823 17143 8857 17177
rect 8983 17143 9017 17177
rect 9143 17143 9177 17177
rect 9303 17143 9337 17177
rect 9463 17143 9497 17177
rect 9623 17143 9657 17177
rect 9783 17143 9817 17177
rect 9943 17143 9977 17177
rect 10103 17143 10137 17177
rect 10263 17143 10297 17177
rect 10423 17143 10457 17177
rect 10583 17143 10617 17177
rect 10743 17143 10777 17177
rect 10903 17143 10937 17177
rect 11063 17143 11097 17177
rect 11223 17143 11257 17177
rect 11383 17143 11417 17177
rect 11543 17143 11577 17177
rect 11703 17143 11737 17177
rect 11863 17143 11897 17177
rect 12023 17143 12057 17177
rect 12183 17143 12217 17177
rect 12343 17143 12377 17177
rect 8503 16983 8537 17017
rect 8663 16983 8697 17017
rect 8823 16983 8857 17017
rect 8983 16983 9017 17017
rect 9143 16983 9177 17017
rect 9303 16983 9337 17017
rect 9463 16983 9497 17017
rect 9623 16983 9657 17017
rect 9783 16983 9817 17017
rect 9943 16983 9977 17017
rect 10103 16983 10137 17017
rect 10263 16983 10297 17017
rect 10423 16983 10457 17017
rect 10583 16983 10617 17017
rect 10743 16983 10777 17017
rect 10903 16983 10937 17017
rect 11063 16983 11097 17017
rect 11223 16983 11257 17017
rect 11383 16983 11417 17017
rect 11543 16983 11577 17017
rect 11703 16983 11737 17017
rect 11863 16983 11897 17017
rect 12023 16983 12057 17017
rect 12183 16983 12217 17017
rect 12343 16983 12377 17017
rect 8503 16823 8537 16857
rect 8663 16823 8697 16857
rect 8823 16823 8857 16857
rect 8983 16823 9017 16857
rect 9143 16823 9177 16857
rect 9303 16823 9337 16857
rect 9463 16823 9497 16857
rect 9623 16823 9657 16857
rect 9783 16823 9817 16857
rect 9943 16823 9977 16857
rect 10103 16823 10137 16857
rect 10263 16823 10297 16857
rect 10423 16823 10457 16857
rect 10583 16823 10617 16857
rect 10743 16823 10777 16857
rect 10903 16823 10937 16857
rect 11063 16823 11097 16857
rect 11223 16823 11257 16857
rect 11383 16823 11417 16857
rect 11543 16823 11577 16857
rect 11703 16823 11737 16857
rect 11863 16823 11897 16857
rect 12023 16823 12057 16857
rect 12183 16823 12217 16857
rect 12343 16823 12377 16857
rect 8503 16663 8537 16697
rect 8663 16663 8697 16697
rect 8823 16663 8857 16697
rect 8983 16663 9017 16697
rect 9143 16663 9177 16697
rect 9303 16663 9337 16697
rect 9463 16663 9497 16697
rect 9623 16663 9657 16697
rect 9783 16663 9817 16697
rect 9943 16663 9977 16697
rect 10103 16663 10137 16697
rect 10263 16663 10297 16697
rect 10423 16663 10457 16697
rect 10583 16663 10617 16697
rect 10743 16663 10777 16697
rect 10903 16663 10937 16697
rect 11063 16663 11097 16697
rect 11223 16663 11257 16697
rect 11383 16663 11417 16697
rect 11543 16663 11577 16697
rect 11703 16663 11737 16697
rect 11863 16663 11897 16697
rect 12023 16663 12057 16697
rect 12183 16663 12217 16697
rect 12343 16663 12377 16697
rect 8503 16503 8537 16537
rect 8663 16503 8697 16537
rect 8823 16503 8857 16537
rect 8983 16503 9017 16537
rect 9143 16503 9177 16537
rect 9303 16503 9337 16537
rect 9463 16503 9497 16537
rect 9623 16503 9657 16537
rect 9783 16503 9817 16537
rect 9943 16503 9977 16537
rect 10103 16503 10137 16537
rect 10263 16503 10297 16537
rect 10423 16503 10457 16537
rect 10583 16503 10617 16537
rect 10743 16503 10777 16537
rect 10903 16503 10937 16537
rect 11063 16503 11097 16537
rect 11223 16503 11257 16537
rect 11383 16503 11417 16537
rect 11543 16503 11577 16537
rect 11703 16503 11737 16537
rect 11863 16503 11897 16537
rect 12023 16503 12057 16537
rect 12183 16503 12217 16537
rect 12343 16503 12377 16537
rect 8503 16343 8537 16377
rect 8663 16343 8697 16377
rect 8823 16343 8857 16377
rect 8983 16343 9017 16377
rect 9143 16343 9177 16377
rect 9303 16343 9337 16377
rect 9463 16343 9497 16377
rect 9623 16343 9657 16377
rect 9783 16343 9817 16377
rect 9943 16343 9977 16377
rect 10103 16343 10137 16377
rect 10263 16343 10297 16377
rect 10423 16343 10457 16377
rect 10583 16343 10617 16377
rect 10743 16343 10777 16377
rect 10903 16343 10937 16377
rect 11063 16343 11097 16377
rect 11223 16343 11257 16377
rect 11383 16343 11417 16377
rect 11543 16343 11577 16377
rect 11703 16343 11737 16377
rect 11863 16343 11897 16377
rect 12023 16343 12057 16377
rect 12183 16343 12217 16377
rect 12343 16343 12377 16377
rect 8503 16183 8537 16217
rect 8663 16183 8697 16217
rect 8823 16183 8857 16217
rect 8983 16183 9017 16217
rect 9143 16183 9177 16217
rect 9303 16183 9337 16217
rect 9463 16183 9497 16217
rect 9623 16183 9657 16217
rect 9783 16183 9817 16217
rect 9943 16183 9977 16217
rect 10103 16183 10137 16217
rect 10263 16183 10297 16217
rect 10423 16183 10457 16217
rect 10583 16183 10617 16217
rect 10743 16183 10777 16217
rect 10903 16183 10937 16217
rect 11063 16183 11097 16217
rect 11223 16183 11257 16217
rect 11383 16183 11417 16217
rect 11543 16183 11577 16217
rect 11703 16183 11737 16217
rect 11863 16183 11897 16217
rect 12023 16183 12057 16217
rect 12183 16183 12217 16217
rect 12343 16183 12377 16217
rect 8503 16023 8537 16057
rect 8663 16023 8697 16057
rect 8823 16023 8857 16057
rect 8983 16023 9017 16057
rect 9143 16023 9177 16057
rect 9303 16023 9337 16057
rect 9463 16023 9497 16057
rect 9623 16023 9657 16057
rect 9783 16023 9817 16057
rect 9943 16023 9977 16057
rect 10103 16023 10137 16057
rect 10263 16023 10297 16057
rect 10423 16023 10457 16057
rect 10583 16023 10617 16057
rect 10743 16023 10777 16057
rect 10903 16023 10937 16057
rect 11063 16023 11097 16057
rect 11223 16023 11257 16057
rect 11383 16023 11417 16057
rect 11543 16023 11577 16057
rect 11703 16023 11737 16057
rect 11863 16023 11897 16057
rect 12023 16023 12057 16057
rect 12183 16023 12217 16057
rect 12343 16023 12377 16057
rect 8503 15863 8537 15897
rect 8663 15863 8697 15897
rect 8823 15863 8857 15897
rect 8983 15863 9017 15897
rect 9143 15863 9177 15897
rect 9303 15863 9337 15897
rect 9463 15863 9497 15897
rect 9623 15863 9657 15897
rect 9783 15863 9817 15897
rect 9943 15863 9977 15897
rect 10103 15863 10137 15897
rect 10263 15863 10297 15897
rect 10423 15863 10457 15897
rect 10583 15863 10617 15897
rect 10743 15863 10777 15897
rect 10903 15863 10937 15897
rect 11063 15863 11097 15897
rect 11223 15863 11257 15897
rect 11383 15863 11417 15897
rect 11543 15863 11577 15897
rect 11703 15863 11737 15897
rect 11863 15863 11897 15897
rect 12023 15863 12057 15897
rect 12183 15863 12217 15897
rect 12343 15863 12377 15897
rect 8503 15703 8537 15737
rect 8663 15703 8697 15737
rect 8823 15703 8857 15737
rect 8983 15703 9017 15737
rect 9143 15703 9177 15737
rect 9303 15703 9337 15737
rect 9463 15703 9497 15737
rect 9623 15703 9657 15737
rect 9783 15703 9817 15737
rect 9943 15703 9977 15737
rect 10103 15703 10137 15737
rect 10263 15703 10297 15737
rect 10423 15703 10457 15737
rect 10583 15703 10617 15737
rect 10743 15703 10777 15737
rect 10903 15703 10937 15737
rect 11063 15703 11097 15737
rect 11223 15703 11257 15737
rect 11383 15703 11417 15737
rect 11543 15703 11577 15737
rect 11703 15703 11737 15737
rect 11863 15703 11897 15737
rect 12023 15703 12057 15737
rect 12183 15703 12217 15737
rect 12343 15703 12377 15737
rect 8503 15543 8537 15577
rect 8663 15543 8697 15577
rect 8823 15543 8857 15577
rect 8983 15543 9017 15577
rect 9143 15543 9177 15577
rect 9303 15543 9337 15577
rect 9463 15543 9497 15577
rect 9623 15543 9657 15577
rect 9783 15543 9817 15577
rect 9943 15543 9977 15577
rect 10103 15543 10137 15577
rect 10263 15543 10297 15577
rect 10423 15543 10457 15577
rect 10583 15543 10617 15577
rect 10743 15543 10777 15577
rect 10903 15543 10937 15577
rect 11063 15543 11097 15577
rect 11223 15543 11257 15577
rect 11383 15543 11417 15577
rect 11543 15543 11577 15577
rect 11703 15543 11737 15577
rect 11863 15543 11897 15577
rect 12023 15543 12057 15577
rect 12183 15543 12217 15577
rect 12343 15543 12377 15577
rect 8503 15383 8537 15417
rect 8663 15383 8697 15417
rect 8823 15383 8857 15417
rect 8983 15383 9017 15417
rect 9143 15383 9177 15417
rect 9303 15383 9337 15417
rect 9463 15383 9497 15417
rect 9623 15383 9657 15417
rect 9783 15383 9817 15417
rect 9943 15383 9977 15417
rect 10103 15383 10137 15417
rect 10263 15383 10297 15417
rect 10423 15383 10457 15417
rect 10583 15383 10617 15417
rect 10743 15383 10777 15417
rect 10903 15383 10937 15417
rect 11063 15383 11097 15417
rect 11223 15383 11257 15417
rect 11383 15383 11417 15417
rect 11543 15383 11577 15417
rect 11703 15383 11737 15417
rect 11863 15383 11897 15417
rect 12023 15383 12057 15417
rect 12183 15383 12217 15417
rect 12343 15383 12377 15417
rect 8503 15223 8537 15257
rect 8663 15223 8697 15257
rect 8823 15223 8857 15257
rect 8983 15223 9017 15257
rect 9143 15223 9177 15257
rect 9303 15223 9337 15257
rect 9463 15223 9497 15257
rect 9623 15223 9657 15257
rect 9783 15223 9817 15257
rect 9943 15223 9977 15257
rect 10103 15223 10137 15257
rect 10263 15223 10297 15257
rect 10423 15223 10457 15257
rect 10583 15223 10617 15257
rect 10743 15223 10777 15257
rect 10903 15223 10937 15257
rect 11063 15223 11097 15257
rect 11223 15223 11257 15257
rect 11383 15223 11417 15257
rect 11543 15223 11577 15257
rect 11703 15223 11737 15257
rect 11863 15223 11897 15257
rect 12023 15223 12057 15257
rect 12183 15223 12217 15257
rect 12343 15223 12377 15257
rect 8503 15063 8537 15097
rect 8663 15063 8697 15097
rect 8823 15063 8857 15097
rect 8983 15063 9017 15097
rect 9143 15063 9177 15097
rect 9303 15063 9337 15097
rect 9463 15063 9497 15097
rect 9623 15063 9657 15097
rect 9783 15063 9817 15097
rect 9943 15063 9977 15097
rect 10103 15063 10137 15097
rect 10263 15063 10297 15097
rect 10423 15063 10457 15097
rect 10583 15063 10617 15097
rect 10743 15063 10777 15097
rect 10903 15063 10937 15097
rect 11063 15063 11097 15097
rect 11223 15063 11257 15097
rect 11383 15063 11417 15097
rect 11543 15063 11577 15097
rect 11703 15063 11737 15097
rect 11863 15063 11897 15097
rect 12023 15063 12057 15097
rect 12183 15063 12217 15097
rect 12343 15063 12377 15097
rect 8503 14903 8537 14937
rect 8663 14903 8697 14937
rect 8823 14903 8857 14937
rect 8983 14903 9017 14937
rect 9143 14903 9177 14937
rect 9303 14903 9337 14937
rect 9463 14903 9497 14937
rect 9623 14903 9657 14937
rect 9783 14903 9817 14937
rect 9943 14903 9977 14937
rect 10103 14903 10137 14937
rect 10263 14903 10297 14937
rect 10423 14903 10457 14937
rect 10583 14903 10617 14937
rect 10743 14903 10777 14937
rect 10903 14903 10937 14937
rect 11063 14903 11097 14937
rect 11223 14903 11257 14937
rect 11383 14903 11417 14937
rect 11543 14903 11577 14937
rect 11703 14903 11737 14937
rect 11863 14903 11897 14937
rect 12023 14903 12057 14937
rect 12183 14903 12217 14937
rect 12343 14903 12377 14937
rect 8503 14743 8537 14777
rect 8663 14743 8697 14777
rect 8823 14743 8857 14777
rect 8983 14743 9017 14777
rect 9143 14743 9177 14777
rect 9303 14743 9337 14777
rect 9463 14743 9497 14777
rect 9623 14743 9657 14777
rect 9783 14743 9817 14777
rect 9943 14743 9977 14777
rect 10103 14743 10137 14777
rect 10263 14743 10297 14777
rect 10423 14743 10457 14777
rect 10583 14743 10617 14777
rect 10743 14743 10777 14777
rect 10903 14743 10937 14777
rect 11063 14743 11097 14777
rect 11223 14743 11257 14777
rect 11383 14743 11417 14777
rect 11543 14743 11577 14777
rect 11703 14743 11737 14777
rect 11863 14743 11897 14777
rect 12023 14743 12057 14777
rect 12183 14743 12217 14777
rect 12343 14743 12377 14777
rect 8503 14583 8537 14617
rect 8663 14583 8697 14617
rect 8823 14583 8857 14617
rect 8983 14583 9017 14617
rect 9143 14583 9177 14617
rect 9303 14583 9337 14617
rect 9463 14583 9497 14617
rect 9623 14583 9657 14617
rect 9783 14583 9817 14617
rect 9943 14583 9977 14617
rect 10103 14583 10137 14617
rect 10263 14583 10297 14617
rect 10423 14583 10457 14617
rect 10583 14583 10617 14617
rect 10743 14583 10777 14617
rect 10903 14583 10937 14617
rect 11063 14583 11097 14617
rect 11223 14583 11257 14617
rect 11383 14583 11417 14617
rect 11543 14583 11577 14617
rect 11703 14583 11737 14617
rect 11863 14583 11897 14617
rect 12023 14583 12057 14617
rect 12183 14583 12217 14617
rect 12343 14583 12377 14617
rect 8503 14423 8537 14457
rect 8663 14423 8697 14457
rect 8823 14423 8857 14457
rect 8983 14423 9017 14457
rect 9143 14423 9177 14457
rect 9303 14423 9337 14457
rect 9463 14423 9497 14457
rect 9623 14423 9657 14457
rect 9783 14423 9817 14457
rect 9943 14423 9977 14457
rect 10103 14423 10137 14457
rect 10263 14423 10297 14457
rect 10423 14423 10457 14457
rect 10583 14423 10617 14457
rect 10743 14423 10777 14457
rect 10903 14423 10937 14457
rect 11063 14423 11097 14457
rect 11223 14423 11257 14457
rect 11383 14423 11417 14457
rect 11543 14423 11577 14457
rect 11703 14423 11737 14457
rect 11863 14423 11897 14457
rect 12023 14423 12057 14457
rect 12183 14423 12217 14457
rect 12343 14423 12377 14457
rect 8503 14263 8537 14297
rect 8663 14263 8697 14297
rect 8823 14263 8857 14297
rect 8983 14263 9017 14297
rect 9143 14263 9177 14297
rect 9303 14263 9337 14297
rect 9463 14263 9497 14297
rect 9623 14263 9657 14297
rect 9783 14263 9817 14297
rect 9943 14263 9977 14297
rect 10103 14263 10137 14297
rect 10263 14263 10297 14297
rect 10423 14263 10457 14297
rect 10583 14263 10617 14297
rect 10743 14263 10777 14297
rect 10903 14263 10937 14297
rect 11063 14263 11097 14297
rect 11223 14263 11257 14297
rect 11383 14263 11417 14297
rect 11543 14263 11577 14297
rect 11703 14263 11737 14297
rect 11863 14263 11897 14297
rect 12023 14263 12057 14297
rect 12183 14263 12217 14297
rect 12343 14263 12377 14297
rect 8503 14103 8537 14137
rect 8663 14103 8697 14137
rect 8823 14103 8857 14137
rect 8983 14103 9017 14137
rect 9143 14103 9177 14137
rect 9303 14103 9337 14137
rect 9463 14103 9497 14137
rect 9623 14103 9657 14137
rect 9783 14103 9817 14137
rect 9943 14103 9977 14137
rect 10103 14103 10137 14137
rect 10263 14103 10297 14137
rect 10423 14103 10457 14137
rect 10583 14103 10617 14137
rect 10743 14103 10777 14137
rect 10903 14103 10937 14137
rect 11063 14103 11097 14137
rect 11223 14103 11257 14137
rect 11383 14103 11417 14137
rect 11543 14103 11577 14137
rect 11703 14103 11737 14137
rect 11863 14103 11897 14137
rect 12023 14103 12057 14137
rect 12183 14103 12217 14137
rect 12343 14103 12377 14137
rect 8503 13943 8537 13977
rect 8663 13943 8697 13977
rect 8823 13943 8857 13977
rect 8983 13943 9017 13977
rect 9143 13943 9177 13977
rect 9303 13943 9337 13977
rect 9463 13943 9497 13977
rect 9623 13943 9657 13977
rect 9783 13943 9817 13977
rect 9943 13943 9977 13977
rect 10103 13943 10137 13977
rect 10263 13943 10297 13977
rect 10423 13943 10457 13977
rect 10583 13943 10617 13977
rect 10743 13943 10777 13977
rect 10903 13943 10937 13977
rect 11063 13943 11097 13977
rect 11223 13943 11257 13977
rect 11383 13943 11417 13977
rect 11543 13943 11577 13977
rect 11703 13943 11737 13977
rect 11863 13943 11897 13977
rect 12023 13943 12057 13977
rect 12183 13943 12217 13977
rect 12343 13943 12377 13977
rect 8503 13783 8537 13817
rect 8663 13783 8697 13817
rect 8823 13783 8857 13817
rect 8983 13783 9017 13817
rect 9143 13783 9177 13817
rect 9303 13783 9337 13817
rect 9463 13783 9497 13817
rect 9623 13783 9657 13817
rect 9783 13783 9817 13817
rect 9943 13783 9977 13817
rect 10103 13783 10137 13817
rect 10263 13783 10297 13817
rect 10423 13783 10457 13817
rect 10583 13783 10617 13817
rect 10743 13783 10777 13817
rect 10903 13783 10937 13817
rect 11063 13783 11097 13817
rect 11223 13783 11257 13817
rect 11383 13783 11417 13817
rect 11543 13783 11577 13817
rect 11703 13783 11737 13817
rect 11863 13783 11897 13817
rect 12023 13783 12057 13817
rect 12183 13783 12217 13817
rect 12343 13783 12377 13817
rect 8503 13623 8537 13657
rect 8663 13623 8697 13657
rect 8823 13623 8857 13657
rect 8983 13623 9017 13657
rect 9143 13623 9177 13657
rect 9303 13623 9337 13657
rect 9463 13623 9497 13657
rect 9623 13623 9657 13657
rect 9783 13623 9817 13657
rect 9943 13623 9977 13657
rect 10103 13623 10137 13657
rect 10263 13623 10297 13657
rect 10423 13623 10457 13657
rect 10583 13623 10617 13657
rect 10743 13623 10777 13657
rect 10903 13623 10937 13657
rect 11063 13623 11097 13657
rect 11223 13623 11257 13657
rect 11383 13623 11417 13657
rect 11543 13623 11577 13657
rect 11703 13623 11737 13657
rect 11863 13623 11897 13657
rect 12023 13623 12057 13657
rect 12183 13623 12217 13657
rect 12343 13623 12377 13657
rect 8503 13463 8537 13497
rect 8663 13463 8697 13497
rect 8823 13463 8857 13497
rect 8983 13463 9017 13497
rect 9143 13463 9177 13497
rect 9303 13463 9337 13497
rect 9463 13463 9497 13497
rect 9623 13463 9657 13497
rect 9783 13463 9817 13497
rect 9943 13463 9977 13497
rect 10103 13463 10137 13497
rect 10263 13463 10297 13497
rect 10423 13463 10457 13497
rect 10583 13463 10617 13497
rect 10743 13463 10777 13497
rect 10903 13463 10937 13497
rect 11063 13463 11097 13497
rect 11223 13463 11257 13497
rect 11383 13463 11417 13497
rect 11543 13463 11577 13497
rect 11703 13463 11737 13497
rect 11863 13463 11897 13497
rect 12023 13463 12057 13497
rect 12183 13463 12217 13497
rect 12343 13463 12377 13497
rect 8503 13303 8537 13337
rect 8663 13303 8697 13337
rect 8823 13303 8857 13337
rect 8983 13303 9017 13337
rect 9143 13303 9177 13337
rect 9303 13303 9337 13337
rect 9463 13303 9497 13337
rect 9623 13303 9657 13337
rect 9783 13303 9817 13337
rect 9943 13303 9977 13337
rect 10103 13303 10137 13337
rect 10263 13303 10297 13337
rect 10423 13303 10457 13337
rect 10583 13303 10617 13337
rect 10743 13303 10777 13337
rect 10903 13303 10937 13337
rect 11063 13303 11097 13337
rect 11223 13303 11257 13337
rect 11383 13303 11417 13337
rect 11543 13303 11577 13337
rect 11703 13303 11737 13337
rect 11863 13303 11897 13337
rect 12023 13303 12057 13337
rect 12183 13303 12217 13337
rect 12343 13303 12377 13337
rect 8503 13143 8537 13177
rect 8663 13143 8697 13177
rect 8823 13143 8857 13177
rect 8983 13143 9017 13177
rect 9143 13143 9177 13177
rect 9303 13143 9337 13177
rect 9463 13143 9497 13177
rect 9623 13143 9657 13177
rect 9783 13143 9817 13177
rect 9943 13143 9977 13177
rect 10103 13143 10137 13177
rect 10263 13143 10297 13177
rect 10423 13143 10457 13177
rect 10583 13143 10617 13177
rect 10743 13143 10777 13177
rect 10903 13143 10937 13177
rect 11063 13143 11097 13177
rect 11223 13143 11257 13177
rect 11383 13143 11417 13177
rect 11543 13143 11577 13177
rect 11703 13143 11737 13177
rect 11863 13143 11897 13177
rect 12023 13143 12057 13177
rect 12183 13143 12217 13177
rect 12343 13143 12377 13177
rect 8503 12983 8537 13017
rect 8663 12983 8697 13017
rect 8823 12983 8857 13017
rect 8983 12983 9017 13017
rect 9143 12983 9177 13017
rect 9303 12983 9337 13017
rect 9463 12983 9497 13017
rect 9623 12983 9657 13017
rect 9783 12983 9817 13017
rect 9943 12983 9977 13017
rect 10103 12983 10137 13017
rect 10263 12983 10297 13017
rect 10423 12983 10457 13017
rect 10583 12983 10617 13017
rect 10743 12983 10777 13017
rect 10903 12983 10937 13017
rect 11063 12983 11097 13017
rect 11223 12983 11257 13017
rect 11383 12983 11417 13017
rect 11543 12983 11577 13017
rect 11703 12983 11737 13017
rect 11863 12983 11897 13017
rect 12023 12983 12057 13017
rect 12183 12983 12217 13017
rect 12343 12983 12377 13017
rect 8503 12823 8537 12857
rect 8663 12823 8697 12857
rect 8823 12823 8857 12857
rect 8983 12823 9017 12857
rect 9143 12823 9177 12857
rect 9303 12823 9337 12857
rect 9463 12823 9497 12857
rect 9623 12823 9657 12857
rect 9783 12823 9817 12857
rect 9943 12823 9977 12857
rect 10103 12823 10137 12857
rect 10263 12823 10297 12857
rect 10423 12823 10457 12857
rect 10583 12823 10617 12857
rect 10743 12823 10777 12857
rect 10903 12823 10937 12857
rect 11063 12823 11097 12857
rect 11223 12823 11257 12857
rect 11383 12823 11417 12857
rect 11543 12823 11577 12857
rect 11703 12823 11737 12857
rect 11863 12823 11897 12857
rect 12023 12823 12057 12857
rect 12183 12823 12217 12857
rect 12343 12823 12377 12857
rect 8503 12663 8537 12697
rect 8663 12663 8697 12697
rect 8823 12663 8857 12697
rect 8983 12663 9017 12697
rect 9143 12663 9177 12697
rect 9303 12663 9337 12697
rect 9463 12663 9497 12697
rect 9623 12663 9657 12697
rect 9783 12663 9817 12697
rect 9943 12663 9977 12697
rect 10103 12663 10137 12697
rect 10263 12663 10297 12697
rect 10423 12663 10457 12697
rect 10583 12663 10617 12697
rect 10743 12663 10777 12697
rect 10903 12663 10937 12697
rect 11063 12663 11097 12697
rect 11223 12663 11257 12697
rect 11383 12663 11417 12697
rect 11543 12663 11577 12697
rect 11703 12663 11737 12697
rect 11863 12663 11897 12697
rect 12023 12663 12057 12697
rect 12183 12663 12217 12697
rect 12343 12663 12377 12697
rect 8503 12503 8537 12537
rect 8663 12503 8697 12537
rect 8823 12503 8857 12537
rect 8983 12503 9017 12537
rect 9143 12503 9177 12537
rect 9303 12503 9337 12537
rect 9463 12503 9497 12537
rect 9623 12503 9657 12537
rect 9783 12503 9817 12537
rect 9943 12503 9977 12537
rect 10103 12503 10137 12537
rect 10263 12503 10297 12537
rect 10423 12503 10457 12537
rect 10583 12503 10617 12537
rect 10743 12503 10777 12537
rect 10903 12503 10937 12537
rect 11063 12503 11097 12537
rect 11223 12503 11257 12537
rect 11383 12503 11417 12537
rect 11543 12503 11577 12537
rect 11703 12503 11737 12537
rect 11863 12503 11897 12537
rect 12023 12503 12057 12537
rect 12183 12503 12217 12537
rect 12343 12503 12377 12537
rect 8503 12343 8537 12377
rect 8663 12343 8697 12377
rect 8823 12343 8857 12377
rect 8983 12343 9017 12377
rect 9143 12343 9177 12377
rect 9303 12343 9337 12377
rect 9463 12343 9497 12377
rect 9623 12343 9657 12377
rect 9783 12343 9817 12377
rect 9943 12343 9977 12377
rect 10103 12343 10137 12377
rect 10263 12343 10297 12377
rect 10423 12343 10457 12377
rect 10583 12343 10617 12377
rect 10743 12343 10777 12377
rect 10903 12343 10937 12377
rect 11063 12343 11097 12377
rect 11223 12343 11257 12377
rect 11383 12343 11417 12377
rect 11543 12343 11577 12377
rect 11703 12343 11737 12377
rect 11863 12343 11897 12377
rect 12023 12343 12057 12377
rect 12183 12343 12217 12377
rect 12343 12343 12377 12377
rect 8503 12183 8537 12217
rect 8663 12183 8697 12217
rect 8823 12183 8857 12217
rect 8983 12183 9017 12217
rect 9143 12183 9177 12217
rect 9303 12183 9337 12217
rect 9463 12183 9497 12217
rect 9623 12183 9657 12217
rect 9783 12183 9817 12217
rect 9943 12183 9977 12217
rect 10103 12183 10137 12217
rect 10263 12183 10297 12217
rect 10423 12183 10457 12217
rect 10583 12183 10617 12217
rect 10743 12183 10777 12217
rect 10903 12183 10937 12217
rect 11063 12183 11097 12217
rect 11223 12183 11257 12217
rect 11383 12183 11417 12217
rect 11543 12183 11577 12217
rect 11703 12183 11737 12217
rect 11863 12183 11897 12217
rect 12023 12183 12057 12217
rect 12183 12183 12217 12217
rect 12343 12183 12377 12217
rect 8503 12023 8537 12057
rect 8663 12023 8697 12057
rect 8823 12023 8857 12057
rect 8983 12023 9017 12057
rect 9143 12023 9177 12057
rect 9303 12023 9337 12057
rect 9463 12023 9497 12057
rect 9623 12023 9657 12057
rect 9783 12023 9817 12057
rect 9943 12023 9977 12057
rect 10103 12023 10137 12057
rect 10263 12023 10297 12057
rect 10423 12023 10457 12057
rect 10583 12023 10617 12057
rect 10743 12023 10777 12057
rect 10903 12023 10937 12057
rect 11063 12023 11097 12057
rect 11223 12023 11257 12057
rect 11383 12023 11417 12057
rect 11543 12023 11577 12057
rect 11703 12023 11737 12057
rect 11863 12023 11897 12057
rect 12023 12023 12057 12057
rect 12183 12023 12217 12057
rect 12343 12023 12377 12057
rect 8503 11863 8537 11897
rect 8663 11863 8697 11897
rect 8823 11863 8857 11897
rect 8983 11863 9017 11897
rect 9143 11863 9177 11897
rect 9303 11863 9337 11897
rect 9463 11863 9497 11897
rect 9623 11863 9657 11897
rect 9783 11863 9817 11897
rect 9943 11863 9977 11897
rect 10103 11863 10137 11897
rect 10263 11863 10297 11897
rect 10423 11863 10457 11897
rect 10583 11863 10617 11897
rect 10743 11863 10777 11897
rect 10903 11863 10937 11897
rect 11063 11863 11097 11897
rect 11223 11863 11257 11897
rect 11383 11863 11417 11897
rect 11543 11863 11577 11897
rect 11703 11863 11737 11897
rect 11863 11863 11897 11897
rect 12023 11863 12057 11897
rect 12183 11863 12217 11897
rect 12343 11863 12377 11897
rect 8503 11703 8537 11737
rect 8663 11703 8697 11737
rect 8823 11703 8857 11737
rect 8983 11703 9017 11737
rect 9143 11703 9177 11737
rect 9303 11703 9337 11737
rect 9463 11703 9497 11737
rect 9623 11703 9657 11737
rect 9783 11703 9817 11737
rect 9943 11703 9977 11737
rect 10103 11703 10137 11737
rect 10263 11703 10297 11737
rect 10423 11703 10457 11737
rect 10583 11703 10617 11737
rect 10743 11703 10777 11737
rect 10903 11703 10937 11737
rect 11063 11703 11097 11737
rect 11223 11703 11257 11737
rect 11383 11703 11417 11737
rect 11543 11703 11577 11737
rect 11703 11703 11737 11737
rect 11863 11703 11897 11737
rect 12023 11703 12057 11737
rect 12183 11703 12217 11737
rect 12343 11703 12377 11737
rect 8503 11543 8537 11577
rect 8663 11543 8697 11577
rect 8823 11543 8857 11577
rect 8983 11543 9017 11577
rect 9143 11543 9177 11577
rect 9303 11543 9337 11577
rect 9463 11543 9497 11577
rect 9623 11543 9657 11577
rect 9783 11543 9817 11577
rect 9943 11543 9977 11577
rect 10103 11543 10137 11577
rect 10263 11543 10297 11577
rect 10423 11543 10457 11577
rect 10583 11543 10617 11577
rect 10743 11543 10777 11577
rect 10903 11543 10937 11577
rect 11063 11543 11097 11577
rect 11223 11543 11257 11577
rect 11383 11543 11417 11577
rect 11543 11543 11577 11577
rect 11703 11543 11737 11577
rect 11863 11543 11897 11577
rect 12023 11543 12057 11577
rect 12183 11543 12217 11577
rect 12343 11543 12377 11577
rect 8503 11383 8537 11417
rect 8663 11383 8697 11417
rect 8823 11383 8857 11417
rect 8983 11383 9017 11417
rect 9143 11383 9177 11417
rect 9303 11383 9337 11417
rect 9463 11383 9497 11417
rect 9623 11383 9657 11417
rect 9783 11383 9817 11417
rect 9943 11383 9977 11417
rect 10103 11383 10137 11417
rect 10263 11383 10297 11417
rect 10423 11383 10457 11417
rect 10583 11383 10617 11417
rect 10743 11383 10777 11417
rect 10903 11383 10937 11417
rect 11063 11383 11097 11417
rect 11223 11383 11257 11417
rect 11383 11383 11417 11417
rect 11543 11383 11577 11417
rect 11703 11383 11737 11417
rect 11863 11383 11897 11417
rect 12023 11383 12057 11417
rect 12183 11383 12217 11417
rect 12343 11383 12377 11417
rect 8503 11223 8537 11257
rect 8663 11223 8697 11257
rect 8823 11223 8857 11257
rect 8983 11223 9017 11257
rect 9143 11223 9177 11257
rect 9303 11223 9337 11257
rect 9463 11223 9497 11257
rect 9623 11223 9657 11257
rect 9783 11223 9817 11257
rect 9943 11223 9977 11257
rect 10103 11223 10137 11257
rect 10263 11223 10297 11257
rect 10423 11223 10457 11257
rect 10583 11223 10617 11257
rect 10743 11223 10777 11257
rect 10903 11223 10937 11257
rect 11063 11223 11097 11257
rect 11223 11223 11257 11257
rect 11383 11223 11417 11257
rect 11543 11223 11577 11257
rect 11703 11223 11737 11257
rect 11863 11223 11897 11257
rect 12023 11223 12057 11257
rect 12183 11223 12217 11257
rect 12343 11223 12377 11257
rect 8503 11063 8537 11097
rect 8663 11063 8697 11097
rect 8823 11063 8857 11097
rect 8983 11063 9017 11097
rect 9143 11063 9177 11097
rect 9303 11063 9337 11097
rect 9463 11063 9497 11097
rect 9623 11063 9657 11097
rect 9783 11063 9817 11097
rect 9943 11063 9977 11097
rect 10103 11063 10137 11097
rect 10263 11063 10297 11097
rect 10423 11063 10457 11097
rect 10583 11063 10617 11097
rect 10743 11063 10777 11097
rect 10903 11063 10937 11097
rect 11063 11063 11097 11097
rect 11223 11063 11257 11097
rect 11383 11063 11417 11097
rect 11543 11063 11577 11097
rect 11703 11063 11737 11097
rect 11863 11063 11897 11097
rect 12023 11063 12057 11097
rect 12183 11063 12217 11097
rect 12343 11063 12377 11097
rect 8503 10903 8537 10937
rect 8663 10903 8697 10937
rect 8823 10903 8857 10937
rect 8983 10903 9017 10937
rect 9143 10903 9177 10937
rect 9303 10903 9337 10937
rect 9463 10903 9497 10937
rect 9623 10903 9657 10937
rect 9783 10903 9817 10937
rect 9943 10903 9977 10937
rect 10103 10903 10137 10937
rect 10263 10903 10297 10937
rect 10423 10903 10457 10937
rect 10583 10903 10617 10937
rect 10743 10903 10777 10937
rect 10903 10903 10937 10937
rect 11063 10903 11097 10937
rect 11223 10903 11257 10937
rect 11383 10903 11417 10937
rect 11543 10903 11577 10937
rect 11703 10903 11737 10937
rect 11863 10903 11897 10937
rect 12023 10903 12057 10937
rect 12183 10903 12217 10937
rect 12343 10903 12377 10937
rect 8503 10743 8537 10777
rect 8663 10743 8697 10777
rect 8823 10743 8857 10777
rect 8983 10743 9017 10777
rect 9143 10743 9177 10777
rect 9303 10743 9337 10777
rect 9463 10743 9497 10777
rect 9623 10743 9657 10777
rect 9783 10743 9817 10777
rect 9943 10743 9977 10777
rect 10103 10743 10137 10777
rect 10263 10743 10297 10777
rect 10423 10743 10457 10777
rect 10583 10743 10617 10777
rect 10743 10743 10777 10777
rect 10903 10743 10937 10777
rect 11063 10743 11097 10777
rect 11223 10743 11257 10777
rect 11383 10743 11417 10777
rect 11543 10743 11577 10777
rect 11703 10743 11737 10777
rect 11863 10743 11897 10777
rect 12023 10743 12057 10777
rect 12183 10743 12217 10777
rect 12343 10743 12377 10777
rect 8503 10583 8537 10617
rect 8663 10583 8697 10617
rect 8823 10583 8857 10617
rect 8983 10583 9017 10617
rect 9143 10583 9177 10617
rect 9303 10583 9337 10617
rect 9463 10583 9497 10617
rect 9623 10583 9657 10617
rect 9783 10583 9817 10617
rect 9943 10583 9977 10617
rect 10103 10583 10137 10617
rect 10263 10583 10297 10617
rect 10423 10583 10457 10617
rect 10583 10583 10617 10617
rect 10743 10583 10777 10617
rect 10903 10583 10937 10617
rect 11063 10583 11097 10617
rect 11223 10583 11257 10617
rect 11383 10583 11417 10617
rect 11543 10583 11577 10617
rect 11703 10583 11737 10617
rect 11863 10583 11897 10617
rect 12023 10583 12057 10617
rect 12183 10583 12217 10617
rect 12343 10583 12377 10617
rect 8503 10423 8537 10457
rect 8663 10423 8697 10457
rect 8823 10423 8857 10457
rect 8983 10423 9017 10457
rect 9143 10423 9177 10457
rect 9303 10423 9337 10457
rect 9463 10423 9497 10457
rect 9623 10423 9657 10457
rect 9783 10423 9817 10457
rect 9943 10423 9977 10457
rect 10103 10423 10137 10457
rect 10263 10423 10297 10457
rect 10423 10423 10457 10457
rect 10583 10423 10617 10457
rect 10743 10423 10777 10457
rect 10903 10423 10937 10457
rect 11063 10423 11097 10457
rect 11223 10423 11257 10457
rect 11383 10423 11417 10457
rect 11543 10423 11577 10457
rect 11703 10423 11737 10457
rect 11863 10423 11897 10457
rect 12023 10423 12057 10457
rect 12183 10423 12217 10457
rect 12343 10423 12377 10457
rect 8503 10263 8537 10297
rect 8663 10263 8697 10297
rect 8823 10263 8857 10297
rect 8983 10263 9017 10297
rect 9143 10263 9177 10297
rect 9303 10263 9337 10297
rect 9463 10263 9497 10297
rect 9623 10263 9657 10297
rect 9783 10263 9817 10297
rect 9943 10263 9977 10297
rect 10103 10263 10137 10297
rect 10263 10263 10297 10297
rect 10423 10263 10457 10297
rect 10583 10263 10617 10297
rect 10743 10263 10777 10297
rect 10903 10263 10937 10297
rect 11063 10263 11097 10297
rect 11223 10263 11257 10297
rect 11383 10263 11417 10297
rect 11543 10263 11577 10297
rect 11703 10263 11737 10297
rect 11863 10263 11897 10297
rect 12023 10263 12057 10297
rect 12183 10263 12217 10297
rect 12343 10263 12377 10297
rect 8503 10103 8537 10137
rect 8663 10103 8697 10137
rect 8823 10103 8857 10137
rect 8983 10103 9017 10137
rect 9143 10103 9177 10137
rect 9303 10103 9337 10137
rect 9463 10103 9497 10137
rect 9623 10103 9657 10137
rect 9783 10103 9817 10137
rect 9943 10103 9977 10137
rect 10103 10103 10137 10137
rect 10263 10103 10297 10137
rect 10423 10103 10457 10137
rect 10583 10103 10617 10137
rect 10743 10103 10777 10137
rect 10903 10103 10937 10137
rect 11063 10103 11097 10137
rect 11223 10103 11257 10137
rect 11383 10103 11417 10137
rect 11543 10103 11577 10137
rect 11703 10103 11737 10137
rect 11863 10103 11897 10137
rect 12023 10103 12057 10137
rect 12183 10103 12217 10137
rect 12343 10103 12377 10137
rect 8503 9943 8537 9977
rect 8663 9943 8697 9977
rect 8823 9943 8857 9977
rect 8983 9943 9017 9977
rect 9143 9943 9177 9977
rect 9303 9943 9337 9977
rect 9463 9943 9497 9977
rect 9623 9943 9657 9977
rect 9783 9943 9817 9977
rect 9943 9943 9977 9977
rect 10103 9943 10137 9977
rect 10263 9943 10297 9977
rect 10423 9943 10457 9977
rect 10583 9943 10617 9977
rect 10743 9943 10777 9977
rect 10903 9943 10937 9977
rect 11063 9943 11097 9977
rect 11223 9943 11257 9977
rect 11383 9943 11417 9977
rect 11543 9943 11577 9977
rect 11703 9943 11737 9977
rect 11863 9943 11897 9977
rect 12023 9943 12057 9977
rect 12183 9943 12217 9977
rect 12343 9943 12377 9977
rect 8503 9783 8537 9817
rect 8663 9783 8697 9817
rect 8823 9783 8857 9817
rect 8983 9783 9017 9817
rect 9143 9783 9177 9817
rect 9303 9783 9337 9817
rect 9463 9783 9497 9817
rect 9623 9783 9657 9817
rect 9783 9783 9817 9817
rect 9943 9783 9977 9817
rect 10103 9783 10137 9817
rect 10263 9783 10297 9817
rect 10423 9783 10457 9817
rect 10583 9783 10617 9817
rect 10743 9783 10777 9817
rect 10903 9783 10937 9817
rect 11063 9783 11097 9817
rect 11223 9783 11257 9817
rect 11383 9783 11417 9817
rect 11543 9783 11577 9817
rect 11703 9783 11737 9817
rect 11863 9783 11897 9817
rect 12023 9783 12057 9817
rect 12183 9783 12217 9817
rect 12343 9783 12377 9817
rect 8503 9623 8537 9657
rect 8663 9623 8697 9657
rect 8823 9623 8857 9657
rect 8983 9623 9017 9657
rect 9143 9623 9177 9657
rect 9303 9623 9337 9657
rect 9463 9623 9497 9657
rect 9623 9623 9657 9657
rect 9783 9623 9817 9657
rect 9943 9623 9977 9657
rect 10103 9623 10137 9657
rect 10263 9623 10297 9657
rect 10423 9623 10457 9657
rect 10583 9623 10617 9657
rect 10743 9623 10777 9657
rect 10903 9623 10937 9657
rect 11063 9623 11097 9657
rect 11223 9623 11257 9657
rect 11383 9623 11417 9657
rect 11543 9623 11577 9657
rect 11703 9623 11737 9657
rect 11863 9623 11897 9657
rect 12023 9623 12057 9657
rect 12183 9623 12217 9657
rect 12343 9623 12377 9657
rect 8503 9463 8537 9497
rect 8663 9463 8697 9497
rect 8823 9463 8857 9497
rect 8983 9463 9017 9497
rect 9143 9463 9177 9497
rect 9303 9463 9337 9497
rect 9463 9463 9497 9497
rect 9623 9463 9657 9497
rect 9783 9463 9817 9497
rect 9943 9463 9977 9497
rect 10103 9463 10137 9497
rect 10263 9463 10297 9497
rect 10423 9463 10457 9497
rect 10583 9463 10617 9497
rect 10743 9463 10777 9497
rect 10903 9463 10937 9497
rect 11063 9463 11097 9497
rect 11223 9463 11257 9497
rect 11383 9463 11417 9497
rect 11543 9463 11577 9497
rect 11703 9463 11737 9497
rect 11863 9463 11897 9497
rect 12023 9463 12057 9497
rect 12183 9463 12217 9497
rect 12343 9463 12377 9497
rect 8503 9303 8537 9337
rect 8663 9303 8697 9337
rect 8823 9303 8857 9337
rect 8983 9303 9017 9337
rect 9143 9303 9177 9337
rect 9303 9303 9337 9337
rect 9463 9303 9497 9337
rect 9623 9303 9657 9337
rect 9783 9303 9817 9337
rect 9943 9303 9977 9337
rect 10103 9303 10137 9337
rect 10263 9303 10297 9337
rect 10423 9303 10457 9337
rect 10583 9303 10617 9337
rect 10743 9303 10777 9337
rect 10903 9303 10937 9337
rect 11063 9303 11097 9337
rect 11223 9303 11257 9337
rect 11383 9303 11417 9337
rect 11543 9303 11577 9337
rect 11703 9303 11737 9337
rect 11863 9303 11897 9337
rect 12023 9303 12057 9337
rect 12183 9303 12217 9337
rect 12343 9303 12377 9337
rect 8503 9143 8537 9177
rect 8663 9143 8697 9177
rect 8823 9143 8857 9177
rect 8983 9143 9017 9177
rect 9143 9143 9177 9177
rect 9303 9143 9337 9177
rect 9463 9143 9497 9177
rect 9623 9143 9657 9177
rect 9783 9143 9817 9177
rect 9943 9143 9977 9177
rect 10103 9143 10137 9177
rect 10263 9143 10297 9177
rect 10423 9143 10457 9177
rect 10583 9143 10617 9177
rect 10743 9143 10777 9177
rect 10903 9143 10937 9177
rect 11063 9143 11097 9177
rect 11223 9143 11257 9177
rect 11383 9143 11417 9177
rect 11543 9143 11577 9177
rect 11703 9143 11737 9177
rect 11863 9143 11897 9177
rect 12023 9143 12057 9177
rect 12183 9143 12217 9177
rect 12343 9143 12377 9177
rect 8503 8983 8537 9017
rect 8663 8983 8697 9017
rect 8823 8983 8857 9017
rect 8983 8983 9017 9017
rect 9143 8983 9177 9017
rect 9303 8983 9337 9017
rect 9463 8983 9497 9017
rect 9623 8983 9657 9017
rect 9783 8983 9817 9017
rect 9943 8983 9977 9017
rect 10103 8983 10137 9017
rect 10263 8983 10297 9017
rect 10423 8983 10457 9017
rect 10583 8983 10617 9017
rect 10743 8983 10777 9017
rect 10903 8983 10937 9017
rect 11063 8983 11097 9017
rect 11223 8983 11257 9017
rect 11383 8983 11417 9017
rect 11543 8983 11577 9017
rect 11703 8983 11737 9017
rect 11863 8983 11897 9017
rect 12023 8983 12057 9017
rect 12183 8983 12217 9017
rect 12343 8983 12377 9017
rect 8503 8823 8537 8857
rect 8663 8823 8697 8857
rect 8823 8823 8857 8857
rect 8983 8823 9017 8857
rect 9143 8823 9177 8857
rect 9303 8823 9337 8857
rect 9463 8823 9497 8857
rect 9623 8823 9657 8857
rect 9783 8823 9817 8857
rect 9943 8823 9977 8857
rect 10103 8823 10137 8857
rect 10263 8823 10297 8857
rect 10423 8823 10457 8857
rect 10583 8823 10617 8857
rect 10743 8823 10777 8857
rect 10903 8823 10937 8857
rect 11063 8823 11097 8857
rect 11223 8823 11257 8857
rect 11383 8823 11417 8857
rect 11543 8823 11577 8857
rect 11703 8823 11737 8857
rect 11863 8823 11897 8857
rect 12023 8823 12057 8857
rect 12183 8823 12217 8857
rect 12343 8823 12377 8857
rect 8503 8663 8537 8697
rect 8663 8663 8697 8697
rect 8823 8663 8857 8697
rect 8983 8663 9017 8697
rect 9143 8663 9177 8697
rect 9303 8663 9337 8697
rect 9463 8663 9497 8697
rect 9623 8663 9657 8697
rect 9783 8663 9817 8697
rect 9943 8663 9977 8697
rect 10103 8663 10137 8697
rect 10263 8663 10297 8697
rect 10423 8663 10457 8697
rect 10583 8663 10617 8697
rect 10743 8663 10777 8697
rect 10903 8663 10937 8697
rect 11063 8663 11097 8697
rect 11223 8663 11257 8697
rect 11383 8663 11417 8697
rect 11543 8663 11577 8697
rect 11703 8663 11737 8697
rect 11863 8663 11897 8697
rect 12023 8663 12057 8697
rect 12183 8663 12217 8697
rect 12343 8663 12377 8697
rect 8503 8503 8537 8537
rect 8663 8503 8697 8537
rect 8823 8503 8857 8537
rect 8983 8503 9017 8537
rect 9143 8503 9177 8537
rect 9303 8503 9337 8537
rect 9463 8503 9497 8537
rect 9623 8503 9657 8537
rect 9783 8503 9817 8537
rect 9943 8503 9977 8537
rect 10103 8503 10137 8537
rect 10263 8503 10297 8537
rect 10423 8503 10457 8537
rect 10583 8503 10617 8537
rect 10743 8503 10777 8537
rect 10903 8503 10937 8537
rect 11063 8503 11097 8537
rect 11223 8503 11257 8537
rect 11383 8503 11417 8537
rect 11543 8503 11577 8537
rect 11703 8503 11737 8537
rect 11863 8503 11897 8537
rect 12023 8503 12057 8537
rect 12183 8503 12217 8537
rect 12343 8503 12377 8537
rect 8503 8343 8537 8377
rect 8663 8343 8697 8377
rect 8823 8343 8857 8377
rect 8983 8343 9017 8377
rect 9143 8343 9177 8377
rect 9303 8343 9337 8377
rect 9463 8343 9497 8377
rect 9623 8343 9657 8377
rect 9783 8343 9817 8377
rect 9943 8343 9977 8377
rect 10103 8343 10137 8377
rect 10263 8343 10297 8377
rect 10423 8343 10457 8377
rect 10583 8343 10617 8377
rect 10743 8343 10777 8377
rect 10903 8343 10937 8377
rect 11063 8343 11097 8377
rect 11223 8343 11257 8377
rect 11383 8343 11417 8377
rect 11543 8343 11577 8377
rect 11703 8343 11737 8377
rect 11863 8343 11897 8377
rect 12023 8343 12057 8377
rect 12183 8343 12217 8377
rect 12343 8343 12377 8377
rect 8503 8183 8537 8217
rect 8663 8183 8697 8217
rect 8823 8183 8857 8217
rect 8983 8183 9017 8217
rect 9143 8183 9177 8217
rect 9303 8183 9337 8217
rect 9463 8183 9497 8217
rect 9623 8183 9657 8217
rect 9783 8183 9817 8217
rect 9943 8183 9977 8217
rect 10103 8183 10137 8217
rect 10263 8183 10297 8217
rect 10423 8183 10457 8217
rect 10583 8183 10617 8217
rect 10743 8183 10777 8217
rect 10903 8183 10937 8217
rect 11063 8183 11097 8217
rect 11223 8183 11257 8217
rect 11383 8183 11417 8217
rect 11543 8183 11577 8217
rect 11703 8183 11737 8217
rect 11863 8183 11897 8217
rect 12023 8183 12057 8217
rect 12183 8183 12217 8217
rect 12343 8183 12377 8217
rect 8503 8023 8537 8057
rect 8663 8023 8697 8057
rect 8823 8023 8857 8057
rect 8983 8023 9017 8057
rect 9143 8023 9177 8057
rect 9303 8023 9337 8057
rect 9463 8023 9497 8057
rect 9623 8023 9657 8057
rect 9783 8023 9817 8057
rect 9943 8023 9977 8057
rect 10103 8023 10137 8057
rect 10263 8023 10297 8057
rect 10423 8023 10457 8057
rect 10583 8023 10617 8057
rect 10743 8023 10777 8057
rect 10903 8023 10937 8057
rect 11063 8023 11097 8057
rect 11223 8023 11257 8057
rect 11383 8023 11417 8057
rect 11543 8023 11577 8057
rect 11703 8023 11737 8057
rect 11863 8023 11897 8057
rect 12023 8023 12057 8057
rect 12183 8023 12217 8057
rect 12343 8023 12377 8057
rect 8503 7863 8537 7897
rect 8663 7863 8697 7897
rect 8823 7863 8857 7897
rect 8983 7863 9017 7897
rect 9143 7863 9177 7897
rect 9303 7863 9337 7897
rect 9463 7863 9497 7897
rect 9623 7863 9657 7897
rect 9783 7863 9817 7897
rect 9943 7863 9977 7897
rect 10103 7863 10137 7897
rect 10263 7863 10297 7897
rect 10423 7863 10457 7897
rect 10583 7863 10617 7897
rect 10743 7863 10777 7897
rect 10903 7863 10937 7897
rect 11063 7863 11097 7897
rect 11223 7863 11257 7897
rect 11383 7863 11417 7897
rect 11543 7863 11577 7897
rect 11703 7863 11737 7897
rect 11863 7863 11897 7897
rect 12023 7863 12057 7897
rect 12183 7863 12217 7897
rect 12343 7863 12377 7897
rect 8503 7703 8537 7737
rect 8663 7703 8697 7737
rect 8823 7703 8857 7737
rect 8983 7703 9017 7737
rect 9143 7703 9177 7737
rect 9303 7703 9337 7737
rect 9463 7703 9497 7737
rect 9623 7703 9657 7737
rect 9783 7703 9817 7737
rect 9943 7703 9977 7737
rect 10103 7703 10137 7737
rect 10263 7703 10297 7737
rect 10423 7703 10457 7737
rect 10583 7703 10617 7737
rect 10743 7703 10777 7737
rect 10903 7703 10937 7737
rect 11063 7703 11097 7737
rect 11223 7703 11257 7737
rect 11383 7703 11417 7737
rect 11543 7703 11577 7737
rect 11703 7703 11737 7737
rect 11863 7703 11897 7737
rect 12023 7703 12057 7737
rect 12183 7703 12217 7737
rect 12343 7703 12377 7737
rect 8503 7543 8537 7577
rect 8663 7543 8697 7577
rect 8823 7543 8857 7577
rect 8983 7543 9017 7577
rect 9143 7543 9177 7577
rect 9303 7543 9337 7577
rect 9463 7543 9497 7577
rect 9623 7543 9657 7577
rect 9783 7543 9817 7577
rect 9943 7543 9977 7577
rect 10103 7543 10137 7577
rect 10263 7543 10297 7577
rect 10423 7543 10457 7577
rect 10583 7543 10617 7577
rect 10743 7543 10777 7577
rect 10903 7543 10937 7577
rect 11063 7543 11097 7577
rect 11223 7543 11257 7577
rect 11383 7543 11417 7577
rect 11543 7543 11577 7577
rect 11703 7543 11737 7577
rect 11863 7543 11897 7577
rect 12023 7543 12057 7577
rect 12183 7543 12217 7577
rect 12343 7543 12377 7577
rect 8503 7383 8537 7417
rect 8663 7383 8697 7417
rect 8823 7383 8857 7417
rect 8983 7383 9017 7417
rect 9143 7383 9177 7417
rect 9303 7383 9337 7417
rect 9463 7383 9497 7417
rect 9623 7383 9657 7417
rect 9783 7383 9817 7417
rect 9943 7383 9977 7417
rect 10103 7383 10137 7417
rect 10263 7383 10297 7417
rect 10423 7383 10457 7417
rect 10583 7383 10617 7417
rect 10743 7383 10777 7417
rect 10903 7383 10937 7417
rect 11063 7383 11097 7417
rect 11223 7383 11257 7417
rect 11383 7383 11417 7417
rect 11543 7383 11577 7417
rect 11703 7383 11737 7417
rect 11863 7383 11897 7417
rect 12023 7383 12057 7417
rect 12183 7383 12217 7417
rect 12343 7383 12377 7417
rect 8503 7223 8537 7257
rect 8663 7223 8697 7257
rect 8823 7223 8857 7257
rect 8983 7223 9017 7257
rect 9143 7223 9177 7257
rect 9303 7223 9337 7257
rect 9463 7223 9497 7257
rect 9623 7223 9657 7257
rect 9783 7223 9817 7257
rect 9943 7223 9977 7257
rect 10103 7223 10137 7257
rect 10263 7223 10297 7257
rect 10423 7223 10457 7257
rect 10583 7223 10617 7257
rect 10743 7223 10777 7257
rect 10903 7223 10937 7257
rect 11063 7223 11097 7257
rect 11223 7223 11257 7257
rect 11383 7223 11417 7257
rect 11543 7223 11577 7257
rect 11703 7223 11737 7257
rect 11863 7223 11897 7257
rect 12023 7223 12057 7257
rect 12183 7223 12217 7257
rect 12343 7223 12377 7257
rect 8503 7063 8537 7097
rect 8663 7063 8697 7097
rect 8823 7063 8857 7097
rect 8983 7063 9017 7097
rect 9143 7063 9177 7097
rect 9303 7063 9337 7097
rect 9463 7063 9497 7097
rect 9623 7063 9657 7097
rect 9783 7063 9817 7097
rect 9943 7063 9977 7097
rect 10103 7063 10137 7097
rect 10263 7063 10297 7097
rect 10423 7063 10457 7097
rect 10583 7063 10617 7097
rect 10743 7063 10777 7097
rect 10903 7063 10937 7097
rect 11063 7063 11097 7097
rect 11223 7063 11257 7097
rect 11383 7063 11417 7097
rect 11543 7063 11577 7097
rect 11703 7063 11737 7097
rect 11863 7063 11897 7097
rect 12023 7063 12057 7097
rect 12183 7063 12217 7097
rect 12343 7063 12377 7097
rect 8503 6903 8537 6937
rect 8663 6903 8697 6937
rect 8823 6903 8857 6937
rect 8983 6903 9017 6937
rect 9143 6903 9177 6937
rect 9303 6903 9337 6937
rect 9463 6903 9497 6937
rect 9623 6903 9657 6937
rect 9783 6903 9817 6937
rect 9943 6903 9977 6937
rect 10103 6903 10137 6937
rect 10263 6903 10297 6937
rect 10423 6903 10457 6937
rect 10583 6903 10617 6937
rect 10743 6903 10777 6937
rect 10903 6903 10937 6937
rect 11063 6903 11097 6937
rect 11223 6903 11257 6937
rect 11383 6903 11417 6937
rect 11543 6903 11577 6937
rect 11703 6903 11737 6937
rect 11863 6903 11897 6937
rect 12023 6903 12057 6937
rect 12183 6903 12217 6937
rect 12343 6903 12377 6937
rect 8503 6743 8537 6777
rect 8663 6743 8697 6777
rect 8823 6743 8857 6777
rect 8983 6743 9017 6777
rect 9143 6743 9177 6777
rect 9303 6743 9337 6777
rect 9463 6743 9497 6777
rect 9623 6743 9657 6777
rect 9783 6743 9817 6777
rect 9943 6743 9977 6777
rect 10103 6743 10137 6777
rect 10263 6743 10297 6777
rect 10423 6743 10457 6777
rect 10583 6743 10617 6777
rect 10743 6743 10777 6777
rect 10903 6743 10937 6777
rect 11063 6743 11097 6777
rect 11223 6743 11257 6777
rect 11383 6743 11417 6777
rect 11543 6743 11577 6777
rect 11703 6743 11737 6777
rect 11863 6743 11897 6777
rect 12023 6743 12057 6777
rect 12183 6743 12217 6777
rect 12343 6743 12377 6777
rect 8503 6583 8537 6617
rect 8663 6583 8697 6617
rect 8823 6583 8857 6617
rect 8983 6583 9017 6617
rect 9143 6583 9177 6617
rect 9303 6583 9337 6617
rect 9463 6583 9497 6617
rect 9623 6583 9657 6617
rect 9783 6583 9817 6617
rect 9943 6583 9977 6617
rect 10103 6583 10137 6617
rect 10263 6583 10297 6617
rect 10423 6583 10457 6617
rect 10583 6583 10617 6617
rect 10743 6583 10777 6617
rect 10903 6583 10937 6617
rect 11063 6583 11097 6617
rect 11223 6583 11257 6617
rect 11383 6583 11417 6617
rect 11543 6583 11577 6617
rect 11703 6583 11737 6617
rect 11863 6583 11897 6617
rect 12023 6583 12057 6617
rect 12183 6583 12217 6617
rect 12343 6583 12377 6617
rect 8503 6423 8537 6457
rect 8663 6423 8697 6457
rect 8823 6423 8857 6457
rect 8983 6423 9017 6457
rect 9143 6423 9177 6457
rect 9303 6423 9337 6457
rect 9463 6423 9497 6457
rect 9623 6423 9657 6457
rect 9783 6423 9817 6457
rect 9943 6423 9977 6457
rect 10103 6423 10137 6457
rect 10263 6423 10297 6457
rect 10423 6423 10457 6457
rect 10583 6423 10617 6457
rect 10743 6423 10777 6457
rect 10903 6423 10937 6457
rect 11063 6423 11097 6457
rect 11223 6423 11257 6457
rect 11383 6423 11417 6457
rect 11543 6423 11577 6457
rect 11703 6423 11737 6457
rect 11863 6423 11897 6457
rect 12023 6423 12057 6457
rect 12183 6423 12217 6457
rect 12343 6423 12377 6457
rect 8503 6263 8537 6297
rect 8663 6263 8697 6297
rect 8823 6263 8857 6297
rect 8983 6263 9017 6297
rect 9143 6263 9177 6297
rect 9303 6263 9337 6297
rect 9463 6263 9497 6297
rect 9623 6263 9657 6297
rect 9783 6263 9817 6297
rect 9943 6263 9977 6297
rect 10103 6263 10137 6297
rect 10263 6263 10297 6297
rect 10423 6263 10457 6297
rect 10583 6263 10617 6297
rect 10743 6263 10777 6297
rect 10903 6263 10937 6297
rect 11063 6263 11097 6297
rect 11223 6263 11257 6297
rect 11383 6263 11417 6297
rect 11543 6263 11577 6297
rect 11703 6263 11737 6297
rect 11863 6263 11897 6297
rect 12023 6263 12057 6297
rect 12183 6263 12217 6297
rect 12343 6263 12377 6297
rect 8503 6103 8537 6137
rect 8663 6103 8697 6137
rect 8823 6103 8857 6137
rect 8983 6103 9017 6137
rect 9143 6103 9177 6137
rect 9303 6103 9337 6137
rect 9463 6103 9497 6137
rect 9623 6103 9657 6137
rect 9783 6103 9817 6137
rect 9943 6103 9977 6137
rect 10103 6103 10137 6137
rect 10263 6103 10297 6137
rect 10423 6103 10457 6137
rect 10583 6103 10617 6137
rect 10743 6103 10777 6137
rect 10903 6103 10937 6137
rect 11063 6103 11097 6137
rect 11223 6103 11257 6137
rect 11383 6103 11417 6137
rect 11543 6103 11577 6137
rect 11703 6103 11737 6137
rect 11863 6103 11897 6137
rect 12023 6103 12057 6137
rect 12183 6103 12217 6137
rect 12343 6103 12377 6137
rect 8503 5943 8537 5977
rect 8663 5943 8697 5977
rect 8823 5943 8857 5977
rect 8983 5943 9017 5977
rect 9143 5943 9177 5977
rect 9303 5943 9337 5977
rect 9463 5943 9497 5977
rect 9623 5943 9657 5977
rect 9783 5943 9817 5977
rect 9943 5943 9977 5977
rect 10103 5943 10137 5977
rect 10263 5943 10297 5977
rect 10423 5943 10457 5977
rect 10583 5943 10617 5977
rect 10743 5943 10777 5977
rect 10903 5943 10937 5977
rect 11063 5943 11097 5977
rect 11223 5943 11257 5977
rect 11383 5943 11417 5977
rect 11543 5943 11577 5977
rect 11703 5943 11737 5977
rect 11863 5943 11897 5977
rect 12023 5943 12057 5977
rect 12183 5943 12217 5977
rect 12343 5943 12377 5977
rect 8503 5783 8537 5817
rect 8663 5783 8697 5817
rect 8823 5783 8857 5817
rect 8983 5783 9017 5817
rect 9143 5783 9177 5817
rect 9303 5783 9337 5817
rect 9463 5783 9497 5817
rect 9623 5783 9657 5817
rect 9783 5783 9817 5817
rect 9943 5783 9977 5817
rect 10103 5783 10137 5817
rect 10263 5783 10297 5817
rect 10423 5783 10457 5817
rect 10583 5783 10617 5817
rect 10743 5783 10777 5817
rect 10903 5783 10937 5817
rect 11063 5783 11097 5817
rect 11223 5783 11257 5817
rect 11383 5783 11417 5817
rect 11543 5783 11577 5817
rect 11703 5783 11737 5817
rect 11863 5783 11897 5817
rect 12023 5783 12057 5817
rect 12183 5783 12217 5817
rect 12343 5783 12377 5817
rect 8503 5623 8537 5657
rect 8663 5623 8697 5657
rect 8823 5623 8857 5657
rect 8983 5623 9017 5657
rect 9143 5623 9177 5657
rect 9303 5623 9337 5657
rect 9463 5623 9497 5657
rect 9623 5623 9657 5657
rect 9783 5623 9817 5657
rect 9943 5623 9977 5657
rect 10103 5623 10137 5657
rect 10263 5623 10297 5657
rect 10423 5623 10457 5657
rect 10583 5623 10617 5657
rect 10743 5623 10777 5657
rect 10903 5623 10937 5657
rect 11063 5623 11097 5657
rect 11223 5623 11257 5657
rect 11383 5623 11417 5657
rect 11543 5623 11577 5657
rect 11703 5623 11737 5657
rect 11863 5623 11897 5657
rect 12023 5623 12057 5657
rect 12183 5623 12217 5657
rect 12343 5623 12377 5657
rect 8503 5463 8537 5497
rect 8663 5463 8697 5497
rect 8823 5463 8857 5497
rect 8983 5463 9017 5497
rect 9143 5463 9177 5497
rect 9303 5463 9337 5497
rect 9463 5463 9497 5497
rect 9623 5463 9657 5497
rect 9783 5463 9817 5497
rect 9943 5463 9977 5497
rect 10103 5463 10137 5497
rect 10263 5463 10297 5497
rect 10423 5463 10457 5497
rect 10583 5463 10617 5497
rect 10743 5463 10777 5497
rect 10903 5463 10937 5497
rect 11063 5463 11097 5497
rect 11223 5463 11257 5497
rect 11383 5463 11417 5497
rect 11543 5463 11577 5497
rect 11703 5463 11737 5497
rect 11863 5463 11897 5497
rect 12023 5463 12057 5497
rect 12183 5463 12217 5497
rect 12343 5463 12377 5497
rect 8503 5303 8537 5337
rect 8663 5303 8697 5337
rect 8823 5303 8857 5337
rect 8983 5303 9017 5337
rect 9143 5303 9177 5337
rect 9303 5303 9337 5337
rect 9463 5303 9497 5337
rect 9623 5303 9657 5337
rect 9783 5303 9817 5337
rect 9943 5303 9977 5337
rect 10103 5303 10137 5337
rect 10263 5303 10297 5337
rect 10423 5303 10457 5337
rect 10583 5303 10617 5337
rect 10743 5303 10777 5337
rect 10903 5303 10937 5337
rect 11063 5303 11097 5337
rect 11223 5303 11257 5337
rect 11383 5303 11417 5337
rect 11543 5303 11577 5337
rect 11703 5303 11737 5337
rect 11863 5303 11897 5337
rect 12023 5303 12057 5337
rect 12183 5303 12217 5337
rect 12343 5303 12377 5337
rect 8503 5143 8537 5177
rect 8663 5143 8697 5177
rect 8823 5143 8857 5177
rect 8983 5143 9017 5177
rect 9143 5143 9177 5177
rect 9303 5143 9337 5177
rect 9463 5143 9497 5177
rect 9623 5143 9657 5177
rect 9783 5143 9817 5177
rect 9943 5143 9977 5177
rect 10103 5143 10137 5177
rect 10263 5143 10297 5177
rect 10423 5143 10457 5177
rect 10583 5143 10617 5177
rect 10743 5143 10777 5177
rect 10903 5143 10937 5177
rect 11063 5143 11097 5177
rect 11223 5143 11257 5177
rect 11383 5143 11417 5177
rect 11543 5143 11577 5177
rect 11703 5143 11737 5177
rect 11863 5143 11897 5177
rect 12023 5143 12057 5177
rect 12183 5143 12217 5177
rect 12343 5143 12377 5177
rect 8503 4983 8537 5017
rect 8663 4983 8697 5017
rect 8823 4983 8857 5017
rect 8983 4983 9017 5017
rect 9143 4983 9177 5017
rect 9303 4983 9337 5017
rect 9463 4983 9497 5017
rect 9623 4983 9657 5017
rect 9783 4983 9817 5017
rect 9943 4983 9977 5017
rect 10103 4983 10137 5017
rect 10263 4983 10297 5017
rect 10423 4983 10457 5017
rect 10583 4983 10617 5017
rect 10743 4983 10777 5017
rect 10903 4983 10937 5017
rect 11063 4983 11097 5017
rect 11223 4983 11257 5017
rect 11383 4983 11417 5017
rect 11543 4983 11577 5017
rect 11703 4983 11737 5017
rect 11863 4983 11897 5017
rect 12023 4983 12057 5017
rect 12183 4983 12217 5017
rect 12343 4983 12377 5017
rect 8503 4823 8537 4857
rect 8663 4823 8697 4857
rect 8823 4823 8857 4857
rect 8983 4823 9017 4857
rect 9143 4823 9177 4857
rect 9303 4823 9337 4857
rect 9463 4823 9497 4857
rect 9623 4823 9657 4857
rect 9783 4823 9817 4857
rect 9943 4823 9977 4857
rect 10103 4823 10137 4857
rect 10263 4823 10297 4857
rect 10423 4823 10457 4857
rect 10583 4823 10617 4857
rect 10743 4823 10777 4857
rect 10903 4823 10937 4857
rect 11063 4823 11097 4857
rect 11223 4823 11257 4857
rect 11383 4823 11417 4857
rect 11543 4823 11577 4857
rect 11703 4823 11737 4857
rect 11863 4823 11897 4857
rect 12023 4823 12057 4857
rect 12183 4823 12217 4857
rect 12343 4823 12377 4857
rect 8503 4663 8537 4697
rect 8663 4663 8697 4697
rect 8823 4663 8857 4697
rect 8983 4663 9017 4697
rect 9143 4663 9177 4697
rect 9303 4663 9337 4697
rect 9463 4663 9497 4697
rect 9623 4663 9657 4697
rect 9783 4663 9817 4697
rect 9943 4663 9977 4697
rect 10103 4663 10137 4697
rect 10263 4663 10297 4697
rect 10423 4663 10457 4697
rect 10583 4663 10617 4697
rect 10743 4663 10777 4697
rect 10903 4663 10937 4697
rect 11063 4663 11097 4697
rect 11223 4663 11257 4697
rect 11383 4663 11417 4697
rect 11543 4663 11577 4697
rect 11703 4663 11737 4697
rect 11863 4663 11897 4697
rect 12023 4663 12057 4697
rect 12183 4663 12217 4697
rect 12343 4663 12377 4697
rect 8503 4503 8537 4537
rect 8663 4503 8697 4537
rect 8823 4503 8857 4537
rect 8983 4503 9017 4537
rect 9143 4503 9177 4537
rect 9303 4503 9337 4537
rect 9463 4503 9497 4537
rect 9623 4503 9657 4537
rect 9783 4503 9817 4537
rect 9943 4503 9977 4537
rect 10103 4503 10137 4537
rect 10263 4503 10297 4537
rect 10423 4503 10457 4537
rect 10583 4503 10617 4537
rect 10743 4503 10777 4537
rect 10903 4503 10937 4537
rect 11063 4503 11097 4537
rect 11223 4503 11257 4537
rect 11383 4503 11417 4537
rect 11543 4503 11577 4537
rect 11703 4503 11737 4537
rect 11863 4503 11897 4537
rect 12023 4503 12057 4537
rect 12183 4503 12217 4537
rect 12343 4503 12377 4537
rect 8503 4343 8537 4377
rect 8663 4343 8697 4377
rect 8823 4343 8857 4377
rect 8983 4343 9017 4377
rect 9143 4343 9177 4377
rect 9303 4343 9337 4377
rect 9463 4343 9497 4377
rect 9623 4343 9657 4377
rect 9783 4343 9817 4377
rect 9943 4343 9977 4377
rect 10103 4343 10137 4377
rect 10263 4343 10297 4377
rect 10423 4343 10457 4377
rect 10583 4343 10617 4377
rect 10743 4343 10777 4377
rect 10903 4343 10937 4377
rect 11063 4343 11097 4377
rect 11223 4343 11257 4377
rect 11383 4343 11417 4377
rect 11543 4343 11577 4377
rect 11703 4343 11737 4377
rect 11863 4343 11897 4377
rect 12023 4343 12057 4377
rect 12183 4343 12217 4377
rect 12343 4343 12377 4377
rect 8503 4183 8537 4217
rect 8663 4183 8697 4217
rect 8823 4183 8857 4217
rect 8983 4183 9017 4217
rect 9143 4183 9177 4217
rect 9303 4183 9337 4217
rect 9463 4183 9497 4217
rect 9623 4183 9657 4217
rect 9783 4183 9817 4217
rect 9943 4183 9977 4217
rect 10103 4183 10137 4217
rect 10263 4183 10297 4217
rect 10423 4183 10457 4217
rect 10583 4183 10617 4217
rect 10743 4183 10777 4217
rect 10903 4183 10937 4217
rect 11063 4183 11097 4217
rect 11223 4183 11257 4217
rect 11383 4183 11417 4217
rect 11543 4183 11577 4217
rect 11703 4183 11737 4217
rect 11863 4183 11897 4217
rect 12023 4183 12057 4217
rect 12183 4183 12217 4217
rect 12343 4183 12377 4217
rect 8503 4023 8537 4057
rect 8663 4023 8697 4057
rect 8823 4023 8857 4057
rect 8983 4023 9017 4057
rect 9143 4023 9177 4057
rect 9303 4023 9337 4057
rect 9463 4023 9497 4057
rect 9623 4023 9657 4057
rect 9783 4023 9817 4057
rect 9943 4023 9977 4057
rect 10103 4023 10137 4057
rect 10263 4023 10297 4057
rect 10423 4023 10457 4057
rect 10583 4023 10617 4057
rect 10743 4023 10777 4057
rect 10903 4023 10937 4057
rect 11063 4023 11097 4057
rect 11223 4023 11257 4057
rect 11383 4023 11417 4057
rect 11543 4023 11577 4057
rect 11703 4023 11737 4057
rect 11863 4023 11897 4057
rect 12023 4023 12057 4057
rect 12183 4023 12217 4057
rect 12343 4023 12377 4057
rect 8503 3863 8537 3897
rect 8663 3863 8697 3897
rect 8823 3863 8857 3897
rect 8983 3863 9017 3897
rect 9143 3863 9177 3897
rect 9303 3863 9337 3897
rect 9463 3863 9497 3897
rect 9623 3863 9657 3897
rect 9783 3863 9817 3897
rect 9943 3863 9977 3897
rect 10103 3863 10137 3897
rect 10263 3863 10297 3897
rect 10423 3863 10457 3897
rect 10583 3863 10617 3897
rect 10743 3863 10777 3897
rect 10903 3863 10937 3897
rect 11063 3863 11097 3897
rect 11223 3863 11257 3897
rect 11383 3863 11417 3897
rect 11543 3863 11577 3897
rect 11703 3863 11737 3897
rect 11863 3863 11897 3897
rect 12023 3863 12057 3897
rect 12183 3863 12217 3897
rect 12343 3863 12377 3897
rect 8503 3703 8537 3737
rect 8663 3703 8697 3737
rect 8823 3703 8857 3737
rect 8983 3703 9017 3737
rect 9143 3703 9177 3737
rect 9303 3703 9337 3737
rect 9463 3703 9497 3737
rect 9623 3703 9657 3737
rect 9783 3703 9817 3737
rect 9943 3703 9977 3737
rect 10103 3703 10137 3737
rect 10263 3703 10297 3737
rect 10423 3703 10457 3737
rect 10583 3703 10617 3737
rect 10743 3703 10777 3737
rect 10903 3703 10937 3737
rect 11063 3703 11097 3737
rect 11223 3703 11257 3737
rect 11383 3703 11417 3737
rect 11543 3703 11577 3737
rect 11703 3703 11737 3737
rect 11863 3703 11897 3737
rect 12023 3703 12057 3737
rect 12183 3703 12217 3737
rect 12343 3703 12377 3737
rect 8503 3543 8537 3577
rect 8663 3543 8697 3577
rect 8823 3543 8857 3577
rect 8983 3543 9017 3577
rect 9143 3543 9177 3577
rect 9303 3543 9337 3577
rect 9463 3543 9497 3577
rect 9623 3543 9657 3577
rect 9783 3543 9817 3577
rect 9943 3543 9977 3577
rect 10103 3543 10137 3577
rect 10263 3543 10297 3577
rect 10423 3543 10457 3577
rect 10583 3543 10617 3577
rect 10743 3543 10777 3577
rect 10903 3543 10937 3577
rect 11063 3543 11097 3577
rect 11223 3543 11257 3577
rect 11383 3543 11417 3577
rect 11543 3543 11577 3577
rect 11703 3543 11737 3577
rect 11863 3543 11897 3577
rect 12023 3543 12057 3577
rect 12183 3543 12217 3577
rect 12343 3543 12377 3577
rect 8503 3383 8537 3417
rect 8663 3383 8697 3417
rect 8823 3383 8857 3417
rect 8983 3383 9017 3417
rect 9143 3383 9177 3417
rect 9303 3383 9337 3417
rect 9463 3383 9497 3417
rect 9623 3383 9657 3417
rect 9783 3383 9817 3417
rect 9943 3383 9977 3417
rect 10103 3383 10137 3417
rect 10263 3383 10297 3417
rect 10423 3383 10457 3417
rect 10583 3383 10617 3417
rect 10743 3383 10777 3417
rect 10903 3383 10937 3417
rect 11063 3383 11097 3417
rect 11223 3383 11257 3417
rect 11383 3383 11417 3417
rect 11543 3383 11577 3417
rect 11703 3383 11737 3417
rect 11863 3383 11897 3417
rect 12023 3383 12057 3417
rect 12183 3383 12217 3417
rect 12343 3383 12377 3417
rect 8503 3223 8537 3257
rect 8663 3223 8697 3257
rect 8823 3223 8857 3257
rect 8983 3223 9017 3257
rect 9143 3223 9177 3257
rect 9303 3223 9337 3257
rect 9463 3223 9497 3257
rect 9623 3223 9657 3257
rect 9783 3223 9817 3257
rect 9943 3223 9977 3257
rect 10103 3223 10137 3257
rect 10263 3223 10297 3257
rect 10423 3223 10457 3257
rect 10583 3223 10617 3257
rect 10743 3223 10777 3257
rect 10903 3223 10937 3257
rect 11063 3223 11097 3257
rect 11223 3223 11257 3257
rect 11383 3223 11417 3257
rect 11543 3223 11577 3257
rect 11703 3223 11737 3257
rect 11863 3223 11897 3257
rect 12023 3223 12057 3257
rect 12183 3223 12217 3257
rect 12343 3223 12377 3257
rect 8503 3063 8537 3097
rect 8663 3063 8697 3097
rect 8823 3063 8857 3097
rect 8983 3063 9017 3097
rect 9143 3063 9177 3097
rect 9303 3063 9337 3097
rect 9463 3063 9497 3097
rect 9623 3063 9657 3097
rect 9783 3063 9817 3097
rect 9943 3063 9977 3097
rect 10103 3063 10137 3097
rect 10263 3063 10297 3097
rect 10423 3063 10457 3097
rect 10583 3063 10617 3097
rect 10743 3063 10777 3097
rect 10903 3063 10937 3097
rect 11063 3063 11097 3097
rect 11223 3063 11257 3097
rect 11383 3063 11417 3097
rect 11543 3063 11577 3097
rect 11703 3063 11737 3097
rect 11863 3063 11897 3097
rect 12023 3063 12057 3097
rect 12183 3063 12217 3097
rect 12343 3063 12377 3097
rect 8503 2903 8537 2937
rect 8663 2903 8697 2937
rect 8823 2903 8857 2937
rect 8983 2903 9017 2937
rect 9143 2903 9177 2937
rect 9303 2903 9337 2937
rect 9463 2903 9497 2937
rect 9623 2903 9657 2937
rect 9783 2903 9817 2937
rect 9943 2903 9977 2937
rect 10103 2903 10137 2937
rect 10263 2903 10297 2937
rect 10423 2903 10457 2937
rect 10583 2903 10617 2937
rect 10743 2903 10777 2937
rect 10903 2903 10937 2937
rect 11063 2903 11097 2937
rect 11223 2903 11257 2937
rect 11383 2903 11417 2937
rect 11543 2903 11577 2937
rect 11703 2903 11737 2937
rect 11863 2903 11897 2937
rect 12023 2903 12057 2937
rect 12183 2903 12217 2937
rect 12343 2903 12377 2937
rect 8503 2743 8537 2777
rect 8663 2743 8697 2777
rect 8823 2743 8857 2777
rect 8983 2743 9017 2777
rect 9143 2743 9177 2777
rect 9303 2743 9337 2777
rect 9463 2743 9497 2777
rect 9623 2743 9657 2777
rect 9783 2743 9817 2777
rect 9943 2743 9977 2777
rect 10103 2743 10137 2777
rect 10263 2743 10297 2777
rect 10423 2743 10457 2777
rect 10583 2743 10617 2777
rect 10743 2743 10777 2777
rect 10903 2743 10937 2777
rect 11063 2743 11097 2777
rect 11223 2743 11257 2777
rect 11383 2743 11417 2777
rect 11543 2743 11577 2777
rect 11703 2743 11737 2777
rect 11863 2743 11897 2777
rect 12023 2743 12057 2777
rect 12183 2743 12217 2777
rect 12343 2743 12377 2777
rect 8503 2583 8537 2617
rect 8663 2583 8697 2617
rect 8823 2583 8857 2617
rect 8983 2583 9017 2617
rect 9143 2583 9177 2617
rect 9303 2583 9337 2617
rect 9463 2583 9497 2617
rect 9623 2583 9657 2617
rect 9783 2583 9817 2617
rect 9943 2583 9977 2617
rect 10103 2583 10137 2617
rect 10263 2583 10297 2617
rect 10423 2583 10457 2617
rect 10583 2583 10617 2617
rect 10743 2583 10777 2617
rect 10903 2583 10937 2617
rect 11063 2583 11097 2617
rect 11223 2583 11257 2617
rect 11383 2583 11417 2617
rect 11543 2583 11577 2617
rect 11703 2583 11737 2617
rect 11863 2583 11897 2617
rect 12023 2583 12057 2617
rect 12183 2583 12217 2617
rect 12343 2583 12377 2617
rect 8503 2423 8537 2457
rect 8663 2423 8697 2457
rect 8823 2423 8857 2457
rect 8983 2423 9017 2457
rect 9143 2423 9177 2457
rect 9303 2423 9337 2457
rect 9463 2423 9497 2457
rect 9623 2423 9657 2457
rect 9783 2423 9817 2457
rect 9943 2423 9977 2457
rect 10103 2423 10137 2457
rect 10263 2423 10297 2457
rect 10423 2423 10457 2457
rect 10583 2423 10617 2457
rect 10743 2423 10777 2457
rect 10903 2423 10937 2457
rect 11063 2423 11097 2457
rect 11223 2423 11257 2457
rect 11383 2423 11417 2457
rect 11543 2423 11577 2457
rect 11703 2423 11737 2457
rect 11863 2423 11897 2457
rect 12023 2423 12057 2457
rect 12183 2423 12217 2457
rect 12343 2423 12377 2457
rect 8503 2263 8537 2297
rect 8663 2263 8697 2297
rect 8823 2263 8857 2297
rect 8983 2263 9017 2297
rect 9143 2263 9177 2297
rect 9303 2263 9337 2297
rect 9463 2263 9497 2297
rect 9623 2263 9657 2297
rect 9783 2263 9817 2297
rect 9943 2263 9977 2297
rect 10103 2263 10137 2297
rect 10263 2263 10297 2297
rect 10423 2263 10457 2297
rect 10583 2263 10617 2297
rect 10743 2263 10777 2297
rect 10903 2263 10937 2297
rect 11063 2263 11097 2297
rect 11223 2263 11257 2297
rect 11383 2263 11417 2297
rect 11543 2263 11577 2297
rect 11703 2263 11737 2297
rect 11863 2263 11897 2297
rect 12023 2263 12057 2297
rect 12183 2263 12217 2297
rect 12343 2263 12377 2297
rect 8503 2103 8537 2137
rect 8663 2103 8697 2137
rect 8823 2103 8857 2137
rect 8983 2103 9017 2137
rect 9143 2103 9177 2137
rect 9303 2103 9337 2137
rect 9463 2103 9497 2137
rect 9623 2103 9657 2137
rect 9783 2103 9817 2137
rect 9943 2103 9977 2137
rect 10103 2103 10137 2137
rect 10263 2103 10297 2137
rect 10423 2103 10457 2137
rect 10583 2103 10617 2137
rect 10743 2103 10777 2137
rect 10903 2103 10937 2137
rect 11063 2103 11097 2137
rect 11223 2103 11257 2137
rect 11383 2103 11417 2137
rect 11543 2103 11577 2137
rect 11703 2103 11737 2137
rect 11863 2103 11897 2137
rect 12023 2103 12057 2137
rect 12183 2103 12217 2137
rect 12343 2103 12377 2137
rect 8503 1943 8537 1977
rect 8663 1943 8697 1977
rect 8823 1943 8857 1977
rect 8983 1943 9017 1977
rect 9143 1943 9177 1977
rect 9303 1943 9337 1977
rect 9463 1943 9497 1977
rect 9623 1943 9657 1977
rect 9783 1943 9817 1977
rect 9943 1943 9977 1977
rect 10103 1943 10137 1977
rect 10263 1943 10297 1977
rect 10423 1943 10457 1977
rect 10583 1943 10617 1977
rect 10743 1943 10777 1977
rect 10903 1943 10937 1977
rect 11063 1943 11097 1977
rect 11223 1943 11257 1977
rect 11383 1943 11417 1977
rect 11543 1943 11577 1977
rect 11703 1943 11737 1977
rect 11863 1943 11897 1977
rect 12023 1943 12057 1977
rect 12183 1943 12217 1977
rect 12343 1943 12377 1977
rect 8503 1783 8537 1817
rect 8663 1783 8697 1817
rect 8823 1783 8857 1817
rect 8983 1783 9017 1817
rect 9143 1783 9177 1817
rect 9303 1783 9337 1817
rect 9463 1783 9497 1817
rect 9623 1783 9657 1817
rect 9783 1783 9817 1817
rect 9943 1783 9977 1817
rect 10103 1783 10137 1817
rect 10263 1783 10297 1817
rect 10423 1783 10457 1817
rect 10583 1783 10617 1817
rect 10743 1783 10777 1817
rect 10903 1783 10937 1817
rect 11063 1783 11097 1817
rect 11223 1783 11257 1817
rect 11383 1783 11417 1817
rect 11543 1783 11577 1817
rect 11703 1783 11737 1817
rect 11863 1783 11897 1817
rect 12023 1783 12057 1817
rect 12183 1783 12217 1817
rect 12343 1783 12377 1817
rect 8503 1623 8537 1657
rect 8663 1623 8697 1657
rect 8823 1623 8857 1657
rect 8983 1623 9017 1657
rect 9143 1623 9177 1657
rect 9303 1623 9337 1657
rect 9463 1623 9497 1657
rect 9623 1623 9657 1657
rect 9783 1623 9817 1657
rect 9943 1623 9977 1657
rect 10103 1623 10137 1657
rect 10263 1623 10297 1657
rect 10423 1623 10457 1657
rect 10583 1623 10617 1657
rect 10743 1623 10777 1657
rect 10903 1623 10937 1657
rect 11063 1623 11097 1657
rect 11223 1623 11257 1657
rect 11383 1623 11417 1657
rect 11543 1623 11577 1657
rect 11703 1623 11737 1657
rect 11863 1623 11897 1657
rect 12023 1623 12057 1657
rect 12183 1623 12217 1657
rect 12343 1623 12377 1657
rect 8503 1463 8537 1497
rect 8663 1463 8697 1497
rect 8823 1463 8857 1497
rect 8983 1463 9017 1497
rect 9143 1463 9177 1497
rect 9303 1463 9337 1497
rect 9463 1463 9497 1497
rect 9623 1463 9657 1497
rect 9783 1463 9817 1497
rect 9943 1463 9977 1497
rect 10103 1463 10137 1497
rect 10263 1463 10297 1497
rect 10423 1463 10457 1497
rect 10583 1463 10617 1497
rect 10743 1463 10777 1497
rect 10903 1463 10937 1497
rect 11063 1463 11097 1497
rect 11223 1463 11257 1497
rect 11383 1463 11417 1497
rect 11543 1463 11577 1497
rect 11703 1463 11737 1497
rect 11863 1463 11897 1497
rect 12023 1463 12057 1497
rect 12183 1463 12217 1497
rect 12343 1463 12377 1497
rect 8503 1303 8537 1337
rect 8663 1303 8697 1337
rect 8823 1303 8857 1337
rect 8983 1303 9017 1337
rect 9143 1303 9177 1337
rect 9303 1303 9337 1337
rect 9463 1303 9497 1337
rect 9623 1303 9657 1337
rect 9783 1303 9817 1337
rect 9943 1303 9977 1337
rect 10103 1303 10137 1337
rect 10263 1303 10297 1337
rect 10423 1303 10457 1337
rect 10583 1303 10617 1337
rect 10743 1303 10777 1337
rect 10903 1303 10937 1337
rect 11063 1303 11097 1337
rect 11223 1303 11257 1337
rect 11383 1303 11417 1337
rect 11543 1303 11577 1337
rect 11703 1303 11737 1337
rect 11863 1303 11897 1337
rect 12023 1303 12057 1337
rect 12183 1303 12217 1337
rect 12343 1303 12377 1337
rect 8503 1143 8537 1177
rect 8663 1143 8697 1177
rect 8823 1143 8857 1177
rect 8983 1143 9017 1177
rect 9143 1143 9177 1177
rect 9303 1143 9337 1177
rect 9463 1143 9497 1177
rect 9623 1143 9657 1177
rect 9783 1143 9817 1177
rect 9943 1143 9977 1177
rect 10103 1143 10137 1177
rect 10263 1143 10297 1177
rect 10423 1143 10457 1177
rect 10583 1143 10617 1177
rect 10743 1143 10777 1177
rect 10903 1143 10937 1177
rect 11063 1143 11097 1177
rect 11223 1143 11257 1177
rect 11383 1143 11417 1177
rect 11543 1143 11577 1177
rect 11703 1143 11737 1177
rect 11863 1143 11897 1177
rect 12023 1143 12057 1177
rect 12183 1143 12217 1177
rect 12343 1143 12377 1177
rect 8503 983 8537 1017
rect 8663 983 8697 1017
rect 8823 983 8857 1017
rect 8983 983 9017 1017
rect 9143 983 9177 1017
rect 9303 983 9337 1017
rect 9463 983 9497 1017
rect 9623 983 9657 1017
rect 9783 983 9817 1017
rect 9943 983 9977 1017
rect 10103 983 10137 1017
rect 10263 983 10297 1017
rect 10423 983 10457 1017
rect 10583 983 10617 1017
rect 10743 983 10777 1017
rect 10903 983 10937 1017
rect 11063 983 11097 1017
rect 11223 983 11257 1017
rect 11383 983 11417 1017
rect 11543 983 11577 1017
rect 11703 983 11737 1017
rect 11863 983 11897 1017
rect 12023 983 12057 1017
rect 12183 983 12217 1017
rect 12343 983 12377 1017
rect 8503 823 8537 857
rect 8663 823 8697 857
rect 8823 823 8857 857
rect 8983 823 9017 857
rect 9143 823 9177 857
rect 9303 823 9337 857
rect 9463 823 9497 857
rect 9623 823 9657 857
rect 9783 823 9817 857
rect 9943 823 9977 857
rect 10103 823 10137 857
rect 10263 823 10297 857
rect 10423 823 10457 857
rect 10583 823 10617 857
rect 10743 823 10777 857
rect 10903 823 10937 857
rect 11063 823 11097 857
rect 11223 823 11257 857
rect 11383 823 11417 857
rect 11543 823 11577 857
rect 11703 823 11737 857
rect 11863 823 11897 857
rect 12023 823 12057 857
rect 12183 823 12217 857
rect 12343 823 12377 857
rect 8503 663 8537 697
rect 8663 663 8697 697
rect 8823 663 8857 697
rect 8983 663 9017 697
rect 9143 663 9177 697
rect 9303 663 9337 697
rect 9463 663 9497 697
rect 9623 663 9657 697
rect 9783 663 9817 697
rect 9943 663 9977 697
rect 10103 663 10137 697
rect 10263 663 10297 697
rect 10423 663 10457 697
rect 10583 663 10617 697
rect 10743 663 10777 697
rect 10903 663 10937 697
rect 11063 663 11097 697
rect 11223 663 11257 697
rect 11383 663 11417 697
rect 11543 663 11577 697
rect 11703 663 11737 697
rect 11863 663 11897 697
rect 12023 663 12057 697
rect 12183 663 12217 697
rect 12343 663 12377 697
rect 8503 503 8537 537
rect 8663 503 8697 537
rect 8823 503 8857 537
rect 8983 503 9017 537
rect 9143 503 9177 537
rect 9303 503 9337 537
rect 9463 503 9497 537
rect 9623 503 9657 537
rect 9783 503 9817 537
rect 9943 503 9977 537
rect 10103 503 10137 537
rect 10263 503 10297 537
rect 10423 503 10457 537
rect 10583 503 10617 537
rect 10743 503 10777 537
rect 10903 503 10937 537
rect 11063 503 11097 537
rect 11223 503 11257 537
rect 11383 503 11417 537
rect 11543 503 11577 537
rect 11703 503 11737 537
rect 11863 503 11897 537
rect 12023 503 12057 537
rect 12183 503 12217 537
rect 12343 503 12377 537
rect 8503 343 8537 377
rect 8663 343 8697 377
rect 8823 343 8857 377
rect 8983 343 9017 377
rect 9143 343 9177 377
rect 9303 343 9337 377
rect 9463 343 9497 377
rect 9623 343 9657 377
rect 9783 343 9817 377
rect 9943 343 9977 377
rect 10103 343 10137 377
rect 10263 343 10297 377
rect 10423 343 10457 377
rect 10583 343 10617 377
rect 10743 343 10777 377
rect 10903 343 10937 377
rect 11063 343 11097 377
rect 11223 343 11257 377
rect 11383 343 11417 377
rect 11543 343 11577 377
rect 11703 343 11737 377
rect 11863 343 11897 377
rect 12023 343 12057 377
rect 12183 343 12217 377
rect 12343 343 12377 377
rect 8503 183 8537 217
rect 8663 183 8697 217
rect 8823 183 8857 217
rect 8983 183 9017 217
rect 9143 183 9177 217
rect 9303 183 9337 217
rect 9463 183 9497 217
rect 9623 183 9657 217
rect 9783 183 9817 217
rect 9943 183 9977 217
rect 10103 183 10137 217
rect 10263 183 10297 217
rect 10423 183 10457 217
rect 10583 183 10617 217
rect 10743 183 10777 217
rect 10903 183 10937 217
rect 11063 183 11097 217
rect 11223 183 11257 217
rect 11383 183 11417 217
rect 11543 183 11577 217
rect 11703 183 11737 217
rect 11863 183 11897 217
rect 12023 183 12057 217
rect 12183 183 12217 217
rect 12343 183 12377 217
rect 8503 23 8537 57
rect 8663 23 8697 57
rect 8823 23 8857 57
rect 8983 23 9017 57
rect 9143 23 9177 57
rect 9303 23 9337 57
rect 9463 23 9497 57
rect 9623 23 9657 57
rect 9783 23 9817 57
rect 9943 23 9977 57
rect 10103 23 10137 57
rect 10263 23 10297 57
rect 10423 23 10457 57
rect 10583 23 10617 57
rect 10743 23 10777 57
rect 10903 23 10937 57
rect 11063 23 11097 57
rect 11223 23 11257 57
rect 11383 23 11417 57
rect 11543 23 11577 57
rect 11703 23 11737 57
rect 11863 23 11897 57
rect 12023 23 12057 57
rect 12183 23 12217 57
rect 12343 23 12377 57
<< metal1 >>
rect 8480 31426 8560 31440
rect 8480 31374 8494 31426
rect 8546 31374 8560 31426
rect 8480 31266 8560 31374
rect 8480 31214 8494 31266
rect 8546 31214 8560 31266
rect 8480 31106 8560 31214
rect 8480 31054 8494 31106
rect 8546 31054 8560 31106
rect 8480 30946 8560 31054
rect 8480 30894 8494 30946
rect 8546 30894 8560 30946
rect 8480 30786 8560 30894
rect 8480 30734 8494 30786
rect 8546 30734 8560 30786
rect 8480 30626 8560 30734
rect 8480 30574 8494 30626
rect 8546 30574 8560 30626
rect 8480 30466 8560 30574
rect 8480 30414 8494 30466
rect 8546 30414 8560 30466
rect 8480 30306 8560 30414
rect 8480 30254 8494 30306
rect 8546 30254 8560 30306
rect 8480 30137 8560 30254
rect 8480 30103 8503 30137
rect 8537 30103 8560 30137
rect 8480 29986 8560 30103
rect 8480 29934 8494 29986
rect 8546 29934 8560 29986
rect 8480 29826 8560 29934
rect 8480 29774 8494 29826
rect 8546 29774 8560 29826
rect 8480 29666 8560 29774
rect 8480 29614 8494 29666
rect 8546 29614 8560 29666
rect 8480 29506 8560 29614
rect 8480 29454 8494 29506
rect 8546 29454 8560 29506
rect 8480 29346 8560 29454
rect 8480 29294 8494 29346
rect 8546 29294 8560 29346
rect 8480 29186 8560 29294
rect 8480 29134 8494 29186
rect 8546 29134 8560 29186
rect 8480 29026 8560 29134
rect 8480 28974 8494 29026
rect 8546 28974 8560 29026
rect 8480 28866 8560 28974
rect 8480 28814 8494 28866
rect 8546 28814 8560 28866
rect 8480 28697 8560 28814
rect 8480 28663 8503 28697
rect 8537 28663 8560 28697
rect 8480 28537 8560 28663
rect 8480 28503 8503 28537
rect 8537 28503 8560 28537
rect 8480 28377 8560 28503
rect 8480 28343 8503 28377
rect 8537 28343 8560 28377
rect 8480 28217 8560 28343
rect 8480 28183 8503 28217
rect 8537 28183 8560 28217
rect 8480 28066 8560 28183
rect 8480 28014 8494 28066
rect 8546 28014 8560 28066
rect 8480 27906 8560 28014
rect 8480 27854 8494 27906
rect 8546 27854 8560 27906
rect 8480 27746 8560 27854
rect 8480 27694 8494 27746
rect 8546 27694 8560 27746
rect 8480 27586 8560 27694
rect 8480 27534 8494 27586
rect 8546 27534 8560 27586
rect 8480 27426 8560 27534
rect 8480 27374 8494 27426
rect 8546 27374 8560 27426
rect 8480 27266 8560 27374
rect 8480 27214 8494 27266
rect 8546 27214 8560 27266
rect 8480 27106 8560 27214
rect 8480 27054 8494 27106
rect 8546 27054 8560 27106
rect 8480 26946 8560 27054
rect 8480 26894 8494 26946
rect 8546 26894 8560 26946
rect 8480 26777 8560 26894
rect 8480 26743 8503 26777
rect 8537 26743 8560 26777
rect 8480 26617 8560 26743
rect 8480 26583 8503 26617
rect 8537 26583 8560 26617
rect 8480 26457 8560 26583
rect 8480 26423 8503 26457
rect 8537 26423 8560 26457
rect 8480 26297 8560 26423
rect 8480 26263 8503 26297
rect 8537 26263 8560 26297
rect 8480 26146 8560 26263
rect 8480 26094 8494 26146
rect 8546 26094 8560 26146
rect 8480 25986 8560 26094
rect 8480 25934 8494 25986
rect 8546 25934 8560 25986
rect 8480 25826 8560 25934
rect 8480 25774 8494 25826
rect 8546 25774 8560 25826
rect 8480 25666 8560 25774
rect 8480 25614 8494 25666
rect 8546 25614 8560 25666
rect 8480 25506 8560 25614
rect 8480 25454 8494 25506
rect 8546 25454 8560 25506
rect 8480 25346 8560 25454
rect 8480 25294 8494 25346
rect 8546 25294 8560 25346
rect 8480 25186 8560 25294
rect 8480 25134 8494 25186
rect 8546 25134 8560 25186
rect 8480 25026 8560 25134
rect 8480 24974 8494 25026
rect 8546 24974 8560 25026
rect 8480 24857 8560 24974
rect 8480 24823 8503 24857
rect 8537 24823 8560 24857
rect 8480 24706 8560 24823
rect 8480 24654 8494 24706
rect 8546 24654 8560 24706
rect 8480 24546 8560 24654
rect 8480 24494 8494 24546
rect 8546 24494 8560 24546
rect 8480 24386 8560 24494
rect 8480 24334 8494 24386
rect 8546 24334 8560 24386
rect 8480 24226 8560 24334
rect 8480 24174 8494 24226
rect 8546 24174 8560 24226
rect 8480 24066 8560 24174
rect 8480 24014 8494 24066
rect 8546 24014 8560 24066
rect 8480 23906 8560 24014
rect 8480 23854 8494 23906
rect 8546 23854 8560 23906
rect 8480 23746 8560 23854
rect 8480 23694 8494 23746
rect 8546 23694 8560 23746
rect 8480 23586 8560 23694
rect 8480 23534 8494 23586
rect 8546 23534 8560 23586
rect 8480 23426 8560 23534
rect 8480 23374 8494 23426
rect 8546 23374 8560 23426
rect 8480 23266 8560 23374
rect 8480 23214 8494 23266
rect 8546 23214 8560 23266
rect 8480 23106 8560 23214
rect 8480 23054 8494 23106
rect 8546 23054 8560 23106
rect 8480 22946 8560 23054
rect 8480 22894 8494 22946
rect 8546 22894 8560 22946
rect 8480 22786 8560 22894
rect 8480 22734 8494 22786
rect 8546 22734 8560 22786
rect 8480 22626 8560 22734
rect 8480 22574 8494 22626
rect 8546 22574 8560 22626
rect 8480 22466 8560 22574
rect 8480 22414 8494 22466
rect 8546 22414 8560 22466
rect 8480 22306 8560 22414
rect 8480 22254 8494 22306
rect 8546 22254 8560 22306
rect 8480 22146 8560 22254
rect 8480 22094 8494 22146
rect 8546 22094 8560 22146
rect 8480 21977 8560 22094
rect 8480 21943 8503 21977
rect 8537 21943 8560 21977
rect 8480 21826 8560 21943
rect 8480 21774 8494 21826
rect 8546 21774 8560 21826
rect 8480 21666 8560 21774
rect 8480 21614 8494 21666
rect 8546 21614 8560 21666
rect 8480 21506 8560 21614
rect 8480 21454 8494 21506
rect 8546 21454 8560 21506
rect 8480 21346 8560 21454
rect 8480 21294 8494 21346
rect 8546 21294 8560 21346
rect 8480 21186 8560 21294
rect 8480 21134 8494 21186
rect 8546 21134 8560 21186
rect 8480 21026 8560 21134
rect 8480 20974 8494 21026
rect 8546 20974 8560 21026
rect 8480 20866 8560 20974
rect 8480 20814 8494 20866
rect 8546 20814 8560 20866
rect 8480 20706 8560 20814
rect 8480 20654 8494 20706
rect 8546 20654 8560 20706
rect 8480 20537 8560 20654
rect 8480 20503 8503 20537
rect 8537 20503 8560 20537
rect 8480 20377 8560 20503
rect 8480 20343 8503 20377
rect 8537 20343 8560 20377
rect 8480 20217 8560 20343
rect 8480 20183 8503 20217
rect 8537 20183 8560 20217
rect 8480 20057 8560 20183
rect 8480 20023 8503 20057
rect 8537 20023 8560 20057
rect 8480 19906 8560 20023
rect 8480 19854 8494 19906
rect 8546 19854 8560 19906
rect 8480 19746 8560 19854
rect 8480 19694 8494 19746
rect 8546 19694 8560 19746
rect 8480 19586 8560 19694
rect 8480 19534 8494 19586
rect 8546 19534 8560 19586
rect 8480 19426 8560 19534
rect 8480 19374 8494 19426
rect 8546 19374 8560 19426
rect 8480 19266 8560 19374
rect 8480 19214 8494 19266
rect 8546 19214 8560 19266
rect 8480 19106 8560 19214
rect 8480 19054 8494 19106
rect 8546 19054 8560 19106
rect 8480 18946 8560 19054
rect 8480 18894 8494 18946
rect 8546 18894 8560 18946
rect 8480 18786 8560 18894
rect 8480 18734 8494 18786
rect 8546 18734 8560 18786
rect 8480 18617 8560 18734
rect 8480 18583 8503 18617
rect 8537 18583 8560 18617
rect 8480 18457 8560 18583
rect 8480 18423 8503 18457
rect 8537 18423 8560 18457
rect 8480 18297 8560 18423
rect 8480 18263 8503 18297
rect 8537 18263 8560 18297
rect 8480 18137 8560 18263
rect 8480 18103 8503 18137
rect 8537 18103 8560 18137
rect 8480 17986 8560 18103
rect 8480 17934 8494 17986
rect 8546 17934 8560 17986
rect 8480 17826 8560 17934
rect 8480 17774 8494 17826
rect 8546 17774 8560 17826
rect 8480 17666 8560 17774
rect 8480 17614 8494 17666
rect 8546 17614 8560 17666
rect 8480 17506 8560 17614
rect 8480 17454 8494 17506
rect 8546 17454 8560 17506
rect 8480 17346 8560 17454
rect 8480 17294 8494 17346
rect 8546 17294 8560 17346
rect 8480 17186 8560 17294
rect 8480 17134 8494 17186
rect 8546 17134 8560 17186
rect 8480 17026 8560 17134
rect 8480 16974 8494 17026
rect 8546 16974 8560 17026
rect 8480 16866 8560 16974
rect 8480 16814 8494 16866
rect 8546 16814 8560 16866
rect 8480 16697 8560 16814
rect 8480 16663 8503 16697
rect 8537 16663 8560 16697
rect 8480 16546 8560 16663
rect 8480 16494 8494 16546
rect 8546 16494 8560 16546
rect 8480 16386 8560 16494
rect 8480 16334 8494 16386
rect 8546 16334 8560 16386
rect 8480 16226 8560 16334
rect 8480 16174 8494 16226
rect 8546 16174 8560 16226
rect 8480 16066 8560 16174
rect 8480 16014 8494 16066
rect 8546 16014 8560 16066
rect 8480 15906 8560 16014
rect 8480 15854 8494 15906
rect 8546 15854 8560 15906
rect 8480 15746 8560 15854
rect 8480 15694 8494 15746
rect 8546 15694 8560 15746
rect 8480 15586 8560 15694
rect 8480 15534 8494 15586
rect 8546 15534 8560 15586
rect 8480 15426 8560 15534
rect 8480 15374 8494 15426
rect 8546 15374 8560 15426
rect 8480 15266 8560 15374
rect 8480 15214 8494 15266
rect 8546 15214 8560 15266
rect 8480 15106 8560 15214
rect 8480 15054 8494 15106
rect 8546 15054 8560 15106
rect 8480 14946 8560 15054
rect 8480 14894 8494 14946
rect 8546 14894 8560 14946
rect 8480 14786 8560 14894
rect 8480 14734 8494 14786
rect 8546 14734 8560 14786
rect 8480 14626 8560 14734
rect 8480 14574 8494 14626
rect 8546 14574 8560 14626
rect 8480 14466 8560 14574
rect 8480 14414 8494 14466
rect 8546 14414 8560 14466
rect 8480 14306 8560 14414
rect 8480 14254 8494 14306
rect 8546 14254 8560 14306
rect 8480 14146 8560 14254
rect 8480 14094 8494 14146
rect 8546 14094 8560 14146
rect 8480 13986 8560 14094
rect 8480 13934 8494 13986
rect 8546 13934 8560 13986
rect 8480 13817 8560 13934
rect 8480 13783 8503 13817
rect 8537 13783 8560 13817
rect 8480 13666 8560 13783
rect 8480 13614 8494 13666
rect 8546 13614 8560 13666
rect 8480 13506 8560 13614
rect 8480 13454 8494 13506
rect 8546 13454 8560 13506
rect 8480 13346 8560 13454
rect 8480 13294 8494 13346
rect 8546 13294 8560 13346
rect 8480 13186 8560 13294
rect 8480 13134 8494 13186
rect 8546 13134 8560 13186
rect 8480 13026 8560 13134
rect 8480 12974 8494 13026
rect 8546 12974 8560 13026
rect 8480 12866 8560 12974
rect 8480 12814 8494 12866
rect 8546 12814 8560 12866
rect 8480 12706 8560 12814
rect 8480 12654 8494 12706
rect 8546 12654 8560 12706
rect 8480 12546 8560 12654
rect 8480 12494 8494 12546
rect 8546 12494 8560 12546
rect 8480 12377 8560 12494
rect 8480 12343 8503 12377
rect 8537 12343 8560 12377
rect 8480 12217 8560 12343
rect 8480 12183 8503 12217
rect 8537 12183 8560 12217
rect 8480 12057 8560 12183
rect 8480 12023 8503 12057
rect 8537 12023 8560 12057
rect 8480 11897 8560 12023
rect 8480 11863 8503 11897
rect 8537 11863 8560 11897
rect 8480 11746 8560 11863
rect 8480 11694 8494 11746
rect 8546 11694 8560 11746
rect 8480 11586 8560 11694
rect 8480 11534 8494 11586
rect 8546 11534 8560 11586
rect 8480 11426 8560 11534
rect 8480 11374 8494 11426
rect 8546 11374 8560 11426
rect 8480 11266 8560 11374
rect 8480 11214 8494 11266
rect 8546 11214 8560 11266
rect 8480 11106 8560 11214
rect 8480 11054 8494 11106
rect 8546 11054 8560 11106
rect 8480 10946 8560 11054
rect 8480 10894 8494 10946
rect 8546 10894 8560 10946
rect 8480 10786 8560 10894
rect 8480 10734 8494 10786
rect 8546 10734 8560 10786
rect 8480 10626 8560 10734
rect 8480 10574 8494 10626
rect 8546 10574 8560 10626
rect 8480 10466 8560 10574
rect 8480 10414 8494 10466
rect 8546 10414 8560 10466
rect 8480 10306 8560 10414
rect 8480 10254 8494 10306
rect 8546 10254 8560 10306
rect 8480 10146 8560 10254
rect 8480 10094 8494 10146
rect 8546 10094 8560 10146
rect 8480 9986 8560 10094
rect 8480 9934 8494 9986
rect 8546 9934 8560 9986
rect 8480 9826 8560 9934
rect 8480 9774 8494 9826
rect 8546 9774 8560 9826
rect 8480 9657 8560 9774
rect 8480 9623 8503 9657
rect 8537 9623 8560 9657
rect 8480 9506 8560 9623
rect 8480 9454 8494 9506
rect 8546 9454 8560 9506
rect 8480 9346 8560 9454
rect 8480 9294 8494 9346
rect 8546 9294 8560 9346
rect 8480 9177 8560 9294
rect 8480 9143 8503 9177
rect 8537 9143 8560 9177
rect 8480 9026 8560 9143
rect 8480 8974 8494 9026
rect 8546 8974 8560 9026
rect 8480 8866 8560 8974
rect 8480 8814 8494 8866
rect 8546 8814 8560 8866
rect 8480 8706 8560 8814
rect 8480 8654 8494 8706
rect 8546 8654 8560 8706
rect 8480 8546 8560 8654
rect 8480 8494 8494 8546
rect 8546 8494 8560 8546
rect 8480 8386 8560 8494
rect 8480 8334 8494 8386
rect 8546 8334 8560 8386
rect 8480 8226 8560 8334
rect 8480 8174 8494 8226
rect 8546 8174 8560 8226
rect 8480 8066 8560 8174
rect 8480 8014 8494 8066
rect 8546 8014 8560 8066
rect 8480 7906 8560 8014
rect 8480 7854 8494 7906
rect 8546 7854 8560 7906
rect 8480 7746 8560 7854
rect 8480 7694 8494 7746
rect 8546 7694 8560 7746
rect 8480 7577 8560 7694
rect 8480 7543 8503 7577
rect 8537 7543 8560 7577
rect 8480 7426 8560 7543
rect 8480 7374 8494 7426
rect 8546 7374 8560 7426
rect 8480 7266 8560 7374
rect 8480 7214 8494 7266
rect 8546 7214 8560 7266
rect 8480 7097 8560 7214
rect 8480 7063 8503 7097
rect 8537 7063 8560 7097
rect 8480 6946 8560 7063
rect 8480 6894 8494 6946
rect 8546 6894 8560 6946
rect 8480 6786 8560 6894
rect 8480 6734 8494 6786
rect 8546 6734 8560 6786
rect 8480 6617 8560 6734
rect 8480 6583 8503 6617
rect 8537 6583 8560 6617
rect 8480 6466 8560 6583
rect 8480 6414 8494 6466
rect 8546 6414 8560 6466
rect 8480 6306 8560 6414
rect 8480 6254 8494 6306
rect 8546 6254 8560 6306
rect 8480 6146 8560 6254
rect 8480 6094 8494 6146
rect 8546 6094 8560 6146
rect 8480 5986 8560 6094
rect 8480 5934 8494 5986
rect 8546 5934 8560 5986
rect 8480 5826 8560 5934
rect 8480 5774 8494 5826
rect 8546 5774 8560 5826
rect 8480 5666 8560 5774
rect 8480 5614 8494 5666
rect 8546 5614 8560 5666
rect 8480 5506 8560 5614
rect 8480 5454 8494 5506
rect 8546 5454 8560 5506
rect 8480 5346 8560 5454
rect 8480 5294 8494 5346
rect 8546 5294 8560 5346
rect 8480 5186 8560 5294
rect 8480 5134 8494 5186
rect 8546 5134 8560 5186
rect 8480 5026 8560 5134
rect 8480 4974 8494 5026
rect 8546 4974 8560 5026
rect 8480 4866 8560 4974
rect 8480 4814 8494 4866
rect 8546 4814 8560 4866
rect 8480 4706 8560 4814
rect 8480 4654 8494 4706
rect 8546 4654 8560 4706
rect 8480 4546 8560 4654
rect 8480 4494 8494 4546
rect 8546 4494 8560 4546
rect 8480 4386 8560 4494
rect 8480 4334 8494 4386
rect 8546 4334 8560 4386
rect 8480 4226 8560 4334
rect 8480 4174 8494 4226
rect 8546 4174 8560 4226
rect 8480 4066 8560 4174
rect 8480 4014 8494 4066
rect 8546 4014 8560 4066
rect 8480 3906 8560 4014
rect 8480 3854 8494 3906
rect 8546 3854 8560 3906
rect 8480 3737 8560 3854
rect 8480 3703 8503 3737
rect 8537 3703 8560 3737
rect 8480 3577 8560 3703
rect 8480 3543 8503 3577
rect 8537 3543 8560 3577
rect 8480 3426 8560 3543
rect 8480 3374 8494 3426
rect 8546 3374 8560 3426
rect 8480 3266 8560 3374
rect 8480 3214 8494 3266
rect 8546 3214 8560 3266
rect 8480 3106 8560 3214
rect 8480 3054 8494 3106
rect 8546 3054 8560 3106
rect 8480 2946 8560 3054
rect 8480 2894 8494 2946
rect 8546 2894 8560 2946
rect 8480 2786 8560 2894
rect 8480 2734 8494 2786
rect 8546 2734 8560 2786
rect 8480 2626 8560 2734
rect 8480 2574 8494 2626
rect 8546 2574 8560 2626
rect 8480 2466 8560 2574
rect 8480 2414 8494 2466
rect 8546 2414 8560 2466
rect 8480 2306 8560 2414
rect 8480 2254 8494 2306
rect 8546 2254 8560 2306
rect 8480 2146 8560 2254
rect 8480 2094 8494 2146
rect 8546 2094 8560 2146
rect 8480 1986 8560 2094
rect 8480 1934 8494 1986
rect 8546 1934 8560 1986
rect 8480 1817 8560 1934
rect 8480 1783 8503 1817
rect 8537 1783 8560 1817
rect 8480 1666 8560 1783
rect 8480 1614 8494 1666
rect 8546 1614 8560 1666
rect 8480 1506 8560 1614
rect 8480 1454 8494 1506
rect 8546 1454 8560 1506
rect 8480 1346 8560 1454
rect 8480 1294 8494 1346
rect 8546 1294 8560 1346
rect 8480 1186 8560 1294
rect 8480 1134 8494 1186
rect 8546 1134 8560 1186
rect 8480 1026 8560 1134
rect 8480 974 8494 1026
rect 8546 974 8560 1026
rect 8480 857 8560 974
rect 8480 823 8503 857
rect 8537 823 8560 857
rect 8480 697 8560 823
rect 8480 663 8503 697
rect 8537 663 8560 697
rect 8480 546 8560 663
rect 8480 494 8494 546
rect 8546 494 8560 546
rect 8480 386 8560 494
rect 8480 334 8494 386
rect 8546 334 8560 386
rect 8480 226 8560 334
rect 8480 174 8494 226
rect 8546 174 8560 226
rect 8480 66 8560 174
rect 8480 14 8494 66
rect 8546 14 8560 66
rect 8480 0 8560 14
rect 8640 31417 8720 31440
rect 8640 31383 8663 31417
rect 8697 31383 8720 31417
rect 8640 31257 8720 31383
rect 8640 31223 8663 31257
rect 8697 31223 8720 31257
rect 8640 31097 8720 31223
rect 8640 31063 8663 31097
rect 8697 31063 8720 31097
rect 8640 30937 8720 31063
rect 8640 30903 8663 30937
rect 8697 30903 8720 30937
rect 8640 30777 8720 30903
rect 8640 30743 8663 30777
rect 8697 30743 8720 30777
rect 8640 30617 8720 30743
rect 8640 30583 8663 30617
rect 8697 30583 8720 30617
rect 8640 30457 8720 30583
rect 8640 30423 8663 30457
rect 8697 30423 8720 30457
rect 8640 30297 8720 30423
rect 8640 30263 8663 30297
rect 8697 30263 8720 30297
rect 8640 30137 8720 30263
rect 8640 30103 8663 30137
rect 8697 30103 8720 30137
rect 8640 29977 8720 30103
rect 8640 29943 8663 29977
rect 8697 29943 8720 29977
rect 8640 29817 8720 29943
rect 8640 29783 8663 29817
rect 8697 29783 8720 29817
rect 8640 29657 8720 29783
rect 8640 29623 8663 29657
rect 8697 29623 8720 29657
rect 8640 29497 8720 29623
rect 8640 29463 8663 29497
rect 8697 29463 8720 29497
rect 8640 29337 8720 29463
rect 8640 29303 8663 29337
rect 8697 29303 8720 29337
rect 8640 29177 8720 29303
rect 8640 29143 8663 29177
rect 8697 29143 8720 29177
rect 8640 29017 8720 29143
rect 8640 28983 8663 29017
rect 8697 28983 8720 29017
rect 8640 28857 8720 28983
rect 8640 28823 8663 28857
rect 8697 28823 8720 28857
rect 8640 28697 8720 28823
rect 8640 28663 8663 28697
rect 8697 28663 8720 28697
rect 8640 28537 8720 28663
rect 8640 28503 8663 28537
rect 8697 28503 8720 28537
rect 8640 28377 8720 28503
rect 8640 28343 8663 28377
rect 8697 28343 8720 28377
rect 8640 28217 8720 28343
rect 8640 28183 8663 28217
rect 8697 28183 8720 28217
rect 8640 28057 8720 28183
rect 8640 28023 8663 28057
rect 8697 28023 8720 28057
rect 8640 27897 8720 28023
rect 8640 27863 8663 27897
rect 8697 27863 8720 27897
rect 8640 27737 8720 27863
rect 8640 27703 8663 27737
rect 8697 27703 8720 27737
rect 8640 27577 8720 27703
rect 8640 27543 8663 27577
rect 8697 27543 8720 27577
rect 8640 27417 8720 27543
rect 8640 27383 8663 27417
rect 8697 27383 8720 27417
rect 8640 27257 8720 27383
rect 8640 27223 8663 27257
rect 8697 27223 8720 27257
rect 8640 27097 8720 27223
rect 8640 27063 8663 27097
rect 8697 27063 8720 27097
rect 8640 26937 8720 27063
rect 8640 26903 8663 26937
rect 8697 26903 8720 26937
rect 8640 26777 8720 26903
rect 8640 26743 8663 26777
rect 8697 26743 8720 26777
rect 8640 26617 8720 26743
rect 8640 26583 8663 26617
rect 8697 26583 8720 26617
rect 8640 26457 8720 26583
rect 8640 26423 8663 26457
rect 8697 26423 8720 26457
rect 8640 26297 8720 26423
rect 8640 26263 8663 26297
rect 8697 26263 8720 26297
rect 8640 26137 8720 26263
rect 8640 26103 8663 26137
rect 8697 26103 8720 26137
rect 8640 25977 8720 26103
rect 8640 25943 8663 25977
rect 8697 25943 8720 25977
rect 8640 25817 8720 25943
rect 8640 25783 8663 25817
rect 8697 25783 8720 25817
rect 8640 25657 8720 25783
rect 8640 25623 8663 25657
rect 8697 25623 8720 25657
rect 8640 25497 8720 25623
rect 8640 25463 8663 25497
rect 8697 25463 8720 25497
rect 8640 25337 8720 25463
rect 8640 25303 8663 25337
rect 8697 25303 8720 25337
rect 8640 25177 8720 25303
rect 8640 25143 8663 25177
rect 8697 25143 8720 25177
rect 8640 25017 8720 25143
rect 8640 24983 8663 25017
rect 8697 24983 8720 25017
rect 8640 24857 8720 24983
rect 8640 24823 8663 24857
rect 8697 24823 8720 24857
rect 8640 24697 8720 24823
rect 8640 24663 8663 24697
rect 8697 24663 8720 24697
rect 8640 24537 8720 24663
rect 8640 24503 8663 24537
rect 8697 24503 8720 24537
rect 8640 24377 8720 24503
rect 8640 24343 8663 24377
rect 8697 24343 8720 24377
rect 8640 24217 8720 24343
rect 8640 24183 8663 24217
rect 8697 24183 8720 24217
rect 8640 24057 8720 24183
rect 8640 24023 8663 24057
rect 8697 24023 8720 24057
rect 8640 23897 8720 24023
rect 8640 23863 8663 23897
rect 8697 23863 8720 23897
rect 8640 23737 8720 23863
rect 8640 23703 8663 23737
rect 8697 23703 8720 23737
rect 8640 23577 8720 23703
rect 8640 23543 8663 23577
rect 8697 23543 8720 23577
rect 8640 23417 8720 23543
rect 8640 23383 8663 23417
rect 8697 23383 8720 23417
rect 8640 23257 8720 23383
rect 8640 23223 8663 23257
rect 8697 23223 8720 23257
rect 8640 23097 8720 23223
rect 8640 23063 8663 23097
rect 8697 23063 8720 23097
rect 8640 22937 8720 23063
rect 8640 22903 8663 22937
rect 8697 22903 8720 22937
rect 8640 22777 8720 22903
rect 8640 22743 8663 22777
rect 8697 22743 8720 22777
rect 8640 22617 8720 22743
rect 8640 22583 8663 22617
rect 8697 22583 8720 22617
rect 8640 22457 8720 22583
rect 8640 22423 8663 22457
rect 8697 22423 8720 22457
rect 8640 22297 8720 22423
rect 8640 22263 8663 22297
rect 8697 22263 8720 22297
rect 8640 22137 8720 22263
rect 8640 22103 8663 22137
rect 8697 22103 8720 22137
rect 8640 21977 8720 22103
rect 8640 21943 8663 21977
rect 8697 21943 8720 21977
rect 8640 21817 8720 21943
rect 8640 21783 8663 21817
rect 8697 21783 8720 21817
rect 8640 21657 8720 21783
rect 8640 21623 8663 21657
rect 8697 21623 8720 21657
rect 8640 21497 8720 21623
rect 8640 21463 8663 21497
rect 8697 21463 8720 21497
rect 8640 21337 8720 21463
rect 8640 21303 8663 21337
rect 8697 21303 8720 21337
rect 8640 21177 8720 21303
rect 8640 21143 8663 21177
rect 8697 21143 8720 21177
rect 8640 21017 8720 21143
rect 8640 20983 8663 21017
rect 8697 20983 8720 21017
rect 8640 20857 8720 20983
rect 8640 20823 8663 20857
rect 8697 20823 8720 20857
rect 8640 20697 8720 20823
rect 8640 20663 8663 20697
rect 8697 20663 8720 20697
rect 8640 20537 8720 20663
rect 8640 20503 8663 20537
rect 8697 20503 8720 20537
rect 8640 20377 8720 20503
rect 8640 20343 8663 20377
rect 8697 20343 8720 20377
rect 8640 20217 8720 20343
rect 8640 20183 8663 20217
rect 8697 20183 8720 20217
rect 8640 20057 8720 20183
rect 8640 20023 8663 20057
rect 8697 20023 8720 20057
rect 8640 19897 8720 20023
rect 8640 19863 8663 19897
rect 8697 19863 8720 19897
rect 8640 19737 8720 19863
rect 8640 19703 8663 19737
rect 8697 19703 8720 19737
rect 8640 19577 8720 19703
rect 8640 19543 8663 19577
rect 8697 19543 8720 19577
rect 8640 19417 8720 19543
rect 8640 19383 8663 19417
rect 8697 19383 8720 19417
rect 8640 19257 8720 19383
rect 8640 19223 8663 19257
rect 8697 19223 8720 19257
rect 8640 19097 8720 19223
rect 8640 19063 8663 19097
rect 8697 19063 8720 19097
rect 8640 18937 8720 19063
rect 8640 18903 8663 18937
rect 8697 18903 8720 18937
rect 8640 18777 8720 18903
rect 8640 18743 8663 18777
rect 8697 18743 8720 18777
rect 8640 18617 8720 18743
rect 8640 18583 8663 18617
rect 8697 18583 8720 18617
rect 8640 18457 8720 18583
rect 8640 18423 8663 18457
rect 8697 18423 8720 18457
rect 8640 18297 8720 18423
rect 8640 18263 8663 18297
rect 8697 18263 8720 18297
rect 8640 18137 8720 18263
rect 8640 18103 8663 18137
rect 8697 18103 8720 18137
rect 8640 17977 8720 18103
rect 8640 17943 8663 17977
rect 8697 17943 8720 17977
rect 8640 17817 8720 17943
rect 8640 17783 8663 17817
rect 8697 17783 8720 17817
rect 8640 17657 8720 17783
rect 8640 17623 8663 17657
rect 8697 17623 8720 17657
rect 8640 17497 8720 17623
rect 8640 17463 8663 17497
rect 8697 17463 8720 17497
rect 8640 17337 8720 17463
rect 8640 17303 8663 17337
rect 8697 17303 8720 17337
rect 8640 17177 8720 17303
rect 8640 17143 8663 17177
rect 8697 17143 8720 17177
rect 8640 17017 8720 17143
rect 8640 16983 8663 17017
rect 8697 16983 8720 17017
rect 8640 16857 8720 16983
rect 8640 16823 8663 16857
rect 8697 16823 8720 16857
rect 8640 16697 8720 16823
rect 8640 16663 8663 16697
rect 8697 16663 8720 16697
rect 8640 16537 8720 16663
rect 8640 16503 8663 16537
rect 8697 16503 8720 16537
rect 8640 16377 8720 16503
rect 8640 16343 8663 16377
rect 8697 16343 8720 16377
rect 8640 16217 8720 16343
rect 8640 16183 8663 16217
rect 8697 16183 8720 16217
rect 8640 16057 8720 16183
rect 8640 16023 8663 16057
rect 8697 16023 8720 16057
rect 8640 15897 8720 16023
rect 8640 15863 8663 15897
rect 8697 15863 8720 15897
rect 8640 15737 8720 15863
rect 8640 15703 8663 15737
rect 8697 15703 8720 15737
rect 8640 15577 8720 15703
rect 8640 15543 8663 15577
rect 8697 15543 8720 15577
rect 8640 15417 8720 15543
rect 8640 15383 8663 15417
rect 8697 15383 8720 15417
rect 8640 15257 8720 15383
rect 8640 15223 8663 15257
rect 8697 15223 8720 15257
rect 8640 15097 8720 15223
rect 8640 15063 8663 15097
rect 8697 15063 8720 15097
rect 8640 14937 8720 15063
rect 8640 14903 8663 14937
rect 8697 14903 8720 14937
rect 8640 14777 8720 14903
rect 8640 14743 8663 14777
rect 8697 14743 8720 14777
rect 8640 14617 8720 14743
rect 8640 14583 8663 14617
rect 8697 14583 8720 14617
rect 8640 14457 8720 14583
rect 8640 14423 8663 14457
rect 8697 14423 8720 14457
rect 8640 14297 8720 14423
rect 8640 14263 8663 14297
rect 8697 14263 8720 14297
rect 8640 14137 8720 14263
rect 8640 14103 8663 14137
rect 8697 14103 8720 14137
rect 8640 13977 8720 14103
rect 8640 13943 8663 13977
rect 8697 13943 8720 13977
rect 8640 13817 8720 13943
rect 8640 13783 8663 13817
rect 8697 13783 8720 13817
rect 8640 13657 8720 13783
rect 8640 13623 8663 13657
rect 8697 13623 8720 13657
rect 8640 13497 8720 13623
rect 8640 13463 8663 13497
rect 8697 13463 8720 13497
rect 8640 13337 8720 13463
rect 8640 13303 8663 13337
rect 8697 13303 8720 13337
rect 8640 13177 8720 13303
rect 8640 13143 8663 13177
rect 8697 13143 8720 13177
rect 8640 13017 8720 13143
rect 8640 12983 8663 13017
rect 8697 12983 8720 13017
rect 8640 12857 8720 12983
rect 8640 12823 8663 12857
rect 8697 12823 8720 12857
rect 8640 12697 8720 12823
rect 8640 12663 8663 12697
rect 8697 12663 8720 12697
rect 8640 12537 8720 12663
rect 8640 12503 8663 12537
rect 8697 12503 8720 12537
rect 8640 12377 8720 12503
rect 8640 12343 8663 12377
rect 8697 12343 8720 12377
rect 8640 12217 8720 12343
rect 8640 12183 8663 12217
rect 8697 12183 8720 12217
rect 8640 12057 8720 12183
rect 8640 12023 8663 12057
rect 8697 12023 8720 12057
rect 8640 11897 8720 12023
rect 8640 11863 8663 11897
rect 8697 11863 8720 11897
rect 8640 11737 8720 11863
rect 8640 11703 8663 11737
rect 8697 11703 8720 11737
rect 8640 11577 8720 11703
rect 8640 11543 8663 11577
rect 8697 11543 8720 11577
rect 8640 11417 8720 11543
rect 8640 11383 8663 11417
rect 8697 11383 8720 11417
rect 8640 11257 8720 11383
rect 8640 11223 8663 11257
rect 8697 11223 8720 11257
rect 8640 11097 8720 11223
rect 8640 11063 8663 11097
rect 8697 11063 8720 11097
rect 8640 10937 8720 11063
rect 8640 10903 8663 10937
rect 8697 10903 8720 10937
rect 8640 10777 8720 10903
rect 8640 10743 8663 10777
rect 8697 10743 8720 10777
rect 8640 10617 8720 10743
rect 8640 10583 8663 10617
rect 8697 10583 8720 10617
rect 8640 10457 8720 10583
rect 8640 10423 8663 10457
rect 8697 10423 8720 10457
rect 8640 10297 8720 10423
rect 8640 10263 8663 10297
rect 8697 10263 8720 10297
rect 8640 10137 8720 10263
rect 8640 10103 8663 10137
rect 8697 10103 8720 10137
rect 8640 9977 8720 10103
rect 8640 9943 8663 9977
rect 8697 9943 8720 9977
rect 8640 9817 8720 9943
rect 8640 9783 8663 9817
rect 8697 9783 8720 9817
rect 8640 9657 8720 9783
rect 8640 9623 8663 9657
rect 8697 9623 8720 9657
rect 8640 9497 8720 9623
rect 8640 9463 8663 9497
rect 8697 9463 8720 9497
rect 8640 9337 8720 9463
rect 8640 9303 8663 9337
rect 8697 9303 8720 9337
rect 8640 9177 8720 9303
rect 8640 9143 8663 9177
rect 8697 9143 8720 9177
rect 8640 9017 8720 9143
rect 8640 8983 8663 9017
rect 8697 8983 8720 9017
rect 8640 8857 8720 8983
rect 8640 8823 8663 8857
rect 8697 8823 8720 8857
rect 8640 8697 8720 8823
rect 8640 8663 8663 8697
rect 8697 8663 8720 8697
rect 8640 8537 8720 8663
rect 8640 8503 8663 8537
rect 8697 8503 8720 8537
rect 8640 8377 8720 8503
rect 8640 8343 8663 8377
rect 8697 8343 8720 8377
rect 8640 8217 8720 8343
rect 8640 8183 8663 8217
rect 8697 8183 8720 8217
rect 8640 8057 8720 8183
rect 8640 8023 8663 8057
rect 8697 8023 8720 8057
rect 8640 7897 8720 8023
rect 8640 7863 8663 7897
rect 8697 7863 8720 7897
rect 8640 7737 8720 7863
rect 8640 7703 8663 7737
rect 8697 7703 8720 7737
rect 8640 7577 8720 7703
rect 8640 7543 8663 7577
rect 8697 7543 8720 7577
rect 8640 7417 8720 7543
rect 8640 7383 8663 7417
rect 8697 7383 8720 7417
rect 8640 7257 8720 7383
rect 8640 7223 8663 7257
rect 8697 7223 8720 7257
rect 8640 7097 8720 7223
rect 8640 7063 8663 7097
rect 8697 7063 8720 7097
rect 8640 6937 8720 7063
rect 8640 6903 8663 6937
rect 8697 6903 8720 6937
rect 8640 6777 8720 6903
rect 8640 6743 8663 6777
rect 8697 6743 8720 6777
rect 8640 6617 8720 6743
rect 8640 6583 8663 6617
rect 8697 6583 8720 6617
rect 8640 6457 8720 6583
rect 8640 6423 8663 6457
rect 8697 6423 8720 6457
rect 8640 6297 8720 6423
rect 8640 6263 8663 6297
rect 8697 6263 8720 6297
rect 8640 6137 8720 6263
rect 8640 6103 8663 6137
rect 8697 6103 8720 6137
rect 8640 5977 8720 6103
rect 8640 5943 8663 5977
rect 8697 5943 8720 5977
rect 8640 5817 8720 5943
rect 8640 5783 8663 5817
rect 8697 5783 8720 5817
rect 8640 5657 8720 5783
rect 8640 5623 8663 5657
rect 8697 5623 8720 5657
rect 8640 5497 8720 5623
rect 8640 5463 8663 5497
rect 8697 5463 8720 5497
rect 8640 5337 8720 5463
rect 8640 5303 8663 5337
rect 8697 5303 8720 5337
rect 8640 5177 8720 5303
rect 8640 5143 8663 5177
rect 8697 5143 8720 5177
rect 8640 5017 8720 5143
rect 8640 4983 8663 5017
rect 8697 4983 8720 5017
rect 8640 4857 8720 4983
rect 8640 4823 8663 4857
rect 8697 4823 8720 4857
rect 8640 4697 8720 4823
rect 8640 4663 8663 4697
rect 8697 4663 8720 4697
rect 8640 4537 8720 4663
rect 8640 4503 8663 4537
rect 8697 4503 8720 4537
rect 8640 4377 8720 4503
rect 8640 4343 8663 4377
rect 8697 4343 8720 4377
rect 8640 4217 8720 4343
rect 8640 4183 8663 4217
rect 8697 4183 8720 4217
rect 8640 4057 8720 4183
rect 8640 4023 8663 4057
rect 8697 4023 8720 4057
rect 8640 3897 8720 4023
rect 8640 3863 8663 3897
rect 8697 3863 8720 3897
rect 8640 3737 8720 3863
rect 8640 3703 8663 3737
rect 8697 3703 8720 3737
rect 8640 3577 8720 3703
rect 8640 3543 8663 3577
rect 8697 3543 8720 3577
rect 8640 3417 8720 3543
rect 8640 3383 8663 3417
rect 8697 3383 8720 3417
rect 8640 3257 8720 3383
rect 8640 3223 8663 3257
rect 8697 3223 8720 3257
rect 8640 3097 8720 3223
rect 8640 3063 8663 3097
rect 8697 3063 8720 3097
rect 8640 2937 8720 3063
rect 8640 2903 8663 2937
rect 8697 2903 8720 2937
rect 8640 2777 8720 2903
rect 8640 2743 8663 2777
rect 8697 2743 8720 2777
rect 8640 2617 8720 2743
rect 8640 2583 8663 2617
rect 8697 2583 8720 2617
rect 8640 2457 8720 2583
rect 8640 2423 8663 2457
rect 8697 2423 8720 2457
rect 8640 2297 8720 2423
rect 8640 2263 8663 2297
rect 8697 2263 8720 2297
rect 8640 2137 8720 2263
rect 8640 2103 8663 2137
rect 8697 2103 8720 2137
rect 8640 1977 8720 2103
rect 8640 1943 8663 1977
rect 8697 1943 8720 1977
rect 8640 1817 8720 1943
rect 8640 1783 8663 1817
rect 8697 1783 8720 1817
rect 8640 1657 8720 1783
rect 8640 1623 8663 1657
rect 8697 1623 8720 1657
rect 8640 1497 8720 1623
rect 8640 1463 8663 1497
rect 8697 1463 8720 1497
rect 8640 1337 8720 1463
rect 8640 1303 8663 1337
rect 8697 1303 8720 1337
rect 8640 1177 8720 1303
rect 8640 1143 8663 1177
rect 8697 1143 8720 1177
rect 8640 1017 8720 1143
rect 8640 983 8663 1017
rect 8697 983 8720 1017
rect 8640 857 8720 983
rect 8640 823 8663 857
rect 8697 823 8720 857
rect 8640 697 8720 823
rect 8640 663 8663 697
rect 8697 663 8720 697
rect 8640 537 8720 663
rect 8640 503 8663 537
rect 8697 503 8720 537
rect 8640 377 8720 503
rect 8640 343 8663 377
rect 8697 343 8720 377
rect 8640 217 8720 343
rect 8640 183 8663 217
rect 8697 183 8720 217
rect 8640 57 8720 183
rect 8640 23 8663 57
rect 8697 23 8720 57
rect 8640 0 8720 23
rect 8800 31426 8880 31440
rect 8800 31374 8814 31426
rect 8866 31374 8880 31426
rect 8800 31266 8880 31374
rect 8800 31214 8814 31266
rect 8866 31214 8880 31266
rect 8800 31106 8880 31214
rect 8800 31054 8814 31106
rect 8866 31054 8880 31106
rect 8800 30946 8880 31054
rect 8800 30894 8814 30946
rect 8866 30894 8880 30946
rect 8800 30786 8880 30894
rect 8800 30734 8814 30786
rect 8866 30734 8880 30786
rect 8800 30626 8880 30734
rect 8800 30574 8814 30626
rect 8866 30574 8880 30626
rect 8800 30466 8880 30574
rect 8800 30414 8814 30466
rect 8866 30414 8880 30466
rect 8800 30306 8880 30414
rect 8800 30254 8814 30306
rect 8866 30254 8880 30306
rect 8800 30137 8880 30254
rect 8800 30103 8823 30137
rect 8857 30103 8880 30137
rect 8800 29986 8880 30103
rect 8800 29934 8814 29986
rect 8866 29934 8880 29986
rect 8800 29826 8880 29934
rect 8800 29774 8814 29826
rect 8866 29774 8880 29826
rect 8800 29666 8880 29774
rect 8800 29614 8814 29666
rect 8866 29614 8880 29666
rect 8800 29506 8880 29614
rect 8800 29454 8814 29506
rect 8866 29454 8880 29506
rect 8800 29346 8880 29454
rect 8800 29294 8814 29346
rect 8866 29294 8880 29346
rect 8800 29186 8880 29294
rect 8800 29134 8814 29186
rect 8866 29134 8880 29186
rect 8800 29026 8880 29134
rect 8800 28974 8814 29026
rect 8866 28974 8880 29026
rect 8800 28866 8880 28974
rect 8800 28814 8814 28866
rect 8866 28814 8880 28866
rect 8800 28697 8880 28814
rect 8800 28663 8823 28697
rect 8857 28663 8880 28697
rect 8800 28537 8880 28663
rect 8800 28503 8823 28537
rect 8857 28503 8880 28537
rect 8800 28377 8880 28503
rect 8800 28343 8823 28377
rect 8857 28343 8880 28377
rect 8800 28217 8880 28343
rect 8800 28183 8823 28217
rect 8857 28183 8880 28217
rect 8800 28066 8880 28183
rect 8800 28014 8814 28066
rect 8866 28014 8880 28066
rect 8800 27906 8880 28014
rect 8800 27854 8814 27906
rect 8866 27854 8880 27906
rect 8800 27746 8880 27854
rect 8800 27694 8814 27746
rect 8866 27694 8880 27746
rect 8800 27586 8880 27694
rect 8800 27534 8814 27586
rect 8866 27534 8880 27586
rect 8800 27426 8880 27534
rect 8800 27374 8814 27426
rect 8866 27374 8880 27426
rect 8800 27266 8880 27374
rect 8800 27214 8814 27266
rect 8866 27214 8880 27266
rect 8800 27106 8880 27214
rect 8800 27054 8814 27106
rect 8866 27054 8880 27106
rect 8800 26946 8880 27054
rect 8800 26894 8814 26946
rect 8866 26894 8880 26946
rect 8800 26777 8880 26894
rect 8800 26743 8823 26777
rect 8857 26743 8880 26777
rect 8800 26617 8880 26743
rect 8800 26583 8823 26617
rect 8857 26583 8880 26617
rect 8800 26457 8880 26583
rect 8800 26423 8823 26457
rect 8857 26423 8880 26457
rect 8800 26297 8880 26423
rect 8800 26263 8823 26297
rect 8857 26263 8880 26297
rect 8800 26146 8880 26263
rect 8800 26094 8814 26146
rect 8866 26094 8880 26146
rect 8800 25986 8880 26094
rect 8800 25934 8814 25986
rect 8866 25934 8880 25986
rect 8800 25826 8880 25934
rect 8800 25774 8814 25826
rect 8866 25774 8880 25826
rect 8800 25666 8880 25774
rect 8800 25614 8814 25666
rect 8866 25614 8880 25666
rect 8800 25506 8880 25614
rect 8800 25454 8814 25506
rect 8866 25454 8880 25506
rect 8800 25346 8880 25454
rect 8800 25294 8814 25346
rect 8866 25294 8880 25346
rect 8800 25186 8880 25294
rect 8800 25134 8814 25186
rect 8866 25134 8880 25186
rect 8800 25026 8880 25134
rect 8800 24974 8814 25026
rect 8866 24974 8880 25026
rect 8800 24857 8880 24974
rect 8800 24823 8823 24857
rect 8857 24823 8880 24857
rect 8800 24706 8880 24823
rect 8800 24654 8814 24706
rect 8866 24654 8880 24706
rect 8800 24546 8880 24654
rect 8800 24494 8814 24546
rect 8866 24494 8880 24546
rect 8800 24386 8880 24494
rect 8800 24334 8814 24386
rect 8866 24334 8880 24386
rect 8800 24226 8880 24334
rect 8800 24174 8814 24226
rect 8866 24174 8880 24226
rect 8800 24066 8880 24174
rect 8800 24014 8814 24066
rect 8866 24014 8880 24066
rect 8800 23906 8880 24014
rect 8800 23854 8814 23906
rect 8866 23854 8880 23906
rect 8800 23746 8880 23854
rect 8800 23694 8814 23746
rect 8866 23694 8880 23746
rect 8800 23586 8880 23694
rect 8800 23534 8814 23586
rect 8866 23534 8880 23586
rect 8800 23426 8880 23534
rect 8800 23374 8814 23426
rect 8866 23374 8880 23426
rect 8800 23266 8880 23374
rect 8800 23214 8814 23266
rect 8866 23214 8880 23266
rect 8800 23106 8880 23214
rect 8800 23054 8814 23106
rect 8866 23054 8880 23106
rect 8800 22946 8880 23054
rect 8800 22894 8814 22946
rect 8866 22894 8880 22946
rect 8800 22786 8880 22894
rect 8800 22734 8814 22786
rect 8866 22734 8880 22786
rect 8800 22626 8880 22734
rect 8800 22574 8814 22626
rect 8866 22574 8880 22626
rect 8800 22466 8880 22574
rect 8800 22414 8814 22466
rect 8866 22414 8880 22466
rect 8800 22306 8880 22414
rect 8800 22254 8814 22306
rect 8866 22254 8880 22306
rect 8800 22146 8880 22254
rect 8800 22094 8814 22146
rect 8866 22094 8880 22146
rect 8800 21977 8880 22094
rect 8800 21943 8823 21977
rect 8857 21943 8880 21977
rect 8800 21826 8880 21943
rect 8800 21774 8814 21826
rect 8866 21774 8880 21826
rect 8800 21666 8880 21774
rect 8800 21614 8814 21666
rect 8866 21614 8880 21666
rect 8800 21506 8880 21614
rect 8800 21454 8814 21506
rect 8866 21454 8880 21506
rect 8800 21346 8880 21454
rect 8800 21294 8814 21346
rect 8866 21294 8880 21346
rect 8800 21186 8880 21294
rect 8800 21134 8814 21186
rect 8866 21134 8880 21186
rect 8800 21026 8880 21134
rect 8800 20974 8814 21026
rect 8866 20974 8880 21026
rect 8800 20866 8880 20974
rect 8800 20814 8814 20866
rect 8866 20814 8880 20866
rect 8800 20706 8880 20814
rect 8800 20654 8814 20706
rect 8866 20654 8880 20706
rect 8800 20537 8880 20654
rect 8800 20503 8823 20537
rect 8857 20503 8880 20537
rect 8800 20377 8880 20503
rect 8800 20343 8823 20377
rect 8857 20343 8880 20377
rect 8800 20217 8880 20343
rect 8800 20183 8823 20217
rect 8857 20183 8880 20217
rect 8800 20057 8880 20183
rect 8800 20023 8823 20057
rect 8857 20023 8880 20057
rect 8800 19906 8880 20023
rect 8800 19854 8814 19906
rect 8866 19854 8880 19906
rect 8800 19746 8880 19854
rect 8800 19694 8814 19746
rect 8866 19694 8880 19746
rect 8800 19586 8880 19694
rect 8800 19534 8814 19586
rect 8866 19534 8880 19586
rect 8800 19426 8880 19534
rect 8800 19374 8814 19426
rect 8866 19374 8880 19426
rect 8800 19266 8880 19374
rect 8800 19214 8814 19266
rect 8866 19214 8880 19266
rect 8800 19106 8880 19214
rect 8800 19054 8814 19106
rect 8866 19054 8880 19106
rect 8800 18946 8880 19054
rect 8800 18894 8814 18946
rect 8866 18894 8880 18946
rect 8800 18786 8880 18894
rect 8800 18734 8814 18786
rect 8866 18734 8880 18786
rect 8800 18617 8880 18734
rect 8800 18583 8823 18617
rect 8857 18583 8880 18617
rect 8800 18457 8880 18583
rect 8800 18423 8823 18457
rect 8857 18423 8880 18457
rect 8800 18297 8880 18423
rect 8800 18263 8823 18297
rect 8857 18263 8880 18297
rect 8800 18137 8880 18263
rect 8800 18103 8823 18137
rect 8857 18103 8880 18137
rect 8800 17986 8880 18103
rect 8800 17934 8814 17986
rect 8866 17934 8880 17986
rect 8800 17826 8880 17934
rect 8800 17774 8814 17826
rect 8866 17774 8880 17826
rect 8800 17666 8880 17774
rect 8800 17614 8814 17666
rect 8866 17614 8880 17666
rect 8800 17506 8880 17614
rect 8800 17454 8814 17506
rect 8866 17454 8880 17506
rect 8800 17346 8880 17454
rect 8800 17294 8814 17346
rect 8866 17294 8880 17346
rect 8800 17186 8880 17294
rect 8800 17134 8814 17186
rect 8866 17134 8880 17186
rect 8800 17026 8880 17134
rect 8800 16974 8814 17026
rect 8866 16974 8880 17026
rect 8800 16866 8880 16974
rect 8800 16814 8814 16866
rect 8866 16814 8880 16866
rect 8800 16697 8880 16814
rect 8800 16663 8823 16697
rect 8857 16663 8880 16697
rect 8800 16546 8880 16663
rect 8800 16494 8814 16546
rect 8866 16494 8880 16546
rect 8800 16386 8880 16494
rect 8800 16334 8814 16386
rect 8866 16334 8880 16386
rect 8800 16226 8880 16334
rect 8800 16174 8814 16226
rect 8866 16174 8880 16226
rect 8800 16066 8880 16174
rect 8800 16014 8814 16066
rect 8866 16014 8880 16066
rect 8800 15906 8880 16014
rect 8800 15854 8814 15906
rect 8866 15854 8880 15906
rect 8800 15746 8880 15854
rect 8800 15694 8814 15746
rect 8866 15694 8880 15746
rect 8800 15586 8880 15694
rect 8800 15534 8814 15586
rect 8866 15534 8880 15586
rect 8800 15426 8880 15534
rect 8800 15374 8814 15426
rect 8866 15374 8880 15426
rect 8800 15266 8880 15374
rect 8800 15214 8814 15266
rect 8866 15214 8880 15266
rect 8800 15106 8880 15214
rect 8800 15054 8814 15106
rect 8866 15054 8880 15106
rect 8800 14946 8880 15054
rect 8800 14894 8814 14946
rect 8866 14894 8880 14946
rect 8800 14786 8880 14894
rect 8800 14734 8814 14786
rect 8866 14734 8880 14786
rect 8800 14626 8880 14734
rect 8800 14574 8814 14626
rect 8866 14574 8880 14626
rect 8800 14466 8880 14574
rect 8800 14414 8814 14466
rect 8866 14414 8880 14466
rect 8800 14306 8880 14414
rect 8800 14254 8814 14306
rect 8866 14254 8880 14306
rect 8800 14146 8880 14254
rect 8800 14094 8814 14146
rect 8866 14094 8880 14146
rect 8800 13986 8880 14094
rect 8800 13934 8814 13986
rect 8866 13934 8880 13986
rect 8800 13817 8880 13934
rect 8800 13783 8823 13817
rect 8857 13783 8880 13817
rect 8800 13666 8880 13783
rect 8800 13614 8814 13666
rect 8866 13614 8880 13666
rect 8800 13506 8880 13614
rect 8800 13454 8814 13506
rect 8866 13454 8880 13506
rect 8800 13346 8880 13454
rect 8800 13294 8814 13346
rect 8866 13294 8880 13346
rect 8800 13186 8880 13294
rect 8800 13134 8814 13186
rect 8866 13134 8880 13186
rect 8800 13026 8880 13134
rect 8800 12974 8814 13026
rect 8866 12974 8880 13026
rect 8800 12866 8880 12974
rect 8800 12814 8814 12866
rect 8866 12814 8880 12866
rect 8800 12706 8880 12814
rect 8800 12654 8814 12706
rect 8866 12654 8880 12706
rect 8800 12546 8880 12654
rect 8800 12494 8814 12546
rect 8866 12494 8880 12546
rect 8800 12377 8880 12494
rect 8800 12343 8823 12377
rect 8857 12343 8880 12377
rect 8800 12217 8880 12343
rect 8800 12183 8823 12217
rect 8857 12183 8880 12217
rect 8800 12057 8880 12183
rect 8800 12023 8823 12057
rect 8857 12023 8880 12057
rect 8800 11897 8880 12023
rect 8800 11863 8823 11897
rect 8857 11863 8880 11897
rect 8800 11746 8880 11863
rect 8800 11694 8814 11746
rect 8866 11694 8880 11746
rect 8800 11586 8880 11694
rect 8800 11534 8814 11586
rect 8866 11534 8880 11586
rect 8800 11426 8880 11534
rect 8800 11374 8814 11426
rect 8866 11374 8880 11426
rect 8800 11266 8880 11374
rect 8800 11214 8814 11266
rect 8866 11214 8880 11266
rect 8800 11106 8880 11214
rect 8800 11054 8814 11106
rect 8866 11054 8880 11106
rect 8800 10946 8880 11054
rect 8800 10894 8814 10946
rect 8866 10894 8880 10946
rect 8800 10786 8880 10894
rect 8800 10734 8814 10786
rect 8866 10734 8880 10786
rect 8800 10626 8880 10734
rect 8800 10574 8814 10626
rect 8866 10574 8880 10626
rect 8800 10466 8880 10574
rect 8800 10414 8814 10466
rect 8866 10414 8880 10466
rect 8800 10306 8880 10414
rect 8800 10254 8814 10306
rect 8866 10254 8880 10306
rect 8800 10146 8880 10254
rect 8800 10094 8814 10146
rect 8866 10094 8880 10146
rect 8800 9986 8880 10094
rect 8800 9934 8814 9986
rect 8866 9934 8880 9986
rect 8800 9826 8880 9934
rect 8800 9774 8814 9826
rect 8866 9774 8880 9826
rect 8800 9657 8880 9774
rect 8800 9623 8823 9657
rect 8857 9623 8880 9657
rect 8800 9506 8880 9623
rect 8800 9454 8814 9506
rect 8866 9454 8880 9506
rect 8800 9346 8880 9454
rect 8800 9294 8814 9346
rect 8866 9294 8880 9346
rect 8800 9177 8880 9294
rect 8800 9143 8823 9177
rect 8857 9143 8880 9177
rect 8800 9026 8880 9143
rect 8800 8974 8814 9026
rect 8866 8974 8880 9026
rect 8800 8866 8880 8974
rect 8800 8814 8814 8866
rect 8866 8814 8880 8866
rect 8800 8706 8880 8814
rect 8800 8654 8814 8706
rect 8866 8654 8880 8706
rect 8800 8546 8880 8654
rect 8800 8494 8814 8546
rect 8866 8494 8880 8546
rect 8800 8386 8880 8494
rect 8800 8334 8814 8386
rect 8866 8334 8880 8386
rect 8800 8226 8880 8334
rect 8800 8174 8814 8226
rect 8866 8174 8880 8226
rect 8800 8066 8880 8174
rect 8800 8014 8814 8066
rect 8866 8014 8880 8066
rect 8800 7906 8880 8014
rect 8800 7854 8814 7906
rect 8866 7854 8880 7906
rect 8800 7746 8880 7854
rect 8800 7694 8814 7746
rect 8866 7694 8880 7746
rect 8800 7577 8880 7694
rect 8800 7543 8823 7577
rect 8857 7543 8880 7577
rect 8800 7426 8880 7543
rect 8800 7374 8814 7426
rect 8866 7374 8880 7426
rect 8800 7266 8880 7374
rect 8800 7214 8814 7266
rect 8866 7214 8880 7266
rect 8800 7097 8880 7214
rect 8800 7063 8823 7097
rect 8857 7063 8880 7097
rect 8800 6946 8880 7063
rect 8800 6894 8814 6946
rect 8866 6894 8880 6946
rect 8800 6786 8880 6894
rect 8800 6734 8814 6786
rect 8866 6734 8880 6786
rect 8800 6617 8880 6734
rect 8800 6583 8823 6617
rect 8857 6583 8880 6617
rect 8800 6466 8880 6583
rect 8800 6414 8814 6466
rect 8866 6414 8880 6466
rect 8800 6306 8880 6414
rect 8800 6254 8814 6306
rect 8866 6254 8880 6306
rect 8800 6146 8880 6254
rect 8800 6094 8814 6146
rect 8866 6094 8880 6146
rect 8800 5986 8880 6094
rect 8800 5934 8814 5986
rect 8866 5934 8880 5986
rect 8800 5826 8880 5934
rect 8800 5774 8814 5826
rect 8866 5774 8880 5826
rect 8800 5666 8880 5774
rect 8800 5614 8814 5666
rect 8866 5614 8880 5666
rect 8800 5506 8880 5614
rect 8800 5454 8814 5506
rect 8866 5454 8880 5506
rect 8800 5346 8880 5454
rect 8800 5294 8814 5346
rect 8866 5294 8880 5346
rect 8800 5186 8880 5294
rect 8800 5134 8814 5186
rect 8866 5134 8880 5186
rect 8800 5026 8880 5134
rect 8800 4974 8814 5026
rect 8866 4974 8880 5026
rect 8800 4866 8880 4974
rect 8800 4814 8814 4866
rect 8866 4814 8880 4866
rect 8800 4706 8880 4814
rect 8800 4654 8814 4706
rect 8866 4654 8880 4706
rect 8800 4546 8880 4654
rect 8800 4494 8814 4546
rect 8866 4494 8880 4546
rect 8800 4386 8880 4494
rect 8800 4334 8814 4386
rect 8866 4334 8880 4386
rect 8800 4226 8880 4334
rect 8800 4174 8814 4226
rect 8866 4174 8880 4226
rect 8800 4066 8880 4174
rect 8800 4014 8814 4066
rect 8866 4014 8880 4066
rect 8800 3906 8880 4014
rect 8800 3854 8814 3906
rect 8866 3854 8880 3906
rect 8800 3737 8880 3854
rect 8800 3703 8823 3737
rect 8857 3703 8880 3737
rect 8800 3577 8880 3703
rect 8800 3543 8823 3577
rect 8857 3543 8880 3577
rect 8800 3426 8880 3543
rect 8800 3374 8814 3426
rect 8866 3374 8880 3426
rect 8800 3266 8880 3374
rect 8800 3214 8814 3266
rect 8866 3214 8880 3266
rect 8800 3106 8880 3214
rect 8800 3054 8814 3106
rect 8866 3054 8880 3106
rect 8800 2946 8880 3054
rect 8800 2894 8814 2946
rect 8866 2894 8880 2946
rect 8800 2786 8880 2894
rect 8800 2734 8814 2786
rect 8866 2734 8880 2786
rect 8800 2626 8880 2734
rect 8800 2574 8814 2626
rect 8866 2574 8880 2626
rect 8800 2466 8880 2574
rect 8800 2414 8814 2466
rect 8866 2414 8880 2466
rect 8800 2306 8880 2414
rect 8800 2254 8814 2306
rect 8866 2254 8880 2306
rect 8800 2146 8880 2254
rect 8800 2094 8814 2146
rect 8866 2094 8880 2146
rect 8800 1986 8880 2094
rect 8800 1934 8814 1986
rect 8866 1934 8880 1986
rect 8800 1817 8880 1934
rect 8800 1783 8823 1817
rect 8857 1783 8880 1817
rect 8800 1666 8880 1783
rect 8800 1614 8814 1666
rect 8866 1614 8880 1666
rect 8800 1506 8880 1614
rect 8800 1454 8814 1506
rect 8866 1454 8880 1506
rect 8800 1346 8880 1454
rect 8800 1294 8814 1346
rect 8866 1294 8880 1346
rect 8800 1186 8880 1294
rect 8800 1134 8814 1186
rect 8866 1134 8880 1186
rect 8800 1026 8880 1134
rect 8800 974 8814 1026
rect 8866 974 8880 1026
rect 8800 857 8880 974
rect 8800 823 8823 857
rect 8857 823 8880 857
rect 8800 697 8880 823
rect 8800 663 8823 697
rect 8857 663 8880 697
rect 8800 546 8880 663
rect 8800 494 8814 546
rect 8866 494 8880 546
rect 8800 386 8880 494
rect 8800 334 8814 386
rect 8866 334 8880 386
rect 8800 226 8880 334
rect 8800 174 8814 226
rect 8866 174 8880 226
rect 8800 66 8880 174
rect 8800 14 8814 66
rect 8866 14 8880 66
rect 8800 0 8880 14
rect 8960 31426 9040 31440
rect 8960 31374 8974 31426
rect 9026 31374 9040 31426
rect 8960 31266 9040 31374
rect 8960 31214 8974 31266
rect 9026 31214 9040 31266
rect 8960 31106 9040 31214
rect 8960 31054 8974 31106
rect 9026 31054 9040 31106
rect 8960 30946 9040 31054
rect 8960 30894 8974 30946
rect 9026 30894 9040 30946
rect 8960 30786 9040 30894
rect 8960 30734 8974 30786
rect 9026 30734 9040 30786
rect 8960 30626 9040 30734
rect 8960 30574 8974 30626
rect 9026 30574 9040 30626
rect 8960 30466 9040 30574
rect 8960 30414 8974 30466
rect 9026 30414 9040 30466
rect 8960 30306 9040 30414
rect 8960 30254 8974 30306
rect 9026 30254 9040 30306
rect 8960 30137 9040 30254
rect 8960 30103 8983 30137
rect 9017 30103 9040 30137
rect 8960 29986 9040 30103
rect 8960 29934 8974 29986
rect 9026 29934 9040 29986
rect 8960 29826 9040 29934
rect 8960 29774 8974 29826
rect 9026 29774 9040 29826
rect 8960 29666 9040 29774
rect 8960 29614 8974 29666
rect 9026 29614 9040 29666
rect 8960 29506 9040 29614
rect 8960 29454 8974 29506
rect 9026 29454 9040 29506
rect 8960 29346 9040 29454
rect 8960 29294 8974 29346
rect 9026 29294 9040 29346
rect 8960 29186 9040 29294
rect 8960 29134 8974 29186
rect 9026 29134 9040 29186
rect 8960 29026 9040 29134
rect 8960 28974 8974 29026
rect 9026 28974 9040 29026
rect 8960 28866 9040 28974
rect 8960 28814 8974 28866
rect 9026 28814 9040 28866
rect 8960 28697 9040 28814
rect 8960 28663 8983 28697
rect 9017 28663 9040 28697
rect 8960 28537 9040 28663
rect 8960 28503 8983 28537
rect 9017 28503 9040 28537
rect 8960 28377 9040 28503
rect 8960 28343 8983 28377
rect 9017 28343 9040 28377
rect 8960 28217 9040 28343
rect 8960 28183 8983 28217
rect 9017 28183 9040 28217
rect 8960 28066 9040 28183
rect 8960 28014 8974 28066
rect 9026 28014 9040 28066
rect 8960 27906 9040 28014
rect 8960 27854 8974 27906
rect 9026 27854 9040 27906
rect 8960 27746 9040 27854
rect 8960 27694 8974 27746
rect 9026 27694 9040 27746
rect 8960 27586 9040 27694
rect 8960 27534 8974 27586
rect 9026 27534 9040 27586
rect 8960 27426 9040 27534
rect 8960 27374 8974 27426
rect 9026 27374 9040 27426
rect 8960 27266 9040 27374
rect 8960 27214 8974 27266
rect 9026 27214 9040 27266
rect 8960 27106 9040 27214
rect 8960 27054 8974 27106
rect 9026 27054 9040 27106
rect 8960 26946 9040 27054
rect 8960 26894 8974 26946
rect 9026 26894 9040 26946
rect 8960 26777 9040 26894
rect 8960 26743 8983 26777
rect 9017 26743 9040 26777
rect 8960 26617 9040 26743
rect 8960 26583 8983 26617
rect 9017 26583 9040 26617
rect 8960 26457 9040 26583
rect 8960 26423 8983 26457
rect 9017 26423 9040 26457
rect 8960 26297 9040 26423
rect 8960 26263 8983 26297
rect 9017 26263 9040 26297
rect 8960 26146 9040 26263
rect 8960 26094 8974 26146
rect 9026 26094 9040 26146
rect 8960 25986 9040 26094
rect 8960 25934 8974 25986
rect 9026 25934 9040 25986
rect 8960 25826 9040 25934
rect 8960 25774 8974 25826
rect 9026 25774 9040 25826
rect 8960 25666 9040 25774
rect 8960 25614 8974 25666
rect 9026 25614 9040 25666
rect 8960 25506 9040 25614
rect 8960 25454 8974 25506
rect 9026 25454 9040 25506
rect 8960 25346 9040 25454
rect 8960 25294 8974 25346
rect 9026 25294 9040 25346
rect 8960 25186 9040 25294
rect 8960 25134 8974 25186
rect 9026 25134 9040 25186
rect 8960 25026 9040 25134
rect 8960 24974 8974 25026
rect 9026 24974 9040 25026
rect 8960 24857 9040 24974
rect 8960 24823 8983 24857
rect 9017 24823 9040 24857
rect 8960 24706 9040 24823
rect 8960 24654 8974 24706
rect 9026 24654 9040 24706
rect 8960 24546 9040 24654
rect 8960 24494 8974 24546
rect 9026 24494 9040 24546
rect 8960 24386 9040 24494
rect 8960 24334 8974 24386
rect 9026 24334 9040 24386
rect 8960 24226 9040 24334
rect 8960 24174 8974 24226
rect 9026 24174 9040 24226
rect 8960 24066 9040 24174
rect 8960 24014 8974 24066
rect 9026 24014 9040 24066
rect 8960 23906 9040 24014
rect 8960 23854 8974 23906
rect 9026 23854 9040 23906
rect 8960 23746 9040 23854
rect 8960 23694 8974 23746
rect 9026 23694 9040 23746
rect 8960 23586 9040 23694
rect 8960 23534 8974 23586
rect 9026 23534 9040 23586
rect 8960 23426 9040 23534
rect 8960 23374 8974 23426
rect 9026 23374 9040 23426
rect 8960 23266 9040 23374
rect 8960 23214 8974 23266
rect 9026 23214 9040 23266
rect 8960 23106 9040 23214
rect 8960 23054 8974 23106
rect 9026 23054 9040 23106
rect 8960 22946 9040 23054
rect 8960 22894 8974 22946
rect 9026 22894 9040 22946
rect 8960 22786 9040 22894
rect 8960 22734 8974 22786
rect 9026 22734 9040 22786
rect 8960 22626 9040 22734
rect 8960 22574 8974 22626
rect 9026 22574 9040 22626
rect 8960 22466 9040 22574
rect 8960 22414 8974 22466
rect 9026 22414 9040 22466
rect 8960 22306 9040 22414
rect 8960 22254 8974 22306
rect 9026 22254 9040 22306
rect 8960 22146 9040 22254
rect 8960 22094 8974 22146
rect 9026 22094 9040 22146
rect 8960 21977 9040 22094
rect 8960 21943 8983 21977
rect 9017 21943 9040 21977
rect 8960 21826 9040 21943
rect 8960 21774 8974 21826
rect 9026 21774 9040 21826
rect 8960 21666 9040 21774
rect 8960 21614 8974 21666
rect 9026 21614 9040 21666
rect 8960 21506 9040 21614
rect 8960 21454 8974 21506
rect 9026 21454 9040 21506
rect 8960 21346 9040 21454
rect 8960 21294 8974 21346
rect 9026 21294 9040 21346
rect 8960 21186 9040 21294
rect 8960 21134 8974 21186
rect 9026 21134 9040 21186
rect 8960 21026 9040 21134
rect 8960 20974 8974 21026
rect 9026 20974 9040 21026
rect 8960 20866 9040 20974
rect 8960 20814 8974 20866
rect 9026 20814 9040 20866
rect 8960 20706 9040 20814
rect 8960 20654 8974 20706
rect 9026 20654 9040 20706
rect 8960 20537 9040 20654
rect 8960 20503 8983 20537
rect 9017 20503 9040 20537
rect 8960 20377 9040 20503
rect 8960 20343 8983 20377
rect 9017 20343 9040 20377
rect 8960 20217 9040 20343
rect 8960 20183 8983 20217
rect 9017 20183 9040 20217
rect 8960 20057 9040 20183
rect 8960 20023 8983 20057
rect 9017 20023 9040 20057
rect 8960 19906 9040 20023
rect 8960 19854 8974 19906
rect 9026 19854 9040 19906
rect 8960 19746 9040 19854
rect 8960 19694 8974 19746
rect 9026 19694 9040 19746
rect 8960 19586 9040 19694
rect 8960 19534 8974 19586
rect 9026 19534 9040 19586
rect 8960 19426 9040 19534
rect 8960 19374 8974 19426
rect 9026 19374 9040 19426
rect 8960 19266 9040 19374
rect 8960 19214 8974 19266
rect 9026 19214 9040 19266
rect 8960 19106 9040 19214
rect 8960 19054 8974 19106
rect 9026 19054 9040 19106
rect 8960 18946 9040 19054
rect 8960 18894 8974 18946
rect 9026 18894 9040 18946
rect 8960 18786 9040 18894
rect 8960 18734 8974 18786
rect 9026 18734 9040 18786
rect 8960 18617 9040 18734
rect 8960 18583 8983 18617
rect 9017 18583 9040 18617
rect 8960 18457 9040 18583
rect 8960 18423 8983 18457
rect 9017 18423 9040 18457
rect 8960 18297 9040 18423
rect 8960 18263 8983 18297
rect 9017 18263 9040 18297
rect 8960 18137 9040 18263
rect 8960 18103 8983 18137
rect 9017 18103 9040 18137
rect 8960 17986 9040 18103
rect 8960 17934 8974 17986
rect 9026 17934 9040 17986
rect 8960 17826 9040 17934
rect 8960 17774 8974 17826
rect 9026 17774 9040 17826
rect 8960 17666 9040 17774
rect 8960 17614 8974 17666
rect 9026 17614 9040 17666
rect 8960 17506 9040 17614
rect 8960 17454 8974 17506
rect 9026 17454 9040 17506
rect 8960 17346 9040 17454
rect 8960 17294 8974 17346
rect 9026 17294 9040 17346
rect 8960 17186 9040 17294
rect 8960 17134 8974 17186
rect 9026 17134 9040 17186
rect 8960 17026 9040 17134
rect 8960 16974 8974 17026
rect 9026 16974 9040 17026
rect 8960 16866 9040 16974
rect 8960 16814 8974 16866
rect 9026 16814 9040 16866
rect 8960 16697 9040 16814
rect 8960 16663 8983 16697
rect 9017 16663 9040 16697
rect 8960 16546 9040 16663
rect 8960 16494 8974 16546
rect 9026 16494 9040 16546
rect 8960 16386 9040 16494
rect 8960 16334 8974 16386
rect 9026 16334 9040 16386
rect 8960 16226 9040 16334
rect 8960 16174 8974 16226
rect 9026 16174 9040 16226
rect 8960 16066 9040 16174
rect 8960 16014 8974 16066
rect 9026 16014 9040 16066
rect 8960 15906 9040 16014
rect 8960 15854 8974 15906
rect 9026 15854 9040 15906
rect 8960 15746 9040 15854
rect 8960 15694 8974 15746
rect 9026 15694 9040 15746
rect 8960 15586 9040 15694
rect 8960 15534 8974 15586
rect 9026 15534 9040 15586
rect 8960 15426 9040 15534
rect 8960 15374 8974 15426
rect 9026 15374 9040 15426
rect 8960 15266 9040 15374
rect 8960 15214 8974 15266
rect 9026 15214 9040 15266
rect 8960 15106 9040 15214
rect 8960 15054 8974 15106
rect 9026 15054 9040 15106
rect 8960 14946 9040 15054
rect 8960 14894 8974 14946
rect 9026 14894 9040 14946
rect 8960 14786 9040 14894
rect 8960 14734 8974 14786
rect 9026 14734 9040 14786
rect 8960 14626 9040 14734
rect 8960 14574 8974 14626
rect 9026 14574 9040 14626
rect 8960 14466 9040 14574
rect 8960 14414 8974 14466
rect 9026 14414 9040 14466
rect 8960 14306 9040 14414
rect 8960 14254 8974 14306
rect 9026 14254 9040 14306
rect 8960 14146 9040 14254
rect 8960 14094 8974 14146
rect 9026 14094 9040 14146
rect 8960 13986 9040 14094
rect 8960 13934 8974 13986
rect 9026 13934 9040 13986
rect 8960 13817 9040 13934
rect 8960 13783 8983 13817
rect 9017 13783 9040 13817
rect 8960 13666 9040 13783
rect 8960 13614 8974 13666
rect 9026 13614 9040 13666
rect 8960 13506 9040 13614
rect 8960 13454 8974 13506
rect 9026 13454 9040 13506
rect 8960 13346 9040 13454
rect 8960 13294 8974 13346
rect 9026 13294 9040 13346
rect 8960 13186 9040 13294
rect 8960 13134 8974 13186
rect 9026 13134 9040 13186
rect 8960 13026 9040 13134
rect 8960 12974 8974 13026
rect 9026 12974 9040 13026
rect 8960 12866 9040 12974
rect 8960 12814 8974 12866
rect 9026 12814 9040 12866
rect 8960 12706 9040 12814
rect 8960 12654 8974 12706
rect 9026 12654 9040 12706
rect 8960 12546 9040 12654
rect 8960 12494 8974 12546
rect 9026 12494 9040 12546
rect 8960 12377 9040 12494
rect 8960 12343 8983 12377
rect 9017 12343 9040 12377
rect 8960 12217 9040 12343
rect 8960 12183 8983 12217
rect 9017 12183 9040 12217
rect 8960 12057 9040 12183
rect 8960 12023 8983 12057
rect 9017 12023 9040 12057
rect 8960 11897 9040 12023
rect 8960 11863 8983 11897
rect 9017 11863 9040 11897
rect 8960 11746 9040 11863
rect 8960 11694 8974 11746
rect 9026 11694 9040 11746
rect 8960 11586 9040 11694
rect 8960 11534 8974 11586
rect 9026 11534 9040 11586
rect 8960 11426 9040 11534
rect 8960 11374 8974 11426
rect 9026 11374 9040 11426
rect 8960 11266 9040 11374
rect 8960 11214 8974 11266
rect 9026 11214 9040 11266
rect 8960 11106 9040 11214
rect 8960 11054 8974 11106
rect 9026 11054 9040 11106
rect 8960 10946 9040 11054
rect 8960 10894 8974 10946
rect 9026 10894 9040 10946
rect 8960 10786 9040 10894
rect 8960 10734 8974 10786
rect 9026 10734 9040 10786
rect 8960 10626 9040 10734
rect 8960 10574 8974 10626
rect 9026 10574 9040 10626
rect 8960 10466 9040 10574
rect 8960 10414 8974 10466
rect 9026 10414 9040 10466
rect 8960 10306 9040 10414
rect 8960 10254 8974 10306
rect 9026 10254 9040 10306
rect 8960 10146 9040 10254
rect 8960 10094 8974 10146
rect 9026 10094 9040 10146
rect 8960 9986 9040 10094
rect 8960 9934 8974 9986
rect 9026 9934 9040 9986
rect 8960 9826 9040 9934
rect 8960 9774 8974 9826
rect 9026 9774 9040 9826
rect 8960 9657 9040 9774
rect 8960 9623 8983 9657
rect 9017 9623 9040 9657
rect 8960 9506 9040 9623
rect 8960 9454 8974 9506
rect 9026 9454 9040 9506
rect 8960 9346 9040 9454
rect 8960 9294 8974 9346
rect 9026 9294 9040 9346
rect 8960 9177 9040 9294
rect 8960 9143 8983 9177
rect 9017 9143 9040 9177
rect 8960 9026 9040 9143
rect 8960 8974 8974 9026
rect 9026 8974 9040 9026
rect 8960 8866 9040 8974
rect 8960 8814 8974 8866
rect 9026 8814 9040 8866
rect 8960 8706 9040 8814
rect 8960 8654 8974 8706
rect 9026 8654 9040 8706
rect 8960 8546 9040 8654
rect 8960 8494 8974 8546
rect 9026 8494 9040 8546
rect 8960 8386 9040 8494
rect 8960 8334 8974 8386
rect 9026 8334 9040 8386
rect 8960 8226 9040 8334
rect 8960 8174 8974 8226
rect 9026 8174 9040 8226
rect 8960 8066 9040 8174
rect 8960 8014 8974 8066
rect 9026 8014 9040 8066
rect 8960 7906 9040 8014
rect 8960 7854 8974 7906
rect 9026 7854 9040 7906
rect 8960 7746 9040 7854
rect 8960 7694 8974 7746
rect 9026 7694 9040 7746
rect 8960 7577 9040 7694
rect 8960 7543 8983 7577
rect 9017 7543 9040 7577
rect 8960 7426 9040 7543
rect 8960 7374 8974 7426
rect 9026 7374 9040 7426
rect 8960 7266 9040 7374
rect 8960 7214 8974 7266
rect 9026 7214 9040 7266
rect 8960 7097 9040 7214
rect 8960 7063 8983 7097
rect 9017 7063 9040 7097
rect 8960 6946 9040 7063
rect 8960 6894 8974 6946
rect 9026 6894 9040 6946
rect 8960 6786 9040 6894
rect 8960 6734 8974 6786
rect 9026 6734 9040 6786
rect 8960 6617 9040 6734
rect 8960 6583 8983 6617
rect 9017 6583 9040 6617
rect 8960 6466 9040 6583
rect 8960 6414 8974 6466
rect 9026 6414 9040 6466
rect 8960 6306 9040 6414
rect 8960 6254 8974 6306
rect 9026 6254 9040 6306
rect 8960 6146 9040 6254
rect 8960 6094 8974 6146
rect 9026 6094 9040 6146
rect 8960 5986 9040 6094
rect 8960 5934 8974 5986
rect 9026 5934 9040 5986
rect 8960 5826 9040 5934
rect 8960 5774 8974 5826
rect 9026 5774 9040 5826
rect 8960 5666 9040 5774
rect 8960 5614 8974 5666
rect 9026 5614 9040 5666
rect 8960 5506 9040 5614
rect 8960 5454 8974 5506
rect 9026 5454 9040 5506
rect 8960 5346 9040 5454
rect 8960 5294 8974 5346
rect 9026 5294 9040 5346
rect 8960 5186 9040 5294
rect 8960 5134 8974 5186
rect 9026 5134 9040 5186
rect 8960 5026 9040 5134
rect 8960 4974 8974 5026
rect 9026 4974 9040 5026
rect 8960 4866 9040 4974
rect 8960 4814 8974 4866
rect 9026 4814 9040 4866
rect 8960 4706 9040 4814
rect 8960 4654 8974 4706
rect 9026 4654 9040 4706
rect 8960 4546 9040 4654
rect 8960 4494 8974 4546
rect 9026 4494 9040 4546
rect 8960 4386 9040 4494
rect 8960 4334 8974 4386
rect 9026 4334 9040 4386
rect 8960 4226 9040 4334
rect 8960 4174 8974 4226
rect 9026 4174 9040 4226
rect 8960 4066 9040 4174
rect 8960 4014 8974 4066
rect 9026 4014 9040 4066
rect 8960 3906 9040 4014
rect 8960 3854 8974 3906
rect 9026 3854 9040 3906
rect 8960 3737 9040 3854
rect 8960 3703 8983 3737
rect 9017 3703 9040 3737
rect 8960 3577 9040 3703
rect 8960 3543 8983 3577
rect 9017 3543 9040 3577
rect 8960 3426 9040 3543
rect 8960 3374 8974 3426
rect 9026 3374 9040 3426
rect 8960 3266 9040 3374
rect 8960 3214 8974 3266
rect 9026 3214 9040 3266
rect 8960 3106 9040 3214
rect 8960 3054 8974 3106
rect 9026 3054 9040 3106
rect 8960 2946 9040 3054
rect 8960 2894 8974 2946
rect 9026 2894 9040 2946
rect 8960 2786 9040 2894
rect 8960 2734 8974 2786
rect 9026 2734 9040 2786
rect 8960 2626 9040 2734
rect 8960 2574 8974 2626
rect 9026 2574 9040 2626
rect 8960 2466 9040 2574
rect 8960 2414 8974 2466
rect 9026 2414 9040 2466
rect 8960 2306 9040 2414
rect 8960 2254 8974 2306
rect 9026 2254 9040 2306
rect 8960 2146 9040 2254
rect 8960 2094 8974 2146
rect 9026 2094 9040 2146
rect 8960 1986 9040 2094
rect 8960 1934 8974 1986
rect 9026 1934 9040 1986
rect 8960 1817 9040 1934
rect 8960 1783 8983 1817
rect 9017 1783 9040 1817
rect 8960 1666 9040 1783
rect 8960 1614 8974 1666
rect 9026 1614 9040 1666
rect 8960 1506 9040 1614
rect 8960 1454 8974 1506
rect 9026 1454 9040 1506
rect 8960 1346 9040 1454
rect 8960 1294 8974 1346
rect 9026 1294 9040 1346
rect 8960 1186 9040 1294
rect 8960 1134 8974 1186
rect 9026 1134 9040 1186
rect 8960 1026 9040 1134
rect 8960 974 8974 1026
rect 9026 974 9040 1026
rect 8960 857 9040 974
rect 8960 823 8983 857
rect 9017 823 9040 857
rect 8960 697 9040 823
rect 8960 663 8983 697
rect 9017 663 9040 697
rect 8960 546 9040 663
rect 8960 494 8974 546
rect 9026 494 9040 546
rect 8960 386 9040 494
rect 8960 334 8974 386
rect 9026 334 9040 386
rect 8960 226 9040 334
rect 8960 174 8974 226
rect 9026 174 9040 226
rect 8960 66 9040 174
rect 8960 14 8974 66
rect 9026 14 9040 66
rect 8960 0 9040 14
rect 9120 31417 9200 31440
rect 9120 31383 9143 31417
rect 9177 31383 9200 31417
rect 9120 31257 9200 31383
rect 9120 31223 9143 31257
rect 9177 31223 9200 31257
rect 9120 31097 9200 31223
rect 9120 31063 9143 31097
rect 9177 31063 9200 31097
rect 9120 30937 9200 31063
rect 9120 30903 9143 30937
rect 9177 30903 9200 30937
rect 9120 30777 9200 30903
rect 9120 30743 9143 30777
rect 9177 30743 9200 30777
rect 9120 30617 9200 30743
rect 9120 30583 9143 30617
rect 9177 30583 9200 30617
rect 9120 30457 9200 30583
rect 9120 30423 9143 30457
rect 9177 30423 9200 30457
rect 9120 30297 9200 30423
rect 9120 30263 9143 30297
rect 9177 30263 9200 30297
rect 9120 30137 9200 30263
rect 9120 30103 9143 30137
rect 9177 30103 9200 30137
rect 9120 29977 9200 30103
rect 9120 29943 9143 29977
rect 9177 29943 9200 29977
rect 9120 29817 9200 29943
rect 9120 29783 9143 29817
rect 9177 29783 9200 29817
rect 9120 29657 9200 29783
rect 9120 29623 9143 29657
rect 9177 29623 9200 29657
rect 9120 29497 9200 29623
rect 9120 29463 9143 29497
rect 9177 29463 9200 29497
rect 9120 29337 9200 29463
rect 9120 29303 9143 29337
rect 9177 29303 9200 29337
rect 9120 29177 9200 29303
rect 9120 29143 9143 29177
rect 9177 29143 9200 29177
rect 9120 29017 9200 29143
rect 9120 28983 9143 29017
rect 9177 28983 9200 29017
rect 9120 28857 9200 28983
rect 9120 28823 9143 28857
rect 9177 28823 9200 28857
rect 9120 28697 9200 28823
rect 9120 28663 9143 28697
rect 9177 28663 9200 28697
rect 9120 28537 9200 28663
rect 9120 28503 9143 28537
rect 9177 28503 9200 28537
rect 9120 28377 9200 28503
rect 9120 28343 9143 28377
rect 9177 28343 9200 28377
rect 9120 28217 9200 28343
rect 9120 28183 9143 28217
rect 9177 28183 9200 28217
rect 9120 28057 9200 28183
rect 9120 28023 9143 28057
rect 9177 28023 9200 28057
rect 9120 27897 9200 28023
rect 9120 27863 9143 27897
rect 9177 27863 9200 27897
rect 9120 27737 9200 27863
rect 9120 27703 9143 27737
rect 9177 27703 9200 27737
rect 9120 27577 9200 27703
rect 9120 27543 9143 27577
rect 9177 27543 9200 27577
rect 9120 27417 9200 27543
rect 9120 27383 9143 27417
rect 9177 27383 9200 27417
rect 9120 27257 9200 27383
rect 9120 27223 9143 27257
rect 9177 27223 9200 27257
rect 9120 27097 9200 27223
rect 9120 27063 9143 27097
rect 9177 27063 9200 27097
rect 9120 26937 9200 27063
rect 9120 26903 9143 26937
rect 9177 26903 9200 26937
rect 9120 26777 9200 26903
rect 9120 26743 9143 26777
rect 9177 26743 9200 26777
rect 9120 26617 9200 26743
rect 9120 26583 9143 26617
rect 9177 26583 9200 26617
rect 9120 26457 9200 26583
rect 9120 26423 9143 26457
rect 9177 26423 9200 26457
rect 9120 26297 9200 26423
rect 9120 26263 9143 26297
rect 9177 26263 9200 26297
rect 9120 26137 9200 26263
rect 9120 26103 9143 26137
rect 9177 26103 9200 26137
rect 9120 25977 9200 26103
rect 9120 25943 9143 25977
rect 9177 25943 9200 25977
rect 9120 25817 9200 25943
rect 9120 25783 9143 25817
rect 9177 25783 9200 25817
rect 9120 25657 9200 25783
rect 9120 25623 9143 25657
rect 9177 25623 9200 25657
rect 9120 25497 9200 25623
rect 9120 25463 9143 25497
rect 9177 25463 9200 25497
rect 9120 25337 9200 25463
rect 9120 25303 9143 25337
rect 9177 25303 9200 25337
rect 9120 25177 9200 25303
rect 9120 25143 9143 25177
rect 9177 25143 9200 25177
rect 9120 25017 9200 25143
rect 9120 24983 9143 25017
rect 9177 24983 9200 25017
rect 9120 24857 9200 24983
rect 9120 24823 9143 24857
rect 9177 24823 9200 24857
rect 9120 24697 9200 24823
rect 9120 24663 9143 24697
rect 9177 24663 9200 24697
rect 9120 24537 9200 24663
rect 9120 24503 9143 24537
rect 9177 24503 9200 24537
rect 9120 24377 9200 24503
rect 9120 24343 9143 24377
rect 9177 24343 9200 24377
rect 9120 24217 9200 24343
rect 9120 24183 9143 24217
rect 9177 24183 9200 24217
rect 9120 24057 9200 24183
rect 9120 24023 9143 24057
rect 9177 24023 9200 24057
rect 9120 23897 9200 24023
rect 9120 23863 9143 23897
rect 9177 23863 9200 23897
rect 9120 23737 9200 23863
rect 9120 23703 9143 23737
rect 9177 23703 9200 23737
rect 9120 23577 9200 23703
rect 9120 23543 9143 23577
rect 9177 23543 9200 23577
rect 9120 23417 9200 23543
rect 9120 23383 9143 23417
rect 9177 23383 9200 23417
rect 9120 23257 9200 23383
rect 9120 23223 9143 23257
rect 9177 23223 9200 23257
rect 9120 23097 9200 23223
rect 9120 23063 9143 23097
rect 9177 23063 9200 23097
rect 9120 22937 9200 23063
rect 9120 22903 9143 22937
rect 9177 22903 9200 22937
rect 9120 22777 9200 22903
rect 9120 22743 9143 22777
rect 9177 22743 9200 22777
rect 9120 22617 9200 22743
rect 9120 22583 9143 22617
rect 9177 22583 9200 22617
rect 9120 22457 9200 22583
rect 9120 22423 9143 22457
rect 9177 22423 9200 22457
rect 9120 22297 9200 22423
rect 9120 22263 9143 22297
rect 9177 22263 9200 22297
rect 9120 22137 9200 22263
rect 9120 22103 9143 22137
rect 9177 22103 9200 22137
rect 9120 21977 9200 22103
rect 9120 21943 9143 21977
rect 9177 21943 9200 21977
rect 9120 21817 9200 21943
rect 9120 21783 9143 21817
rect 9177 21783 9200 21817
rect 9120 21657 9200 21783
rect 9120 21623 9143 21657
rect 9177 21623 9200 21657
rect 9120 21497 9200 21623
rect 9120 21463 9143 21497
rect 9177 21463 9200 21497
rect 9120 21337 9200 21463
rect 9120 21303 9143 21337
rect 9177 21303 9200 21337
rect 9120 21177 9200 21303
rect 9120 21143 9143 21177
rect 9177 21143 9200 21177
rect 9120 21017 9200 21143
rect 9120 20983 9143 21017
rect 9177 20983 9200 21017
rect 9120 20857 9200 20983
rect 9120 20823 9143 20857
rect 9177 20823 9200 20857
rect 9120 20697 9200 20823
rect 9120 20663 9143 20697
rect 9177 20663 9200 20697
rect 9120 20537 9200 20663
rect 9120 20503 9143 20537
rect 9177 20503 9200 20537
rect 9120 20377 9200 20503
rect 9120 20343 9143 20377
rect 9177 20343 9200 20377
rect 9120 20217 9200 20343
rect 9120 20183 9143 20217
rect 9177 20183 9200 20217
rect 9120 20057 9200 20183
rect 9120 20023 9143 20057
rect 9177 20023 9200 20057
rect 9120 19897 9200 20023
rect 9120 19863 9143 19897
rect 9177 19863 9200 19897
rect 9120 19737 9200 19863
rect 9120 19703 9143 19737
rect 9177 19703 9200 19737
rect 9120 19577 9200 19703
rect 9120 19543 9143 19577
rect 9177 19543 9200 19577
rect 9120 19417 9200 19543
rect 9120 19383 9143 19417
rect 9177 19383 9200 19417
rect 9120 19257 9200 19383
rect 9120 19223 9143 19257
rect 9177 19223 9200 19257
rect 9120 19097 9200 19223
rect 9120 19063 9143 19097
rect 9177 19063 9200 19097
rect 9120 18937 9200 19063
rect 9120 18903 9143 18937
rect 9177 18903 9200 18937
rect 9120 18777 9200 18903
rect 9120 18743 9143 18777
rect 9177 18743 9200 18777
rect 9120 18617 9200 18743
rect 9120 18583 9143 18617
rect 9177 18583 9200 18617
rect 9120 18457 9200 18583
rect 9120 18423 9143 18457
rect 9177 18423 9200 18457
rect 9120 18297 9200 18423
rect 9120 18263 9143 18297
rect 9177 18263 9200 18297
rect 9120 18137 9200 18263
rect 9120 18103 9143 18137
rect 9177 18103 9200 18137
rect 9120 17977 9200 18103
rect 9120 17943 9143 17977
rect 9177 17943 9200 17977
rect 9120 17817 9200 17943
rect 9120 17783 9143 17817
rect 9177 17783 9200 17817
rect 9120 17657 9200 17783
rect 9120 17623 9143 17657
rect 9177 17623 9200 17657
rect 9120 17497 9200 17623
rect 9120 17463 9143 17497
rect 9177 17463 9200 17497
rect 9120 17337 9200 17463
rect 9120 17303 9143 17337
rect 9177 17303 9200 17337
rect 9120 17177 9200 17303
rect 9120 17143 9143 17177
rect 9177 17143 9200 17177
rect 9120 17017 9200 17143
rect 9120 16983 9143 17017
rect 9177 16983 9200 17017
rect 9120 16857 9200 16983
rect 9120 16823 9143 16857
rect 9177 16823 9200 16857
rect 9120 16697 9200 16823
rect 9120 16663 9143 16697
rect 9177 16663 9200 16697
rect 9120 16537 9200 16663
rect 9120 16503 9143 16537
rect 9177 16503 9200 16537
rect 9120 16377 9200 16503
rect 9120 16343 9143 16377
rect 9177 16343 9200 16377
rect 9120 16217 9200 16343
rect 9120 16183 9143 16217
rect 9177 16183 9200 16217
rect 9120 16057 9200 16183
rect 9120 16023 9143 16057
rect 9177 16023 9200 16057
rect 9120 15897 9200 16023
rect 9120 15863 9143 15897
rect 9177 15863 9200 15897
rect 9120 15737 9200 15863
rect 9120 15703 9143 15737
rect 9177 15703 9200 15737
rect 9120 15577 9200 15703
rect 9120 15543 9143 15577
rect 9177 15543 9200 15577
rect 9120 15417 9200 15543
rect 9120 15383 9143 15417
rect 9177 15383 9200 15417
rect 9120 15257 9200 15383
rect 9120 15223 9143 15257
rect 9177 15223 9200 15257
rect 9120 15097 9200 15223
rect 9120 15063 9143 15097
rect 9177 15063 9200 15097
rect 9120 14937 9200 15063
rect 9120 14903 9143 14937
rect 9177 14903 9200 14937
rect 9120 14777 9200 14903
rect 9120 14743 9143 14777
rect 9177 14743 9200 14777
rect 9120 14617 9200 14743
rect 9120 14583 9143 14617
rect 9177 14583 9200 14617
rect 9120 14457 9200 14583
rect 9120 14423 9143 14457
rect 9177 14423 9200 14457
rect 9120 14297 9200 14423
rect 9120 14263 9143 14297
rect 9177 14263 9200 14297
rect 9120 14137 9200 14263
rect 9120 14103 9143 14137
rect 9177 14103 9200 14137
rect 9120 13977 9200 14103
rect 9120 13943 9143 13977
rect 9177 13943 9200 13977
rect 9120 13817 9200 13943
rect 9120 13783 9143 13817
rect 9177 13783 9200 13817
rect 9120 13657 9200 13783
rect 9120 13623 9143 13657
rect 9177 13623 9200 13657
rect 9120 13497 9200 13623
rect 9120 13463 9143 13497
rect 9177 13463 9200 13497
rect 9120 13337 9200 13463
rect 9120 13303 9143 13337
rect 9177 13303 9200 13337
rect 9120 13177 9200 13303
rect 9120 13143 9143 13177
rect 9177 13143 9200 13177
rect 9120 13017 9200 13143
rect 9120 12983 9143 13017
rect 9177 12983 9200 13017
rect 9120 12857 9200 12983
rect 9120 12823 9143 12857
rect 9177 12823 9200 12857
rect 9120 12697 9200 12823
rect 9120 12663 9143 12697
rect 9177 12663 9200 12697
rect 9120 12537 9200 12663
rect 9120 12503 9143 12537
rect 9177 12503 9200 12537
rect 9120 12377 9200 12503
rect 9120 12343 9143 12377
rect 9177 12343 9200 12377
rect 9120 12217 9200 12343
rect 9120 12183 9143 12217
rect 9177 12183 9200 12217
rect 9120 12057 9200 12183
rect 9120 12023 9143 12057
rect 9177 12023 9200 12057
rect 9120 11897 9200 12023
rect 9120 11863 9143 11897
rect 9177 11863 9200 11897
rect 9120 11737 9200 11863
rect 9120 11703 9143 11737
rect 9177 11703 9200 11737
rect 9120 11577 9200 11703
rect 9120 11543 9143 11577
rect 9177 11543 9200 11577
rect 9120 11417 9200 11543
rect 9120 11383 9143 11417
rect 9177 11383 9200 11417
rect 9120 11257 9200 11383
rect 9120 11223 9143 11257
rect 9177 11223 9200 11257
rect 9120 11097 9200 11223
rect 9120 11063 9143 11097
rect 9177 11063 9200 11097
rect 9120 10937 9200 11063
rect 9120 10903 9143 10937
rect 9177 10903 9200 10937
rect 9120 10777 9200 10903
rect 9120 10743 9143 10777
rect 9177 10743 9200 10777
rect 9120 10617 9200 10743
rect 9120 10583 9143 10617
rect 9177 10583 9200 10617
rect 9120 10457 9200 10583
rect 9120 10423 9143 10457
rect 9177 10423 9200 10457
rect 9120 10297 9200 10423
rect 9120 10263 9143 10297
rect 9177 10263 9200 10297
rect 9120 10137 9200 10263
rect 9120 10103 9143 10137
rect 9177 10103 9200 10137
rect 9120 9977 9200 10103
rect 9120 9943 9143 9977
rect 9177 9943 9200 9977
rect 9120 9817 9200 9943
rect 9120 9783 9143 9817
rect 9177 9783 9200 9817
rect 9120 9657 9200 9783
rect 9120 9623 9143 9657
rect 9177 9623 9200 9657
rect 9120 9497 9200 9623
rect 9120 9463 9143 9497
rect 9177 9463 9200 9497
rect 9120 9337 9200 9463
rect 9120 9303 9143 9337
rect 9177 9303 9200 9337
rect 9120 9177 9200 9303
rect 9120 9143 9143 9177
rect 9177 9143 9200 9177
rect 9120 9017 9200 9143
rect 9120 8983 9143 9017
rect 9177 8983 9200 9017
rect 9120 8857 9200 8983
rect 9120 8823 9143 8857
rect 9177 8823 9200 8857
rect 9120 8697 9200 8823
rect 9120 8663 9143 8697
rect 9177 8663 9200 8697
rect 9120 8537 9200 8663
rect 9120 8503 9143 8537
rect 9177 8503 9200 8537
rect 9120 8377 9200 8503
rect 9120 8343 9143 8377
rect 9177 8343 9200 8377
rect 9120 8217 9200 8343
rect 9120 8183 9143 8217
rect 9177 8183 9200 8217
rect 9120 8057 9200 8183
rect 9120 8023 9143 8057
rect 9177 8023 9200 8057
rect 9120 7897 9200 8023
rect 9120 7863 9143 7897
rect 9177 7863 9200 7897
rect 9120 7737 9200 7863
rect 9120 7703 9143 7737
rect 9177 7703 9200 7737
rect 9120 7577 9200 7703
rect 9120 7543 9143 7577
rect 9177 7543 9200 7577
rect 9120 7417 9200 7543
rect 9120 7383 9143 7417
rect 9177 7383 9200 7417
rect 9120 7257 9200 7383
rect 9120 7223 9143 7257
rect 9177 7223 9200 7257
rect 9120 7097 9200 7223
rect 9120 7063 9143 7097
rect 9177 7063 9200 7097
rect 9120 6937 9200 7063
rect 9120 6903 9143 6937
rect 9177 6903 9200 6937
rect 9120 6777 9200 6903
rect 9120 6743 9143 6777
rect 9177 6743 9200 6777
rect 9120 6617 9200 6743
rect 9120 6583 9143 6617
rect 9177 6583 9200 6617
rect 9120 6457 9200 6583
rect 9120 6423 9143 6457
rect 9177 6423 9200 6457
rect 9120 6297 9200 6423
rect 9120 6263 9143 6297
rect 9177 6263 9200 6297
rect 9120 6137 9200 6263
rect 9120 6103 9143 6137
rect 9177 6103 9200 6137
rect 9120 5977 9200 6103
rect 9120 5943 9143 5977
rect 9177 5943 9200 5977
rect 9120 5817 9200 5943
rect 9120 5783 9143 5817
rect 9177 5783 9200 5817
rect 9120 5657 9200 5783
rect 9120 5623 9143 5657
rect 9177 5623 9200 5657
rect 9120 5497 9200 5623
rect 9120 5463 9143 5497
rect 9177 5463 9200 5497
rect 9120 5337 9200 5463
rect 9120 5303 9143 5337
rect 9177 5303 9200 5337
rect 9120 5177 9200 5303
rect 9120 5143 9143 5177
rect 9177 5143 9200 5177
rect 9120 5017 9200 5143
rect 9120 4983 9143 5017
rect 9177 4983 9200 5017
rect 9120 4857 9200 4983
rect 9120 4823 9143 4857
rect 9177 4823 9200 4857
rect 9120 4697 9200 4823
rect 9120 4663 9143 4697
rect 9177 4663 9200 4697
rect 9120 4537 9200 4663
rect 9120 4503 9143 4537
rect 9177 4503 9200 4537
rect 9120 4377 9200 4503
rect 9120 4343 9143 4377
rect 9177 4343 9200 4377
rect 9120 4217 9200 4343
rect 9120 4183 9143 4217
rect 9177 4183 9200 4217
rect 9120 4057 9200 4183
rect 9120 4023 9143 4057
rect 9177 4023 9200 4057
rect 9120 3897 9200 4023
rect 9120 3863 9143 3897
rect 9177 3863 9200 3897
rect 9120 3737 9200 3863
rect 9120 3703 9143 3737
rect 9177 3703 9200 3737
rect 9120 3577 9200 3703
rect 9120 3543 9143 3577
rect 9177 3543 9200 3577
rect 9120 3417 9200 3543
rect 9120 3383 9143 3417
rect 9177 3383 9200 3417
rect 9120 3257 9200 3383
rect 9120 3223 9143 3257
rect 9177 3223 9200 3257
rect 9120 3097 9200 3223
rect 9120 3063 9143 3097
rect 9177 3063 9200 3097
rect 9120 2937 9200 3063
rect 9120 2903 9143 2937
rect 9177 2903 9200 2937
rect 9120 2777 9200 2903
rect 9120 2743 9143 2777
rect 9177 2743 9200 2777
rect 9120 2617 9200 2743
rect 9120 2583 9143 2617
rect 9177 2583 9200 2617
rect 9120 2457 9200 2583
rect 9120 2423 9143 2457
rect 9177 2423 9200 2457
rect 9120 2297 9200 2423
rect 9120 2263 9143 2297
rect 9177 2263 9200 2297
rect 9120 2137 9200 2263
rect 9120 2103 9143 2137
rect 9177 2103 9200 2137
rect 9120 1977 9200 2103
rect 9120 1943 9143 1977
rect 9177 1943 9200 1977
rect 9120 1817 9200 1943
rect 9120 1783 9143 1817
rect 9177 1783 9200 1817
rect 9120 1657 9200 1783
rect 9120 1623 9143 1657
rect 9177 1623 9200 1657
rect 9120 1497 9200 1623
rect 9120 1463 9143 1497
rect 9177 1463 9200 1497
rect 9120 1337 9200 1463
rect 9120 1303 9143 1337
rect 9177 1303 9200 1337
rect 9120 1177 9200 1303
rect 9120 1143 9143 1177
rect 9177 1143 9200 1177
rect 9120 1017 9200 1143
rect 9120 983 9143 1017
rect 9177 983 9200 1017
rect 9120 857 9200 983
rect 9120 823 9143 857
rect 9177 823 9200 857
rect 9120 697 9200 823
rect 9120 663 9143 697
rect 9177 663 9200 697
rect 9120 537 9200 663
rect 9120 503 9143 537
rect 9177 503 9200 537
rect 9120 377 9200 503
rect 9120 343 9143 377
rect 9177 343 9200 377
rect 9120 217 9200 343
rect 9120 183 9143 217
rect 9177 183 9200 217
rect 9120 57 9200 183
rect 9120 23 9143 57
rect 9177 23 9200 57
rect 9120 0 9200 23
rect 9280 31426 9360 31440
rect 9280 31374 9294 31426
rect 9346 31374 9360 31426
rect 9280 31266 9360 31374
rect 9280 31214 9294 31266
rect 9346 31214 9360 31266
rect 9280 31106 9360 31214
rect 9280 31054 9294 31106
rect 9346 31054 9360 31106
rect 9280 30946 9360 31054
rect 9280 30894 9294 30946
rect 9346 30894 9360 30946
rect 9280 30786 9360 30894
rect 9280 30734 9294 30786
rect 9346 30734 9360 30786
rect 9280 30626 9360 30734
rect 9280 30574 9294 30626
rect 9346 30574 9360 30626
rect 9280 30466 9360 30574
rect 9280 30414 9294 30466
rect 9346 30414 9360 30466
rect 9280 30306 9360 30414
rect 9280 30254 9294 30306
rect 9346 30254 9360 30306
rect 9280 30137 9360 30254
rect 9280 30103 9303 30137
rect 9337 30103 9360 30137
rect 9280 29986 9360 30103
rect 9280 29934 9294 29986
rect 9346 29934 9360 29986
rect 9280 29826 9360 29934
rect 9280 29774 9294 29826
rect 9346 29774 9360 29826
rect 9280 29666 9360 29774
rect 9280 29614 9294 29666
rect 9346 29614 9360 29666
rect 9280 29506 9360 29614
rect 9280 29454 9294 29506
rect 9346 29454 9360 29506
rect 9280 29346 9360 29454
rect 9280 29294 9294 29346
rect 9346 29294 9360 29346
rect 9280 29186 9360 29294
rect 9280 29134 9294 29186
rect 9346 29134 9360 29186
rect 9280 29026 9360 29134
rect 9280 28974 9294 29026
rect 9346 28974 9360 29026
rect 9280 28866 9360 28974
rect 9280 28814 9294 28866
rect 9346 28814 9360 28866
rect 9280 28697 9360 28814
rect 9280 28663 9303 28697
rect 9337 28663 9360 28697
rect 9280 28537 9360 28663
rect 9280 28503 9303 28537
rect 9337 28503 9360 28537
rect 9280 28377 9360 28503
rect 9280 28343 9303 28377
rect 9337 28343 9360 28377
rect 9280 28217 9360 28343
rect 9280 28183 9303 28217
rect 9337 28183 9360 28217
rect 9280 28066 9360 28183
rect 9280 28014 9294 28066
rect 9346 28014 9360 28066
rect 9280 27906 9360 28014
rect 9280 27854 9294 27906
rect 9346 27854 9360 27906
rect 9280 27746 9360 27854
rect 9280 27694 9294 27746
rect 9346 27694 9360 27746
rect 9280 27586 9360 27694
rect 9280 27534 9294 27586
rect 9346 27534 9360 27586
rect 9280 27426 9360 27534
rect 9280 27374 9294 27426
rect 9346 27374 9360 27426
rect 9280 27266 9360 27374
rect 9280 27214 9294 27266
rect 9346 27214 9360 27266
rect 9280 27106 9360 27214
rect 9280 27054 9294 27106
rect 9346 27054 9360 27106
rect 9280 26946 9360 27054
rect 9280 26894 9294 26946
rect 9346 26894 9360 26946
rect 9280 26777 9360 26894
rect 9280 26743 9303 26777
rect 9337 26743 9360 26777
rect 9280 26617 9360 26743
rect 9280 26583 9303 26617
rect 9337 26583 9360 26617
rect 9280 26457 9360 26583
rect 9280 26423 9303 26457
rect 9337 26423 9360 26457
rect 9280 26297 9360 26423
rect 9280 26263 9303 26297
rect 9337 26263 9360 26297
rect 9280 26146 9360 26263
rect 9280 26094 9294 26146
rect 9346 26094 9360 26146
rect 9280 25986 9360 26094
rect 9280 25934 9294 25986
rect 9346 25934 9360 25986
rect 9280 25826 9360 25934
rect 9280 25774 9294 25826
rect 9346 25774 9360 25826
rect 9280 25666 9360 25774
rect 9280 25614 9294 25666
rect 9346 25614 9360 25666
rect 9280 25506 9360 25614
rect 9280 25454 9294 25506
rect 9346 25454 9360 25506
rect 9280 25346 9360 25454
rect 9280 25294 9294 25346
rect 9346 25294 9360 25346
rect 9280 25186 9360 25294
rect 9280 25134 9294 25186
rect 9346 25134 9360 25186
rect 9280 25026 9360 25134
rect 9280 24974 9294 25026
rect 9346 24974 9360 25026
rect 9280 24857 9360 24974
rect 9280 24823 9303 24857
rect 9337 24823 9360 24857
rect 9280 24706 9360 24823
rect 9280 24654 9294 24706
rect 9346 24654 9360 24706
rect 9280 24546 9360 24654
rect 9280 24494 9294 24546
rect 9346 24494 9360 24546
rect 9280 24386 9360 24494
rect 9280 24334 9294 24386
rect 9346 24334 9360 24386
rect 9280 24226 9360 24334
rect 9280 24174 9294 24226
rect 9346 24174 9360 24226
rect 9280 24066 9360 24174
rect 9280 24014 9294 24066
rect 9346 24014 9360 24066
rect 9280 23906 9360 24014
rect 9280 23854 9294 23906
rect 9346 23854 9360 23906
rect 9280 23746 9360 23854
rect 9280 23694 9294 23746
rect 9346 23694 9360 23746
rect 9280 23586 9360 23694
rect 9280 23534 9294 23586
rect 9346 23534 9360 23586
rect 9280 23426 9360 23534
rect 9280 23374 9294 23426
rect 9346 23374 9360 23426
rect 9280 23266 9360 23374
rect 9280 23214 9294 23266
rect 9346 23214 9360 23266
rect 9280 23106 9360 23214
rect 9280 23054 9294 23106
rect 9346 23054 9360 23106
rect 9280 22946 9360 23054
rect 9280 22894 9294 22946
rect 9346 22894 9360 22946
rect 9280 22786 9360 22894
rect 9280 22734 9294 22786
rect 9346 22734 9360 22786
rect 9280 22626 9360 22734
rect 9280 22574 9294 22626
rect 9346 22574 9360 22626
rect 9280 22466 9360 22574
rect 9280 22414 9294 22466
rect 9346 22414 9360 22466
rect 9280 22306 9360 22414
rect 9280 22254 9294 22306
rect 9346 22254 9360 22306
rect 9280 22146 9360 22254
rect 9280 22094 9294 22146
rect 9346 22094 9360 22146
rect 9280 21977 9360 22094
rect 9280 21943 9303 21977
rect 9337 21943 9360 21977
rect 9280 21826 9360 21943
rect 9280 21774 9294 21826
rect 9346 21774 9360 21826
rect 9280 21666 9360 21774
rect 9280 21614 9294 21666
rect 9346 21614 9360 21666
rect 9280 21506 9360 21614
rect 9280 21454 9294 21506
rect 9346 21454 9360 21506
rect 9280 21346 9360 21454
rect 9280 21294 9294 21346
rect 9346 21294 9360 21346
rect 9280 21186 9360 21294
rect 9280 21134 9294 21186
rect 9346 21134 9360 21186
rect 9280 21026 9360 21134
rect 9280 20974 9294 21026
rect 9346 20974 9360 21026
rect 9280 20866 9360 20974
rect 9280 20814 9294 20866
rect 9346 20814 9360 20866
rect 9280 20706 9360 20814
rect 9280 20654 9294 20706
rect 9346 20654 9360 20706
rect 9280 20537 9360 20654
rect 9280 20503 9303 20537
rect 9337 20503 9360 20537
rect 9280 20377 9360 20503
rect 9280 20343 9303 20377
rect 9337 20343 9360 20377
rect 9280 20217 9360 20343
rect 9280 20183 9303 20217
rect 9337 20183 9360 20217
rect 9280 20057 9360 20183
rect 9280 20023 9303 20057
rect 9337 20023 9360 20057
rect 9280 19906 9360 20023
rect 9280 19854 9294 19906
rect 9346 19854 9360 19906
rect 9280 19746 9360 19854
rect 9280 19694 9294 19746
rect 9346 19694 9360 19746
rect 9280 19586 9360 19694
rect 9280 19534 9294 19586
rect 9346 19534 9360 19586
rect 9280 19426 9360 19534
rect 9280 19374 9294 19426
rect 9346 19374 9360 19426
rect 9280 19266 9360 19374
rect 9280 19214 9294 19266
rect 9346 19214 9360 19266
rect 9280 19106 9360 19214
rect 9280 19054 9294 19106
rect 9346 19054 9360 19106
rect 9280 18946 9360 19054
rect 9280 18894 9294 18946
rect 9346 18894 9360 18946
rect 9280 18786 9360 18894
rect 9280 18734 9294 18786
rect 9346 18734 9360 18786
rect 9280 18617 9360 18734
rect 9280 18583 9303 18617
rect 9337 18583 9360 18617
rect 9280 18457 9360 18583
rect 9280 18423 9303 18457
rect 9337 18423 9360 18457
rect 9280 18297 9360 18423
rect 9280 18263 9303 18297
rect 9337 18263 9360 18297
rect 9280 18137 9360 18263
rect 9280 18103 9303 18137
rect 9337 18103 9360 18137
rect 9280 17986 9360 18103
rect 9280 17934 9294 17986
rect 9346 17934 9360 17986
rect 9280 17826 9360 17934
rect 9280 17774 9294 17826
rect 9346 17774 9360 17826
rect 9280 17666 9360 17774
rect 9280 17614 9294 17666
rect 9346 17614 9360 17666
rect 9280 17506 9360 17614
rect 9280 17454 9294 17506
rect 9346 17454 9360 17506
rect 9280 17346 9360 17454
rect 9280 17294 9294 17346
rect 9346 17294 9360 17346
rect 9280 17186 9360 17294
rect 9280 17134 9294 17186
rect 9346 17134 9360 17186
rect 9280 17026 9360 17134
rect 9280 16974 9294 17026
rect 9346 16974 9360 17026
rect 9280 16866 9360 16974
rect 9280 16814 9294 16866
rect 9346 16814 9360 16866
rect 9280 16697 9360 16814
rect 9280 16663 9303 16697
rect 9337 16663 9360 16697
rect 9280 16546 9360 16663
rect 9280 16494 9294 16546
rect 9346 16494 9360 16546
rect 9280 16386 9360 16494
rect 9280 16334 9294 16386
rect 9346 16334 9360 16386
rect 9280 16226 9360 16334
rect 9280 16174 9294 16226
rect 9346 16174 9360 16226
rect 9280 16066 9360 16174
rect 9280 16014 9294 16066
rect 9346 16014 9360 16066
rect 9280 15906 9360 16014
rect 9280 15854 9294 15906
rect 9346 15854 9360 15906
rect 9280 15746 9360 15854
rect 9280 15694 9294 15746
rect 9346 15694 9360 15746
rect 9280 15586 9360 15694
rect 9280 15534 9294 15586
rect 9346 15534 9360 15586
rect 9280 15426 9360 15534
rect 9280 15374 9294 15426
rect 9346 15374 9360 15426
rect 9280 15266 9360 15374
rect 9280 15214 9294 15266
rect 9346 15214 9360 15266
rect 9280 15106 9360 15214
rect 9280 15054 9294 15106
rect 9346 15054 9360 15106
rect 9280 14946 9360 15054
rect 9280 14894 9294 14946
rect 9346 14894 9360 14946
rect 9280 14786 9360 14894
rect 9280 14734 9294 14786
rect 9346 14734 9360 14786
rect 9280 14626 9360 14734
rect 9280 14574 9294 14626
rect 9346 14574 9360 14626
rect 9280 14466 9360 14574
rect 9280 14414 9294 14466
rect 9346 14414 9360 14466
rect 9280 14306 9360 14414
rect 9280 14254 9294 14306
rect 9346 14254 9360 14306
rect 9280 14146 9360 14254
rect 9280 14094 9294 14146
rect 9346 14094 9360 14146
rect 9280 13986 9360 14094
rect 9280 13934 9294 13986
rect 9346 13934 9360 13986
rect 9280 13817 9360 13934
rect 9280 13783 9303 13817
rect 9337 13783 9360 13817
rect 9280 13666 9360 13783
rect 9280 13614 9294 13666
rect 9346 13614 9360 13666
rect 9280 13506 9360 13614
rect 9280 13454 9294 13506
rect 9346 13454 9360 13506
rect 9280 13346 9360 13454
rect 9280 13294 9294 13346
rect 9346 13294 9360 13346
rect 9280 13186 9360 13294
rect 9280 13134 9294 13186
rect 9346 13134 9360 13186
rect 9280 13026 9360 13134
rect 9280 12974 9294 13026
rect 9346 12974 9360 13026
rect 9280 12866 9360 12974
rect 9280 12814 9294 12866
rect 9346 12814 9360 12866
rect 9280 12706 9360 12814
rect 9280 12654 9294 12706
rect 9346 12654 9360 12706
rect 9280 12546 9360 12654
rect 9280 12494 9294 12546
rect 9346 12494 9360 12546
rect 9280 12377 9360 12494
rect 9280 12343 9303 12377
rect 9337 12343 9360 12377
rect 9280 12217 9360 12343
rect 9280 12183 9303 12217
rect 9337 12183 9360 12217
rect 9280 12057 9360 12183
rect 9280 12023 9303 12057
rect 9337 12023 9360 12057
rect 9280 11897 9360 12023
rect 9280 11863 9303 11897
rect 9337 11863 9360 11897
rect 9280 11746 9360 11863
rect 9280 11694 9294 11746
rect 9346 11694 9360 11746
rect 9280 11586 9360 11694
rect 9280 11534 9294 11586
rect 9346 11534 9360 11586
rect 9280 11426 9360 11534
rect 9280 11374 9294 11426
rect 9346 11374 9360 11426
rect 9280 11266 9360 11374
rect 9280 11214 9294 11266
rect 9346 11214 9360 11266
rect 9280 11106 9360 11214
rect 9280 11054 9294 11106
rect 9346 11054 9360 11106
rect 9280 10946 9360 11054
rect 9280 10894 9294 10946
rect 9346 10894 9360 10946
rect 9280 10786 9360 10894
rect 9280 10734 9294 10786
rect 9346 10734 9360 10786
rect 9280 10626 9360 10734
rect 9280 10574 9294 10626
rect 9346 10574 9360 10626
rect 9280 10466 9360 10574
rect 9280 10414 9294 10466
rect 9346 10414 9360 10466
rect 9280 10306 9360 10414
rect 9280 10254 9294 10306
rect 9346 10254 9360 10306
rect 9280 10146 9360 10254
rect 9280 10094 9294 10146
rect 9346 10094 9360 10146
rect 9280 9986 9360 10094
rect 9280 9934 9294 9986
rect 9346 9934 9360 9986
rect 9280 9826 9360 9934
rect 9280 9774 9294 9826
rect 9346 9774 9360 9826
rect 9280 9657 9360 9774
rect 9280 9623 9303 9657
rect 9337 9623 9360 9657
rect 9280 9506 9360 9623
rect 9280 9454 9294 9506
rect 9346 9454 9360 9506
rect 9280 9346 9360 9454
rect 9280 9294 9294 9346
rect 9346 9294 9360 9346
rect 9280 9177 9360 9294
rect 9280 9143 9303 9177
rect 9337 9143 9360 9177
rect 9280 9026 9360 9143
rect 9280 8974 9294 9026
rect 9346 8974 9360 9026
rect 9280 8866 9360 8974
rect 9280 8814 9294 8866
rect 9346 8814 9360 8866
rect 9280 8706 9360 8814
rect 9280 8654 9294 8706
rect 9346 8654 9360 8706
rect 9280 8546 9360 8654
rect 9280 8494 9294 8546
rect 9346 8494 9360 8546
rect 9280 8386 9360 8494
rect 9280 8334 9294 8386
rect 9346 8334 9360 8386
rect 9280 8226 9360 8334
rect 9280 8174 9294 8226
rect 9346 8174 9360 8226
rect 9280 8066 9360 8174
rect 9280 8014 9294 8066
rect 9346 8014 9360 8066
rect 9280 7906 9360 8014
rect 9280 7854 9294 7906
rect 9346 7854 9360 7906
rect 9280 7746 9360 7854
rect 9280 7694 9294 7746
rect 9346 7694 9360 7746
rect 9280 7577 9360 7694
rect 9280 7543 9303 7577
rect 9337 7543 9360 7577
rect 9280 7426 9360 7543
rect 9280 7374 9294 7426
rect 9346 7374 9360 7426
rect 9280 7266 9360 7374
rect 9280 7214 9294 7266
rect 9346 7214 9360 7266
rect 9280 7097 9360 7214
rect 9280 7063 9303 7097
rect 9337 7063 9360 7097
rect 9280 6946 9360 7063
rect 9280 6894 9294 6946
rect 9346 6894 9360 6946
rect 9280 6786 9360 6894
rect 9280 6734 9294 6786
rect 9346 6734 9360 6786
rect 9280 6617 9360 6734
rect 9280 6583 9303 6617
rect 9337 6583 9360 6617
rect 9280 6466 9360 6583
rect 9280 6414 9294 6466
rect 9346 6414 9360 6466
rect 9280 6306 9360 6414
rect 9280 6254 9294 6306
rect 9346 6254 9360 6306
rect 9280 6146 9360 6254
rect 9280 6094 9294 6146
rect 9346 6094 9360 6146
rect 9280 5986 9360 6094
rect 9280 5934 9294 5986
rect 9346 5934 9360 5986
rect 9280 5826 9360 5934
rect 9280 5774 9294 5826
rect 9346 5774 9360 5826
rect 9280 5666 9360 5774
rect 9280 5614 9294 5666
rect 9346 5614 9360 5666
rect 9280 5506 9360 5614
rect 9280 5454 9294 5506
rect 9346 5454 9360 5506
rect 9280 5346 9360 5454
rect 9280 5294 9294 5346
rect 9346 5294 9360 5346
rect 9280 5186 9360 5294
rect 9280 5134 9294 5186
rect 9346 5134 9360 5186
rect 9280 5026 9360 5134
rect 9280 4974 9294 5026
rect 9346 4974 9360 5026
rect 9280 4866 9360 4974
rect 9280 4814 9294 4866
rect 9346 4814 9360 4866
rect 9280 4706 9360 4814
rect 9280 4654 9294 4706
rect 9346 4654 9360 4706
rect 9280 4546 9360 4654
rect 9280 4494 9294 4546
rect 9346 4494 9360 4546
rect 9280 4386 9360 4494
rect 9280 4334 9294 4386
rect 9346 4334 9360 4386
rect 9280 4226 9360 4334
rect 9280 4174 9294 4226
rect 9346 4174 9360 4226
rect 9280 4066 9360 4174
rect 9280 4014 9294 4066
rect 9346 4014 9360 4066
rect 9280 3906 9360 4014
rect 9280 3854 9294 3906
rect 9346 3854 9360 3906
rect 9280 3737 9360 3854
rect 9280 3703 9303 3737
rect 9337 3703 9360 3737
rect 9280 3577 9360 3703
rect 9280 3543 9303 3577
rect 9337 3543 9360 3577
rect 9280 3426 9360 3543
rect 9280 3374 9294 3426
rect 9346 3374 9360 3426
rect 9280 3266 9360 3374
rect 9280 3214 9294 3266
rect 9346 3214 9360 3266
rect 9280 3106 9360 3214
rect 9280 3054 9294 3106
rect 9346 3054 9360 3106
rect 9280 2946 9360 3054
rect 9280 2894 9294 2946
rect 9346 2894 9360 2946
rect 9280 2786 9360 2894
rect 9280 2734 9294 2786
rect 9346 2734 9360 2786
rect 9280 2626 9360 2734
rect 9280 2574 9294 2626
rect 9346 2574 9360 2626
rect 9280 2466 9360 2574
rect 9280 2414 9294 2466
rect 9346 2414 9360 2466
rect 9280 2306 9360 2414
rect 9280 2254 9294 2306
rect 9346 2254 9360 2306
rect 9280 2146 9360 2254
rect 9280 2094 9294 2146
rect 9346 2094 9360 2146
rect 9280 1986 9360 2094
rect 9280 1934 9294 1986
rect 9346 1934 9360 1986
rect 9280 1817 9360 1934
rect 9280 1783 9303 1817
rect 9337 1783 9360 1817
rect 9280 1666 9360 1783
rect 9280 1614 9294 1666
rect 9346 1614 9360 1666
rect 9280 1506 9360 1614
rect 9280 1454 9294 1506
rect 9346 1454 9360 1506
rect 9280 1346 9360 1454
rect 9280 1294 9294 1346
rect 9346 1294 9360 1346
rect 9280 1186 9360 1294
rect 9280 1134 9294 1186
rect 9346 1134 9360 1186
rect 9280 1026 9360 1134
rect 9280 974 9294 1026
rect 9346 974 9360 1026
rect 9280 857 9360 974
rect 9280 823 9303 857
rect 9337 823 9360 857
rect 9280 697 9360 823
rect 9280 663 9303 697
rect 9337 663 9360 697
rect 9280 546 9360 663
rect 9280 494 9294 546
rect 9346 494 9360 546
rect 9280 386 9360 494
rect 9280 334 9294 386
rect 9346 334 9360 386
rect 9280 226 9360 334
rect 9280 174 9294 226
rect 9346 174 9360 226
rect 9280 66 9360 174
rect 9280 14 9294 66
rect 9346 14 9360 66
rect 9280 0 9360 14
rect 9440 31426 9520 31440
rect 9440 31374 9454 31426
rect 9506 31374 9520 31426
rect 9440 31266 9520 31374
rect 9440 31214 9454 31266
rect 9506 31214 9520 31266
rect 9440 31106 9520 31214
rect 9440 31054 9454 31106
rect 9506 31054 9520 31106
rect 9440 30946 9520 31054
rect 9440 30894 9454 30946
rect 9506 30894 9520 30946
rect 9440 30786 9520 30894
rect 9440 30734 9454 30786
rect 9506 30734 9520 30786
rect 9440 30626 9520 30734
rect 9440 30574 9454 30626
rect 9506 30574 9520 30626
rect 9440 30466 9520 30574
rect 9440 30414 9454 30466
rect 9506 30414 9520 30466
rect 9440 30306 9520 30414
rect 9440 30254 9454 30306
rect 9506 30254 9520 30306
rect 9440 30137 9520 30254
rect 9440 30103 9463 30137
rect 9497 30103 9520 30137
rect 9440 29986 9520 30103
rect 9440 29934 9454 29986
rect 9506 29934 9520 29986
rect 9440 29826 9520 29934
rect 9440 29774 9454 29826
rect 9506 29774 9520 29826
rect 9440 29666 9520 29774
rect 9440 29614 9454 29666
rect 9506 29614 9520 29666
rect 9440 29506 9520 29614
rect 9440 29454 9454 29506
rect 9506 29454 9520 29506
rect 9440 29346 9520 29454
rect 9440 29294 9454 29346
rect 9506 29294 9520 29346
rect 9440 29186 9520 29294
rect 9440 29134 9454 29186
rect 9506 29134 9520 29186
rect 9440 29026 9520 29134
rect 9440 28974 9454 29026
rect 9506 28974 9520 29026
rect 9440 28866 9520 28974
rect 9440 28814 9454 28866
rect 9506 28814 9520 28866
rect 9440 28697 9520 28814
rect 9440 28663 9463 28697
rect 9497 28663 9520 28697
rect 9440 28537 9520 28663
rect 9440 28503 9463 28537
rect 9497 28503 9520 28537
rect 9440 28377 9520 28503
rect 9440 28343 9463 28377
rect 9497 28343 9520 28377
rect 9440 28217 9520 28343
rect 9440 28183 9463 28217
rect 9497 28183 9520 28217
rect 9440 28066 9520 28183
rect 9440 28014 9454 28066
rect 9506 28014 9520 28066
rect 9440 27906 9520 28014
rect 9440 27854 9454 27906
rect 9506 27854 9520 27906
rect 9440 27746 9520 27854
rect 9440 27694 9454 27746
rect 9506 27694 9520 27746
rect 9440 27586 9520 27694
rect 9440 27534 9454 27586
rect 9506 27534 9520 27586
rect 9440 27426 9520 27534
rect 9440 27374 9454 27426
rect 9506 27374 9520 27426
rect 9440 27266 9520 27374
rect 9440 27214 9454 27266
rect 9506 27214 9520 27266
rect 9440 27106 9520 27214
rect 9440 27054 9454 27106
rect 9506 27054 9520 27106
rect 9440 26946 9520 27054
rect 9440 26894 9454 26946
rect 9506 26894 9520 26946
rect 9440 26777 9520 26894
rect 9440 26743 9463 26777
rect 9497 26743 9520 26777
rect 9440 26617 9520 26743
rect 9440 26583 9463 26617
rect 9497 26583 9520 26617
rect 9440 26457 9520 26583
rect 9440 26423 9463 26457
rect 9497 26423 9520 26457
rect 9440 26297 9520 26423
rect 9440 26263 9463 26297
rect 9497 26263 9520 26297
rect 9440 26146 9520 26263
rect 9440 26094 9454 26146
rect 9506 26094 9520 26146
rect 9440 25986 9520 26094
rect 9440 25934 9454 25986
rect 9506 25934 9520 25986
rect 9440 25826 9520 25934
rect 9440 25774 9454 25826
rect 9506 25774 9520 25826
rect 9440 25666 9520 25774
rect 9440 25614 9454 25666
rect 9506 25614 9520 25666
rect 9440 25506 9520 25614
rect 9440 25454 9454 25506
rect 9506 25454 9520 25506
rect 9440 25346 9520 25454
rect 9440 25294 9454 25346
rect 9506 25294 9520 25346
rect 9440 25186 9520 25294
rect 9440 25134 9454 25186
rect 9506 25134 9520 25186
rect 9440 25026 9520 25134
rect 9440 24974 9454 25026
rect 9506 24974 9520 25026
rect 9440 24857 9520 24974
rect 9440 24823 9463 24857
rect 9497 24823 9520 24857
rect 9440 24706 9520 24823
rect 9440 24654 9454 24706
rect 9506 24654 9520 24706
rect 9440 24546 9520 24654
rect 9440 24494 9454 24546
rect 9506 24494 9520 24546
rect 9440 24386 9520 24494
rect 9440 24334 9454 24386
rect 9506 24334 9520 24386
rect 9440 24226 9520 24334
rect 9440 24174 9454 24226
rect 9506 24174 9520 24226
rect 9440 24066 9520 24174
rect 9440 24014 9454 24066
rect 9506 24014 9520 24066
rect 9440 23906 9520 24014
rect 9440 23854 9454 23906
rect 9506 23854 9520 23906
rect 9440 23746 9520 23854
rect 9440 23694 9454 23746
rect 9506 23694 9520 23746
rect 9440 23586 9520 23694
rect 9440 23534 9454 23586
rect 9506 23534 9520 23586
rect 9440 23426 9520 23534
rect 9440 23374 9454 23426
rect 9506 23374 9520 23426
rect 9440 23266 9520 23374
rect 9440 23214 9454 23266
rect 9506 23214 9520 23266
rect 9440 23106 9520 23214
rect 9440 23054 9454 23106
rect 9506 23054 9520 23106
rect 9440 22946 9520 23054
rect 9440 22894 9454 22946
rect 9506 22894 9520 22946
rect 9440 22786 9520 22894
rect 9440 22734 9454 22786
rect 9506 22734 9520 22786
rect 9440 22626 9520 22734
rect 9440 22574 9454 22626
rect 9506 22574 9520 22626
rect 9440 22466 9520 22574
rect 9440 22414 9454 22466
rect 9506 22414 9520 22466
rect 9440 22306 9520 22414
rect 9440 22254 9454 22306
rect 9506 22254 9520 22306
rect 9440 22146 9520 22254
rect 9440 22094 9454 22146
rect 9506 22094 9520 22146
rect 9440 21977 9520 22094
rect 9440 21943 9463 21977
rect 9497 21943 9520 21977
rect 9440 21826 9520 21943
rect 9440 21774 9454 21826
rect 9506 21774 9520 21826
rect 9440 21666 9520 21774
rect 9440 21614 9454 21666
rect 9506 21614 9520 21666
rect 9440 21506 9520 21614
rect 9440 21454 9454 21506
rect 9506 21454 9520 21506
rect 9440 21346 9520 21454
rect 9440 21294 9454 21346
rect 9506 21294 9520 21346
rect 9440 21186 9520 21294
rect 9440 21134 9454 21186
rect 9506 21134 9520 21186
rect 9440 21026 9520 21134
rect 9440 20974 9454 21026
rect 9506 20974 9520 21026
rect 9440 20866 9520 20974
rect 9440 20814 9454 20866
rect 9506 20814 9520 20866
rect 9440 20706 9520 20814
rect 9440 20654 9454 20706
rect 9506 20654 9520 20706
rect 9440 20537 9520 20654
rect 9440 20503 9463 20537
rect 9497 20503 9520 20537
rect 9440 20377 9520 20503
rect 9440 20343 9463 20377
rect 9497 20343 9520 20377
rect 9440 20217 9520 20343
rect 9440 20183 9463 20217
rect 9497 20183 9520 20217
rect 9440 20057 9520 20183
rect 9440 20023 9463 20057
rect 9497 20023 9520 20057
rect 9440 19906 9520 20023
rect 9440 19854 9454 19906
rect 9506 19854 9520 19906
rect 9440 19746 9520 19854
rect 9440 19694 9454 19746
rect 9506 19694 9520 19746
rect 9440 19586 9520 19694
rect 9440 19534 9454 19586
rect 9506 19534 9520 19586
rect 9440 19426 9520 19534
rect 9440 19374 9454 19426
rect 9506 19374 9520 19426
rect 9440 19266 9520 19374
rect 9440 19214 9454 19266
rect 9506 19214 9520 19266
rect 9440 19106 9520 19214
rect 9440 19054 9454 19106
rect 9506 19054 9520 19106
rect 9440 18946 9520 19054
rect 9440 18894 9454 18946
rect 9506 18894 9520 18946
rect 9440 18786 9520 18894
rect 9440 18734 9454 18786
rect 9506 18734 9520 18786
rect 9440 18617 9520 18734
rect 9440 18583 9463 18617
rect 9497 18583 9520 18617
rect 9440 18457 9520 18583
rect 9440 18423 9463 18457
rect 9497 18423 9520 18457
rect 9440 18297 9520 18423
rect 9440 18263 9463 18297
rect 9497 18263 9520 18297
rect 9440 18137 9520 18263
rect 9440 18103 9463 18137
rect 9497 18103 9520 18137
rect 9440 17986 9520 18103
rect 9440 17934 9454 17986
rect 9506 17934 9520 17986
rect 9440 17826 9520 17934
rect 9440 17774 9454 17826
rect 9506 17774 9520 17826
rect 9440 17666 9520 17774
rect 9440 17614 9454 17666
rect 9506 17614 9520 17666
rect 9440 17506 9520 17614
rect 9440 17454 9454 17506
rect 9506 17454 9520 17506
rect 9440 17346 9520 17454
rect 9440 17294 9454 17346
rect 9506 17294 9520 17346
rect 9440 17186 9520 17294
rect 9440 17134 9454 17186
rect 9506 17134 9520 17186
rect 9440 17026 9520 17134
rect 9440 16974 9454 17026
rect 9506 16974 9520 17026
rect 9440 16866 9520 16974
rect 9440 16814 9454 16866
rect 9506 16814 9520 16866
rect 9440 16697 9520 16814
rect 9440 16663 9463 16697
rect 9497 16663 9520 16697
rect 9440 16546 9520 16663
rect 9440 16494 9454 16546
rect 9506 16494 9520 16546
rect 9440 16386 9520 16494
rect 9440 16334 9454 16386
rect 9506 16334 9520 16386
rect 9440 16226 9520 16334
rect 9440 16174 9454 16226
rect 9506 16174 9520 16226
rect 9440 16066 9520 16174
rect 9440 16014 9454 16066
rect 9506 16014 9520 16066
rect 9440 15906 9520 16014
rect 9440 15854 9454 15906
rect 9506 15854 9520 15906
rect 9440 15746 9520 15854
rect 9440 15694 9454 15746
rect 9506 15694 9520 15746
rect 9440 15586 9520 15694
rect 9440 15534 9454 15586
rect 9506 15534 9520 15586
rect 9440 15426 9520 15534
rect 9440 15374 9454 15426
rect 9506 15374 9520 15426
rect 9440 15266 9520 15374
rect 9440 15214 9454 15266
rect 9506 15214 9520 15266
rect 9440 15106 9520 15214
rect 9440 15054 9454 15106
rect 9506 15054 9520 15106
rect 9440 14946 9520 15054
rect 9440 14894 9454 14946
rect 9506 14894 9520 14946
rect 9440 14786 9520 14894
rect 9440 14734 9454 14786
rect 9506 14734 9520 14786
rect 9440 14626 9520 14734
rect 9440 14574 9454 14626
rect 9506 14574 9520 14626
rect 9440 14466 9520 14574
rect 9440 14414 9454 14466
rect 9506 14414 9520 14466
rect 9440 14306 9520 14414
rect 9440 14254 9454 14306
rect 9506 14254 9520 14306
rect 9440 14146 9520 14254
rect 9440 14094 9454 14146
rect 9506 14094 9520 14146
rect 9440 13986 9520 14094
rect 9440 13934 9454 13986
rect 9506 13934 9520 13986
rect 9440 13817 9520 13934
rect 9440 13783 9463 13817
rect 9497 13783 9520 13817
rect 9440 13666 9520 13783
rect 9440 13614 9454 13666
rect 9506 13614 9520 13666
rect 9440 13506 9520 13614
rect 9440 13454 9454 13506
rect 9506 13454 9520 13506
rect 9440 13346 9520 13454
rect 9440 13294 9454 13346
rect 9506 13294 9520 13346
rect 9440 13186 9520 13294
rect 9440 13134 9454 13186
rect 9506 13134 9520 13186
rect 9440 13026 9520 13134
rect 9440 12974 9454 13026
rect 9506 12974 9520 13026
rect 9440 12866 9520 12974
rect 9440 12814 9454 12866
rect 9506 12814 9520 12866
rect 9440 12706 9520 12814
rect 9440 12654 9454 12706
rect 9506 12654 9520 12706
rect 9440 12546 9520 12654
rect 9440 12494 9454 12546
rect 9506 12494 9520 12546
rect 9440 12377 9520 12494
rect 9440 12343 9463 12377
rect 9497 12343 9520 12377
rect 9440 12217 9520 12343
rect 9440 12183 9463 12217
rect 9497 12183 9520 12217
rect 9440 12057 9520 12183
rect 9440 12023 9463 12057
rect 9497 12023 9520 12057
rect 9440 11897 9520 12023
rect 9440 11863 9463 11897
rect 9497 11863 9520 11897
rect 9440 11746 9520 11863
rect 9440 11694 9454 11746
rect 9506 11694 9520 11746
rect 9440 11586 9520 11694
rect 9440 11534 9454 11586
rect 9506 11534 9520 11586
rect 9440 11426 9520 11534
rect 9440 11374 9454 11426
rect 9506 11374 9520 11426
rect 9440 11266 9520 11374
rect 9440 11214 9454 11266
rect 9506 11214 9520 11266
rect 9440 11106 9520 11214
rect 9440 11054 9454 11106
rect 9506 11054 9520 11106
rect 9440 10946 9520 11054
rect 9440 10894 9454 10946
rect 9506 10894 9520 10946
rect 9440 10786 9520 10894
rect 9440 10734 9454 10786
rect 9506 10734 9520 10786
rect 9440 10626 9520 10734
rect 9440 10574 9454 10626
rect 9506 10574 9520 10626
rect 9440 10466 9520 10574
rect 9440 10414 9454 10466
rect 9506 10414 9520 10466
rect 9440 10306 9520 10414
rect 9440 10254 9454 10306
rect 9506 10254 9520 10306
rect 9440 10146 9520 10254
rect 9440 10094 9454 10146
rect 9506 10094 9520 10146
rect 9440 9986 9520 10094
rect 9440 9934 9454 9986
rect 9506 9934 9520 9986
rect 9440 9826 9520 9934
rect 9440 9774 9454 9826
rect 9506 9774 9520 9826
rect 9440 9657 9520 9774
rect 9440 9623 9463 9657
rect 9497 9623 9520 9657
rect 9440 9506 9520 9623
rect 9440 9454 9454 9506
rect 9506 9454 9520 9506
rect 9440 9346 9520 9454
rect 9440 9294 9454 9346
rect 9506 9294 9520 9346
rect 9440 9177 9520 9294
rect 9440 9143 9463 9177
rect 9497 9143 9520 9177
rect 9440 9026 9520 9143
rect 9440 8974 9454 9026
rect 9506 8974 9520 9026
rect 9440 8866 9520 8974
rect 9440 8814 9454 8866
rect 9506 8814 9520 8866
rect 9440 8706 9520 8814
rect 9440 8654 9454 8706
rect 9506 8654 9520 8706
rect 9440 8546 9520 8654
rect 9440 8494 9454 8546
rect 9506 8494 9520 8546
rect 9440 8386 9520 8494
rect 9440 8334 9454 8386
rect 9506 8334 9520 8386
rect 9440 8226 9520 8334
rect 9440 8174 9454 8226
rect 9506 8174 9520 8226
rect 9440 8066 9520 8174
rect 9440 8014 9454 8066
rect 9506 8014 9520 8066
rect 9440 7906 9520 8014
rect 9440 7854 9454 7906
rect 9506 7854 9520 7906
rect 9440 7746 9520 7854
rect 9440 7694 9454 7746
rect 9506 7694 9520 7746
rect 9440 7577 9520 7694
rect 9440 7543 9463 7577
rect 9497 7543 9520 7577
rect 9440 7426 9520 7543
rect 9440 7374 9454 7426
rect 9506 7374 9520 7426
rect 9440 7266 9520 7374
rect 9440 7214 9454 7266
rect 9506 7214 9520 7266
rect 9440 7097 9520 7214
rect 9440 7063 9463 7097
rect 9497 7063 9520 7097
rect 9440 6946 9520 7063
rect 9440 6894 9454 6946
rect 9506 6894 9520 6946
rect 9440 6786 9520 6894
rect 9440 6734 9454 6786
rect 9506 6734 9520 6786
rect 9440 6617 9520 6734
rect 9440 6583 9463 6617
rect 9497 6583 9520 6617
rect 9440 6466 9520 6583
rect 9440 6414 9454 6466
rect 9506 6414 9520 6466
rect 9440 6306 9520 6414
rect 9440 6254 9454 6306
rect 9506 6254 9520 6306
rect 9440 6146 9520 6254
rect 9440 6094 9454 6146
rect 9506 6094 9520 6146
rect 9440 5986 9520 6094
rect 9440 5934 9454 5986
rect 9506 5934 9520 5986
rect 9440 5826 9520 5934
rect 9440 5774 9454 5826
rect 9506 5774 9520 5826
rect 9440 5666 9520 5774
rect 9440 5614 9454 5666
rect 9506 5614 9520 5666
rect 9440 5506 9520 5614
rect 9440 5454 9454 5506
rect 9506 5454 9520 5506
rect 9440 5346 9520 5454
rect 9440 5294 9454 5346
rect 9506 5294 9520 5346
rect 9440 5186 9520 5294
rect 9440 5134 9454 5186
rect 9506 5134 9520 5186
rect 9440 5026 9520 5134
rect 9440 4974 9454 5026
rect 9506 4974 9520 5026
rect 9440 4866 9520 4974
rect 9440 4814 9454 4866
rect 9506 4814 9520 4866
rect 9440 4706 9520 4814
rect 9440 4654 9454 4706
rect 9506 4654 9520 4706
rect 9440 4546 9520 4654
rect 9440 4494 9454 4546
rect 9506 4494 9520 4546
rect 9440 4386 9520 4494
rect 9440 4334 9454 4386
rect 9506 4334 9520 4386
rect 9440 4226 9520 4334
rect 9440 4174 9454 4226
rect 9506 4174 9520 4226
rect 9440 4066 9520 4174
rect 9440 4014 9454 4066
rect 9506 4014 9520 4066
rect 9440 3906 9520 4014
rect 9440 3854 9454 3906
rect 9506 3854 9520 3906
rect 9440 3737 9520 3854
rect 9440 3703 9463 3737
rect 9497 3703 9520 3737
rect 9440 3577 9520 3703
rect 9440 3543 9463 3577
rect 9497 3543 9520 3577
rect 9440 3426 9520 3543
rect 9440 3374 9454 3426
rect 9506 3374 9520 3426
rect 9440 3266 9520 3374
rect 9440 3214 9454 3266
rect 9506 3214 9520 3266
rect 9440 3106 9520 3214
rect 9440 3054 9454 3106
rect 9506 3054 9520 3106
rect 9440 2946 9520 3054
rect 9440 2894 9454 2946
rect 9506 2894 9520 2946
rect 9440 2786 9520 2894
rect 9440 2734 9454 2786
rect 9506 2734 9520 2786
rect 9440 2626 9520 2734
rect 9440 2574 9454 2626
rect 9506 2574 9520 2626
rect 9440 2466 9520 2574
rect 9440 2414 9454 2466
rect 9506 2414 9520 2466
rect 9440 2306 9520 2414
rect 9440 2254 9454 2306
rect 9506 2254 9520 2306
rect 9440 2146 9520 2254
rect 9440 2094 9454 2146
rect 9506 2094 9520 2146
rect 9440 1986 9520 2094
rect 9440 1934 9454 1986
rect 9506 1934 9520 1986
rect 9440 1817 9520 1934
rect 9440 1783 9463 1817
rect 9497 1783 9520 1817
rect 9440 1666 9520 1783
rect 9440 1614 9454 1666
rect 9506 1614 9520 1666
rect 9440 1506 9520 1614
rect 9440 1454 9454 1506
rect 9506 1454 9520 1506
rect 9440 1346 9520 1454
rect 9440 1294 9454 1346
rect 9506 1294 9520 1346
rect 9440 1186 9520 1294
rect 9440 1134 9454 1186
rect 9506 1134 9520 1186
rect 9440 1026 9520 1134
rect 9440 974 9454 1026
rect 9506 974 9520 1026
rect 9440 857 9520 974
rect 9440 823 9463 857
rect 9497 823 9520 857
rect 9440 697 9520 823
rect 9440 663 9463 697
rect 9497 663 9520 697
rect 9440 546 9520 663
rect 9440 494 9454 546
rect 9506 494 9520 546
rect 9440 386 9520 494
rect 9440 334 9454 386
rect 9506 334 9520 386
rect 9440 226 9520 334
rect 9440 174 9454 226
rect 9506 174 9520 226
rect 9440 66 9520 174
rect 9440 14 9454 66
rect 9506 14 9520 66
rect 9440 0 9520 14
rect 9600 31417 9680 31440
rect 9600 31383 9623 31417
rect 9657 31383 9680 31417
rect 9600 31257 9680 31383
rect 9600 31223 9623 31257
rect 9657 31223 9680 31257
rect 9600 31097 9680 31223
rect 9600 31063 9623 31097
rect 9657 31063 9680 31097
rect 9600 30937 9680 31063
rect 9600 30903 9623 30937
rect 9657 30903 9680 30937
rect 9600 30777 9680 30903
rect 9600 30743 9623 30777
rect 9657 30743 9680 30777
rect 9600 30617 9680 30743
rect 9600 30583 9623 30617
rect 9657 30583 9680 30617
rect 9600 30457 9680 30583
rect 9600 30423 9623 30457
rect 9657 30423 9680 30457
rect 9600 30297 9680 30423
rect 9600 30263 9623 30297
rect 9657 30263 9680 30297
rect 9600 30137 9680 30263
rect 9600 30103 9623 30137
rect 9657 30103 9680 30137
rect 9600 29977 9680 30103
rect 9600 29943 9623 29977
rect 9657 29943 9680 29977
rect 9600 29817 9680 29943
rect 9600 29783 9623 29817
rect 9657 29783 9680 29817
rect 9600 29657 9680 29783
rect 9600 29623 9623 29657
rect 9657 29623 9680 29657
rect 9600 29497 9680 29623
rect 9600 29463 9623 29497
rect 9657 29463 9680 29497
rect 9600 29337 9680 29463
rect 9600 29303 9623 29337
rect 9657 29303 9680 29337
rect 9600 29177 9680 29303
rect 9600 29143 9623 29177
rect 9657 29143 9680 29177
rect 9600 29017 9680 29143
rect 9600 28983 9623 29017
rect 9657 28983 9680 29017
rect 9600 28857 9680 28983
rect 9600 28823 9623 28857
rect 9657 28823 9680 28857
rect 9600 28697 9680 28823
rect 9600 28663 9623 28697
rect 9657 28663 9680 28697
rect 9600 28537 9680 28663
rect 9600 28503 9623 28537
rect 9657 28503 9680 28537
rect 9600 28377 9680 28503
rect 9600 28343 9623 28377
rect 9657 28343 9680 28377
rect 9600 28217 9680 28343
rect 9600 28183 9623 28217
rect 9657 28183 9680 28217
rect 9600 28057 9680 28183
rect 9600 28023 9623 28057
rect 9657 28023 9680 28057
rect 9600 27897 9680 28023
rect 9600 27863 9623 27897
rect 9657 27863 9680 27897
rect 9600 27737 9680 27863
rect 9600 27703 9623 27737
rect 9657 27703 9680 27737
rect 9600 27577 9680 27703
rect 9600 27543 9623 27577
rect 9657 27543 9680 27577
rect 9600 27417 9680 27543
rect 9600 27383 9623 27417
rect 9657 27383 9680 27417
rect 9600 27257 9680 27383
rect 9600 27223 9623 27257
rect 9657 27223 9680 27257
rect 9600 27097 9680 27223
rect 9600 27063 9623 27097
rect 9657 27063 9680 27097
rect 9600 26937 9680 27063
rect 9600 26903 9623 26937
rect 9657 26903 9680 26937
rect 9600 26777 9680 26903
rect 9600 26743 9623 26777
rect 9657 26743 9680 26777
rect 9600 26617 9680 26743
rect 9600 26583 9623 26617
rect 9657 26583 9680 26617
rect 9600 26457 9680 26583
rect 9600 26423 9623 26457
rect 9657 26423 9680 26457
rect 9600 26297 9680 26423
rect 9600 26263 9623 26297
rect 9657 26263 9680 26297
rect 9600 26137 9680 26263
rect 9600 26103 9623 26137
rect 9657 26103 9680 26137
rect 9600 25977 9680 26103
rect 9600 25943 9623 25977
rect 9657 25943 9680 25977
rect 9600 25817 9680 25943
rect 9600 25783 9623 25817
rect 9657 25783 9680 25817
rect 9600 25657 9680 25783
rect 9600 25623 9623 25657
rect 9657 25623 9680 25657
rect 9600 25497 9680 25623
rect 9600 25463 9623 25497
rect 9657 25463 9680 25497
rect 9600 25337 9680 25463
rect 9600 25303 9623 25337
rect 9657 25303 9680 25337
rect 9600 25177 9680 25303
rect 9600 25143 9623 25177
rect 9657 25143 9680 25177
rect 9600 25017 9680 25143
rect 9600 24983 9623 25017
rect 9657 24983 9680 25017
rect 9600 24857 9680 24983
rect 9600 24823 9623 24857
rect 9657 24823 9680 24857
rect 9600 24697 9680 24823
rect 9600 24663 9623 24697
rect 9657 24663 9680 24697
rect 9600 24537 9680 24663
rect 9600 24503 9623 24537
rect 9657 24503 9680 24537
rect 9600 24377 9680 24503
rect 9600 24343 9623 24377
rect 9657 24343 9680 24377
rect 9600 24217 9680 24343
rect 9600 24183 9623 24217
rect 9657 24183 9680 24217
rect 9600 24057 9680 24183
rect 9600 24023 9623 24057
rect 9657 24023 9680 24057
rect 9600 23897 9680 24023
rect 9600 23863 9623 23897
rect 9657 23863 9680 23897
rect 9600 23737 9680 23863
rect 9600 23703 9623 23737
rect 9657 23703 9680 23737
rect 9600 23577 9680 23703
rect 9600 23543 9623 23577
rect 9657 23543 9680 23577
rect 9600 23417 9680 23543
rect 9600 23383 9623 23417
rect 9657 23383 9680 23417
rect 9600 23257 9680 23383
rect 9600 23223 9623 23257
rect 9657 23223 9680 23257
rect 9600 23097 9680 23223
rect 9600 23063 9623 23097
rect 9657 23063 9680 23097
rect 9600 22937 9680 23063
rect 9600 22903 9623 22937
rect 9657 22903 9680 22937
rect 9600 22777 9680 22903
rect 9600 22743 9623 22777
rect 9657 22743 9680 22777
rect 9600 22617 9680 22743
rect 9600 22583 9623 22617
rect 9657 22583 9680 22617
rect 9600 22457 9680 22583
rect 9600 22423 9623 22457
rect 9657 22423 9680 22457
rect 9600 22297 9680 22423
rect 9600 22263 9623 22297
rect 9657 22263 9680 22297
rect 9600 22137 9680 22263
rect 9600 22103 9623 22137
rect 9657 22103 9680 22137
rect 9600 21977 9680 22103
rect 9600 21943 9623 21977
rect 9657 21943 9680 21977
rect 9600 21817 9680 21943
rect 9600 21783 9623 21817
rect 9657 21783 9680 21817
rect 9600 21657 9680 21783
rect 9600 21623 9623 21657
rect 9657 21623 9680 21657
rect 9600 21497 9680 21623
rect 9600 21463 9623 21497
rect 9657 21463 9680 21497
rect 9600 21337 9680 21463
rect 9600 21303 9623 21337
rect 9657 21303 9680 21337
rect 9600 21177 9680 21303
rect 9600 21143 9623 21177
rect 9657 21143 9680 21177
rect 9600 21017 9680 21143
rect 9600 20983 9623 21017
rect 9657 20983 9680 21017
rect 9600 20857 9680 20983
rect 9600 20823 9623 20857
rect 9657 20823 9680 20857
rect 9600 20697 9680 20823
rect 9600 20663 9623 20697
rect 9657 20663 9680 20697
rect 9600 20537 9680 20663
rect 9600 20503 9623 20537
rect 9657 20503 9680 20537
rect 9600 20377 9680 20503
rect 9600 20343 9623 20377
rect 9657 20343 9680 20377
rect 9600 20217 9680 20343
rect 9600 20183 9623 20217
rect 9657 20183 9680 20217
rect 9600 20057 9680 20183
rect 9600 20023 9623 20057
rect 9657 20023 9680 20057
rect 9600 19897 9680 20023
rect 9600 19863 9623 19897
rect 9657 19863 9680 19897
rect 9600 19737 9680 19863
rect 9600 19703 9623 19737
rect 9657 19703 9680 19737
rect 9600 19577 9680 19703
rect 9600 19543 9623 19577
rect 9657 19543 9680 19577
rect 9600 19417 9680 19543
rect 9600 19383 9623 19417
rect 9657 19383 9680 19417
rect 9600 19257 9680 19383
rect 9600 19223 9623 19257
rect 9657 19223 9680 19257
rect 9600 19097 9680 19223
rect 9600 19063 9623 19097
rect 9657 19063 9680 19097
rect 9600 18937 9680 19063
rect 9600 18903 9623 18937
rect 9657 18903 9680 18937
rect 9600 18777 9680 18903
rect 9600 18743 9623 18777
rect 9657 18743 9680 18777
rect 9600 18617 9680 18743
rect 9600 18583 9623 18617
rect 9657 18583 9680 18617
rect 9600 18457 9680 18583
rect 9600 18423 9623 18457
rect 9657 18423 9680 18457
rect 9600 18297 9680 18423
rect 9600 18263 9623 18297
rect 9657 18263 9680 18297
rect 9600 18137 9680 18263
rect 9600 18103 9623 18137
rect 9657 18103 9680 18137
rect 9600 17977 9680 18103
rect 9600 17943 9623 17977
rect 9657 17943 9680 17977
rect 9600 17817 9680 17943
rect 9600 17783 9623 17817
rect 9657 17783 9680 17817
rect 9600 17657 9680 17783
rect 9600 17623 9623 17657
rect 9657 17623 9680 17657
rect 9600 17497 9680 17623
rect 9600 17463 9623 17497
rect 9657 17463 9680 17497
rect 9600 17337 9680 17463
rect 9600 17303 9623 17337
rect 9657 17303 9680 17337
rect 9600 17177 9680 17303
rect 9600 17143 9623 17177
rect 9657 17143 9680 17177
rect 9600 17017 9680 17143
rect 9600 16983 9623 17017
rect 9657 16983 9680 17017
rect 9600 16857 9680 16983
rect 9600 16823 9623 16857
rect 9657 16823 9680 16857
rect 9600 16697 9680 16823
rect 9600 16663 9623 16697
rect 9657 16663 9680 16697
rect 9600 16537 9680 16663
rect 9600 16503 9623 16537
rect 9657 16503 9680 16537
rect 9600 16377 9680 16503
rect 9600 16343 9623 16377
rect 9657 16343 9680 16377
rect 9600 16217 9680 16343
rect 9600 16183 9623 16217
rect 9657 16183 9680 16217
rect 9600 16057 9680 16183
rect 9600 16023 9623 16057
rect 9657 16023 9680 16057
rect 9600 15897 9680 16023
rect 9600 15863 9623 15897
rect 9657 15863 9680 15897
rect 9600 15737 9680 15863
rect 9600 15703 9623 15737
rect 9657 15703 9680 15737
rect 9600 15577 9680 15703
rect 9600 15543 9623 15577
rect 9657 15543 9680 15577
rect 9600 15417 9680 15543
rect 9600 15383 9623 15417
rect 9657 15383 9680 15417
rect 9600 15257 9680 15383
rect 9600 15223 9623 15257
rect 9657 15223 9680 15257
rect 9600 15097 9680 15223
rect 9600 15063 9623 15097
rect 9657 15063 9680 15097
rect 9600 14937 9680 15063
rect 9600 14903 9623 14937
rect 9657 14903 9680 14937
rect 9600 14777 9680 14903
rect 9600 14743 9623 14777
rect 9657 14743 9680 14777
rect 9600 14617 9680 14743
rect 9600 14583 9623 14617
rect 9657 14583 9680 14617
rect 9600 14457 9680 14583
rect 9600 14423 9623 14457
rect 9657 14423 9680 14457
rect 9600 14297 9680 14423
rect 9600 14263 9623 14297
rect 9657 14263 9680 14297
rect 9600 14137 9680 14263
rect 9600 14103 9623 14137
rect 9657 14103 9680 14137
rect 9600 13977 9680 14103
rect 9600 13943 9623 13977
rect 9657 13943 9680 13977
rect 9600 13817 9680 13943
rect 9600 13783 9623 13817
rect 9657 13783 9680 13817
rect 9600 13657 9680 13783
rect 9600 13623 9623 13657
rect 9657 13623 9680 13657
rect 9600 13497 9680 13623
rect 9600 13463 9623 13497
rect 9657 13463 9680 13497
rect 9600 13337 9680 13463
rect 9600 13303 9623 13337
rect 9657 13303 9680 13337
rect 9600 13177 9680 13303
rect 9600 13143 9623 13177
rect 9657 13143 9680 13177
rect 9600 13017 9680 13143
rect 9600 12983 9623 13017
rect 9657 12983 9680 13017
rect 9600 12857 9680 12983
rect 9600 12823 9623 12857
rect 9657 12823 9680 12857
rect 9600 12697 9680 12823
rect 9600 12663 9623 12697
rect 9657 12663 9680 12697
rect 9600 12537 9680 12663
rect 9600 12503 9623 12537
rect 9657 12503 9680 12537
rect 9600 12377 9680 12503
rect 9600 12343 9623 12377
rect 9657 12343 9680 12377
rect 9600 12217 9680 12343
rect 9600 12183 9623 12217
rect 9657 12183 9680 12217
rect 9600 12057 9680 12183
rect 9600 12023 9623 12057
rect 9657 12023 9680 12057
rect 9600 11897 9680 12023
rect 9600 11863 9623 11897
rect 9657 11863 9680 11897
rect 9600 11737 9680 11863
rect 9600 11703 9623 11737
rect 9657 11703 9680 11737
rect 9600 11577 9680 11703
rect 9600 11543 9623 11577
rect 9657 11543 9680 11577
rect 9600 11417 9680 11543
rect 9600 11383 9623 11417
rect 9657 11383 9680 11417
rect 9600 11257 9680 11383
rect 9600 11223 9623 11257
rect 9657 11223 9680 11257
rect 9600 11097 9680 11223
rect 9600 11063 9623 11097
rect 9657 11063 9680 11097
rect 9600 10937 9680 11063
rect 9600 10903 9623 10937
rect 9657 10903 9680 10937
rect 9600 10777 9680 10903
rect 9600 10743 9623 10777
rect 9657 10743 9680 10777
rect 9600 10617 9680 10743
rect 9600 10583 9623 10617
rect 9657 10583 9680 10617
rect 9600 10457 9680 10583
rect 9600 10423 9623 10457
rect 9657 10423 9680 10457
rect 9600 10297 9680 10423
rect 9600 10263 9623 10297
rect 9657 10263 9680 10297
rect 9600 10137 9680 10263
rect 9600 10103 9623 10137
rect 9657 10103 9680 10137
rect 9600 9977 9680 10103
rect 9600 9943 9623 9977
rect 9657 9943 9680 9977
rect 9600 9817 9680 9943
rect 9600 9783 9623 9817
rect 9657 9783 9680 9817
rect 9600 9657 9680 9783
rect 9600 9623 9623 9657
rect 9657 9623 9680 9657
rect 9600 9497 9680 9623
rect 9600 9463 9623 9497
rect 9657 9463 9680 9497
rect 9600 9337 9680 9463
rect 9600 9303 9623 9337
rect 9657 9303 9680 9337
rect 9600 9177 9680 9303
rect 9600 9143 9623 9177
rect 9657 9143 9680 9177
rect 9600 9017 9680 9143
rect 9600 8983 9623 9017
rect 9657 8983 9680 9017
rect 9600 8857 9680 8983
rect 9600 8823 9623 8857
rect 9657 8823 9680 8857
rect 9600 8697 9680 8823
rect 9600 8663 9623 8697
rect 9657 8663 9680 8697
rect 9600 8537 9680 8663
rect 9600 8503 9623 8537
rect 9657 8503 9680 8537
rect 9600 8377 9680 8503
rect 9600 8343 9623 8377
rect 9657 8343 9680 8377
rect 9600 8217 9680 8343
rect 9600 8183 9623 8217
rect 9657 8183 9680 8217
rect 9600 8057 9680 8183
rect 9600 8023 9623 8057
rect 9657 8023 9680 8057
rect 9600 7897 9680 8023
rect 9600 7863 9623 7897
rect 9657 7863 9680 7897
rect 9600 7737 9680 7863
rect 9600 7703 9623 7737
rect 9657 7703 9680 7737
rect 9600 7577 9680 7703
rect 9600 7543 9623 7577
rect 9657 7543 9680 7577
rect 9600 7417 9680 7543
rect 9600 7383 9623 7417
rect 9657 7383 9680 7417
rect 9600 7257 9680 7383
rect 9600 7223 9623 7257
rect 9657 7223 9680 7257
rect 9600 7097 9680 7223
rect 9600 7063 9623 7097
rect 9657 7063 9680 7097
rect 9600 6937 9680 7063
rect 9600 6903 9623 6937
rect 9657 6903 9680 6937
rect 9600 6777 9680 6903
rect 9600 6743 9623 6777
rect 9657 6743 9680 6777
rect 9600 6617 9680 6743
rect 9600 6583 9623 6617
rect 9657 6583 9680 6617
rect 9600 6457 9680 6583
rect 9600 6423 9623 6457
rect 9657 6423 9680 6457
rect 9600 6297 9680 6423
rect 9600 6263 9623 6297
rect 9657 6263 9680 6297
rect 9600 6137 9680 6263
rect 9600 6103 9623 6137
rect 9657 6103 9680 6137
rect 9600 5977 9680 6103
rect 9600 5943 9623 5977
rect 9657 5943 9680 5977
rect 9600 5817 9680 5943
rect 9600 5783 9623 5817
rect 9657 5783 9680 5817
rect 9600 5657 9680 5783
rect 9600 5623 9623 5657
rect 9657 5623 9680 5657
rect 9600 5497 9680 5623
rect 9600 5463 9623 5497
rect 9657 5463 9680 5497
rect 9600 5337 9680 5463
rect 9600 5303 9623 5337
rect 9657 5303 9680 5337
rect 9600 5177 9680 5303
rect 9600 5143 9623 5177
rect 9657 5143 9680 5177
rect 9600 5017 9680 5143
rect 9600 4983 9623 5017
rect 9657 4983 9680 5017
rect 9600 4857 9680 4983
rect 9600 4823 9623 4857
rect 9657 4823 9680 4857
rect 9600 4697 9680 4823
rect 9600 4663 9623 4697
rect 9657 4663 9680 4697
rect 9600 4537 9680 4663
rect 9600 4503 9623 4537
rect 9657 4503 9680 4537
rect 9600 4377 9680 4503
rect 9600 4343 9623 4377
rect 9657 4343 9680 4377
rect 9600 4217 9680 4343
rect 9600 4183 9623 4217
rect 9657 4183 9680 4217
rect 9600 4057 9680 4183
rect 9600 4023 9623 4057
rect 9657 4023 9680 4057
rect 9600 3897 9680 4023
rect 9600 3863 9623 3897
rect 9657 3863 9680 3897
rect 9600 3737 9680 3863
rect 9600 3703 9623 3737
rect 9657 3703 9680 3737
rect 9600 3577 9680 3703
rect 9600 3543 9623 3577
rect 9657 3543 9680 3577
rect 9600 3417 9680 3543
rect 9600 3383 9623 3417
rect 9657 3383 9680 3417
rect 9600 3257 9680 3383
rect 9600 3223 9623 3257
rect 9657 3223 9680 3257
rect 9600 3097 9680 3223
rect 9600 3063 9623 3097
rect 9657 3063 9680 3097
rect 9600 2937 9680 3063
rect 9600 2903 9623 2937
rect 9657 2903 9680 2937
rect 9600 2777 9680 2903
rect 9600 2743 9623 2777
rect 9657 2743 9680 2777
rect 9600 2617 9680 2743
rect 9600 2583 9623 2617
rect 9657 2583 9680 2617
rect 9600 2457 9680 2583
rect 9600 2423 9623 2457
rect 9657 2423 9680 2457
rect 9600 2297 9680 2423
rect 9600 2263 9623 2297
rect 9657 2263 9680 2297
rect 9600 2137 9680 2263
rect 9600 2103 9623 2137
rect 9657 2103 9680 2137
rect 9600 1977 9680 2103
rect 9600 1943 9623 1977
rect 9657 1943 9680 1977
rect 9600 1817 9680 1943
rect 9600 1783 9623 1817
rect 9657 1783 9680 1817
rect 9600 1657 9680 1783
rect 9600 1623 9623 1657
rect 9657 1623 9680 1657
rect 9600 1497 9680 1623
rect 9600 1463 9623 1497
rect 9657 1463 9680 1497
rect 9600 1337 9680 1463
rect 9600 1303 9623 1337
rect 9657 1303 9680 1337
rect 9600 1177 9680 1303
rect 9600 1143 9623 1177
rect 9657 1143 9680 1177
rect 9600 1017 9680 1143
rect 9600 983 9623 1017
rect 9657 983 9680 1017
rect 9600 857 9680 983
rect 9600 823 9623 857
rect 9657 823 9680 857
rect 9600 697 9680 823
rect 9600 663 9623 697
rect 9657 663 9680 697
rect 9600 537 9680 663
rect 9600 503 9623 537
rect 9657 503 9680 537
rect 9600 377 9680 503
rect 9600 343 9623 377
rect 9657 343 9680 377
rect 9600 217 9680 343
rect 9600 183 9623 217
rect 9657 183 9680 217
rect 9600 57 9680 183
rect 9600 23 9623 57
rect 9657 23 9680 57
rect 9600 0 9680 23
rect 9760 31426 9840 31440
rect 9760 31374 9774 31426
rect 9826 31374 9840 31426
rect 9760 31266 9840 31374
rect 9760 31214 9774 31266
rect 9826 31214 9840 31266
rect 9760 31106 9840 31214
rect 9760 31054 9774 31106
rect 9826 31054 9840 31106
rect 9760 30946 9840 31054
rect 9760 30894 9774 30946
rect 9826 30894 9840 30946
rect 9760 30786 9840 30894
rect 9760 30734 9774 30786
rect 9826 30734 9840 30786
rect 9760 30626 9840 30734
rect 9760 30574 9774 30626
rect 9826 30574 9840 30626
rect 9760 30466 9840 30574
rect 9760 30414 9774 30466
rect 9826 30414 9840 30466
rect 9760 30306 9840 30414
rect 9760 30254 9774 30306
rect 9826 30254 9840 30306
rect 9760 30137 9840 30254
rect 9760 30103 9783 30137
rect 9817 30103 9840 30137
rect 9760 29986 9840 30103
rect 9760 29934 9774 29986
rect 9826 29934 9840 29986
rect 9760 29826 9840 29934
rect 9760 29774 9774 29826
rect 9826 29774 9840 29826
rect 9760 29666 9840 29774
rect 9760 29614 9774 29666
rect 9826 29614 9840 29666
rect 9760 29506 9840 29614
rect 9760 29454 9774 29506
rect 9826 29454 9840 29506
rect 9760 29346 9840 29454
rect 9760 29294 9774 29346
rect 9826 29294 9840 29346
rect 9760 29186 9840 29294
rect 9760 29134 9774 29186
rect 9826 29134 9840 29186
rect 9760 29026 9840 29134
rect 9760 28974 9774 29026
rect 9826 28974 9840 29026
rect 9760 28866 9840 28974
rect 9760 28814 9774 28866
rect 9826 28814 9840 28866
rect 9760 28697 9840 28814
rect 9760 28663 9783 28697
rect 9817 28663 9840 28697
rect 9760 28537 9840 28663
rect 9760 28503 9783 28537
rect 9817 28503 9840 28537
rect 9760 28377 9840 28503
rect 9760 28343 9783 28377
rect 9817 28343 9840 28377
rect 9760 28217 9840 28343
rect 9760 28183 9783 28217
rect 9817 28183 9840 28217
rect 9760 28066 9840 28183
rect 9760 28014 9774 28066
rect 9826 28014 9840 28066
rect 9760 27906 9840 28014
rect 9760 27854 9774 27906
rect 9826 27854 9840 27906
rect 9760 27746 9840 27854
rect 9760 27694 9774 27746
rect 9826 27694 9840 27746
rect 9760 27586 9840 27694
rect 9760 27534 9774 27586
rect 9826 27534 9840 27586
rect 9760 27426 9840 27534
rect 9760 27374 9774 27426
rect 9826 27374 9840 27426
rect 9760 27266 9840 27374
rect 9760 27214 9774 27266
rect 9826 27214 9840 27266
rect 9760 27106 9840 27214
rect 9760 27054 9774 27106
rect 9826 27054 9840 27106
rect 9760 26946 9840 27054
rect 9760 26894 9774 26946
rect 9826 26894 9840 26946
rect 9760 26777 9840 26894
rect 9760 26743 9783 26777
rect 9817 26743 9840 26777
rect 9760 26617 9840 26743
rect 9760 26583 9783 26617
rect 9817 26583 9840 26617
rect 9760 26457 9840 26583
rect 9760 26423 9783 26457
rect 9817 26423 9840 26457
rect 9760 26297 9840 26423
rect 9760 26263 9783 26297
rect 9817 26263 9840 26297
rect 9760 26146 9840 26263
rect 9760 26094 9774 26146
rect 9826 26094 9840 26146
rect 9760 25986 9840 26094
rect 9760 25934 9774 25986
rect 9826 25934 9840 25986
rect 9760 25826 9840 25934
rect 9760 25774 9774 25826
rect 9826 25774 9840 25826
rect 9760 25666 9840 25774
rect 9760 25614 9774 25666
rect 9826 25614 9840 25666
rect 9760 25506 9840 25614
rect 9760 25454 9774 25506
rect 9826 25454 9840 25506
rect 9760 25346 9840 25454
rect 9760 25294 9774 25346
rect 9826 25294 9840 25346
rect 9760 25186 9840 25294
rect 9760 25134 9774 25186
rect 9826 25134 9840 25186
rect 9760 25026 9840 25134
rect 9760 24974 9774 25026
rect 9826 24974 9840 25026
rect 9760 24857 9840 24974
rect 9760 24823 9783 24857
rect 9817 24823 9840 24857
rect 9760 24706 9840 24823
rect 9760 24654 9774 24706
rect 9826 24654 9840 24706
rect 9760 24546 9840 24654
rect 9760 24494 9774 24546
rect 9826 24494 9840 24546
rect 9760 24386 9840 24494
rect 9760 24334 9774 24386
rect 9826 24334 9840 24386
rect 9760 24226 9840 24334
rect 9760 24174 9774 24226
rect 9826 24174 9840 24226
rect 9760 24066 9840 24174
rect 9760 24014 9774 24066
rect 9826 24014 9840 24066
rect 9760 23906 9840 24014
rect 9760 23854 9774 23906
rect 9826 23854 9840 23906
rect 9760 23746 9840 23854
rect 9760 23694 9774 23746
rect 9826 23694 9840 23746
rect 9760 23586 9840 23694
rect 9760 23534 9774 23586
rect 9826 23534 9840 23586
rect 9760 23426 9840 23534
rect 9760 23374 9774 23426
rect 9826 23374 9840 23426
rect 9760 23266 9840 23374
rect 9760 23214 9774 23266
rect 9826 23214 9840 23266
rect 9760 23106 9840 23214
rect 9760 23054 9774 23106
rect 9826 23054 9840 23106
rect 9760 22946 9840 23054
rect 9760 22894 9774 22946
rect 9826 22894 9840 22946
rect 9760 22786 9840 22894
rect 9760 22734 9774 22786
rect 9826 22734 9840 22786
rect 9760 22626 9840 22734
rect 9760 22574 9774 22626
rect 9826 22574 9840 22626
rect 9760 22466 9840 22574
rect 9760 22414 9774 22466
rect 9826 22414 9840 22466
rect 9760 22306 9840 22414
rect 9760 22254 9774 22306
rect 9826 22254 9840 22306
rect 9760 22146 9840 22254
rect 9760 22094 9774 22146
rect 9826 22094 9840 22146
rect 9760 21977 9840 22094
rect 9760 21943 9783 21977
rect 9817 21943 9840 21977
rect 9760 21826 9840 21943
rect 9760 21774 9774 21826
rect 9826 21774 9840 21826
rect 9760 21666 9840 21774
rect 9760 21614 9774 21666
rect 9826 21614 9840 21666
rect 9760 21506 9840 21614
rect 9760 21454 9774 21506
rect 9826 21454 9840 21506
rect 9760 21346 9840 21454
rect 9760 21294 9774 21346
rect 9826 21294 9840 21346
rect 9760 21186 9840 21294
rect 9760 21134 9774 21186
rect 9826 21134 9840 21186
rect 9760 21026 9840 21134
rect 9760 20974 9774 21026
rect 9826 20974 9840 21026
rect 9760 20866 9840 20974
rect 9760 20814 9774 20866
rect 9826 20814 9840 20866
rect 9760 20706 9840 20814
rect 9760 20654 9774 20706
rect 9826 20654 9840 20706
rect 9760 20537 9840 20654
rect 9760 20503 9783 20537
rect 9817 20503 9840 20537
rect 9760 20377 9840 20503
rect 9760 20343 9783 20377
rect 9817 20343 9840 20377
rect 9760 20217 9840 20343
rect 9760 20183 9783 20217
rect 9817 20183 9840 20217
rect 9760 20057 9840 20183
rect 9760 20023 9783 20057
rect 9817 20023 9840 20057
rect 9760 19906 9840 20023
rect 9760 19854 9774 19906
rect 9826 19854 9840 19906
rect 9760 19746 9840 19854
rect 9760 19694 9774 19746
rect 9826 19694 9840 19746
rect 9760 19586 9840 19694
rect 9760 19534 9774 19586
rect 9826 19534 9840 19586
rect 9760 19426 9840 19534
rect 9760 19374 9774 19426
rect 9826 19374 9840 19426
rect 9760 19266 9840 19374
rect 9760 19214 9774 19266
rect 9826 19214 9840 19266
rect 9760 19106 9840 19214
rect 9760 19054 9774 19106
rect 9826 19054 9840 19106
rect 9760 18946 9840 19054
rect 9760 18894 9774 18946
rect 9826 18894 9840 18946
rect 9760 18786 9840 18894
rect 9760 18734 9774 18786
rect 9826 18734 9840 18786
rect 9760 18617 9840 18734
rect 9760 18583 9783 18617
rect 9817 18583 9840 18617
rect 9760 18457 9840 18583
rect 9760 18423 9783 18457
rect 9817 18423 9840 18457
rect 9760 18297 9840 18423
rect 9760 18263 9783 18297
rect 9817 18263 9840 18297
rect 9760 18137 9840 18263
rect 9760 18103 9783 18137
rect 9817 18103 9840 18137
rect 9760 17986 9840 18103
rect 9760 17934 9774 17986
rect 9826 17934 9840 17986
rect 9760 17826 9840 17934
rect 9760 17774 9774 17826
rect 9826 17774 9840 17826
rect 9760 17666 9840 17774
rect 9760 17614 9774 17666
rect 9826 17614 9840 17666
rect 9760 17506 9840 17614
rect 9760 17454 9774 17506
rect 9826 17454 9840 17506
rect 9760 17346 9840 17454
rect 9760 17294 9774 17346
rect 9826 17294 9840 17346
rect 9760 17186 9840 17294
rect 9760 17134 9774 17186
rect 9826 17134 9840 17186
rect 9760 17026 9840 17134
rect 9760 16974 9774 17026
rect 9826 16974 9840 17026
rect 9760 16866 9840 16974
rect 9760 16814 9774 16866
rect 9826 16814 9840 16866
rect 9760 16697 9840 16814
rect 9760 16663 9783 16697
rect 9817 16663 9840 16697
rect 9760 16546 9840 16663
rect 9760 16494 9774 16546
rect 9826 16494 9840 16546
rect 9760 16386 9840 16494
rect 9760 16334 9774 16386
rect 9826 16334 9840 16386
rect 9760 16226 9840 16334
rect 9760 16174 9774 16226
rect 9826 16174 9840 16226
rect 9760 16066 9840 16174
rect 9760 16014 9774 16066
rect 9826 16014 9840 16066
rect 9760 15906 9840 16014
rect 9760 15854 9774 15906
rect 9826 15854 9840 15906
rect 9760 15746 9840 15854
rect 9760 15694 9774 15746
rect 9826 15694 9840 15746
rect 9760 15586 9840 15694
rect 9760 15534 9774 15586
rect 9826 15534 9840 15586
rect 9760 15426 9840 15534
rect 9760 15374 9774 15426
rect 9826 15374 9840 15426
rect 9760 15266 9840 15374
rect 9760 15214 9774 15266
rect 9826 15214 9840 15266
rect 9760 15106 9840 15214
rect 9760 15054 9774 15106
rect 9826 15054 9840 15106
rect 9760 14946 9840 15054
rect 9760 14894 9774 14946
rect 9826 14894 9840 14946
rect 9760 14786 9840 14894
rect 9760 14734 9774 14786
rect 9826 14734 9840 14786
rect 9760 14626 9840 14734
rect 9760 14574 9774 14626
rect 9826 14574 9840 14626
rect 9760 14466 9840 14574
rect 9760 14414 9774 14466
rect 9826 14414 9840 14466
rect 9760 14306 9840 14414
rect 9760 14254 9774 14306
rect 9826 14254 9840 14306
rect 9760 14146 9840 14254
rect 9760 14094 9774 14146
rect 9826 14094 9840 14146
rect 9760 13986 9840 14094
rect 9760 13934 9774 13986
rect 9826 13934 9840 13986
rect 9760 13817 9840 13934
rect 9760 13783 9783 13817
rect 9817 13783 9840 13817
rect 9760 13666 9840 13783
rect 9760 13614 9774 13666
rect 9826 13614 9840 13666
rect 9760 13506 9840 13614
rect 9760 13454 9774 13506
rect 9826 13454 9840 13506
rect 9760 13346 9840 13454
rect 9760 13294 9774 13346
rect 9826 13294 9840 13346
rect 9760 13186 9840 13294
rect 9760 13134 9774 13186
rect 9826 13134 9840 13186
rect 9760 13026 9840 13134
rect 9760 12974 9774 13026
rect 9826 12974 9840 13026
rect 9760 12866 9840 12974
rect 9760 12814 9774 12866
rect 9826 12814 9840 12866
rect 9760 12706 9840 12814
rect 9760 12654 9774 12706
rect 9826 12654 9840 12706
rect 9760 12546 9840 12654
rect 9760 12494 9774 12546
rect 9826 12494 9840 12546
rect 9760 12377 9840 12494
rect 9760 12343 9783 12377
rect 9817 12343 9840 12377
rect 9760 12217 9840 12343
rect 9760 12183 9783 12217
rect 9817 12183 9840 12217
rect 9760 12057 9840 12183
rect 9760 12023 9783 12057
rect 9817 12023 9840 12057
rect 9760 11897 9840 12023
rect 9760 11863 9783 11897
rect 9817 11863 9840 11897
rect 9760 11746 9840 11863
rect 9760 11694 9774 11746
rect 9826 11694 9840 11746
rect 9760 11586 9840 11694
rect 9760 11534 9774 11586
rect 9826 11534 9840 11586
rect 9760 11426 9840 11534
rect 9760 11374 9774 11426
rect 9826 11374 9840 11426
rect 9760 11266 9840 11374
rect 9760 11214 9774 11266
rect 9826 11214 9840 11266
rect 9760 11106 9840 11214
rect 9760 11054 9774 11106
rect 9826 11054 9840 11106
rect 9760 10946 9840 11054
rect 9760 10894 9774 10946
rect 9826 10894 9840 10946
rect 9760 10786 9840 10894
rect 9760 10734 9774 10786
rect 9826 10734 9840 10786
rect 9760 10626 9840 10734
rect 9760 10574 9774 10626
rect 9826 10574 9840 10626
rect 9760 10466 9840 10574
rect 9760 10414 9774 10466
rect 9826 10414 9840 10466
rect 9760 10306 9840 10414
rect 9760 10254 9774 10306
rect 9826 10254 9840 10306
rect 9760 10146 9840 10254
rect 9760 10094 9774 10146
rect 9826 10094 9840 10146
rect 9760 9986 9840 10094
rect 9760 9934 9774 9986
rect 9826 9934 9840 9986
rect 9760 9826 9840 9934
rect 9760 9774 9774 9826
rect 9826 9774 9840 9826
rect 9760 9657 9840 9774
rect 9760 9623 9783 9657
rect 9817 9623 9840 9657
rect 9760 9506 9840 9623
rect 9760 9454 9774 9506
rect 9826 9454 9840 9506
rect 9760 9346 9840 9454
rect 9760 9294 9774 9346
rect 9826 9294 9840 9346
rect 9760 9177 9840 9294
rect 9760 9143 9783 9177
rect 9817 9143 9840 9177
rect 9760 9026 9840 9143
rect 9760 8974 9774 9026
rect 9826 8974 9840 9026
rect 9760 8866 9840 8974
rect 9760 8814 9774 8866
rect 9826 8814 9840 8866
rect 9760 8706 9840 8814
rect 9760 8654 9774 8706
rect 9826 8654 9840 8706
rect 9760 8546 9840 8654
rect 9760 8494 9774 8546
rect 9826 8494 9840 8546
rect 9760 8386 9840 8494
rect 9760 8334 9774 8386
rect 9826 8334 9840 8386
rect 9760 8226 9840 8334
rect 9760 8174 9774 8226
rect 9826 8174 9840 8226
rect 9760 8066 9840 8174
rect 9760 8014 9774 8066
rect 9826 8014 9840 8066
rect 9760 7906 9840 8014
rect 9760 7854 9774 7906
rect 9826 7854 9840 7906
rect 9760 7746 9840 7854
rect 9760 7694 9774 7746
rect 9826 7694 9840 7746
rect 9760 7577 9840 7694
rect 9760 7543 9783 7577
rect 9817 7543 9840 7577
rect 9760 7426 9840 7543
rect 9760 7374 9774 7426
rect 9826 7374 9840 7426
rect 9760 7266 9840 7374
rect 9760 7214 9774 7266
rect 9826 7214 9840 7266
rect 9760 7097 9840 7214
rect 9760 7063 9783 7097
rect 9817 7063 9840 7097
rect 9760 6946 9840 7063
rect 9760 6894 9774 6946
rect 9826 6894 9840 6946
rect 9760 6786 9840 6894
rect 9760 6734 9774 6786
rect 9826 6734 9840 6786
rect 9760 6617 9840 6734
rect 9760 6583 9783 6617
rect 9817 6583 9840 6617
rect 9760 6466 9840 6583
rect 9760 6414 9774 6466
rect 9826 6414 9840 6466
rect 9760 6306 9840 6414
rect 9760 6254 9774 6306
rect 9826 6254 9840 6306
rect 9760 6146 9840 6254
rect 9760 6094 9774 6146
rect 9826 6094 9840 6146
rect 9760 5986 9840 6094
rect 9760 5934 9774 5986
rect 9826 5934 9840 5986
rect 9760 5826 9840 5934
rect 9760 5774 9774 5826
rect 9826 5774 9840 5826
rect 9760 5666 9840 5774
rect 9760 5614 9774 5666
rect 9826 5614 9840 5666
rect 9760 5506 9840 5614
rect 9760 5454 9774 5506
rect 9826 5454 9840 5506
rect 9760 5346 9840 5454
rect 9760 5294 9774 5346
rect 9826 5294 9840 5346
rect 9760 5186 9840 5294
rect 9760 5134 9774 5186
rect 9826 5134 9840 5186
rect 9760 5026 9840 5134
rect 9760 4974 9774 5026
rect 9826 4974 9840 5026
rect 9760 4866 9840 4974
rect 9760 4814 9774 4866
rect 9826 4814 9840 4866
rect 9760 4706 9840 4814
rect 9760 4654 9774 4706
rect 9826 4654 9840 4706
rect 9760 4546 9840 4654
rect 9760 4494 9774 4546
rect 9826 4494 9840 4546
rect 9760 4386 9840 4494
rect 9760 4334 9774 4386
rect 9826 4334 9840 4386
rect 9760 4226 9840 4334
rect 9760 4174 9774 4226
rect 9826 4174 9840 4226
rect 9760 4066 9840 4174
rect 9760 4014 9774 4066
rect 9826 4014 9840 4066
rect 9760 3906 9840 4014
rect 9760 3854 9774 3906
rect 9826 3854 9840 3906
rect 9760 3737 9840 3854
rect 9760 3703 9783 3737
rect 9817 3703 9840 3737
rect 9760 3577 9840 3703
rect 9760 3543 9783 3577
rect 9817 3543 9840 3577
rect 9760 3426 9840 3543
rect 9760 3374 9774 3426
rect 9826 3374 9840 3426
rect 9760 3266 9840 3374
rect 9760 3214 9774 3266
rect 9826 3214 9840 3266
rect 9760 3106 9840 3214
rect 9760 3054 9774 3106
rect 9826 3054 9840 3106
rect 9760 2946 9840 3054
rect 9760 2894 9774 2946
rect 9826 2894 9840 2946
rect 9760 2786 9840 2894
rect 9760 2734 9774 2786
rect 9826 2734 9840 2786
rect 9760 2626 9840 2734
rect 9760 2574 9774 2626
rect 9826 2574 9840 2626
rect 9760 2466 9840 2574
rect 9760 2414 9774 2466
rect 9826 2414 9840 2466
rect 9760 2306 9840 2414
rect 9760 2254 9774 2306
rect 9826 2254 9840 2306
rect 9760 2146 9840 2254
rect 9760 2094 9774 2146
rect 9826 2094 9840 2146
rect 9760 1986 9840 2094
rect 9760 1934 9774 1986
rect 9826 1934 9840 1986
rect 9760 1817 9840 1934
rect 9760 1783 9783 1817
rect 9817 1783 9840 1817
rect 9760 1666 9840 1783
rect 9760 1614 9774 1666
rect 9826 1614 9840 1666
rect 9760 1506 9840 1614
rect 9760 1454 9774 1506
rect 9826 1454 9840 1506
rect 9760 1346 9840 1454
rect 9760 1294 9774 1346
rect 9826 1294 9840 1346
rect 9760 1186 9840 1294
rect 9760 1134 9774 1186
rect 9826 1134 9840 1186
rect 9760 1026 9840 1134
rect 9760 974 9774 1026
rect 9826 974 9840 1026
rect 9760 857 9840 974
rect 9760 823 9783 857
rect 9817 823 9840 857
rect 9760 697 9840 823
rect 9760 663 9783 697
rect 9817 663 9840 697
rect 9760 546 9840 663
rect 9760 494 9774 546
rect 9826 494 9840 546
rect 9760 386 9840 494
rect 9760 334 9774 386
rect 9826 334 9840 386
rect 9760 226 9840 334
rect 9760 174 9774 226
rect 9826 174 9840 226
rect 9760 66 9840 174
rect 9760 14 9774 66
rect 9826 14 9840 66
rect 9760 0 9840 14
rect 9920 31417 10000 31440
rect 9920 31383 9943 31417
rect 9977 31383 10000 31417
rect 9920 31257 10000 31383
rect 9920 31223 9943 31257
rect 9977 31223 10000 31257
rect 9920 31097 10000 31223
rect 9920 31063 9943 31097
rect 9977 31063 10000 31097
rect 9920 30937 10000 31063
rect 9920 30903 9943 30937
rect 9977 30903 10000 30937
rect 9920 30777 10000 30903
rect 9920 30743 9943 30777
rect 9977 30743 10000 30777
rect 9920 30617 10000 30743
rect 9920 30583 9943 30617
rect 9977 30583 10000 30617
rect 9920 30457 10000 30583
rect 9920 30423 9943 30457
rect 9977 30423 10000 30457
rect 9920 30297 10000 30423
rect 9920 30263 9943 30297
rect 9977 30263 10000 30297
rect 9920 30137 10000 30263
rect 9920 30103 9943 30137
rect 9977 30103 10000 30137
rect 9920 29977 10000 30103
rect 9920 29943 9943 29977
rect 9977 29943 10000 29977
rect 9920 29817 10000 29943
rect 9920 29783 9943 29817
rect 9977 29783 10000 29817
rect 9920 29657 10000 29783
rect 9920 29623 9943 29657
rect 9977 29623 10000 29657
rect 9920 29497 10000 29623
rect 9920 29463 9943 29497
rect 9977 29463 10000 29497
rect 9920 29337 10000 29463
rect 9920 29303 9943 29337
rect 9977 29303 10000 29337
rect 9920 29177 10000 29303
rect 9920 29143 9943 29177
rect 9977 29143 10000 29177
rect 9920 29017 10000 29143
rect 9920 28983 9943 29017
rect 9977 28983 10000 29017
rect 9920 28857 10000 28983
rect 9920 28823 9943 28857
rect 9977 28823 10000 28857
rect 9920 28697 10000 28823
rect 9920 28663 9943 28697
rect 9977 28663 10000 28697
rect 9920 28537 10000 28663
rect 9920 28503 9943 28537
rect 9977 28503 10000 28537
rect 9920 28377 10000 28503
rect 9920 28343 9943 28377
rect 9977 28343 10000 28377
rect 9920 28217 10000 28343
rect 9920 28183 9943 28217
rect 9977 28183 10000 28217
rect 9920 28057 10000 28183
rect 9920 28023 9943 28057
rect 9977 28023 10000 28057
rect 9920 27897 10000 28023
rect 9920 27863 9943 27897
rect 9977 27863 10000 27897
rect 9920 27737 10000 27863
rect 9920 27703 9943 27737
rect 9977 27703 10000 27737
rect 9920 27577 10000 27703
rect 9920 27543 9943 27577
rect 9977 27543 10000 27577
rect 9920 27417 10000 27543
rect 9920 27383 9943 27417
rect 9977 27383 10000 27417
rect 9920 27257 10000 27383
rect 9920 27223 9943 27257
rect 9977 27223 10000 27257
rect 9920 27097 10000 27223
rect 9920 27063 9943 27097
rect 9977 27063 10000 27097
rect 9920 26937 10000 27063
rect 9920 26903 9943 26937
rect 9977 26903 10000 26937
rect 9920 26777 10000 26903
rect 9920 26743 9943 26777
rect 9977 26743 10000 26777
rect 9920 26617 10000 26743
rect 9920 26583 9943 26617
rect 9977 26583 10000 26617
rect 9920 26457 10000 26583
rect 9920 26423 9943 26457
rect 9977 26423 10000 26457
rect 9920 26297 10000 26423
rect 9920 26263 9943 26297
rect 9977 26263 10000 26297
rect 9920 26137 10000 26263
rect 9920 26103 9943 26137
rect 9977 26103 10000 26137
rect 9920 25977 10000 26103
rect 9920 25943 9943 25977
rect 9977 25943 10000 25977
rect 9920 25817 10000 25943
rect 9920 25783 9943 25817
rect 9977 25783 10000 25817
rect 9920 25657 10000 25783
rect 9920 25623 9943 25657
rect 9977 25623 10000 25657
rect 9920 25497 10000 25623
rect 9920 25463 9943 25497
rect 9977 25463 10000 25497
rect 9920 25337 10000 25463
rect 9920 25303 9943 25337
rect 9977 25303 10000 25337
rect 9920 25177 10000 25303
rect 9920 25143 9943 25177
rect 9977 25143 10000 25177
rect 9920 25017 10000 25143
rect 9920 24983 9943 25017
rect 9977 24983 10000 25017
rect 9920 24857 10000 24983
rect 9920 24823 9943 24857
rect 9977 24823 10000 24857
rect 9920 24697 10000 24823
rect 9920 24663 9943 24697
rect 9977 24663 10000 24697
rect 9920 24537 10000 24663
rect 9920 24503 9943 24537
rect 9977 24503 10000 24537
rect 9920 24377 10000 24503
rect 9920 24343 9943 24377
rect 9977 24343 10000 24377
rect 9920 24217 10000 24343
rect 9920 24183 9943 24217
rect 9977 24183 10000 24217
rect 9920 24057 10000 24183
rect 9920 24023 9943 24057
rect 9977 24023 10000 24057
rect 9920 23897 10000 24023
rect 9920 23863 9943 23897
rect 9977 23863 10000 23897
rect 9920 23737 10000 23863
rect 9920 23703 9943 23737
rect 9977 23703 10000 23737
rect 9920 23577 10000 23703
rect 9920 23543 9943 23577
rect 9977 23543 10000 23577
rect 9920 23417 10000 23543
rect 9920 23383 9943 23417
rect 9977 23383 10000 23417
rect 9920 23257 10000 23383
rect 9920 23223 9943 23257
rect 9977 23223 10000 23257
rect 9920 23097 10000 23223
rect 9920 23063 9943 23097
rect 9977 23063 10000 23097
rect 9920 22937 10000 23063
rect 9920 22903 9943 22937
rect 9977 22903 10000 22937
rect 9920 22777 10000 22903
rect 9920 22743 9943 22777
rect 9977 22743 10000 22777
rect 9920 22617 10000 22743
rect 9920 22583 9943 22617
rect 9977 22583 10000 22617
rect 9920 22457 10000 22583
rect 9920 22423 9943 22457
rect 9977 22423 10000 22457
rect 9920 22297 10000 22423
rect 9920 22263 9943 22297
rect 9977 22263 10000 22297
rect 9920 22137 10000 22263
rect 9920 22103 9943 22137
rect 9977 22103 10000 22137
rect 9920 21977 10000 22103
rect 9920 21943 9943 21977
rect 9977 21943 10000 21977
rect 9920 21817 10000 21943
rect 9920 21783 9943 21817
rect 9977 21783 10000 21817
rect 9920 21657 10000 21783
rect 9920 21623 9943 21657
rect 9977 21623 10000 21657
rect 9920 21497 10000 21623
rect 9920 21463 9943 21497
rect 9977 21463 10000 21497
rect 9920 21337 10000 21463
rect 9920 21303 9943 21337
rect 9977 21303 10000 21337
rect 9920 21177 10000 21303
rect 9920 21143 9943 21177
rect 9977 21143 10000 21177
rect 9920 21017 10000 21143
rect 9920 20983 9943 21017
rect 9977 20983 10000 21017
rect 9920 20857 10000 20983
rect 9920 20823 9943 20857
rect 9977 20823 10000 20857
rect 9920 20697 10000 20823
rect 9920 20663 9943 20697
rect 9977 20663 10000 20697
rect 9920 20537 10000 20663
rect 9920 20503 9943 20537
rect 9977 20503 10000 20537
rect 9920 20377 10000 20503
rect 9920 20343 9943 20377
rect 9977 20343 10000 20377
rect 9920 20217 10000 20343
rect 9920 20183 9943 20217
rect 9977 20183 10000 20217
rect 9920 20057 10000 20183
rect 9920 20023 9943 20057
rect 9977 20023 10000 20057
rect 9920 19897 10000 20023
rect 9920 19863 9943 19897
rect 9977 19863 10000 19897
rect 9920 19737 10000 19863
rect 9920 19703 9943 19737
rect 9977 19703 10000 19737
rect 9920 19577 10000 19703
rect 9920 19543 9943 19577
rect 9977 19543 10000 19577
rect 9920 19417 10000 19543
rect 9920 19383 9943 19417
rect 9977 19383 10000 19417
rect 9920 19257 10000 19383
rect 9920 19223 9943 19257
rect 9977 19223 10000 19257
rect 9920 19097 10000 19223
rect 9920 19063 9943 19097
rect 9977 19063 10000 19097
rect 9920 18937 10000 19063
rect 9920 18903 9943 18937
rect 9977 18903 10000 18937
rect 9920 18777 10000 18903
rect 9920 18743 9943 18777
rect 9977 18743 10000 18777
rect 9920 18617 10000 18743
rect 9920 18583 9943 18617
rect 9977 18583 10000 18617
rect 9920 18457 10000 18583
rect 9920 18423 9943 18457
rect 9977 18423 10000 18457
rect 9920 18297 10000 18423
rect 9920 18263 9943 18297
rect 9977 18263 10000 18297
rect 9920 18137 10000 18263
rect 9920 18103 9943 18137
rect 9977 18103 10000 18137
rect 9920 17977 10000 18103
rect 9920 17943 9943 17977
rect 9977 17943 10000 17977
rect 9920 17817 10000 17943
rect 9920 17783 9943 17817
rect 9977 17783 10000 17817
rect 9920 17657 10000 17783
rect 9920 17623 9943 17657
rect 9977 17623 10000 17657
rect 9920 17497 10000 17623
rect 9920 17463 9943 17497
rect 9977 17463 10000 17497
rect 9920 17337 10000 17463
rect 9920 17303 9943 17337
rect 9977 17303 10000 17337
rect 9920 17177 10000 17303
rect 9920 17143 9943 17177
rect 9977 17143 10000 17177
rect 9920 17017 10000 17143
rect 9920 16983 9943 17017
rect 9977 16983 10000 17017
rect 9920 16857 10000 16983
rect 9920 16823 9943 16857
rect 9977 16823 10000 16857
rect 9920 16697 10000 16823
rect 9920 16663 9943 16697
rect 9977 16663 10000 16697
rect 9920 16537 10000 16663
rect 9920 16503 9943 16537
rect 9977 16503 10000 16537
rect 9920 16377 10000 16503
rect 9920 16343 9943 16377
rect 9977 16343 10000 16377
rect 9920 16217 10000 16343
rect 9920 16183 9943 16217
rect 9977 16183 10000 16217
rect 9920 16057 10000 16183
rect 9920 16023 9943 16057
rect 9977 16023 10000 16057
rect 9920 15897 10000 16023
rect 9920 15863 9943 15897
rect 9977 15863 10000 15897
rect 9920 15737 10000 15863
rect 9920 15703 9943 15737
rect 9977 15703 10000 15737
rect 9920 15577 10000 15703
rect 9920 15543 9943 15577
rect 9977 15543 10000 15577
rect 9920 15417 10000 15543
rect 9920 15383 9943 15417
rect 9977 15383 10000 15417
rect 9920 15257 10000 15383
rect 9920 15223 9943 15257
rect 9977 15223 10000 15257
rect 9920 15097 10000 15223
rect 9920 15063 9943 15097
rect 9977 15063 10000 15097
rect 9920 14937 10000 15063
rect 9920 14903 9943 14937
rect 9977 14903 10000 14937
rect 9920 14777 10000 14903
rect 9920 14743 9943 14777
rect 9977 14743 10000 14777
rect 9920 14617 10000 14743
rect 9920 14583 9943 14617
rect 9977 14583 10000 14617
rect 9920 14457 10000 14583
rect 9920 14423 9943 14457
rect 9977 14423 10000 14457
rect 9920 14297 10000 14423
rect 9920 14263 9943 14297
rect 9977 14263 10000 14297
rect 9920 14137 10000 14263
rect 9920 14103 9943 14137
rect 9977 14103 10000 14137
rect 9920 13977 10000 14103
rect 9920 13943 9943 13977
rect 9977 13943 10000 13977
rect 9920 13817 10000 13943
rect 9920 13783 9943 13817
rect 9977 13783 10000 13817
rect 9920 13657 10000 13783
rect 9920 13623 9943 13657
rect 9977 13623 10000 13657
rect 9920 13497 10000 13623
rect 9920 13463 9943 13497
rect 9977 13463 10000 13497
rect 9920 13337 10000 13463
rect 9920 13303 9943 13337
rect 9977 13303 10000 13337
rect 9920 13177 10000 13303
rect 9920 13143 9943 13177
rect 9977 13143 10000 13177
rect 9920 13017 10000 13143
rect 9920 12983 9943 13017
rect 9977 12983 10000 13017
rect 9920 12857 10000 12983
rect 9920 12823 9943 12857
rect 9977 12823 10000 12857
rect 9920 12697 10000 12823
rect 9920 12663 9943 12697
rect 9977 12663 10000 12697
rect 9920 12537 10000 12663
rect 9920 12503 9943 12537
rect 9977 12503 10000 12537
rect 9920 12377 10000 12503
rect 9920 12343 9943 12377
rect 9977 12343 10000 12377
rect 9920 12217 10000 12343
rect 9920 12183 9943 12217
rect 9977 12183 10000 12217
rect 9920 12057 10000 12183
rect 9920 12023 9943 12057
rect 9977 12023 10000 12057
rect 9920 11897 10000 12023
rect 9920 11863 9943 11897
rect 9977 11863 10000 11897
rect 9920 11737 10000 11863
rect 9920 11703 9943 11737
rect 9977 11703 10000 11737
rect 9920 11577 10000 11703
rect 9920 11543 9943 11577
rect 9977 11543 10000 11577
rect 9920 11417 10000 11543
rect 9920 11383 9943 11417
rect 9977 11383 10000 11417
rect 9920 11257 10000 11383
rect 9920 11223 9943 11257
rect 9977 11223 10000 11257
rect 9920 11097 10000 11223
rect 9920 11063 9943 11097
rect 9977 11063 10000 11097
rect 9920 10937 10000 11063
rect 9920 10903 9943 10937
rect 9977 10903 10000 10937
rect 9920 10777 10000 10903
rect 9920 10743 9943 10777
rect 9977 10743 10000 10777
rect 9920 10617 10000 10743
rect 9920 10583 9943 10617
rect 9977 10583 10000 10617
rect 9920 10457 10000 10583
rect 9920 10423 9943 10457
rect 9977 10423 10000 10457
rect 9920 10297 10000 10423
rect 9920 10263 9943 10297
rect 9977 10263 10000 10297
rect 9920 10137 10000 10263
rect 9920 10103 9943 10137
rect 9977 10103 10000 10137
rect 9920 9977 10000 10103
rect 9920 9943 9943 9977
rect 9977 9943 10000 9977
rect 9920 9817 10000 9943
rect 9920 9783 9943 9817
rect 9977 9783 10000 9817
rect 9920 9657 10000 9783
rect 9920 9623 9943 9657
rect 9977 9623 10000 9657
rect 9920 9497 10000 9623
rect 9920 9463 9943 9497
rect 9977 9463 10000 9497
rect 9920 9337 10000 9463
rect 9920 9303 9943 9337
rect 9977 9303 10000 9337
rect 9920 9177 10000 9303
rect 9920 9143 9943 9177
rect 9977 9143 10000 9177
rect 9920 9017 10000 9143
rect 9920 8983 9943 9017
rect 9977 8983 10000 9017
rect 9920 8857 10000 8983
rect 9920 8823 9943 8857
rect 9977 8823 10000 8857
rect 9920 8697 10000 8823
rect 9920 8663 9943 8697
rect 9977 8663 10000 8697
rect 9920 8537 10000 8663
rect 9920 8503 9943 8537
rect 9977 8503 10000 8537
rect 9920 8377 10000 8503
rect 9920 8343 9943 8377
rect 9977 8343 10000 8377
rect 9920 8217 10000 8343
rect 9920 8183 9943 8217
rect 9977 8183 10000 8217
rect 9920 8057 10000 8183
rect 9920 8023 9943 8057
rect 9977 8023 10000 8057
rect 9920 7897 10000 8023
rect 9920 7863 9943 7897
rect 9977 7863 10000 7897
rect 9920 7737 10000 7863
rect 9920 7703 9943 7737
rect 9977 7703 10000 7737
rect 9920 7577 10000 7703
rect 9920 7543 9943 7577
rect 9977 7543 10000 7577
rect 9920 7417 10000 7543
rect 9920 7383 9943 7417
rect 9977 7383 10000 7417
rect 9920 7257 10000 7383
rect 9920 7223 9943 7257
rect 9977 7223 10000 7257
rect 9920 7097 10000 7223
rect 9920 7063 9943 7097
rect 9977 7063 10000 7097
rect 9920 6937 10000 7063
rect 9920 6903 9943 6937
rect 9977 6903 10000 6937
rect 9920 6777 10000 6903
rect 9920 6743 9943 6777
rect 9977 6743 10000 6777
rect 9920 6617 10000 6743
rect 9920 6583 9943 6617
rect 9977 6583 10000 6617
rect 9920 6457 10000 6583
rect 9920 6423 9943 6457
rect 9977 6423 10000 6457
rect 9920 6297 10000 6423
rect 9920 6263 9943 6297
rect 9977 6263 10000 6297
rect 9920 6137 10000 6263
rect 9920 6103 9943 6137
rect 9977 6103 10000 6137
rect 9920 5977 10000 6103
rect 9920 5943 9943 5977
rect 9977 5943 10000 5977
rect 9920 5817 10000 5943
rect 9920 5783 9943 5817
rect 9977 5783 10000 5817
rect 9920 5657 10000 5783
rect 9920 5623 9943 5657
rect 9977 5623 10000 5657
rect 9920 5497 10000 5623
rect 9920 5463 9943 5497
rect 9977 5463 10000 5497
rect 9920 5337 10000 5463
rect 9920 5303 9943 5337
rect 9977 5303 10000 5337
rect 9920 5177 10000 5303
rect 9920 5143 9943 5177
rect 9977 5143 10000 5177
rect 9920 5017 10000 5143
rect 9920 4983 9943 5017
rect 9977 4983 10000 5017
rect 9920 4857 10000 4983
rect 9920 4823 9943 4857
rect 9977 4823 10000 4857
rect 9920 4697 10000 4823
rect 9920 4663 9943 4697
rect 9977 4663 10000 4697
rect 9920 4537 10000 4663
rect 9920 4503 9943 4537
rect 9977 4503 10000 4537
rect 9920 4377 10000 4503
rect 9920 4343 9943 4377
rect 9977 4343 10000 4377
rect 9920 4217 10000 4343
rect 9920 4183 9943 4217
rect 9977 4183 10000 4217
rect 9920 4057 10000 4183
rect 9920 4023 9943 4057
rect 9977 4023 10000 4057
rect 9920 3897 10000 4023
rect 9920 3863 9943 3897
rect 9977 3863 10000 3897
rect 9920 3737 10000 3863
rect 9920 3703 9943 3737
rect 9977 3703 10000 3737
rect 9920 3577 10000 3703
rect 9920 3543 9943 3577
rect 9977 3543 10000 3577
rect 9920 3417 10000 3543
rect 9920 3383 9943 3417
rect 9977 3383 10000 3417
rect 9920 3257 10000 3383
rect 9920 3223 9943 3257
rect 9977 3223 10000 3257
rect 9920 3097 10000 3223
rect 9920 3063 9943 3097
rect 9977 3063 10000 3097
rect 9920 2937 10000 3063
rect 9920 2903 9943 2937
rect 9977 2903 10000 2937
rect 9920 2777 10000 2903
rect 9920 2743 9943 2777
rect 9977 2743 10000 2777
rect 9920 2617 10000 2743
rect 9920 2583 9943 2617
rect 9977 2583 10000 2617
rect 9920 2457 10000 2583
rect 9920 2423 9943 2457
rect 9977 2423 10000 2457
rect 9920 2297 10000 2423
rect 9920 2263 9943 2297
rect 9977 2263 10000 2297
rect 9920 2137 10000 2263
rect 9920 2103 9943 2137
rect 9977 2103 10000 2137
rect 9920 1977 10000 2103
rect 9920 1943 9943 1977
rect 9977 1943 10000 1977
rect 9920 1817 10000 1943
rect 9920 1783 9943 1817
rect 9977 1783 10000 1817
rect 9920 1657 10000 1783
rect 9920 1623 9943 1657
rect 9977 1623 10000 1657
rect 9920 1497 10000 1623
rect 9920 1463 9943 1497
rect 9977 1463 10000 1497
rect 9920 1337 10000 1463
rect 9920 1303 9943 1337
rect 9977 1303 10000 1337
rect 9920 1177 10000 1303
rect 9920 1143 9943 1177
rect 9977 1143 10000 1177
rect 9920 1017 10000 1143
rect 9920 983 9943 1017
rect 9977 983 10000 1017
rect 9920 857 10000 983
rect 9920 823 9943 857
rect 9977 823 10000 857
rect 9920 697 10000 823
rect 9920 663 9943 697
rect 9977 663 10000 697
rect 9920 537 10000 663
rect 9920 503 9943 537
rect 9977 503 10000 537
rect 9920 377 10000 503
rect 9920 343 9943 377
rect 9977 343 10000 377
rect 9920 217 10000 343
rect 9920 183 9943 217
rect 9977 183 10000 217
rect 9920 57 10000 183
rect 9920 23 9943 57
rect 9977 23 10000 57
rect 9920 0 10000 23
rect 10080 31426 10160 31440
rect 10080 31374 10094 31426
rect 10146 31374 10160 31426
rect 10080 31266 10160 31374
rect 10080 31214 10094 31266
rect 10146 31214 10160 31266
rect 10080 31106 10160 31214
rect 10080 31054 10094 31106
rect 10146 31054 10160 31106
rect 10080 30946 10160 31054
rect 10080 30894 10094 30946
rect 10146 30894 10160 30946
rect 10080 30786 10160 30894
rect 10080 30734 10094 30786
rect 10146 30734 10160 30786
rect 10080 30626 10160 30734
rect 10080 30574 10094 30626
rect 10146 30574 10160 30626
rect 10080 30466 10160 30574
rect 10080 30414 10094 30466
rect 10146 30414 10160 30466
rect 10080 30306 10160 30414
rect 10080 30254 10094 30306
rect 10146 30254 10160 30306
rect 10080 30137 10160 30254
rect 10080 30103 10103 30137
rect 10137 30103 10160 30137
rect 10080 29986 10160 30103
rect 10080 29934 10094 29986
rect 10146 29934 10160 29986
rect 10080 29826 10160 29934
rect 10080 29774 10094 29826
rect 10146 29774 10160 29826
rect 10080 29666 10160 29774
rect 10080 29614 10094 29666
rect 10146 29614 10160 29666
rect 10080 29506 10160 29614
rect 10080 29454 10094 29506
rect 10146 29454 10160 29506
rect 10080 29346 10160 29454
rect 10080 29294 10094 29346
rect 10146 29294 10160 29346
rect 10080 29186 10160 29294
rect 10080 29134 10094 29186
rect 10146 29134 10160 29186
rect 10080 29026 10160 29134
rect 10080 28974 10094 29026
rect 10146 28974 10160 29026
rect 10080 28866 10160 28974
rect 10080 28814 10094 28866
rect 10146 28814 10160 28866
rect 10080 28697 10160 28814
rect 10080 28663 10103 28697
rect 10137 28663 10160 28697
rect 10080 28537 10160 28663
rect 10080 28503 10103 28537
rect 10137 28503 10160 28537
rect 10080 28377 10160 28503
rect 10080 28343 10103 28377
rect 10137 28343 10160 28377
rect 10080 28217 10160 28343
rect 10080 28183 10103 28217
rect 10137 28183 10160 28217
rect 10080 28066 10160 28183
rect 10080 28014 10094 28066
rect 10146 28014 10160 28066
rect 10080 27906 10160 28014
rect 10080 27854 10094 27906
rect 10146 27854 10160 27906
rect 10080 27746 10160 27854
rect 10080 27694 10094 27746
rect 10146 27694 10160 27746
rect 10080 27586 10160 27694
rect 10080 27534 10094 27586
rect 10146 27534 10160 27586
rect 10080 27426 10160 27534
rect 10080 27374 10094 27426
rect 10146 27374 10160 27426
rect 10080 27266 10160 27374
rect 10080 27214 10094 27266
rect 10146 27214 10160 27266
rect 10080 27106 10160 27214
rect 10080 27054 10094 27106
rect 10146 27054 10160 27106
rect 10080 26946 10160 27054
rect 10080 26894 10094 26946
rect 10146 26894 10160 26946
rect 10080 26777 10160 26894
rect 10080 26743 10103 26777
rect 10137 26743 10160 26777
rect 10080 26617 10160 26743
rect 10080 26583 10103 26617
rect 10137 26583 10160 26617
rect 10080 26457 10160 26583
rect 10080 26423 10103 26457
rect 10137 26423 10160 26457
rect 10080 26297 10160 26423
rect 10080 26263 10103 26297
rect 10137 26263 10160 26297
rect 10080 26146 10160 26263
rect 10080 26094 10094 26146
rect 10146 26094 10160 26146
rect 10080 25986 10160 26094
rect 10080 25934 10094 25986
rect 10146 25934 10160 25986
rect 10080 25826 10160 25934
rect 10080 25774 10094 25826
rect 10146 25774 10160 25826
rect 10080 25666 10160 25774
rect 10080 25614 10094 25666
rect 10146 25614 10160 25666
rect 10080 25506 10160 25614
rect 10080 25454 10094 25506
rect 10146 25454 10160 25506
rect 10080 25346 10160 25454
rect 10080 25294 10094 25346
rect 10146 25294 10160 25346
rect 10080 25186 10160 25294
rect 10080 25134 10094 25186
rect 10146 25134 10160 25186
rect 10080 25026 10160 25134
rect 10080 24974 10094 25026
rect 10146 24974 10160 25026
rect 10080 24857 10160 24974
rect 10080 24823 10103 24857
rect 10137 24823 10160 24857
rect 10080 24706 10160 24823
rect 10080 24654 10094 24706
rect 10146 24654 10160 24706
rect 10080 24546 10160 24654
rect 10080 24494 10094 24546
rect 10146 24494 10160 24546
rect 10080 24386 10160 24494
rect 10080 24334 10094 24386
rect 10146 24334 10160 24386
rect 10080 24226 10160 24334
rect 10080 24174 10094 24226
rect 10146 24174 10160 24226
rect 10080 24066 10160 24174
rect 10080 24014 10094 24066
rect 10146 24014 10160 24066
rect 10080 23906 10160 24014
rect 10080 23854 10094 23906
rect 10146 23854 10160 23906
rect 10080 23746 10160 23854
rect 10080 23694 10094 23746
rect 10146 23694 10160 23746
rect 10080 23586 10160 23694
rect 10080 23534 10094 23586
rect 10146 23534 10160 23586
rect 10080 23426 10160 23534
rect 10080 23374 10094 23426
rect 10146 23374 10160 23426
rect 10080 23266 10160 23374
rect 10080 23214 10094 23266
rect 10146 23214 10160 23266
rect 10080 23106 10160 23214
rect 10080 23054 10094 23106
rect 10146 23054 10160 23106
rect 10080 22946 10160 23054
rect 10080 22894 10094 22946
rect 10146 22894 10160 22946
rect 10080 22786 10160 22894
rect 10080 22734 10094 22786
rect 10146 22734 10160 22786
rect 10080 22626 10160 22734
rect 10080 22574 10094 22626
rect 10146 22574 10160 22626
rect 10080 22466 10160 22574
rect 10080 22414 10094 22466
rect 10146 22414 10160 22466
rect 10080 22306 10160 22414
rect 10080 22254 10094 22306
rect 10146 22254 10160 22306
rect 10080 22146 10160 22254
rect 10080 22094 10094 22146
rect 10146 22094 10160 22146
rect 10080 21977 10160 22094
rect 10080 21943 10103 21977
rect 10137 21943 10160 21977
rect 10080 21826 10160 21943
rect 10080 21774 10094 21826
rect 10146 21774 10160 21826
rect 10080 21666 10160 21774
rect 10080 21614 10094 21666
rect 10146 21614 10160 21666
rect 10080 21506 10160 21614
rect 10080 21454 10094 21506
rect 10146 21454 10160 21506
rect 10080 21346 10160 21454
rect 10080 21294 10094 21346
rect 10146 21294 10160 21346
rect 10080 21186 10160 21294
rect 10080 21134 10094 21186
rect 10146 21134 10160 21186
rect 10080 21026 10160 21134
rect 10080 20974 10094 21026
rect 10146 20974 10160 21026
rect 10080 20866 10160 20974
rect 10080 20814 10094 20866
rect 10146 20814 10160 20866
rect 10080 20706 10160 20814
rect 10080 20654 10094 20706
rect 10146 20654 10160 20706
rect 10080 20537 10160 20654
rect 10080 20503 10103 20537
rect 10137 20503 10160 20537
rect 10080 20377 10160 20503
rect 10080 20343 10103 20377
rect 10137 20343 10160 20377
rect 10080 20217 10160 20343
rect 10080 20183 10103 20217
rect 10137 20183 10160 20217
rect 10080 20057 10160 20183
rect 10080 20023 10103 20057
rect 10137 20023 10160 20057
rect 10080 19906 10160 20023
rect 10080 19854 10094 19906
rect 10146 19854 10160 19906
rect 10080 19746 10160 19854
rect 10080 19694 10094 19746
rect 10146 19694 10160 19746
rect 10080 19586 10160 19694
rect 10080 19534 10094 19586
rect 10146 19534 10160 19586
rect 10080 19426 10160 19534
rect 10080 19374 10094 19426
rect 10146 19374 10160 19426
rect 10080 19266 10160 19374
rect 10080 19214 10094 19266
rect 10146 19214 10160 19266
rect 10080 19106 10160 19214
rect 10080 19054 10094 19106
rect 10146 19054 10160 19106
rect 10080 18946 10160 19054
rect 10080 18894 10094 18946
rect 10146 18894 10160 18946
rect 10080 18786 10160 18894
rect 10080 18734 10094 18786
rect 10146 18734 10160 18786
rect 10080 18617 10160 18734
rect 10080 18583 10103 18617
rect 10137 18583 10160 18617
rect 10080 18457 10160 18583
rect 10080 18423 10103 18457
rect 10137 18423 10160 18457
rect 10080 18297 10160 18423
rect 10080 18263 10103 18297
rect 10137 18263 10160 18297
rect 10080 18137 10160 18263
rect 10080 18103 10103 18137
rect 10137 18103 10160 18137
rect 10080 17986 10160 18103
rect 10080 17934 10094 17986
rect 10146 17934 10160 17986
rect 10080 17826 10160 17934
rect 10080 17774 10094 17826
rect 10146 17774 10160 17826
rect 10080 17666 10160 17774
rect 10080 17614 10094 17666
rect 10146 17614 10160 17666
rect 10080 17506 10160 17614
rect 10080 17454 10094 17506
rect 10146 17454 10160 17506
rect 10080 17346 10160 17454
rect 10080 17294 10094 17346
rect 10146 17294 10160 17346
rect 10080 17186 10160 17294
rect 10080 17134 10094 17186
rect 10146 17134 10160 17186
rect 10080 17026 10160 17134
rect 10080 16974 10094 17026
rect 10146 16974 10160 17026
rect 10080 16866 10160 16974
rect 10080 16814 10094 16866
rect 10146 16814 10160 16866
rect 10080 16697 10160 16814
rect 10080 16663 10103 16697
rect 10137 16663 10160 16697
rect 10080 16546 10160 16663
rect 10080 16494 10094 16546
rect 10146 16494 10160 16546
rect 10080 16386 10160 16494
rect 10080 16334 10094 16386
rect 10146 16334 10160 16386
rect 10080 16226 10160 16334
rect 10080 16174 10094 16226
rect 10146 16174 10160 16226
rect 10080 16066 10160 16174
rect 10080 16014 10094 16066
rect 10146 16014 10160 16066
rect 10080 15906 10160 16014
rect 10080 15854 10094 15906
rect 10146 15854 10160 15906
rect 10080 15746 10160 15854
rect 10080 15694 10094 15746
rect 10146 15694 10160 15746
rect 10080 15586 10160 15694
rect 10080 15534 10094 15586
rect 10146 15534 10160 15586
rect 10080 15426 10160 15534
rect 10080 15374 10094 15426
rect 10146 15374 10160 15426
rect 10080 15266 10160 15374
rect 10080 15214 10094 15266
rect 10146 15214 10160 15266
rect 10080 15106 10160 15214
rect 10080 15054 10094 15106
rect 10146 15054 10160 15106
rect 10080 14946 10160 15054
rect 10080 14894 10094 14946
rect 10146 14894 10160 14946
rect 10080 14786 10160 14894
rect 10080 14734 10094 14786
rect 10146 14734 10160 14786
rect 10080 14626 10160 14734
rect 10080 14574 10094 14626
rect 10146 14574 10160 14626
rect 10080 14466 10160 14574
rect 10080 14414 10094 14466
rect 10146 14414 10160 14466
rect 10080 14306 10160 14414
rect 10080 14254 10094 14306
rect 10146 14254 10160 14306
rect 10080 14146 10160 14254
rect 10080 14094 10094 14146
rect 10146 14094 10160 14146
rect 10080 13986 10160 14094
rect 10080 13934 10094 13986
rect 10146 13934 10160 13986
rect 10080 13817 10160 13934
rect 10080 13783 10103 13817
rect 10137 13783 10160 13817
rect 10080 13666 10160 13783
rect 10080 13614 10094 13666
rect 10146 13614 10160 13666
rect 10080 13506 10160 13614
rect 10080 13454 10094 13506
rect 10146 13454 10160 13506
rect 10080 13346 10160 13454
rect 10080 13294 10094 13346
rect 10146 13294 10160 13346
rect 10080 13186 10160 13294
rect 10080 13134 10094 13186
rect 10146 13134 10160 13186
rect 10080 13026 10160 13134
rect 10080 12974 10094 13026
rect 10146 12974 10160 13026
rect 10080 12866 10160 12974
rect 10080 12814 10094 12866
rect 10146 12814 10160 12866
rect 10080 12706 10160 12814
rect 10080 12654 10094 12706
rect 10146 12654 10160 12706
rect 10080 12546 10160 12654
rect 10080 12494 10094 12546
rect 10146 12494 10160 12546
rect 10080 12377 10160 12494
rect 10080 12343 10103 12377
rect 10137 12343 10160 12377
rect 10080 12217 10160 12343
rect 10080 12183 10103 12217
rect 10137 12183 10160 12217
rect 10080 12057 10160 12183
rect 10080 12023 10103 12057
rect 10137 12023 10160 12057
rect 10080 11897 10160 12023
rect 10080 11863 10103 11897
rect 10137 11863 10160 11897
rect 10080 11746 10160 11863
rect 10080 11694 10094 11746
rect 10146 11694 10160 11746
rect 10080 11586 10160 11694
rect 10080 11534 10094 11586
rect 10146 11534 10160 11586
rect 10080 11426 10160 11534
rect 10080 11374 10094 11426
rect 10146 11374 10160 11426
rect 10080 11266 10160 11374
rect 10080 11214 10094 11266
rect 10146 11214 10160 11266
rect 10080 11106 10160 11214
rect 10080 11054 10094 11106
rect 10146 11054 10160 11106
rect 10080 10946 10160 11054
rect 10080 10894 10094 10946
rect 10146 10894 10160 10946
rect 10080 10786 10160 10894
rect 10080 10734 10094 10786
rect 10146 10734 10160 10786
rect 10080 10626 10160 10734
rect 10080 10574 10094 10626
rect 10146 10574 10160 10626
rect 10080 10466 10160 10574
rect 10080 10414 10094 10466
rect 10146 10414 10160 10466
rect 10080 10306 10160 10414
rect 10080 10254 10094 10306
rect 10146 10254 10160 10306
rect 10080 10146 10160 10254
rect 10080 10094 10094 10146
rect 10146 10094 10160 10146
rect 10080 9986 10160 10094
rect 10080 9934 10094 9986
rect 10146 9934 10160 9986
rect 10080 9826 10160 9934
rect 10080 9774 10094 9826
rect 10146 9774 10160 9826
rect 10080 9657 10160 9774
rect 10080 9623 10103 9657
rect 10137 9623 10160 9657
rect 10080 9506 10160 9623
rect 10080 9454 10094 9506
rect 10146 9454 10160 9506
rect 10080 9346 10160 9454
rect 10080 9294 10094 9346
rect 10146 9294 10160 9346
rect 10080 9177 10160 9294
rect 10080 9143 10103 9177
rect 10137 9143 10160 9177
rect 10080 9026 10160 9143
rect 10080 8974 10094 9026
rect 10146 8974 10160 9026
rect 10080 8866 10160 8974
rect 10080 8814 10094 8866
rect 10146 8814 10160 8866
rect 10080 8706 10160 8814
rect 10080 8654 10094 8706
rect 10146 8654 10160 8706
rect 10080 8546 10160 8654
rect 10080 8494 10094 8546
rect 10146 8494 10160 8546
rect 10080 8386 10160 8494
rect 10080 8334 10094 8386
rect 10146 8334 10160 8386
rect 10080 8226 10160 8334
rect 10080 8174 10094 8226
rect 10146 8174 10160 8226
rect 10080 8066 10160 8174
rect 10080 8014 10094 8066
rect 10146 8014 10160 8066
rect 10080 7906 10160 8014
rect 10080 7854 10094 7906
rect 10146 7854 10160 7906
rect 10080 7746 10160 7854
rect 10080 7694 10094 7746
rect 10146 7694 10160 7746
rect 10080 7577 10160 7694
rect 10080 7543 10103 7577
rect 10137 7543 10160 7577
rect 10080 7426 10160 7543
rect 10080 7374 10094 7426
rect 10146 7374 10160 7426
rect 10080 7266 10160 7374
rect 10080 7214 10094 7266
rect 10146 7214 10160 7266
rect 10080 7097 10160 7214
rect 10080 7063 10103 7097
rect 10137 7063 10160 7097
rect 10080 6946 10160 7063
rect 10080 6894 10094 6946
rect 10146 6894 10160 6946
rect 10080 6786 10160 6894
rect 10080 6734 10094 6786
rect 10146 6734 10160 6786
rect 10080 6617 10160 6734
rect 10080 6583 10103 6617
rect 10137 6583 10160 6617
rect 10080 6466 10160 6583
rect 10080 6414 10094 6466
rect 10146 6414 10160 6466
rect 10080 6306 10160 6414
rect 10080 6254 10094 6306
rect 10146 6254 10160 6306
rect 10080 6146 10160 6254
rect 10080 6094 10094 6146
rect 10146 6094 10160 6146
rect 10080 5986 10160 6094
rect 10080 5934 10094 5986
rect 10146 5934 10160 5986
rect 10080 5826 10160 5934
rect 10080 5774 10094 5826
rect 10146 5774 10160 5826
rect 10080 5666 10160 5774
rect 10080 5614 10094 5666
rect 10146 5614 10160 5666
rect 10080 5506 10160 5614
rect 10080 5454 10094 5506
rect 10146 5454 10160 5506
rect 10080 5346 10160 5454
rect 10080 5294 10094 5346
rect 10146 5294 10160 5346
rect 10080 5186 10160 5294
rect 10080 5134 10094 5186
rect 10146 5134 10160 5186
rect 10080 5026 10160 5134
rect 10080 4974 10094 5026
rect 10146 4974 10160 5026
rect 10080 4866 10160 4974
rect 10080 4814 10094 4866
rect 10146 4814 10160 4866
rect 10080 4706 10160 4814
rect 10080 4654 10094 4706
rect 10146 4654 10160 4706
rect 10080 4546 10160 4654
rect 10080 4494 10094 4546
rect 10146 4494 10160 4546
rect 10080 4386 10160 4494
rect 10080 4334 10094 4386
rect 10146 4334 10160 4386
rect 10080 4226 10160 4334
rect 10080 4174 10094 4226
rect 10146 4174 10160 4226
rect 10080 4066 10160 4174
rect 10080 4014 10094 4066
rect 10146 4014 10160 4066
rect 10080 3906 10160 4014
rect 10080 3854 10094 3906
rect 10146 3854 10160 3906
rect 10080 3737 10160 3854
rect 10080 3703 10103 3737
rect 10137 3703 10160 3737
rect 10080 3577 10160 3703
rect 10080 3543 10103 3577
rect 10137 3543 10160 3577
rect 10080 3426 10160 3543
rect 10080 3374 10094 3426
rect 10146 3374 10160 3426
rect 10080 3266 10160 3374
rect 10080 3214 10094 3266
rect 10146 3214 10160 3266
rect 10080 3106 10160 3214
rect 10080 3054 10094 3106
rect 10146 3054 10160 3106
rect 10080 2946 10160 3054
rect 10080 2894 10094 2946
rect 10146 2894 10160 2946
rect 10080 2786 10160 2894
rect 10080 2734 10094 2786
rect 10146 2734 10160 2786
rect 10080 2626 10160 2734
rect 10080 2574 10094 2626
rect 10146 2574 10160 2626
rect 10080 2466 10160 2574
rect 10080 2414 10094 2466
rect 10146 2414 10160 2466
rect 10080 2306 10160 2414
rect 10080 2254 10094 2306
rect 10146 2254 10160 2306
rect 10080 2146 10160 2254
rect 10080 2094 10094 2146
rect 10146 2094 10160 2146
rect 10080 1986 10160 2094
rect 10080 1934 10094 1986
rect 10146 1934 10160 1986
rect 10080 1817 10160 1934
rect 10080 1783 10103 1817
rect 10137 1783 10160 1817
rect 10080 1666 10160 1783
rect 10080 1614 10094 1666
rect 10146 1614 10160 1666
rect 10080 1506 10160 1614
rect 10080 1454 10094 1506
rect 10146 1454 10160 1506
rect 10080 1346 10160 1454
rect 10080 1294 10094 1346
rect 10146 1294 10160 1346
rect 10080 1186 10160 1294
rect 10080 1134 10094 1186
rect 10146 1134 10160 1186
rect 10080 1026 10160 1134
rect 10080 974 10094 1026
rect 10146 974 10160 1026
rect 10080 857 10160 974
rect 10080 823 10103 857
rect 10137 823 10160 857
rect 10080 697 10160 823
rect 10080 663 10103 697
rect 10137 663 10160 697
rect 10080 546 10160 663
rect 10080 494 10094 546
rect 10146 494 10160 546
rect 10080 386 10160 494
rect 10080 334 10094 386
rect 10146 334 10160 386
rect 10080 226 10160 334
rect 10080 174 10094 226
rect 10146 174 10160 226
rect 10080 66 10160 174
rect 10080 14 10094 66
rect 10146 14 10160 66
rect 10080 0 10160 14
rect 10240 31417 10320 31440
rect 10240 31383 10263 31417
rect 10297 31383 10320 31417
rect 10240 31257 10320 31383
rect 10240 31223 10263 31257
rect 10297 31223 10320 31257
rect 10240 31097 10320 31223
rect 10240 31063 10263 31097
rect 10297 31063 10320 31097
rect 10240 30937 10320 31063
rect 10240 30903 10263 30937
rect 10297 30903 10320 30937
rect 10240 30777 10320 30903
rect 10240 30743 10263 30777
rect 10297 30743 10320 30777
rect 10240 30617 10320 30743
rect 10240 30583 10263 30617
rect 10297 30583 10320 30617
rect 10240 30457 10320 30583
rect 10240 30423 10263 30457
rect 10297 30423 10320 30457
rect 10240 30297 10320 30423
rect 10240 30263 10263 30297
rect 10297 30263 10320 30297
rect 10240 30137 10320 30263
rect 10240 30103 10263 30137
rect 10297 30103 10320 30137
rect 10240 29977 10320 30103
rect 10240 29943 10263 29977
rect 10297 29943 10320 29977
rect 10240 29817 10320 29943
rect 10240 29783 10263 29817
rect 10297 29783 10320 29817
rect 10240 29657 10320 29783
rect 10240 29623 10263 29657
rect 10297 29623 10320 29657
rect 10240 29497 10320 29623
rect 10240 29463 10263 29497
rect 10297 29463 10320 29497
rect 10240 29337 10320 29463
rect 10240 29303 10263 29337
rect 10297 29303 10320 29337
rect 10240 29177 10320 29303
rect 10240 29143 10263 29177
rect 10297 29143 10320 29177
rect 10240 29017 10320 29143
rect 10240 28983 10263 29017
rect 10297 28983 10320 29017
rect 10240 28857 10320 28983
rect 10240 28823 10263 28857
rect 10297 28823 10320 28857
rect 10240 28697 10320 28823
rect 10240 28663 10263 28697
rect 10297 28663 10320 28697
rect 10240 28537 10320 28663
rect 10240 28503 10263 28537
rect 10297 28503 10320 28537
rect 10240 28377 10320 28503
rect 10240 28343 10263 28377
rect 10297 28343 10320 28377
rect 10240 28217 10320 28343
rect 10240 28183 10263 28217
rect 10297 28183 10320 28217
rect 10240 28057 10320 28183
rect 10240 28023 10263 28057
rect 10297 28023 10320 28057
rect 10240 27897 10320 28023
rect 10240 27863 10263 27897
rect 10297 27863 10320 27897
rect 10240 27737 10320 27863
rect 10240 27703 10263 27737
rect 10297 27703 10320 27737
rect 10240 27577 10320 27703
rect 10240 27543 10263 27577
rect 10297 27543 10320 27577
rect 10240 27417 10320 27543
rect 10240 27383 10263 27417
rect 10297 27383 10320 27417
rect 10240 27257 10320 27383
rect 10240 27223 10263 27257
rect 10297 27223 10320 27257
rect 10240 27097 10320 27223
rect 10240 27063 10263 27097
rect 10297 27063 10320 27097
rect 10240 26937 10320 27063
rect 10240 26903 10263 26937
rect 10297 26903 10320 26937
rect 10240 26777 10320 26903
rect 10240 26743 10263 26777
rect 10297 26743 10320 26777
rect 10240 26617 10320 26743
rect 10240 26583 10263 26617
rect 10297 26583 10320 26617
rect 10240 26457 10320 26583
rect 10240 26423 10263 26457
rect 10297 26423 10320 26457
rect 10240 26297 10320 26423
rect 10240 26263 10263 26297
rect 10297 26263 10320 26297
rect 10240 26137 10320 26263
rect 10240 26103 10263 26137
rect 10297 26103 10320 26137
rect 10240 25977 10320 26103
rect 10240 25943 10263 25977
rect 10297 25943 10320 25977
rect 10240 25817 10320 25943
rect 10240 25783 10263 25817
rect 10297 25783 10320 25817
rect 10240 25657 10320 25783
rect 10240 25623 10263 25657
rect 10297 25623 10320 25657
rect 10240 25497 10320 25623
rect 10240 25463 10263 25497
rect 10297 25463 10320 25497
rect 10240 25337 10320 25463
rect 10240 25303 10263 25337
rect 10297 25303 10320 25337
rect 10240 25177 10320 25303
rect 10240 25143 10263 25177
rect 10297 25143 10320 25177
rect 10240 25017 10320 25143
rect 10240 24983 10263 25017
rect 10297 24983 10320 25017
rect 10240 24857 10320 24983
rect 10240 24823 10263 24857
rect 10297 24823 10320 24857
rect 10240 24697 10320 24823
rect 10240 24663 10263 24697
rect 10297 24663 10320 24697
rect 10240 24537 10320 24663
rect 10240 24503 10263 24537
rect 10297 24503 10320 24537
rect 10240 24377 10320 24503
rect 10240 24343 10263 24377
rect 10297 24343 10320 24377
rect 10240 24217 10320 24343
rect 10240 24183 10263 24217
rect 10297 24183 10320 24217
rect 10240 24057 10320 24183
rect 10240 24023 10263 24057
rect 10297 24023 10320 24057
rect 10240 23897 10320 24023
rect 10240 23863 10263 23897
rect 10297 23863 10320 23897
rect 10240 23737 10320 23863
rect 10240 23703 10263 23737
rect 10297 23703 10320 23737
rect 10240 23577 10320 23703
rect 10240 23543 10263 23577
rect 10297 23543 10320 23577
rect 10240 23417 10320 23543
rect 10240 23383 10263 23417
rect 10297 23383 10320 23417
rect 10240 23257 10320 23383
rect 10240 23223 10263 23257
rect 10297 23223 10320 23257
rect 10240 23097 10320 23223
rect 10240 23063 10263 23097
rect 10297 23063 10320 23097
rect 10240 22937 10320 23063
rect 10240 22903 10263 22937
rect 10297 22903 10320 22937
rect 10240 22777 10320 22903
rect 10240 22743 10263 22777
rect 10297 22743 10320 22777
rect 10240 22617 10320 22743
rect 10240 22583 10263 22617
rect 10297 22583 10320 22617
rect 10240 22457 10320 22583
rect 10240 22423 10263 22457
rect 10297 22423 10320 22457
rect 10240 22297 10320 22423
rect 10240 22263 10263 22297
rect 10297 22263 10320 22297
rect 10240 22137 10320 22263
rect 10240 22103 10263 22137
rect 10297 22103 10320 22137
rect 10240 21977 10320 22103
rect 10240 21943 10263 21977
rect 10297 21943 10320 21977
rect 10240 21817 10320 21943
rect 10240 21783 10263 21817
rect 10297 21783 10320 21817
rect 10240 21657 10320 21783
rect 10240 21623 10263 21657
rect 10297 21623 10320 21657
rect 10240 21497 10320 21623
rect 10240 21463 10263 21497
rect 10297 21463 10320 21497
rect 10240 21337 10320 21463
rect 10240 21303 10263 21337
rect 10297 21303 10320 21337
rect 10240 21177 10320 21303
rect 10240 21143 10263 21177
rect 10297 21143 10320 21177
rect 10240 21017 10320 21143
rect 10240 20983 10263 21017
rect 10297 20983 10320 21017
rect 10240 20857 10320 20983
rect 10240 20823 10263 20857
rect 10297 20823 10320 20857
rect 10240 20697 10320 20823
rect 10240 20663 10263 20697
rect 10297 20663 10320 20697
rect 10240 20537 10320 20663
rect 10240 20503 10263 20537
rect 10297 20503 10320 20537
rect 10240 20377 10320 20503
rect 10240 20343 10263 20377
rect 10297 20343 10320 20377
rect 10240 20217 10320 20343
rect 10240 20183 10263 20217
rect 10297 20183 10320 20217
rect 10240 20057 10320 20183
rect 10240 20023 10263 20057
rect 10297 20023 10320 20057
rect 10240 19897 10320 20023
rect 10240 19863 10263 19897
rect 10297 19863 10320 19897
rect 10240 19737 10320 19863
rect 10240 19703 10263 19737
rect 10297 19703 10320 19737
rect 10240 19577 10320 19703
rect 10240 19543 10263 19577
rect 10297 19543 10320 19577
rect 10240 19417 10320 19543
rect 10240 19383 10263 19417
rect 10297 19383 10320 19417
rect 10240 19257 10320 19383
rect 10240 19223 10263 19257
rect 10297 19223 10320 19257
rect 10240 19097 10320 19223
rect 10240 19063 10263 19097
rect 10297 19063 10320 19097
rect 10240 18937 10320 19063
rect 10240 18903 10263 18937
rect 10297 18903 10320 18937
rect 10240 18777 10320 18903
rect 10240 18743 10263 18777
rect 10297 18743 10320 18777
rect 10240 18617 10320 18743
rect 10240 18583 10263 18617
rect 10297 18583 10320 18617
rect 10240 18457 10320 18583
rect 10240 18423 10263 18457
rect 10297 18423 10320 18457
rect 10240 18297 10320 18423
rect 10240 18263 10263 18297
rect 10297 18263 10320 18297
rect 10240 18137 10320 18263
rect 10240 18103 10263 18137
rect 10297 18103 10320 18137
rect 10240 17977 10320 18103
rect 10240 17943 10263 17977
rect 10297 17943 10320 17977
rect 10240 17817 10320 17943
rect 10240 17783 10263 17817
rect 10297 17783 10320 17817
rect 10240 17657 10320 17783
rect 10240 17623 10263 17657
rect 10297 17623 10320 17657
rect 10240 17497 10320 17623
rect 10240 17463 10263 17497
rect 10297 17463 10320 17497
rect 10240 17337 10320 17463
rect 10240 17303 10263 17337
rect 10297 17303 10320 17337
rect 10240 17177 10320 17303
rect 10240 17143 10263 17177
rect 10297 17143 10320 17177
rect 10240 17017 10320 17143
rect 10240 16983 10263 17017
rect 10297 16983 10320 17017
rect 10240 16857 10320 16983
rect 10240 16823 10263 16857
rect 10297 16823 10320 16857
rect 10240 16697 10320 16823
rect 10240 16663 10263 16697
rect 10297 16663 10320 16697
rect 10240 16537 10320 16663
rect 10240 16503 10263 16537
rect 10297 16503 10320 16537
rect 10240 16377 10320 16503
rect 10240 16343 10263 16377
rect 10297 16343 10320 16377
rect 10240 16217 10320 16343
rect 10240 16183 10263 16217
rect 10297 16183 10320 16217
rect 10240 16057 10320 16183
rect 10240 16023 10263 16057
rect 10297 16023 10320 16057
rect 10240 15897 10320 16023
rect 10240 15863 10263 15897
rect 10297 15863 10320 15897
rect 10240 15737 10320 15863
rect 10240 15703 10263 15737
rect 10297 15703 10320 15737
rect 10240 15577 10320 15703
rect 10240 15543 10263 15577
rect 10297 15543 10320 15577
rect 10240 15417 10320 15543
rect 10240 15383 10263 15417
rect 10297 15383 10320 15417
rect 10240 15257 10320 15383
rect 10240 15223 10263 15257
rect 10297 15223 10320 15257
rect 10240 15097 10320 15223
rect 10240 15063 10263 15097
rect 10297 15063 10320 15097
rect 10240 14937 10320 15063
rect 10240 14903 10263 14937
rect 10297 14903 10320 14937
rect 10240 14777 10320 14903
rect 10240 14743 10263 14777
rect 10297 14743 10320 14777
rect 10240 14617 10320 14743
rect 10240 14583 10263 14617
rect 10297 14583 10320 14617
rect 10240 14457 10320 14583
rect 10240 14423 10263 14457
rect 10297 14423 10320 14457
rect 10240 14297 10320 14423
rect 10240 14263 10263 14297
rect 10297 14263 10320 14297
rect 10240 14137 10320 14263
rect 10240 14103 10263 14137
rect 10297 14103 10320 14137
rect 10240 13977 10320 14103
rect 10240 13943 10263 13977
rect 10297 13943 10320 13977
rect 10240 13817 10320 13943
rect 10240 13783 10263 13817
rect 10297 13783 10320 13817
rect 10240 13657 10320 13783
rect 10240 13623 10263 13657
rect 10297 13623 10320 13657
rect 10240 13497 10320 13623
rect 10240 13463 10263 13497
rect 10297 13463 10320 13497
rect 10240 13337 10320 13463
rect 10240 13303 10263 13337
rect 10297 13303 10320 13337
rect 10240 13177 10320 13303
rect 10240 13143 10263 13177
rect 10297 13143 10320 13177
rect 10240 13017 10320 13143
rect 10240 12983 10263 13017
rect 10297 12983 10320 13017
rect 10240 12857 10320 12983
rect 10240 12823 10263 12857
rect 10297 12823 10320 12857
rect 10240 12697 10320 12823
rect 10240 12663 10263 12697
rect 10297 12663 10320 12697
rect 10240 12537 10320 12663
rect 10240 12503 10263 12537
rect 10297 12503 10320 12537
rect 10240 12377 10320 12503
rect 10240 12343 10263 12377
rect 10297 12343 10320 12377
rect 10240 12217 10320 12343
rect 10240 12183 10263 12217
rect 10297 12183 10320 12217
rect 10240 12057 10320 12183
rect 10240 12023 10263 12057
rect 10297 12023 10320 12057
rect 10240 11897 10320 12023
rect 10240 11863 10263 11897
rect 10297 11863 10320 11897
rect 10240 11737 10320 11863
rect 10240 11703 10263 11737
rect 10297 11703 10320 11737
rect 10240 11577 10320 11703
rect 10240 11543 10263 11577
rect 10297 11543 10320 11577
rect 10240 11417 10320 11543
rect 10240 11383 10263 11417
rect 10297 11383 10320 11417
rect 10240 11257 10320 11383
rect 10240 11223 10263 11257
rect 10297 11223 10320 11257
rect 10240 11097 10320 11223
rect 10240 11063 10263 11097
rect 10297 11063 10320 11097
rect 10240 10937 10320 11063
rect 10240 10903 10263 10937
rect 10297 10903 10320 10937
rect 10240 10777 10320 10903
rect 10240 10743 10263 10777
rect 10297 10743 10320 10777
rect 10240 10617 10320 10743
rect 10240 10583 10263 10617
rect 10297 10583 10320 10617
rect 10240 10457 10320 10583
rect 10240 10423 10263 10457
rect 10297 10423 10320 10457
rect 10240 10297 10320 10423
rect 10240 10263 10263 10297
rect 10297 10263 10320 10297
rect 10240 10137 10320 10263
rect 10240 10103 10263 10137
rect 10297 10103 10320 10137
rect 10240 9977 10320 10103
rect 10240 9943 10263 9977
rect 10297 9943 10320 9977
rect 10240 9817 10320 9943
rect 10240 9783 10263 9817
rect 10297 9783 10320 9817
rect 10240 9657 10320 9783
rect 10240 9623 10263 9657
rect 10297 9623 10320 9657
rect 10240 9497 10320 9623
rect 10240 9463 10263 9497
rect 10297 9463 10320 9497
rect 10240 9337 10320 9463
rect 10240 9303 10263 9337
rect 10297 9303 10320 9337
rect 10240 9177 10320 9303
rect 10240 9143 10263 9177
rect 10297 9143 10320 9177
rect 10240 9017 10320 9143
rect 10240 8983 10263 9017
rect 10297 8983 10320 9017
rect 10240 8857 10320 8983
rect 10240 8823 10263 8857
rect 10297 8823 10320 8857
rect 10240 8697 10320 8823
rect 10240 8663 10263 8697
rect 10297 8663 10320 8697
rect 10240 8537 10320 8663
rect 10240 8503 10263 8537
rect 10297 8503 10320 8537
rect 10240 8377 10320 8503
rect 10240 8343 10263 8377
rect 10297 8343 10320 8377
rect 10240 8217 10320 8343
rect 10240 8183 10263 8217
rect 10297 8183 10320 8217
rect 10240 8057 10320 8183
rect 10240 8023 10263 8057
rect 10297 8023 10320 8057
rect 10240 7897 10320 8023
rect 10240 7863 10263 7897
rect 10297 7863 10320 7897
rect 10240 7737 10320 7863
rect 10240 7703 10263 7737
rect 10297 7703 10320 7737
rect 10240 7577 10320 7703
rect 10240 7543 10263 7577
rect 10297 7543 10320 7577
rect 10240 7417 10320 7543
rect 10240 7383 10263 7417
rect 10297 7383 10320 7417
rect 10240 7257 10320 7383
rect 10240 7223 10263 7257
rect 10297 7223 10320 7257
rect 10240 7097 10320 7223
rect 10240 7063 10263 7097
rect 10297 7063 10320 7097
rect 10240 6937 10320 7063
rect 10240 6903 10263 6937
rect 10297 6903 10320 6937
rect 10240 6777 10320 6903
rect 10240 6743 10263 6777
rect 10297 6743 10320 6777
rect 10240 6617 10320 6743
rect 10240 6583 10263 6617
rect 10297 6583 10320 6617
rect 10240 6457 10320 6583
rect 10240 6423 10263 6457
rect 10297 6423 10320 6457
rect 10240 6297 10320 6423
rect 10240 6263 10263 6297
rect 10297 6263 10320 6297
rect 10240 6137 10320 6263
rect 10240 6103 10263 6137
rect 10297 6103 10320 6137
rect 10240 5977 10320 6103
rect 10240 5943 10263 5977
rect 10297 5943 10320 5977
rect 10240 5817 10320 5943
rect 10240 5783 10263 5817
rect 10297 5783 10320 5817
rect 10240 5657 10320 5783
rect 10240 5623 10263 5657
rect 10297 5623 10320 5657
rect 10240 5497 10320 5623
rect 10240 5463 10263 5497
rect 10297 5463 10320 5497
rect 10240 5337 10320 5463
rect 10240 5303 10263 5337
rect 10297 5303 10320 5337
rect 10240 5177 10320 5303
rect 10240 5143 10263 5177
rect 10297 5143 10320 5177
rect 10240 5017 10320 5143
rect 10240 4983 10263 5017
rect 10297 4983 10320 5017
rect 10240 4857 10320 4983
rect 10240 4823 10263 4857
rect 10297 4823 10320 4857
rect 10240 4697 10320 4823
rect 10240 4663 10263 4697
rect 10297 4663 10320 4697
rect 10240 4537 10320 4663
rect 10240 4503 10263 4537
rect 10297 4503 10320 4537
rect 10240 4377 10320 4503
rect 10240 4343 10263 4377
rect 10297 4343 10320 4377
rect 10240 4217 10320 4343
rect 10240 4183 10263 4217
rect 10297 4183 10320 4217
rect 10240 4057 10320 4183
rect 10240 4023 10263 4057
rect 10297 4023 10320 4057
rect 10240 3897 10320 4023
rect 10240 3863 10263 3897
rect 10297 3863 10320 3897
rect 10240 3737 10320 3863
rect 10240 3703 10263 3737
rect 10297 3703 10320 3737
rect 10240 3577 10320 3703
rect 10240 3543 10263 3577
rect 10297 3543 10320 3577
rect 10240 3417 10320 3543
rect 10240 3383 10263 3417
rect 10297 3383 10320 3417
rect 10240 3257 10320 3383
rect 10240 3223 10263 3257
rect 10297 3223 10320 3257
rect 10240 3097 10320 3223
rect 10240 3063 10263 3097
rect 10297 3063 10320 3097
rect 10240 2937 10320 3063
rect 10240 2903 10263 2937
rect 10297 2903 10320 2937
rect 10240 2777 10320 2903
rect 10240 2743 10263 2777
rect 10297 2743 10320 2777
rect 10240 2617 10320 2743
rect 10240 2583 10263 2617
rect 10297 2583 10320 2617
rect 10240 2457 10320 2583
rect 10240 2423 10263 2457
rect 10297 2423 10320 2457
rect 10240 2297 10320 2423
rect 10240 2263 10263 2297
rect 10297 2263 10320 2297
rect 10240 2137 10320 2263
rect 10240 2103 10263 2137
rect 10297 2103 10320 2137
rect 10240 1977 10320 2103
rect 10240 1943 10263 1977
rect 10297 1943 10320 1977
rect 10240 1817 10320 1943
rect 10240 1783 10263 1817
rect 10297 1783 10320 1817
rect 10240 1657 10320 1783
rect 10240 1623 10263 1657
rect 10297 1623 10320 1657
rect 10240 1497 10320 1623
rect 10240 1463 10263 1497
rect 10297 1463 10320 1497
rect 10240 1337 10320 1463
rect 10240 1303 10263 1337
rect 10297 1303 10320 1337
rect 10240 1177 10320 1303
rect 10240 1143 10263 1177
rect 10297 1143 10320 1177
rect 10240 1017 10320 1143
rect 10240 983 10263 1017
rect 10297 983 10320 1017
rect 10240 857 10320 983
rect 10240 823 10263 857
rect 10297 823 10320 857
rect 10240 697 10320 823
rect 10240 663 10263 697
rect 10297 663 10320 697
rect 10240 537 10320 663
rect 10240 503 10263 537
rect 10297 503 10320 537
rect 10240 377 10320 503
rect 10240 343 10263 377
rect 10297 343 10320 377
rect 10240 217 10320 343
rect 10240 183 10263 217
rect 10297 183 10320 217
rect 10240 57 10320 183
rect 10240 23 10263 57
rect 10297 23 10320 57
rect 10240 0 10320 23
rect 10400 31426 10480 31440
rect 10400 31374 10414 31426
rect 10466 31374 10480 31426
rect 10400 31266 10480 31374
rect 10400 31214 10414 31266
rect 10466 31214 10480 31266
rect 10400 31106 10480 31214
rect 10400 31054 10414 31106
rect 10466 31054 10480 31106
rect 10400 30946 10480 31054
rect 10400 30894 10414 30946
rect 10466 30894 10480 30946
rect 10400 30786 10480 30894
rect 10400 30734 10414 30786
rect 10466 30734 10480 30786
rect 10400 30626 10480 30734
rect 10400 30574 10414 30626
rect 10466 30574 10480 30626
rect 10400 30466 10480 30574
rect 10400 30414 10414 30466
rect 10466 30414 10480 30466
rect 10400 30306 10480 30414
rect 10400 30254 10414 30306
rect 10466 30254 10480 30306
rect 10400 30137 10480 30254
rect 10400 30103 10423 30137
rect 10457 30103 10480 30137
rect 10400 29986 10480 30103
rect 10400 29934 10414 29986
rect 10466 29934 10480 29986
rect 10400 29826 10480 29934
rect 10400 29774 10414 29826
rect 10466 29774 10480 29826
rect 10400 29666 10480 29774
rect 10400 29614 10414 29666
rect 10466 29614 10480 29666
rect 10400 29506 10480 29614
rect 10400 29454 10414 29506
rect 10466 29454 10480 29506
rect 10400 29346 10480 29454
rect 10400 29294 10414 29346
rect 10466 29294 10480 29346
rect 10400 29186 10480 29294
rect 10400 29134 10414 29186
rect 10466 29134 10480 29186
rect 10400 29026 10480 29134
rect 10400 28974 10414 29026
rect 10466 28974 10480 29026
rect 10400 28866 10480 28974
rect 10400 28814 10414 28866
rect 10466 28814 10480 28866
rect 10400 28697 10480 28814
rect 10400 28663 10423 28697
rect 10457 28663 10480 28697
rect 10400 28537 10480 28663
rect 10400 28503 10423 28537
rect 10457 28503 10480 28537
rect 10400 28377 10480 28503
rect 10400 28343 10423 28377
rect 10457 28343 10480 28377
rect 10400 28217 10480 28343
rect 10400 28183 10423 28217
rect 10457 28183 10480 28217
rect 10400 28066 10480 28183
rect 10400 28014 10414 28066
rect 10466 28014 10480 28066
rect 10400 27906 10480 28014
rect 10400 27854 10414 27906
rect 10466 27854 10480 27906
rect 10400 27746 10480 27854
rect 10400 27694 10414 27746
rect 10466 27694 10480 27746
rect 10400 27586 10480 27694
rect 10400 27534 10414 27586
rect 10466 27534 10480 27586
rect 10400 27426 10480 27534
rect 10400 27374 10414 27426
rect 10466 27374 10480 27426
rect 10400 27266 10480 27374
rect 10400 27214 10414 27266
rect 10466 27214 10480 27266
rect 10400 27106 10480 27214
rect 10400 27054 10414 27106
rect 10466 27054 10480 27106
rect 10400 26946 10480 27054
rect 10400 26894 10414 26946
rect 10466 26894 10480 26946
rect 10400 26777 10480 26894
rect 10400 26743 10423 26777
rect 10457 26743 10480 26777
rect 10400 26617 10480 26743
rect 10400 26583 10423 26617
rect 10457 26583 10480 26617
rect 10400 26457 10480 26583
rect 10400 26423 10423 26457
rect 10457 26423 10480 26457
rect 10400 26297 10480 26423
rect 10400 26263 10423 26297
rect 10457 26263 10480 26297
rect 10400 26146 10480 26263
rect 10400 26094 10414 26146
rect 10466 26094 10480 26146
rect 10400 25986 10480 26094
rect 10400 25934 10414 25986
rect 10466 25934 10480 25986
rect 10400 25826 10480 25934
rect 10400 25774 10414 25826
rect 10466 25774 10480 25826
rect 10400 25666 10480 25774
rect 10400 25614 10414 25666
rect 10466 25614 10480 25666
rect 10400 25506 10480 25614
rect 10400 25454 10414 25506
rect 10466 25454 10480 25506
rect 10400 25346 10480 25454
rect 10400 25294 10414 25346
rect 10466 25294 10480 25346
rect 10400 25186 10480 25294
rect 10400 25134 10414 25186
rect 10466 25134 10480 25186
rect 10400 25026 10480 25134
rect 10400 24974 10414 25026
rect 10466 24974 10480 25026
rect 10400 24857 10480 24974
rect 10400 24823 10423 24857
rect 10457 24823 10480 24857
rect 10400 24706 10480 24823
rect 10400 24654 10414 24706
rect 10466 24654 10480 24706
rect 10400 24546 10480 24654
rect 10400 24494 10414 24546
rect 10466 24494 10480 24546
rect 10400 24386 10480 24494
rect 10400 24334 10414 24386
rect 10466 24334 10480 24386
rect 10400 24226 10480 24334
rect 10400 24174 10414 24226
rect 10466 24174 10480 24226
rect 10400 24066 10480 24174
rect 10400 24014 10414 24066
rect 10466 24014 10480 24066
rect 10400 23906 10480 24014
rect 10400 23854 10414 23906
rect 10466 23854 10480 23906
rect 10400 23746 10480 23854
rect 10400 23694 10414 23746
rect 10466 23694 10480 23746
rect 10400 23586 10480 23694
rect 10400 23534 10414 23586
rect 10466 23534 10480 23586
rect 10400 23426 10480 23534
rect 10400 23374 10414 23426
rect 10466 23374 10480 23426
rect 10400 23266 10480 23374
rect 10400 23214 10414 23266
rect 10466 23214 10480 23266
rect 10400 23106 10480 23214
rect 10400 23054 10414 23106
rect 10466 23054 10480 23106
rect 10400 22946 10480 23054
rect 10400 22894 10414 22946
rect 10466 22894 10480 22946
rect 10400 22786 10480 22894
rect 10400 22734 10414 22786
rect 10466 22734 10480 22786
rect 10400 22626 10480 22734
rect 10400 22574 10414 22626
rect 10466 22574 10480 22626
rect 10400 22466 10480 22574
rect 10400 22414 10414 22466
rect 10466 22414 10480 22466
rect 10400 22306 10480 22414
rect 10400 22254 10414 22306
rect 10466 22254 10480 22306
rect 10400 22146 10480 22254
rect 10400 22094 10414 22146
rect 10466 22094 10480 22146
rect 10400 21977 10480 22094
rect 10400 21943 10423 21977
rect 10457 21943 10480 21977
rect 10400 21826 10480 21943
rect 10400 21774 10414 21826
rect 10466 21774 10480 21826
rect 10400 21666 10480 21774
rect 10400 21614 10414 21666
rect 10466 21614 10480 21666
rect 10400 21506 10480 21614
rect 10400 21454 10414 21506
rect 10466 21454 10480 21506
rect 10400 21346 10480 21454
rect 10400 21294 10414 21346
rect 10466 21294 10480 21346
rect 10400 21186 10480 21294
rect 10400 21134 10414 21186
rect 10466 21134 10480 21186
rect 10400 21026 10480 21134
rect 10400 20974 10414 21026
rect 10466 20974 10480 21026
rect 10400 20866 10480 20974
rect 10400 20814 10414 20866
rect 10466 20814 10480 20866
rect 10400 20706 10480 20814
rect 10400 20654 10414 20706
rect 10466 20654 10480 20706
rect 10400 20537 10480 20654
rect 10400 20503 10423 20537
rect 10457 20503 10480 20537
rect 10400 20377 10480 20503
rect 10400 20343 10423 20377
rect 10457 20343 10480 20377
rect 10400 20217 10480 20343
rect 10400 20183 10423 20217
rect 10457 20183 10480 20217
rect 10400 20057 10480 20183
rect 10400 20023 10423 20057
rect 10457 20023 10480 20057
rect 10400 19906 10480 20023
rect 10400 19854 10414 19906
rect 10466 19854 10480 19906
rect 10400 19746 10480 19854
rect 10400 19694 10414 19746
rect 10466 19694 10480 19746
rect 10400 19586 10480 19694
rect 10400 19534 10414 19586
rect 10466 19534 10480 19586
rect 10400 19426 10480 19534
rect 10400 19374 10414 19426
rect 10466 19374 10480 19426
rect 10400 19266 10480 19374
rect 10400 19214 10414 19266
rect 10466 19214 10480 19266
rect 10400 19106 10480 19214
rect 10400 19054 10414 19106
rect 10466 19054 10480 19106
rect 10400 18946 10480 19054
rect 10400 18894 10414 18946
rect 10466 18894 10480 18946
rect 10400 18786 10480 18894
rect 10400 18734 10414 18786
rect 10466 18734 10480 18786
rect 10400 18617 10480 18734
rect 10400 18583 10423 18617
rect 10457 18583 10480 18617
rect 10400 18457 10480 18583
rect 10400 18423 10423 18457
rect 10457 18423 10480 18457
rect 10400 18297 10480 18423
rect 10400 18263 10423 18297
rect 10457 18263 10480 18297
rect 10400 18137 10480 18263
rect 10400 18103 10423 18137
rect 10457 18103 10480 18137
rect 10400 17986 10480 18103
rect 10400 17934 10414 17986
rect 10466 17934 10480 17986
rect 10400 17826 10480 17934
rect 10400 17774 10414 17826
rect 10466 17774 10480 17826
rect 10400 17666 10480 17774
rect 10400 17614 10414 17666
rect 10466 17614 10480 17666
rect 10400 17506 10480 17614
rect 10400 17454 10414 17506
rect 10466 17454 10480 17506
rect 10400 17346 10480 17454
rect 10400 17294 10414 17346
rect 10466 17294 10480 17346
rect 10400 17186 10480 17294
rect 10400 17134 10414 17186
rect 10466 17134 10480 17186
rect 10400 17026 10480 17134
rect 10400 16974 10414 17026
rect 10466 16974 10480 17026
rect 10400 16866 10480 16974
rect 10400 16814 10414 16866
rect 10466 16814 10480 16866
rect 10400 16697 10480 16814
rect 10400 16663 10423 16697
rect 10457 16663 10480 16697
rect 10400 16546 10480 16663
rect 10400 16494 10414 16546
rect 10466 16494 10480 16546
rect 10400 16386 10480 16494
rect 10400 16334 10414 16386
rect 10466 16334 10480 16386
rect 10400 16226 10480 16334
rect 10400 16174 10414 16226
rect 10466 16174 10480 16226
rect 10400 16066 10480 16174
rect 10400 16014 10414 16066
rect 10466 16014 10480 16066
rect 10400 15906 10480 16014
rect 10400 15854 10414 15906
rect 10466 15854 10480 15906
rect 10400 15746 10480 15854
rect 10400 15694 10414 15746
rect 10466 15694 10480 15746
rect 10400 15586 10480 15694
rect 10400 15534 10414 15586
rect 10466 15534 10480 15586
rect 10400 15426 10480 15534
rect 10400 15374 10414 15426
rect 10466 15374 10480 15426
rect 10400 15266 10480 15374
rect 10400 15214 10414 15266
rect 10466 15214 10480 15266
rect 10400 15106 10480 15214
rect 10400 15054 10414 15106
rect 10466 15054 10480 15106
rect 10400 14946 10480 15054
rect 10400 14894 10414 14946
rect 10466 14894 10480 14946
rect 10400 14786 10480 14894
rect 10400 14734 10414 14786
rect 10466 14734 10480 14786
rect 10400 14626 10480 14734
rect 10400 14574 10414 14626
rect 10466 14574 10480 14626
rect 10400 14466 10480 14574
rect 10400 14414 10414 14466
rect 10466 14414 10480 14466
rect 10400 14306 10480 14414
rect 10400 14254 10414 14306
rect 10466 14254 10480 14306
rect 10400 14146 10480 14254
rect 10400 14094 10414 14146
rect 10466 14094 10480 14146
rect 10400 13986 10480 14094
rect 10400 13934 10414 13986
rect 10466 13934 10480 13986
rect 10400 13817 10480 13934
rect 10400 13783 10423 13817
rect 10457 13783 10480 13817
rect 10400 13666 10480 13783
rect 10400 13614 10414 13666
rect 10466 13614 10480 13666
rect 10400 13506 10480 13614
rect 10400 13454 10414 13506
rect 10466 13454 10480 13506
rect 10400 13346 10480 13454
rect 10400 13294 10414 13346
rect 10466 13294 10480 13346
rect 10400 13186 10480 13294
rect 10400 13134 10414 13186
rect 10466 13134 10480 13186
rect 10400 13026 10480 13134
rect 10400 12974 10414 13026
rect 10466 12974 10480 13026
rect 10400 12866 10480 12974
rect 10400 12814 10414 12866
rect 10466 12814 10480 12866
rect 10400 12706 10480 12814
rect 10400 12654 10414 12706
rect 10466 12654 10480 12706
rect 10400 12546 10480 12654
rect 10400 12494 10414 12546
rect 10466 12494 10480 12546
rect 10400 12377 10480 12494
rect 10400 12343 10423 12377
rect 10457 12343 10480 12377
rect 10400 12217 10480 12343
rect 10400 12183 10423 12217
rect 10457 12183 10480 12217
rect 10400 12057 10480 12183
rect 10400 12023 10423 12057
rect 10457 12023 10480 12057
rect 10400 11897 10480 12023
rect 10400 11863 10423 11897
rect 10457 11863 10480 11897
rect 10400 11746 10480 11863
rect 10400 11694 10414 11746
rect 10466 11694 10480 11746
rect 10400 11586 10480 11694
rect 10400 11534 10414 11586
rect 10466 11534 10480 11586
rect 10400 11426 10480 11534
rect 10400 11374 10414 11426
rect 10466 11374 10480 11426
rect 10400 11266 10480 11374
rect 10400 11214 10414 11266
rect 10466 11214 10480 11266
rect 10400 11106 10480 11214
rect 10400 11054 10414 11106
rect 10466 11054 10480 11106
rect 10400 10946 10480 11054
rect 10400 10894 10414 10946
rect 10466 10894 10480 10946
rect 10400 10786 10480 10894
rect 10400 10734 10414 10786
rect 10466 10734 10480 10786
rect 10400 10626 10480 10734
rect 10400 10574 10414 10626
rect 10466 10574 10480 10626
rect 10400 10466 10480 10574
rect 10400 10414 10414 10466
rect 10466 10414 10480 10466
rect 10400 10306 10480 10414
rect 10400 10254 10414 10306
rect 10466 10254 10480 10306
rect 10400 10146 10480 10254
rect 10400 10094 10414 10146
rect 10466 10094 10480 10146
rect 10400 9986 10480 10094
rect 10400 9934 10414 9986
rect 10466 9934 10480 9986
rect 10400 9826 10480 9934
rect 10400 9774 10414 9826
rect 10466 9774 10480 9826
rect 10400 9657 10480 9774
rect 10400 9623 10423 9657
rect 10457 9623 10480 9657
rect 10400 9506 10480 9623
rect 10400 9454 10414 9506
rect 10466 9454 10480 9506
rect 10400 9346 10480 9454
rect 10400 9294 10414 9346
rect 10466 9294 10480 9346
rect 10400 9177 10480 9294
rect 10400 9143 10423 9177
rect 10457 9143 10480 9177
rect 10400 9026 10480 9143
rect 10400 8974 10414 9026
rect 10466 8974 10480 9026
rect 10400 8866 10480 8974
rect 10400 8814 10414 8866
rect 10466 8814 10480 8866
rect 10400 8706 10480 8814
rect 10400 8654 10414 8706
rect 10466 8654 10480 8706
rect 10400 8546 10480 8654
rect 10400 8494 10414 8546
rect 10466 8494 10480 8546
rect 10400 8386 10480 8494
rect 10400 8334 10414 8386
rect 10466 8334 10480 8386
rect 10400 8226 10480 8334
rect 10400 8174 10414 8226
rect 10466 8174 10480 8226
rect 10400 8066 10480 8174
rect 10400 8014 10414 8066
rect 10466 8014 10480 8066
rect 10400 7906 10480 8014
rect 10400 7854 10414 7906
rect 10466 7854 10480 7906
rect 10400 7746 10480 7854
rect 10400 7694 10414 7746
rect 10466 7694 10480 7746
rect 10400 7577 10480 7694
rect 10400 7543 10423 7577
rect 10457 7543 10480 7577
rect 10400 7426 10480 7543
rect 10400 7374 10414 7426
rect 10466 7374 10480 7426
rect 10400 7266 10480 7374
rect 10400 7214 10414 7266
rect 10466 7214 10480 7266
rect 10400 7097 10480 7214
rect 10400 7063 10423 7097
rect 10457 7063 10480 7097
rect 10400 6946 10480 7063
rect 10400 6894 10414 6946
rect 10466 6894 10480 6946
rect 10400 6786 10480 6894
rect 10400 6734 10414 6786
rect 10466 6734 10480 6786
rect 10400 6617 10480 6734
rect 10400 6583 10423 6617
rect 10457 6583 10480 6617
rect 10400 6466 10480 6583
rect 10400 6414 10414 6466
rect 10466 6414 10480 6466
rect 10400 6306 10480 6414
rect 10400 6254 10414 6306
rect 10466 6254 10480 6306
rect 10400 6146 10480 6254
rect 10400 6094 10414 6146
rect 10466 6094 10480 6146
rect 10400 5986 10480 6094
rect 10400 5934 10414 5986
rect 10466 5934 10480 5986
rect 10400 5826 10480 5934
rect 10400 5774 10414 5826
rect 10466 5774 10480 5826
rect 10400 5666 10480 5774
rect 10400 5614 10414 5666
rect 10466 5614 10480 5666
rect 10400 5506 10480 5614
rect 10400 5454 10414 5506
rect 10466 5454 10480 5506
rect 10400 5346 10480 5454
rect 10400 5294 10414 5346
rect 10466 5294 10480 5346
rect 10400 5186 10480 5294
rect 10400 5134 10414 5186
rect 10466 5134 10480 5186
rect 10400 5026 10480 5134
rect 10400 4974 10414 5026
rect 10466 4974 10480 5026
rect 10400 4866 10480 4974
rect 10400 4814 10414 4866
rect 10466 4814 10480 4866
rect 10400 4706 10480 4814
rect 10400 4654 10414 4706
rect 10466 4654 10480 4706
rect 10400 4546 10480 4654
rect 10400 4494 10414 4546
rect 10466 4494 10480 4546
rect 10400 4386 10480 4494
rect 10400 4334 10414 4386
rect 10466 4334 10480 4386
rect 10400 4226 10480 4334
rect 10400 4174 10414 4226
rect 10466 4174 10480 4226
rect 10400 4066 10480 4174
rect 10400 4014 10414 4066
rect 10466 4014 10480 4066
rect 10400 3906 10480 4014
rect 10400 3854 10414 3906
rect 10466 3854 10480 3906
rect 10400 3737 10480 3854
rect 10400 3703 10423 3737
rect 10457 3703 10480 3737
rect 10400 3577 10480 3703
rect 10400 3543 10423 3577
rect 10457 3543 10480 3577
rect 10400 3426 10480 3543
rect 10400 3374 10414 3426
rect 10466 3374 10480 3426
rect 10400 3266 10480 3374
rect 10400 3214 10414 3266
rect 10466 3214 10480 3266
rect 10400 3106 10480 3214
rect 10400 3054 10414 3106
rect 10466 3054 10480 3106
rect 10400 2946 10480 3054
rect 10400 2894 10414 2946
rect 10466 2894 10480 2946
rect 10400 2786 10480 2894
rect 10400 2734 10414 2786
rect 10466 2734 10480 2786
rect 10400 2626 10480 2734
rect 10400 2574 10414 2626
rect 10466 2574 10480 2626
rect 10400 2466 10480 2574
rect 10400 2414 10414 2466
rect 10466 2414 10480 2466
rect 10400 2306 10480 2414
rect 10400 2254 10414 2306
rect 10466 2254 10480 2306
rect 10400 2146 10480 2254
rect 10400 2094 10414 2146
rect 10466 2094 10480 2146
rect 10400 1986 10480 2094
rect 10400 1934 10414 1986
rect 10466 1934 10480 1986
rect 10400 1817 10480 1934
rect 10400 1783 10423 1817
rect 10457 1783 10480 1817
rect 10400 1666 10480 1783
rect 10400 1614 10414 1666
rect 10466 1614 10480 1666
rect 10400 1506 10480 1614
rect 10400 1454 10414 1506
rect 10466 1454 10480 1506
rect 10400 1346 10480 1454
rect 10400 1294 10414 1346
rect 10466 1294 10480 1346
rect 10400 1186 10480 1294
rect 10400 1134 10414 1186
rect 10466 1134 10480 1186
rect 10400 1026 10480 1134
rect 10400 974 10414 1026
rect 10466 974 10480 1026
rect 10400 857 10480 974
rect 10400 823 10423 857
rect 10457 823 10480 857
rect 10400 697 10480 823
rect 10400 663 10423 697
rect 10457 663 10480 697
rect 10400 546 10480 663
rect 10400 494 10414 546
rect 10466 494 10480 546
rect 10400 386 10480 494
rect 10400 334 10414 386
rect 10466 334 10480 386
rect 10400 226 10480 334
rect 10400 174 10414 226
rect 10466 174 10480 226
rect 10400 66 10480 174
rect 10400 14 10414 66
rect 10466 14 10480 66
rect 10400 0 10480 14
rect 10560 31417 10640 31440
rect 10560 31383 10583 31417
rect 10617 31383 10640 31417
rect 10560 31257 10640 31383
rect 10560 31223 10583 31257
rect 10617 31223 10640 31257
rect 10560 31097 10640 31223
rect 10560 31063 10583 31097
rect 10617 31063 10640 31097
rect 10560 30937 10640 31063
rect 10560 30903 10583 30937
rect 10617 30903 10640 30937
rect 10560 30777 10640 30903
rect 10560 30743 10583 30777
rect 10617 30743 10640 30777
rect 10560 30617 10640 30743
rect 10560 30583 10583 30617
rect 10617 30583 10640 30617
rect 10560 30457 10640 30583
rect 10560 30423 10583 30457
rect 10617 30423 10640 30457
rect 10560 30297 10640 30423
rect 10560 30263 10583 30297
rect 10617 30263 10640 30297
rect 10560 30137 10640 30263
rect 10560 30103 10583 30137
rect 10617 30103 10640 30137
rect 10560 29977 10640 30103
rect 10560 29943 10583 29977
rect 10617 29943 10640 29977
rect 10560 29817 10640 29943
rect 10560 29783 10583 29817
rect 10617 29783 10640 29817
rect 10560 29657 10640 29783
rect 10560 29623 10583 29657
rect 10617 29623 10640 29657
rect 10560 29497 10640 29623
rect 10560 29463 10583 29497
rect 10617 29463 10640 29497
rect 10560 29337 10640 29463
rect 10560 29303 10583 29337
rect 10617 29303 10640 29337
rect 10560 29177 10640 29303
rect 10560 29143 10583 29177
rect 10617 29143 10640 29177
rect 10560 29017 10640 29143
rect 10560 28983 10583 29017
rect 10617 28983 10640 29017
rect 10560 28857 10640 28983
rect 10560 28823 10583 28857
rect 10617 28823 10640 28857
rect 10560 28697 10640 28823
rect 10560 28663 10583 28697
rect 10617 28663 10640 28697
rect 10560 28537 10640 28663
rect 10560 28503 10583 28537
rect 10617 28503 10640 28537
rect 10560 28377 10640 28503
rect 10560 28343 10583 28377
rect 10617 28343 10640 28377
rect 10560 28217 10640 28343
rect 10560 28183 10583 28217
rect 10617 28183 10640 28217
rect 10560 28057 10640 28183
rect 10560 28023 10583 28057
rect 10617 28023 10640 28057
rect 10560 27897 10640 28023
rect 10560 27863 10583 27897
rect 10617 27863 10640 27897
rect 10560 27737 10640 27863
rect 10560 27703 10583 27737
rect 10617 27703 10640 27737
rect 10560 27577 10640 27703
rect 10560 27543 10583 27577
rect 10617 27543 10640 27577
rect 10560 27417 10640 27543
rect 10560 27383 10583 27417
rect 10617 27383 10640 27417
rect 10560 27257 10640 27383
rect 10560 27223 10583 27257
rect 10617 27223 10640 27257
rect 10560 27097 10640 27223
rect 10560 27063 10583 27097
rect 10617 27063 10640 27097
rect 10560 26937 10640 27063
rect 10560 26903 10583 26937
rect 10617 26903 10640 26937
rect 10560 26777 10640 26903
rect 10560 26743 10583 26777
rect 10617 26743 10640 26777
rect 10560 26617 10640 26743
rect 10560 26583 10583 26617
rect 10617 26583 10640 26617
rect 10560 26457 10640 26583
rect 10560 26423 10583 26457
rect 10617 26423 10640 26457
rect 10560 26297 10640 26423
rect 10560 26263 10583 26297
rect 10617 26263 10640 26297
rect 10560 26137 10640 26263
rect 10560 26103 10583 26137
rect 10617 26103 10640 26137
rect 10560 25977 10640 26103
rect 10560 25943 10583 25977
rect 10617 25943 10640 25977
rect 10560 25817 10640 25943
rect 10560 25783 10583 25817
rect 10617 25783 10640 25817
rect 10560 25657 10640 25783
rect 10560 25623 10583 25657
rect 10617 25623 10640 25657
rect 10560 25497 10640 25623
rect 10560 25463 10583 25497
rect 10617 25463 10640 25497
rect 10560 25337 10640 25463
rect 10560 25303 10583 25337
rect 10617 25303 10640 25337
rect 10560 25177 10640 25303
rect 10560 25143 10583 25177
rect 10617 25143 10640 25177
rect 10560 25017 10640 25143
rect 10560 24983 10583 25017
rect 10617 24983 10640 25017
rect 10560 24857 10640 24983
rect 10560 24823 10583 24857
rect 10617 24823 10640 24857
rect 10560 24697 10640 24823
rect 10560 24663 10583 24697
rect 10617 24663 10640 24697
rect 10560 24537 10640 24663
rect 10560 24503 10583 24537
rect 10617 24503 10640 24537
rect 10560 24377 10640 24503
rect 10560 24343 10583 24377
rect 10617 24343 10640 24377
rect 10560 24217 10640 24343
rect 10560 24183 10583 24217
rect 10617 24183 10640 24217
rect 10560 24057 10640 24183
rect 10560 24023 10583 24057
rect 10617 24023 10640 24057
rect 10560 23897 10640 24023
rect 10560 23863 10583 23897
rect 10617 23863 10640 23897
rect 10560 23737 10640 23863
rect 10560 23703 10583 23737
rect 10617 23703 10640 23737
rect 10560 23577 10640 23703
rect 10560 23543 10583 23577
rect 10617 23543 10640 23577
rect 10560 23417 10640 23543
rect 10560 23383 10583 23417
rect 10617 23383 10640 23417
rect 10560 23257 10640 23383
rect 10560 23223 10583 23257
rect 10617 23223 10640 23257
rect 10560 23097 10640 23223
rect 10560 23063 10583 23097
rect 10617 23063 10640 23097
rect 10560 22937 10640 23063
rect 10560 22903 10583 22937
rect 10617 22903 10640 22937
rect 10560 22777 10640 22903
rect 10560 22743 10583 22777
rect 10617 22743 10640 22777
rect 10560 22617 10640 22743
rect 10560 22583 10583 22617
rect 10617 22583 10640 22617
rect 10560 22457 10640 22583
rect 10560 22423 10583 22457
rect 10617 22423 10640 22457
rect 10560 22297 10640 22423
rect 10560 22263 10583 22297
rect 10617 22263 10640 22297
rect 10560 22137 10640 22263
rect 10560 22103 10583 22137
rect 10617 22103 10640 22137
rect 10560 21977 10640 22103
rect 10560 21943 10583 21977
rect 10617 21943 10640 21977
rect 10560 21817 10640 21943
rect 10560 21783 10583 21817
rect 10617 21783 10640 21817
rect 10560 21657 10640 21783
rect 10560 21623 10583 21657
rect 10617 21623 10640 21657
rect 10560 21497 10640 21623
rect 10560 21463 10583 21497
rect 10617 21463 10640 21497
rect 10560 21337 10640 21463
rect 10560 21303 10583 21337
rect 10617 21303 10640 21337
rect 10560 21177 10640 21303
rect 10560 21143 10583 21177
rect 10617 21143 10640 21177
rect 10560 21017 10640 21143
rect 10560 20983 10583 21017
rect 10617 20983 10640 21017
rect 10560 20857 10640 20983
rect 10560 20823 10583 20857
rect 10617 20823 10640 20857
rect 10560 20697 10640 20823
rect 10560 20663 10583 20697
rect 10617 20663 10640 20697
rect 10560 20537 10640 20663
rect 10560 20503 10583 20537
rect 10617 20503 10640 20537
rect 10560 20377 10640 20503
rect 10560 20343 10583 20377
rect 10617 20343 10640 20377
rect 10560 20217 10640 20343
rect 10560 20183 10583 20217
rect 10617 20183 10640 20217
rect 10560 20057 10640 20183
rect 10560 20023 10583 20057
rect 10617 20023 10640 20057
rect 10560 19897 10640 20023
rect 10560 19863 10583 19897
rect 10617 19863 10640 19897
rect 10560 19737 10640 19863
rect 10560 19703 10583 19737
rect 10617 19703 10640 19737
rect 10560 19577 10640 19703
rect 10560 19543 10583 19577
rect 10617 19543 10640 19577
rect 10560 19417 10640 19543
rect 10560 19383 10583 19417
rect 10617 19383 10640 19417
rect 10560 19257 10640 19383
rect 10560 19223 10583 19257
rect 10617 19223 10640 19257
rect 10560 19097 10640 19223
rect 10560 19063 10583 19097
rect 10617 19063 10640 19097
rect 10560 18937 10640 19063
rect 10560 18903 10583 18937
rect 10617 18903 10640 18937
rect 10560 18777 10640 18903
rect 10560 18743 10583 18777
rect 10617 18743 10640 18777
rect 10560 18617 10640 18743
rect 10560 18583 10583 18617
rect 10617 18583 10640 18617
rect 10560 18457 10640 18583
rect 10560 18423 10583 18457
rect 10617 18423 10640 18457
rect 10560 18297 10640 18423
rect 10560 18263 10583 18297
rect 10617 18263 10640 18297
rect 10560 18137 10640 18263
rect 10560 18103 10583 18137
rect 10617 18103 10640 18137
rect 10560 17977 10640 18103
rect 10560 17943 10583 17977
rect 10617 17943 10640 17977
rect 10560 17817 10640 17943
rect 10560 17783 10583 17817
rect 10617 17783 10640 17817
rect 10560 17657 10640 17783
rect 10560 17623 10583 17657
rect 10617 17623 10640 17657
rect 10560 17497 10640 17623
rect 10560 17463 10583 17497
rect 10617 17463 10640 17497
rect 10560 17337 10640 17463
rect 10560 17303 10583 17337
rect 10617 17303 10640 17337
rect 10560 17177 10640 17303
rect 10560 17143 10583 17177
rect 10617 17143 10640 17177
rect 10560 17017 10640 17143
rect 10560 16983 10583 17017
rect 10617 16983 10640 17017
rect 10560 16857 10640 16983
rect 10560 16823 10583 16857
rect 10617 16823 10640 16857
rect 10560 16697 10640 16823
rect 10560 16663 10583 16697
rect 10617 16663 10640 16697
rect 10560 16537 10640 16663
rect 10560 16503 10583 16537
rect 10617 16503 10640 16537
rect 10560 16377 10640 16503
rect 10560 16343 10583 16377
rect 10617 16343 10640 16377
rect 10560 16217 10640 16343
rect 10560 16183 10583 16217
rect 10617 16183 10640 16217
rect 10560 16057 10640 16183
rect 10560 16023 10583 16057
rect 10617 16023 10640 16057
rect 10560 15897 10640 16023
rect 10560 15863 10583 15897
rect 10617 15863 10640 15897
rect 10560 15737 10640 15863
rect 10560 15703 10583 15737
rect 10617 15703 10640 15737
rect 10560 15577 10640 15703
rect 10560 15543 10583 15577
rect 10617 15543 10640 15577
rect 10560 15417 10640 15543
rect 10560 15383 10583 15417
rect 10617 15383 10640 15417
rect 10560 15257 10640 15383
rect 10560 15223 10583 15257
rect 10617 15223 10640 15257
rect 10560 15097 10640 15223
rect 10560 15063 10583 15097
rect 10617 15063 10640 15097
rect 10560 14937 10640 15063
rect 10560 14903 10583 14937
rect 10617 14903 10640 14937
rect 10560 14777 10640 14903
rect 10560 14743 10583 14777
rect 10617 14743 10640 14777
rect 10560 14617 10640 14743
rect 10560 14583 10583 14617
rect 10617 14583 10640 14617
rect 10560 14457 10640 14583
rect 10560 14423 10583 14457
rect 10617 14423 10640 14457
rect 10560 14297 10640 14423
rect 10560 14263 10583 14297
rect 10617 14263 10640 14297
rect 10560 14137 10640 14263
rect 10560 14103 10583 14137
rect 10617 14103 10640 14137
rect 10560 13977 10640 14103
rect 10560 13943 10583 13977
rect 10617 13943 10640 13977
rect 10560 13817 10640 13943
rect 10560 13783 10583 13817
rect 10617 13783 10640 13817
rect 10560 13657 10640 13783
rect 10560 13623 10583 13657
rect 10617 13623 10640 13657
rect 10560 13497 10640 13623
rect 10560 13463 10583 13497
rect 10617 13463 10640 13497
rect 10560 13337 10640 13463
rect 10560 13303 10583 13337
rect 10617 13303 10640 13337
rect 10560 13177 10640 13303
rect 10560 13143 10583 13177
rect 10617 13143 10640 13177
rect 10560 13017 10640 13143
rect 10560 12983 10583 13017
rect 10617 12983 10640 13017
rect 10560 12857 10640 12983
rect 10560 12823 10583 12857
rect 10617 12823 10640 12857
rect 10560 12697 10640 12823
rect 10560 12663 10583 12697
rect 10617 12663 10640 12697
rect 10560 12537 10640 12663
rect 10560 12503 10583 12537
rect 10617 12503 10640 12537
rect 10560 12377 10640 12503
rect 10560 12343 10583 12377
rect 10617 12343 10640 12377
rect 10560 12217 10640 12343
rect 10560 12183 10583 12217
rect 10617 12183 10640 12217
rect 10560 12057 10640 12183
rect 10560 12023 10583 12057
rect 10617 12023 10640 12057
rect 10560 11897 10640 12023
rect 10560 11863 10583 11897
rect 10617 11863 10640 11897
rect 10560 11737 10640 11863
rect 10560 11703 10583 11737
rect 10617 11703 10640 11737
rect 10560 11577 10640 11703
rect 10560 11543 10583 11577
rect 10617 11543 10640 11577
rect 10560 11417 10640 11543
rect 10560 11383 10583 11417
rect 10617 11383 10640 11417
rect 10560 11257 10640 11383
rect 10560 11223 10583 11257
rect 10617 11223 10640 11257
rect 10560 11097 10640 11223
rect 10560 11063 10583 11097
rect 10617 11063 10640 11097
rect 10560 10937 10640 11063
rect 10560 10903 10583 10937
rect 10617 10903 10640 10937
rect 10560 10777 10640 10903
rect 10560 10743 10583 10777
rect 10617 10743 10640 10777
rect 10560 10617 10640 10743
rect 10560 10583 10583 10617
rect 10617 10583 10640 10617
rect 10560 10457 10640 10583
rect 10560 10423 10583 10457
rect 10617 10423 10640 10457
rect 10560 10297 10640 10423
rect 10560 10263 10583 10297
rect 10617 10263 10640 10297
rect 10560 10137 10640 10263
rect 10560 10103 10583 10137
rect 10617 10103 10640 10137
rect 10560 9977 10640 10103
rect 10560 9943 10583 9977
rect 10617 9943 10640 9977
rect 10560 9817 10640 9943
rect 10560 9783 10583 9817
rect 10617 9783 10640 9817
rect 10560 9657 10640 9783
rect 10560 9623 10583 9657
rect 10617 9623 10640 9657
rect 10560 9497 10640 9623
rect 10560 9463 10583 9497
rect 10617 9463 10640 9497
rect 10560 9337 10640 9463
rect 10560 9303 10583 9337
rect 10617 9303 10640 9337
rect 10560 9177 10640 9303
rect 10560 9143 10583 9177
rect 10617 9143 10640 9177
rect 10560 9017 10640 9143
rect 10560 8983 10583 9017
rect 10617 8983 10640 9017
rect 10560 8857 10640 8983
rect 10560 8823 10583 8857
rect 10617 8823 10640 8857
rect 10560 8697 10640 8823
rect 10560 8663 10583 8697
rect 10617 8663 10640 8697
rect 10560 8537 10640 8663
rect 10560 8503 10583 8537
rect 10617 8503 10640 8537
rect 10560 8377 10640 8503
rect 10560 8343 10583 8377
rect 10617 8343 10640 8377
rect 10560 8217 10640 8343
rect 10560 8183 10583 8217
rect 10617 8183 10640 8217
rect 10560 8057 10640 8183
rect 10560 8023 10583 8057
rect 10617 8023 10640 8057
rect 10560 7897 10640 8023
rect 10560 7863 10583 7897
rect 10617 7863 10640 7897
rect 10560 7737 10640 7863
rect 10560 7703 10583 7737
rect 10617 7703 10640 7737
rect 10560 7577 10640 7703
rect 10560 7543 10583 7577
rect 10617 7543 10640 7577
rect 10560 7417 10640 7543
rect 10560 7383 10583 7417
rect 10617 7383 10640 7417
rect 10560 7257 10640 7383
rect 10560 7223 10583 7257
rect 10617 7223 10640 7257
rect 10560 7097 10640 7223
rect 10560 7063 10583 7097
rect 10617 7063 10640 7097
rect 10560 6937 10640 7063
rect 10560 6903 10583 6937
rect 10617 6903 10640 6937
rect 10560 6777 10640 6903
rect 10560 6743 10583 6777
rect 10617 6743 10640 6777
rect 10560 6617 10640 6743
rect 10560 6583 10583 6617
rect 10617 6583 10640 6617
rect 10560 6457 10640 6583
rect 10560 6423 10583 6457
rect 10617 6423 10640 6457
rect 10560 6297 10640 6423
rect 10560 6263 10583 6297
rect 10617 6263 10640 6297
rect 10560 6137 10640 6263
rect 10560 6103 10583 6137
rect 10617 6103 10640 6137
rect 10560 5977 10640 6103
rect 10560 5943 10583 5977
rect 10617 5943 10640 5977
rect 10560 5817 10640 5943
rect 10560 5783 10583 5817
rect 10617 5783 10640 5817
rect 10560 5657 10640 5783
rect 10560 5623 10583 5657
rect 10617 5623 10640 5657
rect 10560 5497 10640 5623
rect 10560 5463 10583 5497
rect 10617 5463 10640 5497
rect 10560 5337 10640 5463
rect 10560 5303 10583 5337
rect 10617 5303 10640 5337
rect 10560 5177 10640 5303
rect 10560 5143 10583 5177
rect 10617 5143 10640 5177
rect 10560 5017 10640 5143
rect 10560 4983 10583 5017
rect 10617 4983 10640 5017
rect 10560 4857 10640 4983
rect 10560 4823 10583 4857
rect 10617 4823 10640 4857
rect 10560 4697 10640 4823
rect 10560 4663 10583 4697
rect 10617 4663 10640 4697
rect 10560 4537 10640 4663
rect 10560 4503 10583 4537
rect 10617 4503 10640 4537
rect 10560 4377 10640 4503
rect 10560 4343 10583 4377
rect 10617 4343 10640 4377
rect 10560 4217 10640 4343
rect 10560 4183 10583 4217
rect 10617 4183 10640 4217
rect 10560 4057 10640 4183
rect 10560 4023 10583 4057
rect 10617 4023 10640 4057
rect 10560 3897 10640 4023
rect 10560 3863 10583 3897
rect 10617 3863 10640 3897
rect 10560 3737 10640 3863
rect 10560 3703 10583 3737
rect 10617 3703 10640 3737
rect 10560 3577 10640 3703
rect 10560 3543 10583 3577
rect 10617 3543 10640 3577
rect 10560 3417 10640 3543
rect 10560 3383 10583 3417
rect 10617 3383 10640 3417
rect 10560 3257 10640 3383
rect 10560 3223 10583 3257
rect 10617 3223 10640 3257
rect 10560 3097 10640 3223
rect 10560 3063 10583 3097
rect 10617 3063 10640 3097
rect 10560 2937 10640 3063
rect 10560 2903 10583 2937
rect 10617 2903 10640 2937
rect 10560 2777 10640 2903
rect 10560 2743 10583 2777
rect 10617 2743 10640 2777
rect 10560 2617 10640 2743
rect 10560 2583 10583 2617
rect 10617 2583 10640 2617
rect 10560 2457 10640 2583
rect 10560 2423 10583 2457
rect 10617 2423 10640 2457
rect 10560 2297 10640 2423
rect 10560 2263 10583 2297
rect 10617 2263 10640 2297
rect 10560 2137 10640 2263
rect 10560 2103 10583 2137
rect 10617 2103 10640 2137
rect 10560 1977 10640 2103
rect 10560 1943 10583 1977
rect 10617 1943 10640 1977
rect 10560 1817 10640 1943
rect 10560 1783 10583 1817
rect 10617 1783 10640 1817
rect 10560 1657 10640 1783
rect 10560 1623 10583 1657
rect 10617 1623 10640 1657
rect 10560 1497 10640 1623
rect 10560 1463 10583 1497
rect 10617 1463 10640 1497
rect 10560 1337 10640 1463
rect 10560 1303 10583 1337
rect 10617 1303 10640 1337
rect 10560 1177 10640 1303
rect 10560 1143 10583 1177
rect 10617 1143 10640 1177
rect 10560 1017 10640 1143
rect 10560 983 10583 1017
rect 10617 983 10640 1017
rect 10560 857 10640 983
rect 10560 823 10583 857
rect 10617 823 10640 857
rect 10560 697 10640 823
rect 10560 663 10583 697
rect 10617 663 10640 697
rect 10560 537 10640 663
rect 10560 503 10583 537
rect 10617 503 10640 537
rect 10560 377 10640 503
rect 10560 343 10583 377
rect 10617 343 10640 377
rect 10560 217 10640 343
rect 10560 183 10583 217
rect 10617 183 10640 217
rect 10560 57 10640 183
rect 10560 23 10583 57
rect 10617 23 10640 57
rect 10560 0 10640 23
rect 10720 31426 10800 31440
rect 10720 31374 10734 31426
rect 10786 31374 10800 31426
rect 10720 31266 10800 31374
rect 10720 31214 10734 31266
rect 10786 31214 10800 31266
rect 10720 31106 10800 31214
rect 10720 31054 10734 31106
rect 10786 31054 10800 31106
rect 10720 30946 10800 31054
rect 10720 30894 10734 30946
rect 10786 30894 10800 30946
rect 10720 30786 10800 30894
rect 10720 30734 10734 30786
rect 10786 30734 10800 30786
rect 10720 30626 10800 30734
rect 10720 30574 10734 30626
rect 10786 30574 10800 30626
rect 10720 30466 10800 30574
rect 10720 30414 10734 30466
rect 10786 30414 10800 30466
rect 10720 30306 10800 30414
rect 10720 30254 10734 30306
rect 10786 30254 10800 30306
rect 10720 30137 10800 30254
rect 10720 30103 10743 30137
rect 10777 30103 10800 30137
rect 10720 29986 10800 30103
rect 10720 29934 10734 29986
rect 10786 29934 10800 29986
rect 10720 29826 10800 29934
rect 10720 29774 10734 29826
rect 10786 29774 10800 29826
rect 10720 29666 10800 29774
rect 10720 29614 10734 29666
rect 10786 29614 10800 29666
rect 10720 29506 10800 29614
rect 10720 29454 10734 29506
rect 10786 29454 10800 29506
rect 10720 29346 10800 29454
rect 10720 29294 10734 29346
rect 10786 29294 10800 29346
rect 10720 29186 10800 29294
rect 10720 29134 10734 29186
rect 10786 29134 10800 29186
rect 10720 29026 10800 29134
rect 10720 28974 10734 29026
rect 10786 28974 10800 29026
rect 10720 28866 10800 28974
rect 10720 28814 10734 28866
rect 10786 28814 10800 28866
rect 10720 28697 10800 28814
rect 10720 28663 10743 28697
rect 10777 28663 10800 28697
rect 10720 28537 10800 28663
rect 10720 28503 10743 28537
rect 10777 28503 10800 28537
rect 10720 28377 10800 28503
rect 10720 28343 10743 28377
rect 10777 28343 10800 28377
rect 10720 28217 10800 28343
rect 10720 28183 10743 28217
rect 10777 28183 10800 28217
rect 10720 28066 10800 28183
rect 10720 28014 10734 28066
rect 10786 28014 10800 28066
rect 10720 27906 10800 28014
rect 10720 27854 10734 27906
rect 10786 27854 10800 27906
rect 10720 27746 10800 27854
rect 10720 27694 10734 27746
rect 10786 27694 10800 27746
rect 10720 27586 10800 27694
rect 10720 27534 10734 27586
rect 10786 27534 10800 27586
rect 10720 27426 10800 27534
rect 10720 27374 10734 27426
rect 10786 27374 10800 27426
rect 10720 27266 10800 27374
rect 10720 27214 10734 27266
rect 10786 27214 10800 27266
rect 10720 27106 10800 27214
rect 10720 27054 10734 27106
rect 10786 27054 10800 27106
rect 10720 26946 10800 27054
rect 10720 26894 10734 26946
rect 10786 26894 10800 26946
rect 10720 26777 10800 26894
rect 10720 26743 10743 26777
rect 10777 26743 10800 26777
rect 10720 26617 10800 26743
rect 10720 26583 10743 26617
rect 10777 26583 10800 26617
rect 10720 26457 10800 26583
rect 10720 26423 10743 26457
rect 10777 26423 10800 26457
rect 10720 26297 10800 26423
rect 10720 26263 10743 26297
rect 10777 26263 10800 26297
rect 10720 26146 10800 26263
rect 10720 26094 10734 26146
rect 10786 26094 10800 26146
rect 10720 25986 10800 26094
rect 10720 25934 10734 25986
rect 10786 25934 10800 25986
rect 10720 25826 10800 25934
rect 10720 25774 10734 25826
rect 10786 25774 10800 25826
rect 10720 25666 10800 25774
rect 10720 25614 10734 25666
rect 10786 25614 10800 25666
rect 10720 25506 10800 25614
rect 10720 25454 10734 25506
rect 10786 25454 10800 25506
rect 10720 25346 10800 25454
rect 10720 25294 10734 25346
rect 10786 25294 10800 25346
rect 10720 25186 10800 25294
rect 10720 25134 10734 25186
rect 10786 25134 10800 25186
rect 10720 25026 10800 25134
rect 10720 24974 10734 25026
rect 10786 24974 10800 25026
rect 10720 24857 10800 24974
rect 10720 24823 10743 24857
rect 10777 24823 10800 24857
rect 10720 24706 10800 24823
rect 10720 24654 10734 24706
rect 10786 24654 10800 24706
rect 10720 24546 10800 24654
rect 10720 24494 10734 24546
rect 10786 24494 10800 24546
rect 10720 24386 10800 24494
rect 10720 24334 10734 24386
rect 10786 24334 10800 24386
rect 10720 24226 10800 24334
rect 10720 24174 10734 24226
rect 10786 24174 10800 24226
rect 10720 24066 10800 24174
rect 10720 24014 10734 24066
rect 10786 24014 10800 24066
rect 10720 23906 10800 24014
rect 10720 23854 10734 23906
rect 10786 23854 10800 23906
rect 10720 23746 10800 23854
rect 10720 23694 10734 23746
rect 10786 23694 10800 23746
rect 10720 23586 10800 23694
rect 10720 23534 10734 23586
rect 10786 23534 10800 23586
rect 10720 23426 10800 23534
rect 10720 23374 10734 23426
rect 10786 23374 10800 23426
rect 10720 23266 10800 23374
rect 10720 23214 10734 23266
rect 10786 23214 10800 23266
rect 10720 23106 10800 23214
rect 10720 23054 10734 23106
rect 10786 23054 10800 23106
rect 10720 22946 10800 23054
rect 10720 22894 10734 22946
rect 10786 22894 10800 22946
rect 10720 22786 10800 22894
rect 10720 22734 10734 22786
rect 10786 22734 10800 22786
rect 10720 22626 10800 22734
rect 10720 22574 10734 22626
rect 10786 22574 10800 22626
rect 10720 22466 10800 22574
rect 10720 22414 10734 22466
rect 10786 22414 10800 22466
rect 10720 22306 10800 22414
rect 10720 22254 10734 22306
rect 10786 22254 10800 22306
rect 10720 22146 10800 22254
rect 10720 22094 10734 22146
rect 10786 22094 10800 22146
rect 10720 21977 10800 22094
rect 10720 21943 10743 21977
rect 10777 21943 10800 21977
rect 10720 21826 10800 21943
rect 10720 21774 10734 21826
rect 10786 21774 10800 21826
rect 10720 21666 10800 21774
rect 10720 21614 10734 21666
rect 10786 21614 10800 21666
rect 10720 21506 10800 21614
rect 10720 21454 10734 21506
rect 10786 21454 10800 21506
rect 10720 21346 10800 21454
rect 10720 21294 10734 21346
rect 10786 21294 10800 21346
rect 10720 21186 10800 21294
rect 10720 21134 10734 21186
rect 10786 21134 10800 21186
rect 10720 21026 10800 21134
rect 10720 20974 10734 21026
rect 10786 20974 10800 21026
rect 10720 20866 10800 20974
rect 10720 20814 10734 20866
rect 10786 20814 10800 20866
rect 10720 20706 10800 20814
rect 10720 20654 10734 20706
rect 10786 20654 10800 20706
rect 10720 20537 10800 20654
rect 10720 20503 10743 20537
rect 10777 20503 10800 20537
rect 10720 20377 10800 20503
rect 10720 20343 10743 20377
rect 10777 20343 10800 20377
rect 10720 20217 10800 20343
rect 10720 20183 10743 20217
rect 10777 20183 10800 20217
rect 10720 20057 10800 20183
rect 10720 20023 10743 20057
rect 10777 20023 10800 20057
rect 10720 19906 10800 20023
rect 10720 19854 10734 19906
rect 10786 19854 10800 19906
rect 10720 19746 10800 19854
rect 10720 19694 10734 19746
rect 10786 19694 10800 19746
rect 10720 19586 10800 19694
rect 10720 19534 10734 19586
rect 10786 19534 10800 19586
rect 10720 19426 10800 19534
rect 10720 19374 10734 19426
rect 10786 19374 10800 19426
rect 10720 19266 10800 19374
rect 10720 19214 10734 19266
rect 10786 19214 10800 19266
rect 10720 19106 10800 19214
rect 10720 19054 10734 19106
rect 10786 19054 10800 19106
rect 10720 18946 10800 19054
rect 10720 18894 10734 18946
rect 10786 18894 10800 18946
rect 10720 18786 10800 18894
rect 10720 18734 10734 18786
rect 10786 18734 10800 18786
rect 10720 18617 10800 18734
rect 10720 18583 10743 18617
rect 10777 18583 10800 18617
rect 10720 18457 10800 18583
rect 10720 18423 10743 18457
rect 10777 18423 10800 18457
rect 10720 18297 10800 18423
rect 10720 18263 10743 18297
rect 10777 18263 10800 18297
rect 10720 18137 10800 18263
rect 10720 18103 10743 18137
rect 10777 18103 10800 18137
rect 10720 17986 10800 18103
rect 10720 17934 10734 17986
rect 10786 17934 10800 17986
rect 10720 17826 10800 17934
rect 10720 17774 10734 17826
rect 10786 17774 10800 17826
rect 10720 17666 10800 17774
rect 10720 17614 10734 17666
rect 10786 17614 10800 17666
rect 10720 17506 10800 17614
rect 10720 17454 10734 17506
rect 10786 17454 10800 17506
rect 10720 17346 10800 17454
rect 10720 17294 10734 17346
rect 10786 17294 10800 17346
rect 10720 17186 10800 17294
rect 10720 17134 10734 17186
rect 10786 17134 10800 17186
rect 10720 17026 10800 17134
rect 10720 16974 10734 17026
rect 10786 16974 10800 17026
rect 10720 16866 10800 16974
rect 10720 16814 10734 16866
rect 10786 16814 10800 16866
rect 10720 16697 10800 16814
rect 10720 16663 10743 16697
rect 10777 16663 10800 16697
rect 10720 16546 10800 16663
rect 10720 16494 10734 16546
rect 10786 16494 10800 16546
rect 10720 16386 10800 16494
rect 10720 16334 10734 16386
rect 10786 16334 10800 16386
rect 10720 16226 10800 16334
rect 10720 16174 10734 16226
rect 10786 16174 10800 16226
rect 10720 16066 10800 16174
rect 10720 16014 10734 16066
rect 10786 16014 10800 16066
rect 10720 15906 10800 16014
rect 10720 15854 10734 15906
rect 10786 15854 10800 15906
rect 10720 15746 10800 15854
rect 10720 15694 10734 15746
rect 10786 15694 10800 15746
rect 10720 15586 10800 15694
rect 10720 15534 10734 15586
rect 10786 15534 10800 15586
rect 10720 15426 10800 15534
rect 10720 15374 10734 15426
rect 10786 15374 10800 15426
rect 10720 15266 10800 15374
rect 10720 15214 10734 15266
rect 10786 15214 10800 15266
rect 10720 15106 10800 15214
rect 10720 15054 10734 15106
rect 10786 15054 10800 15106
rect 10720 14946 10800 15054
rect 10720 14894 10734 14946
rect 10786 14894 10800 14946
rect 10720 14786 10800 14894
rect 10720 14734 10734 14786
rect 10786 14734 10800 14786
rect 10720 14626 10800 14734
rect 10720 14574 10734 14626
rect 10786 14574 10800 14626
rect 10720 14466 10800 14574
rect 10720 14414 10734 14466
rect 10786 14414 10800 14466
rect 10720 14306 10800 14414
rect 10720 14254 10734 14306
rect 10786 14254 10800 14306
rect 10720 14146 10800 14254
rect 10720 14094 10734 14146
rect 10786 14094 10800 14146
rect 10720 13986 10800 14094
rect 10720 13934 10734 13986
rect 10786 13934 10800 13986
rect 10720 13817 10800 13934
rect 10720 13783 10743 13817
rect 10777 13783 10800 13817
rect 10720 13666 10800 13783
rect 10720 13614 10734 13666
rect 10786 13614 10800 13666
rect 10720 13506 10800 13614
rect 10720 13454 10734 13506
rect 10786 13454 10800 13506
rect 10720 13346 10800 13454
rect 10720 13294 10734 13346
rect 10786 13294 10800 13346
rect 10720 13186 10800 13294
rect 10720 13134 10734 13186
rect 10786 13134 10800 13186
rect 10720 13026 10800 13134
rect 10720 12974 10734 13026
rect 10786 12974 10800 13026
rect 10720 12866 10800 12974
rect 10720 12814 10734 12866
rect 10786 12814 10800 12866
rect 10720 12706 10800 12814
rect 10720 12654 10734 12706
rect 10786 12654 10800 12706
rect 10720 12546 10800 12654
rect 10720 12494 10734 12546
rect 10786 12494 10800 12546
rect 10720 12377 10800 12494
rect 10720 12343 10743 12377
rect 10777 12343 10800 12377
rect 10720 12217 10800 12343
rect 10720 12183 10743 12217
rect 10777 12183 10800 12217
rect 10720 12057 10800 12183
rect 10720 12023 10743 12057
rect 10777 12023 10800 12057
rect 10720 11897 10800 12023
rect 10720 11863 10743 11897
rect 10777 11863 10800 11897
rect 10720 11746 10800 11863
rect 10720 11694 10734 11746
rect 10786 11694 10800 11746
rect 10720 11586 10800 11694
rect 10720 11534 10734 11586
rect 10786 11534 10800 11586
rect 10720 11426 10800 11534
rect 10720 11374 10734 11426
rect 10786 11374 10800 11426
rect 10720 11266 10800 11374
rect 10720 11214 10734 11266
rect 10786 11214 10800 11266
rect 10720 11106 10800 11214
rect 10720 11054 10734 11106
rect 10786 11054 10800 11106
rect 10720 10946 10800 11054
rect 10720 10894 10734 10946
rect 10786 10894 10800 10946
rect 10720 10786 10800 10894
rect 10720 10734 10734 10786
rect 10786 10734 10800 10786
rect 10720 10626 10800 10734
rect 10720 10574 10734 10626
rect 10786 10574 10800 10626
rect 10720 10466 10800 10574
rect 10720 10414 10734 10466
rect 10786 10414 10800 10466
rect 10720 10306 10800 10414
rect 10720 10254 10734 10306
rect 10786 10254 10800 10306
rect 10720 10146 10800 10254
rect 10720 10094 10734 10146
rect 10786 10094 10800 10146
rect 10720 9986 10800 10094
rect 10720 9934 10734 9986
rect 10786 9934 10800 9986
rect 10720 9826 10800 9934
rect 10720 9774 10734 9826
rect 10786 9774 10800 9826
rect 10720 9657 10800 9774
rect 10720 9623 10743 9657
rect 10777 9623 10800 9657
rect 10720 9506 10800 9623
rect 10720 9454 10734 9506
rect 10786 9454 10800 9506
rect 10720 9346 10800 9454
rect 10720 9294 10734 9346
rect 10786 9294 10800 9346
rect 10720 9177 10800 9294
rect 10720 9143 10743 9177
rect 10777 9143 10800 9177
rect 10720 9026 10800 9143
rect 10720 8974 10734 9026
rect 10786 8974 10800 9026
rect 10720 8866 10800 8974
rect 10720 8814 10734 8866
rect 10786 8814 10800 8866
rect 10720 8706 10800 8814
rect 10720 8654 10734 8706
rect 10786 8654 10800 8706
rect 10720 8546 10800 8654
rect 10720 8494 10734 8546
rect 10786 8494 10800 8546
rect 10720 8386 10800 8494
rect 10720 8334 10734 8386
rect 10786 8334 10800 8386
rect 10720 8226 10800 8334
rect 10720 8174 10734 8226
rect 10786 8174 10800 8226
rect 10720 8066 10800 8174
rect 10720 8014 10734 8066
rect 10786 8014 10800 8066
rect 10720 7906 10800 8014
rect 10720 7854 10734 7906
rect 10786 7854 10800 7906
rect 10720 7746 10800 7854
rect 10720 7694 10734 7746
rect 10786 7694 10800 7746
rect 10720 7577 10800 7694
rect 10720 7543 10743 7577
rect 10777 7543 10800 7577
rect 10720 7426 10800 7543
rect 10720 7374 10734 7426
rect 10786 7374 10800 7426
rect 10720 7266 10800 7374
rect 10720 7214 10734 7266
rect 10786 7214 10800 7266
rect 10720 7097 10800 7214
rect 10720 7063 10743 7097
rect 10777 7063 10800 7097
rect 10720 6946 10800 7063
rect 10720 6894 10734 6946
rect 10786 6894 10800 6946
rect 10720 6786 10800 6894
rect 10720 6734 10734 6786
rect 10786 6734 10800 6786
rect 10720 6617 10800 6734
rect 10720 6583 10743 6617
rect 10777 6583 10800 6617
rect 10720 6466 10800 6583
rect 10720 6414 10734 6466
rect 10786 6414 10800 6466
rect 10720 6306 10800 6414
rect 10720 6254 10734 6306
rect 10786 6254 10800 6306
rect 10720 6146 10800 6254
rect 10720 6094 10734 6146
rect 10786 6094 10800 6146
rect 10720 5986 10800 6094
rect 10720 5934 10734 5986
rect 10786 5934 10800 5986
rect 10720 5826 10800 5934
rect 10720 5774 10734 5826
rect 10786 5774 10800 5826
rect 10720 5666 10800 5774
rect 10720 5614 10734 5666
rect 10786 5614 10800 5666
rect 10720 5506 10800 5614
rect 10720 5454 10734 5506
rect 10786 5454 10800 5506
rect 10720 5346 10800 5454
rect 10720 5294 10734 5346
rect 10786 5294 10800 5346
rect 10720 5186 10800 5294
rect 10720 5134 10734 5186
rect 10786 5134 10800 5186
rect 10720 5026 10800 5134
rect 10720 4974 10734 5026
rect 10786 4974 10800 5026
rect 10720 4866 10800 4974
rect 10720 4814 10734 4866
rect 10786 4814 10800 4866
rect 10720 4706 10800 4814
rect 10720 4654 10734 4706
rect 10786 4654 10800 4706
rect 10720 4546 10800 4654
rect 10720 4494 10734 4546
rect 10786 4494 10800 4546
rect 10720 4386 10800 4494
rect 10720 4334 10734 4386
rect 10786 4334 10800 4386
rect 10720 4226 10800 4334
rect 10720 4174 10734 4226
rect 10786 4174 10800 4226
rect 10720 4066 10800 4174
rect 10720 4014 10734 4066
rect 10786 4014 10800 4066
rect 10720 3906 10800 4014
rect 10720 3854 10734 3906
rect 10786 3854 10800 3906
rect 10720 3737 10800 3854
rect 10720 3703 10743 3737
rect 10777 3703 10800 3737
rect 10720 3577 10800 3703
rect 10720 3543 10743 3577
rect 10777 3543 10800 3577
rect 10720 3426 10800 3543
rect 10720 3374 10734 3426
rect 10786 3374 10800 3426
rect 10720 3266 10800 3374
rect 10720 3214 10734 3266
rect 10786 3214 10800 3266
rect 10720 3106 10800 3214
rect 10720 3054 10734 3106
rect 10786 3054 10800 3106
rect 10720 2946 10800 3054
rect 10720 2894 10734 2946
rect 10786 2894 10800 2946
rect 10720 2786 10800 2894
rect 10720 2734 10734 2786
rect 10786 2734 10800 2786
rect 10720 2626 10800 2734
rect 10720 2574 10734 2626
rect 10786 2574 10800 2626
rect 10720 2466 10800 2574
rect 10720 2414 10734 2466
rect 10786 2414 10800 2466
rect 10720 2306 10800 2414
rect 10720 2254 10734 2306
rect 10786 2254 10800 2306
rect 10720 2146 10800 2254
rect 10720 2094 10734 2146
rect 10786 2094 10800 2146
rect 10720 1986 10800 2094
rect 10720 1934 10734 1986
rect 10786 1934 10800 1986
rect 10720 1817 10800 1934
rect 10720 1783 10743 1817
rect 10777 1783 10800 1817
rect 10720 1666 10800 1783
rect 10720 1614 10734 1666
rect 10786 1614 10800 1666
rect 10720 1506 10800 1614
rect 10720 1454 10734 1506
rect 10786 1454 10800 1506
rect 10720 1346 10800 1454
rect 10720 1294 10734 1346
rect 10786 1294 10800 1346
rect 10720 1186 10800 1294
rect 10720 1134 10734 1186
rect 10786 1134 10800 1186
rect 10720 1026 10800 1134
rect 10720 974 10734 1026
rect 10786 974 10800 1026
rect 10720 857 10800 974
rect 10720 823 10743 857
rect 10777 823 10800 857
rect 10720 697 10800 823
rect 10720 663 10743 697
rect 10777 663 10800 697
rect 10720 546 10800 663
rect 10720 494 10734 546
rect 10786 494 10800 546
rect 10720 386 10800 494
rect 10720 334 10734 386
rect 10786 334 10800 386
rect 10720 226 10800 334
rect 10720 174 10734 226
rect 10786 174 10800 226
rect 10720 66 10800 174
rect 10720 14 10734 66
rect 10786 14 10800 66
rect 10720 0 10800 14
rect 10880 31417 10960 31440
rect 10880 31383 10903 31417
rect 10937 31383 10960 31417
rect 10880 31257 10960 31383
rect 10880 31223 10903 31257
rect 10937 31223 10960 31257
rect 10880 31097 10960 31223
rect 10880 31063 10903 31097
rect 10937 31063 10960 31097
rect 10880 30937 10960 31063
rect 10880 30903 10903 30937
rect 10937 30903 10960 30937
rect 10880 30777 10960 30903
rect 10880 30743 10903 30777
rect 10937 30743 10960 30777
rect 10880 30617 10960 30743
rect 10880 30583 10903 30617
rect 10937 30583 10960 30617
rect 10880 30457 10960 30583
rect 10880 30423 10903 30457
rect 10937 30423 10960 30457
rect 10880 30297 10960 30423
rect 10880 30263 10903 30297
rect 10937 30263 10960 30297
rect 10880 30137 10960 30263
rect 10880 30103 10903 30137
rect 10937 30103 10960 30137
rect 10880 29977 10960 30103
rect 10880 29943 10903 29977
rect 10937 29943 10960 29977
rect 10880 29817 10960 29943
rect 10880 29783 10903 29817
rect 10937 29783 10960 29817
rect 10880 29657 10960 29783
rect 10880 29623 10903 29657
rect 10937 29623 10960 29657
rect 10880 29497 10960 29623
rect 10880 29463 10903 29497
rect 10937 29463 10960 29497
rect 10880 29337 10960 29463
rect 10880 29303 10903 29337
rect 10937 29303 10960 29337
rect 10880 29177 10960 29303
rect 10880 29143 10903 29177
rect 10937 29143 10960 29177
rect 10880 29017 10960 29143
rect 10880 28983 10903 29017
rect 10937 28983 10960 29017
rect 10880 28857 10960 28983
rect 10880 28823 10903 28857
rect 10937 28823 10960 28857
rect 10880 28697 10960 28823
rect 10880 28663 10903 28697
rect 10937 28663 10960 28697
rect 10880 28537 10960 28663
rect 10880 28503 10903 28537
rect 10937 28503 10960 28537
rect 10880 28377 10960 28503
rect 10880 28343 10903 28377
rect 10937 28343 10960 28377
rect 10880 28217 10960 28343
rect 10880 28183 10903 28217
rect 10937 28183 10960 28217
rect 10880 28057 10960 28183
rect 10880 28023 10903 28057
rect 10937 28023 10960 28057
rect 10880 27897 10960 28023
rect 10880 27863 10903 27897
rect 10937 27863 10960 27897
rect 10880 27737 10960 27863
rect 10880 27703 10903 27737
rect 10937 27703 10960 27737
rect 10880 27577 10960 27703
rect 10880 27543 10903 27577
rect 10937 27543 10960 27577
rect 10880 27417 10960 27543
rect 10880 27383 10903 27417
rect 10937 27383 10960 27417
rect 10880 27257 10960 27383
rect 10880 27223 10903 27257
rect 10937 27223 10960 27257
rect 10880 27097 10960 27223
rect 10880 27063 10903 27097
rect 10937 27063 10960 27097
rect 10880 26937 10960 27063
rect 10880 26903 10903 26937
rect 10937 26903 10960 26937
rect 10880 26777 10960 26903
rect 10880 26743 10903 26777
rect 10937 26743 10960 26777
rect 10880 26617 10960 26743
rect 10880 26583 10903 26617
rect 10937 26583 10960 26617
rect 10880 26457 10960 26583
rect 10880 26423 10903 26457
rect 10937 26423 10960 26457
rect 10880 26297 10960 26423
rect 10880 26263 10903 26297
rect 10937 26263 10960 26297
rect 10880 26137 10960 26263
rect 10880 26103 10903 26137
rect 10937 26103 10960 26137
rect 10880 25977 10960 26103
rect 10880 25943 10903 25977
rect 10937 25943 10960 25977
rect 10880 25817 10960 25943
rect 10880 25783 10903 25817
rect 10937 25783 10960 25817
rect 10880 25657 10960 25783
rect 10880 25623 10903 25657
rect 10937 25623 10960 25657
rect 10880 25497 10960 25623
rect 10880 25463 10903 25497
rect 10937 25463 10960 25497
rect 10880 25337 10960 25463
rect 10880 25303 10903 25337
rect 10937 25303 10960 25337
rect 10880 25177 10960 25303
rect 10880 25143 10903 25177
rect 10937 25143 10960 25177
rect 10880 25017 10960 25143
rect 10880 24983 10903 25017
rect 10937 24983 10960 25017
rect 10880 24857 10960 24983
rect 10880 24823 10903 24857
rect 10937 24823 10960 24857
rect 10880 24697 10960 24823
rect 10880 24663 10903 24697
rect 10937 24663 10960 24697
rect 10880 24537 10960 24663
rect 10880 24503 10903 24537
rect 10937 24503 10960 24537
rect 10880 24377 10960 24503
rect 10880 24343 10903 24377
rect 10937 24343 10960 24377
rect 10880 24217 10960 24343
rect 10880 24183 10903 24217
rect 10937 24183 10960 24217
rect 10880 24057 10960 24183
rect 10880 24023 10903 24057
rect 10937 24023 10960 24057
rect 10880 23897 10960 24023
rect 10880 23863 10903 23897
rect 10937 23863 10960 23897
rect 10880 23737 10960 23863
rect 10880 23703 10903 23737
rect 10937 23703 10960 23737
rect 10880 23577 10960 23703
rect 10880 23543 10903 23577
rect 10937 23543 10960 23577
rect 10880 23417 10960 23543
rect 10880 23383 10903 23417
rect 10937 23383 10960 23417
rect 10880 23257 10960 23383
rect 10880 23223 10903 23257
rect 10937 23223 10960 23257
rect 10880 23097 10960 23223
rect 10880 23063 10903 23097
rect 10937 23063 10960 23097
rect 10880 22937 10960 23063
rect 10880 22903 10903 22937
rect 10937 22903 10960 22937
rect 10880 22777 10960 22903
rect 10880 22743 10903 22777
rect 10937 22743 10960 22777
rect 10880 22617 10960 22743
rect 10880 22583 10903 22617
rect 10937 22583 10960 22617
rect 10880 22457 10960 22583
rect 10880 22423 10903 22457
rect 10937 22423 10960 22457
rect 10880 22297 10960 22423
rect 10880 22263 10903 22297
rect 10937 22263 10960 22297
rect 10880 22137 10960 22263
rect 10880 22103 10903 22137
rect 10937 22103 10960 22137
rect 10880 21977 10960 22103
rect 10880 21943 10903 21977
rect 10937 21943 10960 21977
rect 10880 21817 10960 21943
rect 10880 21783 10903 21817
rect 10937 21783 10960 21817
rect 10880 21657 10960 21783
rect 10880 21623 10903 21657
rect 10937 21623 10960 21657
rect 10880 21497 10960 21623
rect 10880 21463 10903 21497
rect 10937 21463 10960 21497
rect 10880 21337 10960 21463
rect 10880 21303 10903 21337
rect 10937 21303 10960 21337
rect 10880 21177 10960 21303
rect 10880 21143 10903 21177
rect 10937 21143 10960 21177
rect 10880 21017 10960 21143
rect 10880 20983 10903 21017
rect 10937 20983 10960 21017
rect 10880 20857 10960 20983
rect 10880 20823 10903 20857
rect 10937 20823 10960 20857
rect 10880 20697 10960 20823
rect 10880 20663 10903 20697
rect 10937 20663 10960 20697
rect 10880 20537 10960 20663
rect 10880 20503 10903 20537
rect 10937 20503 10960 20537
rect 10880 20377 10960 20503
rect 10880 20343 10903 20377
rect 10937 20343 10960 20377
rect 10880 20217 10960 20343
rect 10880 20183 10903 20217
rect 10937 20183 10960 20217
rect 10880 20057 10960 20183
rect 10880 20023 10903 20057
rect 10937 20023 10960 20057
rect 10880 19897 10960 20023
rect 10880 19863 10903 19897
rect 10937 19863 10960 19897
rect 10880 19737 10960 19863
rect 10880 19703 10903 19737
rect 10937 19703 10960 19737
rect 10880 19577 10960 19703
rect 10880 19543 10903 19577
rect 10937 19543 10960 19577
rect 10880 19417 10960 19543
rect 10880 19383 10903 19417
rect 10937 19383 10960 19417
rect 10880 19257 10960 19383
rect 10880 19223 10903 19257
rect 10937 19223 10960 19257
rect 10880 19097 10960 19223
rect 10880 19063 10903 19097
rect 10937 19063 10960 19097
rect 10880 18937 10960 19063
rect 10880 18903 10903 18937
rect 10937 18903 10960 18937
rect 10880 18777 10960 18903
rect 10880 18743 10903 18777
rect 10937 18743 10960 18777
rect 10880 18617 10960 18743
rect 10880 18583 10903 18617
rect 10937 18583 10960 18617
rect 10880 18457 10960 18583
rect 10880 18423 10903 18457
rect 10937 18423 10960 18457
rect 10880 18297 10960 18423
rect 10880 18263 10903 18297
rect 10937 18263 10960 18297
rect 10880 18137 10960 18263
rect 10880 18103 10903 18137
rect 10937 18103 10960 18137
rect 10880 17977 10960 18103
rect 10880 17943 10903 17977
rect 10937 17943 10960 17977
rect 10880 17817 10960 17943
rect 10880 17783 10903 17817
rect 10937 17783 10960 17817
rect 10880 17657 10960 17783
rect 10880 17623 10903 17657
rect 10937 17623 10960 17657
rect 10880 17497 10960 17623
rect 10880 17463 10903 17497
rect 10937 17463 10960 17497
rect 10880 17337 10960 17463
rect 10880 17303 10903 17337
rect 10937 17303 10960 17337
rect 10880 17177 10960 17303
rect 10880 17143 10903 17177
rect 10937 17143 10960 17177
rect 10880 17017 10960 17143
rect 10880 16983 10903 17017
rect 10937 16983 10960 17017
rect 10880 16857 10960 16983
rect 10880 16823 10903 16857
rect 10937 16823 10960 16857
rect 10880 16697 10960 16823
rect 10880 16663 10903 16697
rect 10937 16663 10960 16697
rect 10880 16537 10960 16663
rect 10880 16503 10903 16537
rect 10937 16503 10960 16537
rect 10880 16377 10960 16503
rect 10880 16343 10903 16377
rect 10937 16343 10960 16377
rect 10880 16217 10960 16343
rect 10880 16183 10903 16217
rect 10937 16183 10960 16217
rect 10880 16057 10960 16183
rect 10880 16023 10903 16057
rect 10937 16023 10960 16057
rect 10880 15897 10960 16023
rect 10880 15863 10903 15897
rect 10937 15863 10960 15897
rect 10880 15737 10960 15863
rect 10880 15703 10903 15737
rect 10937 15703 10960 15737
rect 10880 15577 10960 15703
rect 10880 15543 10903 15577
rect 10937 15543 10960 15577
rect 10880 15417 10960 15543
rect 10880 15383 10903 15417
rect 10937 15383 10960 15417
rect 10880 15257 10960 15383
rect 10880 15223 10903 15257
rect 10937 15223 10960 15257
rect 10880 15097 10960 15223
rect 10880 15063 10903 15097
rect 10937 15063 10960 15097
rect 10880 14937 10960 15063
rect 10880 14903 10903 14937
rect 10937 14903 10960 14937
rect 10880 14777 10960 14903
rect 10880 14743 10903 14777
rect 10937 14743 10960 14777
rect 10880 14617 10960 14743
rect 10880 14583 10903 14617
rect 10937 14583 10960 14617
rect 10880 14457 10960 14583
rect 10880 14423 10903 14457
rect 10937 14423 10960 14457
rect 10880 14297 10960 14423
rect 10880 14263 10903 14297
rect 10937 14263 10960 14297
rect 10880 14137 10960 14263
rect 10880 14103 10903 14137
rect 10937 14103 10960 14137
rect 10880 13977 10960 14103
rect 10880 13943 10903 13977
rect 10937 13943 10960 13977
rect 10880 13817 10960 13943
rect 10880 13783 10903 13817
rect 10937 13783 10960 13817
rect 10880 13657 10960 13783
rect 10880 13623 10903 13657
rect 10937 13623 10960 13657
rect 10880 13497 10960 13623
rect 10880 13463 10903 13497
rect 10937 13463 10960 13497
rect 10880 13337 10960 13463
rect 10880 13303 10903 13337
rect 10937 13303 10960 13337
rect 10880 13177 10960 13303
rect 10880 13143 10903 13177
rect 10937 13143 10960 13177
rect 10880 13017 10960 13143
rect 10880 12983 10903 13017
rect 10937 12983 10960 13017
rect 10880 12857 10960 12983
rect 10880 12823 10903 12857
rect 10937 12823 10960 12857
rect 10880 12697 10960 12823
rect 10880 12663 10903 12697
rect 10937 12663 10960 12697
rect 10880 12537 10960 12663
rect 10880 12503 10903 12537
rect 10937 12503 10960 12537
rect 10880 12377 10960 12503
rect 10880 12343 10903 12377
rect 10937 12343 10960 12377
rect 10880 12217 10960 12343
rect 10880 12183 10903 12217
rect 10937 12183 10960 12217
rect 10880 12057 10960 12183
rect 10880 12023 10903 12057
rect 10937 12023 10960 12057
rect 10880 11897 10960 12023
rect 10880 11863 10903 11897
rect 10937 11863 10960 11897
rect 10880 11737 10960 11863
rect 10880 11703 10903 11737
rect 10937 11703 10960 11737
rect 10880 11577 10960 11703
rect 10880 11543 10903 11577
rect 10937 11543 10960 11577
rect 10880 11417 10960 11543
rect 10880 11383 10903 11417
rect 10937 11383 10960 11417
rect 10880 11257 10960 11383
rect 10880 11223 10903 11257
rect 10937 11223 10960 11257
rect 10880 11097 10960 11223
rect 10880 11063 10903 11097
rect 10937 11063 10960 11097
rect 10880 10937 10960 11063
rect 10880 10903 10903 10937
rect 10937 10903 10960 10937
rect 10880 10777 10960 10903
rect 10880 10743 10903 10777
rect 10937 10743 10960 10777
rect 10880 10617 10960 10743
rect 10880 10583 10903 10617
rect 10937 10583 10960 10617
rect 10880 10457 10960 10583
rect 10880 10423 10903 10457
rect 10937 10423 10960 10457
rect 10880 10297 10960 10423
rect 10880 10263 10903 10297
rect 10937 10263 10960 10297
rect 10880 10137 10960 10263
rect 10880 10103 10903 10137
rect 10937 10103 10960 10137
rect 10880 9977 10960 10103
rect 10880 9943 10903 9977
rect 10937 9943 10960 9977
rect 10880 9817 10960 9943
rect 10880 9783 10903 9817
rect 10937 9783 10960 9817
rect 10880 9657 10960 9783
rect 10880 9623 10903 9657
rect 10937 9623 10960 9657
rect 10880 9497 10960 9623
rect 10880 9463 10903 9497
rect 10937 9463 10960 9497
rect 10880 9337 10960 9463
rect 10880 9303 10903 9337
rect 10937 9303 10960 9337
rect 10880 9177 10960 9303
rect 10880 9143 10903 9177
rect 10937 9143 10960 9177
rect 10880 9017 10960 9143
rect 10880 8983 10903 9017
rect 10937 8983 10960 9017
rect 10880 8857 10960 8983
rect 10880 8823 10903 8857
rect 10937 8823 10960 8857
rect 10880 8697 10960 8823
rect 10880 8663 10903 8697
rect 10937 8663 10960 8697
rect 10880 8537 10960 8663
rect 10880 8503 10903 8537
rect 10937 8503 10960 8537
rect 10880 8377 10960 8503
rect 10880 8343 10903 8377
rect 10937 8343 10960 8377
rect 10880 8217 10960 8343
rect 10880 8183 10903 8217
rect 10937 8183 10960 8217
rect 10880 8057 10960 8183
rect 10880 8023 10903 8057
rect 10937 8023 10960 8057
rect 10880 7897 10960 8023
rect 10880 7863 10903 7897
rect 10937 7863 10960 7897
rect 10880 7737 10960 7863
rect 10880 7703 10903 7737
rect 10937 7703 10960 7737
rect 10880 7577 10960 7703
rect 10880 7543 10903 7577
rect 10937 7543 10960 7577
rect 10880 7417 10960 7543
rect 10880 7383 10903 7417
rect 10937 7383 10960 7417
rect 10880 7257 10960 7383
rect 10880 7223 10903 7257
rect 10937 7223 10960 7257
rect 10880 7097 10960 7223
rect 10880 7063 10903 7097
rect 10937 7063 10960 7097
rect 10880 6937 10960 7063
rect 10880 6903 10903 6937
rect 10937 6903 10960 6937
rect 10880 6777 10960 6903
rect 10880 6743 10903 6777
rect 10937 6743 10960 6777
rect 10880 6617 10960 6743
rect 10880 6583 10903 6617
rect 10937 6583 10960 6617
rect 10880 6457 10960 6583
rect 10880 6423 10903 6457
rect 10937 6423 10960 6457
rect 10880 6297 10960 6423
rect 10880 6263 10903 6297
rect 10937 6263 10960 6297
rect 10880 6137 10960 6263
rect 10880 6103 10903 6137
rect 10937 6103 10960 6137
rect 10880 5977 10960 6103
rect 10880 5943 10903 5977
rect 10937 5943 10960 5977
rect 10880 5817 10960 5943
rect 10880 5783 10903 5817
rect 10937 5783 10960 5817
rect 10880 5657 10960 5783
rect 10880 5623 10903 5657
rect 10937 5623 10960 5657
rect 10880 5497 10960 5623
rect 10880 5463 10903 5497
rect 10937 5463 10960 5497
rect 10880 5337 10960 5463
rect 10880 5303 10903 5337
rect 10937 5303 10960 5337
rect 10880 5177 10960 5303
rect 10880 5143 10903 5177
rect 10937 5143 10960 5177
rect 10880 5017 10960 5143
rect 10880 4983 10903 5017
rect 10937 4983 10960 5017
rect 10880 4857 10960 4983
rect 10880 4823 10903 4857
rect 10937 4823 10960 4857
rect 10880 4697 10960 4823
rect 10880 4663 10903 4697
rect 10937 4663 10960 4697
rect 10880 4537 10960 4663
rect 10880 4503 10903 4537
rect 10937 4503 10960 4537
rect 10880 4377 10960 4503
rect 10880 4343 10903 4377
rect 10937 4343 10960 4377
rect 10880 4217 10960 4343
rect 10880 4183 10903 4217
rect 10937 4183 10960 4217
rect 10880 4057 10960 4183
rect 10880 4023 10903 4057
rect 10937 4023 10960 4057
rect 10880 3897 10960 4023
rect 10880 3863 10903 3897
rect 10937 3863 10960 3897
rect 10880 3737 10960 3863
rect 10880 3703 10903 3737
rect 10937 3703 10960 3737
rect 10880 3577 10960 3703
rect 10880 3543 10903 3577
rect 10937 3543 10960 3577
rect 10880 3417 10960 3543
rect 10880 3383 10903 3417
rect 10937 3383 10960 3417
rect 10880 3257 10960 3383
rect 10880 3223 10903 3257
rect 10937 3223 10960 3257
rect 10880 3097 10960 3223
rect 10880 3063 10903 3097
rect 10937 3063 10960 3097
rect 10880 2937 10960 3063
rect 10880 2903 10903 2937
rect 10937 2903 10960 2937
rect 10880 2777 10960 2903
rect 10880 2743 10903 2777
rect 10937 2743 10960 2777
rect 10880 2617 10960 2743
rect 10880 2583 10903 2617
rect 10937 2583 10960 2617
rect 10880 2457 10960 2583
rect 10880 2423 10903 2457
rect 10937 2423 10960 2457
rect 10880 2297 10960 2423
rect 10880 2263 10903 2297
rect 10937 2263 10960 2297
rect 10880 2137 10960 2263
rect 10880 2103 10903 2137
rect 10937 2103 10960 2137
rect 10880 1977 10960 2103
rect 10880 1943 10903 1977
rect 10937 1943 10960 1977
rect 10880 1817 10960 1943
rect 10880 1783 10903 1817
rect 10937 1783 10960 1817
rect 10880 1657 10960 1783
rect 10880 1623 10903 1657
rect 10937 1623 10960 1657
rect 10880 1497 10960 1623
rect 10880 1463 10903 1497
rect 10937 1463 10960 1497
rect 10880 1337 10960 1463
rect 10880 1303 10903 1337
rect 10937 1303 10960 1337
rect 10880 1177 10960 1303
rect 10880 1143 10903 1177
rect 10937 1143 10960 1177
rect 10880 1017 10960 1143
rect 10880 983 10903 1017
rect 10937 983 10960 1017
rect 10880 857 10960 983
rect 10880 823 10903 857
rect 10937 823 10960 857
rect 10880 697 10960 823
rect 10880 663 10903 697
rect 10937 663 10960 697
rect 10880 537 10960 663
rect 10880 503 10903 537
rect 10937 503 10960 537
rect 10880 377 10960 503
rect 10880 343 10903 377
rect 10937 343 10960 377
rect 10880 217 10960 343
rect 10880 183 10903 217
rect 10937 183 10960 217
rect 10880 57 10960 183
rect 10880 23 10903 57
rect 10937 23 10960 57
rect 10880 0 10960 23
rect 11040 31426 11120 31440
rect 11040 31374 11054 31426
rect 11106 31374 11120 31426
rect 11040 31266 11120 31374
rect 11040 31214 11054 31266
rect 11106 31214 11120 31266
rect 11040 31106 11120 31214
rect 11040 31054 11054 31106
rect 11106 31054 11120 31106
rect 11040 30946 11120 31054
rect 11040 30894 11054 30946
rect 11106 30894 11120 30946
rect 11040 30786 11120 30894
rect 11040 30734 11054 30786
rect 11106 30734 11120 30786
rect 11040 30626 11120 30734
rect 11040 30574 11054 30626
rect 11106 30574 11120 30626
rect 11040 30466 11120 30574
rect 11040 30414 11054 30466
rect 11106 30414 11120 30466
rect 11040 30306 11120 30414
rect 11040 30254 11054 30306
rect 11106 30254 11120 30306
rect 11040 30137 11120 30254
rect 11040 30103 11063 30137
rect 11097 30103 11120 30137
rect 11040 29986 11120 30103
rect 11040 29934 11054 29986
rect 11106 29934 11120 29986
rect 11040 29826 11120 29934
rect 11040 29774 11054 29826
rect 11106 29774 11120 29826
rect 11040 29666 11120 29774
rect 11040 29614 11054 29666
rect 11106 29614 11120 29666
rect 11040 29506 11120 29614
rect 11040 29454 11054 29506
rect 11106 29454 11120 29506
rect 11040 29346 11120 29454
rect 11040 29294 11054 29346
rect 11106 29294 11120 29346
rect 11040 29186 11120 29294
rect 11040 29134 11054 29186
rect 11106 29134 11120 29186
rect 11040 29026 11120 29134
rect 11040 28974 11054 29026
rect 11106 28974 11120 29026
rect 11040 28866 11120 28974
rect 11040 28814 11054 28866
rect 11106 28814 11120 28866
rect 11040 28697 11120 28814
rect 11040 28663 11063 28697
rect 11097 28663 11120 28697
rect 11040 28537 11120 28663
rect 11040 28503 11063 28537
rect 11097 28503 11120 28537
rect 11040 28377 11120 28503
rect 11040 28343 11063 28377
rect 11097 28343 11120 28377
rect 11040 28217 11120 28343
rect 11040 28183 11063 28217
rect 11097 28183 11120 28217
rect 11040 28066 11120 28183
rect 11040 28014 11054 28066
rect 11106 28014 11120 28066
rect 11040 27906 11120 28014
rect 11040 27854 11054 27906
rect 11106 27854 11120 27906
rect 11040 27746 11120 27854
rect 11040 27694 11054 27746
rect 11106 27694 11120 27746
rect 11040 27586 11120 27694
rect 11040 27534 11054 27586
rect 11106 27534 11120 27586
rect 11040 27426 11120 27534
rect 11040 27374 11054 27426
rect 11106 27374 11120 27426
rect 11040 27266 11120 27374
rect 11040 27214 11054 27266
rect 11106 27214 11120 27266
rect 11040 27106 11120 27214
rect 11040 27054 11054 27106
rect 11106 27054 11120 27106
rect 11040 26946 11120 27054
rect 11040 26894 11054 26946
rect 11106 26894 11120 26946
rect 11040 26777 11120 26894
rect 11040 26743 11063 26777
rect 11097 26743 11120 26777
rect 11040 26617 11120 26743
rect 11040 26583 11063 26617
rect 11097 26583 11120 26617
rect 11040 26457 11120 26583
rect 11040 26423 11063 26457
rect 11097 26423 11120 26457
rect 11040 26297 11120 26423
rect 11040 26263 11063 26297
rect 11097 26263 11120 26297
rect 11040 26146 11120 26263
rect 11040 26094 11054 26146
rect 11106 26094 11120 26146
rect 11040 25986 11120 26094
rect 11040 25934 11054 25986
rect 11106 25934 11120 25986
rect 11040 25826 11120 25934
rect 11040 25774 11054 25826
rect 11106 25774 11120 25826
rect 11040 25666 11120 25774
rect 11040 25614 11054 25666
rect 11106 25614 11120 25666
rect 11040 25506 11120 25614
rect 11040 25454 11054 25506
rect 11106 25454 11120 25506
rect 11040 25346 11120 25454
rect 11040 25294 11054 25346
rect 11106 25294 11120 25346
rect 11040 25186 11120 25294
rect 11040 25134 11054 25186
rect 11106 25134 11120 25186
rect 11040 25026 11120 25134
rect 11040 24974 11054 25026
rect 11106 24974 11120 25026
rect 11040 24857 11120 24974
rect 11040 24823 11063 24857
rect 11097 24823 11120 24857
rect 11040 24706 11120 24823
rect 11040 24654 11054 24706
rect 11106 24654 11120 24706
rect 11040 24546 11120 24654
rect 11040 24494 11054 24546
rect 11106 24494 11120 24546
rect 11040 24386 11120 24494
rect 11040 24334 11054 24386
rect 11106 24334 11120 24386
rect 11040 24226 11120 24334
rect 11040 24174 11054 24226
rect 11106 24174 11120 24226
rect 11040 24066 11120 24174
rect 11040 24014 11054 24066
rect 11106 24014 11120 24066
rect 11040 23906 11120 24014
rect 11040 23854 11054 23906
rect 11106 23854 11120 23906
rect 11040 23746 11120 23854
rect 11040 23694 11054 23746
rect 11106 23694 11120 23746
rect 11040 23586 11120 23694
rect 11040 23534 11054 23586
rect 11106 23534 11120 23586
rect 11040 23426 11120 23534
rect 11040 23374 11054 23426
rect 11106 23374 11120 23426
rect 11040 23266 11120 23374
rect 11040 23214 11054 23266
rect 11106 23214 11120 23266
rect 11040 23106 11120 23214
rect 11040 23054 11054 23106
rect 11106 23054 11120 23106
rect 11040 22946 11120 23054
rect 11040 22894 11054 22946
rect 11106 22894 11120 22946
rect 11040 22786 11120 22894
rect 11040 22734 11054 22786
rect 11106 22734 11120 22786
rect 11040 22626 11120 22734
rect 11040 22574 11054 22626
rect 11106 22574 11120 22626
rect 11040 22466 11120 22574
rect 11040 22414 11054 22466
rect 11106 22414 11120 22466
rect 11040 22306 11120 22414
rect 11040 22254 11054 22306
rect 11106 22254 11120 22306
rect 11040 22146 11120 22254
rect 11040 22094 11054 22146
rect 11106 22094 11120 22146
rect 11040 21977 11120 22094
rect 11040 21943 11063 21977
rect 11097 21943 11120 21977
rect 11040 21826 11120 21943
rect 11040 21774 11054 21826
rect 11106 21774 11120 21826
rect 11040 21666 11120 21774
rect 11040 21614 11054 21666
rect 11106 21614 11120 21666
rect 11040 21506 11120 21614
rect 11040 21454 11054 21506
rect 11106 21454 11120 21506
rect 11040 21346 11120 21454
rect 11040 21294 11054 21346
rect 11106 21294 11120 21346
rect 11040 21186 11120 21294
rect 11040 21134 11054 21186
rect 11106 21134 11120 21186
rect 11040 21026 11120 21134
rect 11040 20974 11054 21026
rect 11106 20974 11120 21026
rect 11040 20866 11120 20974
rect 11040 20814 11054 20866
rect 11106 20814 11120 20866
rect 11040 20706 11120 20814
rect 11040 20654 11054 20706
rect 11106 20654 11120 20706
rect 11040 20537 11120 20654
rect 11040 20503 11063 20537
rect 11097 20503 11120 20537
rect 11040 20377 11120 20503
rect 11040 20343 11063 20377
rect 11097 20343 11120 20377
rect 11040 20217 11120 20343
rect 11040 20183 11063 20217
rect 11097 20183 11120 20217
rect 11040 20057 11120 20183
rect 11040 20023 11063 20057
rect 11097 20023 11120 20057
rect 11040 19906 11120 20023
rect 11040 19854 11054 19906
rect 11106 19854 11120 19906
rect 11040 19746 11120 19854
rect 11040 19694 11054 19746
rect 11106 19694 11120 19746
rect 11040 19586 11120 19694
rect 11040 19534 11054 19586
rect 11106 19534 11120 19586
rect 11040 19426 11120 19534
rect 11040 19374 11054 19426
rect 11106 19374 11120 19426
rect 11040 19266 11120 19374
rect 11040 19214 11054 19266
rect 11106 19214 11120 19266
rect 11040 19106 11120 19214
rect 11040 19054 11054 19106
rect 11106 19054 11120 19106
rect 11040 18946 11120 19054
rect 11040 18894 11054 18946
rect 11106 18894 11120 18946
rect 11040 18786 11120 18894
rect 11040 18734 11054 18786
rect 11106 18734 11120 18786
rect 11040 18617 11120 18734
rect 11040 18583 11063 18617
rect 11097 18583 11120 18617
rect 11040 18457 11120 18583
rect 11040 18423 11063 18457
rect 11097 18423 11120 18457
rect 11040 18297 11120 18423
rect 11040 18263 11063 18297
rect 11097 18263 11120 18297
rect 11040 18137 11120 18263
rect 11040 18103 11063 18137
rect 11097 18103 11120 18137
rect 11040 17986 11120 18103
rect 11040 17934 11054 17986
rect 11106 17934 11120 17986
rect 11040 17826 11120 17934
rect 11040 17774 11054 17826
rect 11106 17774 11120 17826
rect 11040 17666 11120 17774
rect 11040 17614 11054 17666
rect 11106 17614 11120 17666
rect 11040 17506 11120 17614
rect 11040 17454 11054 17506
rect 11106 17454 11120 17506
rect 11040 17346 11120 17454
rect 11040 17294 11054 17346
rect 11106 17294 11120 17346
rect 11040 17186 11120 17294
rect 11040 17134 11054 17186
rect 11106 17134 11120 17186
rect 11040 17026 11120 17134
rect 11040 16974 11054 17026
rect 11106 16974 11120 17026
rect 11040 16866 11120 16974
rect 11040 16814 11054 16866
rect 11106 16814 11120 16866
rect 11040 16697 11120 16814
rect 11040 16663 11063 16697
rect 11097 16663 11120 16697
rect 11040 16546 11120 16663
rect 11040 16494 11054 16546
rect 11106 16494 11120 16546
rect 11040 16386 11120 16494
rect 11040 16334 11054 16386
rect 11106 16334 11120 16386
rect 11040 16226 11120 16334
rect 11040 16174 11054 16226
rect 11106 16174 11120 16226
rect 11040 16066 11120 16174
rect 11040 16014 11054 16066
rect 11106 16014 11120 16066
rect 11040 15906 11120 16014
rect 11040 15854 11054 15906
rect 11106 15854 11120 15906
rect 11040 15746 11120 15854
rect 11040 15694 11054 15746
rect 11106 15694 11120 15746
rect 11040 15586 11120 15694
rect 11040 15534 11054 15586
rect 11106 15534 11120 15586
rect 11040 15426 11120 15534
rect 11040 15374 11054 15426
rect 11106 15374 11120 15426
rect 11040 15266 11120 15374
rect 11040 15214 11054 15266
rect 11106 15214 11120 15266
rect 11040 15106 11120 15214
rect 11040 15054 11054 15106
rect 11106 15054 11120 15106
rect 11040 14946 11120 15054
rect 11040 14894 11054 14946
rect 11106 14894 11120 14946
rect 11040 14786 11120 14894
rect 11040 14734 11054 14786
rect 11106 14734 11120 14786
rect 11040 14626 11120 14734
rect 11040 14574 11054 14626
rect 11106 14574 11120 14626
rect 11040 14466 11120 14574
rect 11040 14414 11054 14466
rect 11106 14414 11120 14466
rect 11040 14306 11120 14414
rect 11040 14254 11054 14306
rect 11106 14254 11120 14306
rect 11040 14146 11120 14254
rect 11040 14094 11054 14146
rect 11106 14094 11120 14146
rect 11040 13986 11120 14094
rect 11040 13934 11054 13986
rect 11106 13934 11120 13986
rect 11040 13817 11120 13934
rect 11040 13783 11063 13817
rect 11097 13783 11120 13817
rect 11040 13666 11120 13783
rect 11040 13614 11054 13666
rect 11106 13614 11120 13666
rect 11040 13506 11120 13614
rect 11040 13454 11054 13506
rect 11106 13454 11120 13506
rect 11040 13346 11120 13454
rect 11040 13294 11054 13346
rect 11106 13294 11120 13346
rect 11040 13186 11120 13294
rect 11040 13134 11054 13186
rect 11106 13134 11120 13186
rect 11040 13026 11120 13134
rect 11040 12974 11054 13026
rect 11106 12974 11120 13026
rect 11040 12866 11120 12974
rect 11040 12814 11054 12866
rect 11106 12814 11120 12866
rect 11040 12706 11120 12814
rect 11040 12654 11054 12706
rect 11106 12654 11120 12706
rect 11040 12546 11120 12654
rect 11040 12494 11054 12546
rect 11106 12494 11120 12546
rect 11040 12377 11120 12494
rect 11040 12343 11063 12377
rect 11097 12343 11120 12377
rect 11040 12217 11120 12343
rect 11040 12183 11063 12217
rect 11097 12183 11120 12217
rect 11040 12057 11120 12183
rect 11040 12023 11063 12057
rect 11097 12023 11120 12057
rect 11040 11897 11120 12023
rect 11040 11863 11063 11897
rect 11097 11863 11120 11897
rect 11040 11746 11120 11863
rect 11040 11694 11054 11746
rect 11106 11694 11120 11746
rect 11040 11586 11120 11694
rect 11040 11534 11054 11586
rect 11106 11534 11120 11586
rect 11040 11426 11120 11534
rect 11040 11374 11054 11426
rect 11106 11374 11120 11426
rect 11040 11266 11120 11374
rect 11040 11214 11054 11266
rect 11106 11214 11120 11266
rect 11040 11106 11120 11214
rect 11040 11054 11054 11106
rect 11106 11054 11120 11106
rect 11040 10946 11120 11054
rect 11040 10894 11054 10946
rect 11106 10894 11120 10946
rect 11040 10786 11120 10894
rect 11040 10734 11054 10786
rect 11106 10734 11120 10786
rect 11040 10626 11120 10734
rect 11040 10574 11054 10626
rect 11106 10574 11120 10626
rect 11040 10466 11120 10574
rect 11040 10414 11054 10466
rect 11106 10414 11120 10466
rect 11040 10306 11120 10414
rect 11040 10254 11054 10306
rect 11106 10254 11120 10306
rect 11040 10146 11120 10254
rect 11040 10094 11054 10146
rect 11106 10094 11120 10146
rect 11040 9986 11120 10094
rect 11040 9934 11054 9986
rect 11106 9934 11120 9986
rect 11040 9826 11120 9934
rect 11040 9774 11054 9826
rect 11106 9774 11120 9826
rect 11040 9657 11120 9774
rect 11040 9623 11063 9657
rect 11097 9623 11120 9657
rect 11040 9506 11120 9623
rect 11040 9454 11054 9506
rect 11106 9454 11120 9506
rect 11040 9346 11120 9454
rect 11040 9294 11054 9346
rect 11106 9294 11120 9346
rect 11040 9177 11120 9294
rect 11040 9143 11063 9177
rect 11097 9143 11120 9177
rect 11040 9026 11120 9143
rect 11040 8974 11054 9026
rect 11106 8974 11120 9026
rect 11040 8866 11120 8974
rect 11040 8814 11054 8866
rect 11106 8814 11120 8866
rect 11040 8706 11120 8814
rect 11040 8654 11054 8706
rect 11106 8654 11120 8706
rect 11040 8546 11120 8654
rect 11040 8494 11054 8546
rect 11106 8494 11120 8546
rect 11040 8386 11120 8494
rect 11040 8334 11054 8386
rect 11106 8334 11120 8386
rect 11040 8226 11120 8334
rect 11040 8174 11054 8226
rect 11106 8174 11120 8226
rect 11040 8066 11120 8174
rect 11040 8014 11054 8066
rect 11106 8014 11120 8066
rect 11040 7906 11120 8014
rect 11040 7854 11054 7906
rect 11106 7854 11120 7906
rect 11040 7746 11120 7854
rect 11040 7694 11054 7746
rect 11106 7694 11120 7746
rect 11040 7577 11120 7694
rect 11040 7543 11063 7577
rect 11097 7543 11120 7577
rect 11040 7426 11120 7543
rect 11040 7374 11054 7426
rect 11106 7374 11120 7426
rect 11040 7266 11120 7374
rect 11040 7214 11054 7266
rect 11106 7214 11120 7266
rect 11040 7097 11120 7214
rect 11040 7063 11063 7097
rect 11097 7063 11120 7097
rect 11040 6946 11120 7063
rect 11040 6894 11054 6946
rect 11106 6894 11120 6946
rect 11040 6786 11120 6894
rect 11040 6734 11054 6786
rect 11106 6734 11120 6786
rect 11040 6617 11120 6734
rect 11040 6583 11063 6617
rect 11097 6583 11120 6617
rect 11040 6466 11120 6583
rect 11040 6414 11054 6466
rect 11106 6414 11120 6466
rect 11040 6306 11120 6414
rect 11040 6254 11054 6306
rect 11106 6254 11120 6306
rect 11040 6146 11120 6254
rect 11040 6094 11054 6146
rect 11106 6094 11120 6146
rect 11040 5986 11120 6094
rect 11040 5934 11054 5986
rect 11106 5934 11120 5986
rect 11040 5826 11120 5934
rect 11040 5774 11054 5826
rect 11106 5774 11120 5826
rect 11040 5666 11120 5774
rect 11040 5614 11054 5666
rect 11106 5614 11120 5666
rect 11040 5506 11120 5614
rect 11040 5454 11054 5506
rect 11106 5454 11120 5506
rect 11040 5346 11120 5454
rect 11040 5294 11054 5346
rect 11106 5294 11120 5346
rect 11040 5186 11120 5294
rect 11040 5134 11054 5186
rect 11106 5134 11120 5186
rect 11040 5026 11120 5134
rect 11040 4974 11054 5026
rect 11106 4974 11120 5026
rect 11040 4866 11120 4974
rect 11040 4814 11054 4866
rect 11106 4814 11120 4866
rect 11040 4706 11120 4814
rect 11040 4654 11054 4706
rect 11106 4654 11120 4706
rect 11040 4546 11120 4654
rect 11040 4494 11054 4546
rect 11106 4494 11120 4546
rect 11040 4386 11120 4494
rect 11040 4334 11054 4386
rect 11106 4334 11120 4386
rect 11040 4226 11120 4334
rect 11040 4174 11054 4226
rect 11106 4174 11120 4226
rect 11040 4066 11120 4174
rect 11040 4014 11054 4066
rect 11106 4014 11120 4066
rect 11040 3906 11120 4014
rect 11040 3854 11054 3906
rect 11106 3854 11120 3906
rect 11040 3737 11120 3854
rect 11040 3703 11063 3737
rect 11097 3703 11120 3737
rect 11040 3577 11120 3703
rect 11040 3543 11063 3577
rect 11097 3543 11120 3577
rect 11040 3426 11120 3543
rect 11040 3374 11054 3426
rect 11106 3374 11120 3426
rect 11040 3266 11120 3374
rect 11040 3214 11054 3266
rect 11106 3214 11120 3266
rect 11040 3106 11120 3214
rect 11040 3054 11054 3106
rect 11106 3054 11120 3106
rect 11040 2946 11120 3054
rect 11040 2894 11054 2946
rect 11106 2894 11120 2946
rect 11040 2786 11120 2894
rect 11040 2734 11054 2786
rect 11106 2734 11120 2786
rect 11040 2626 11120 2734
rect 11040 2574 11054 2626
rect 11106 2574 11120 2626
rect 11040 2466 11120 2574
rect 11040 2414 11054 2466
rect 11106 2414 11120 2466
rect 11040 2306 11120 2414
rect 11040 2254 11054 2306
rect 11106 2254 11120 2306
rect 11040 2146 11120 2254
rect 11040 2094 11054 2146
rect 11106 2094 11120 2146
rect 11040 1986 11120 2094
rect 11040 1934 11054 1986
rect 11106 1934 11120 1986
rect 11040 1817 11120 1934
rect 11040 1783 11063 1817
rect 11097 1783 11120 1817
rect 11040 1666 11120 1783
rect 11040 1614 11054 1666
rect 11106 1614 11120 1666
rect 11040 1506 11120 1614
rect 11040 1454 11054 1506
rect 11106 1454 11120 1506
rect 11040 1346 11120 1454
rect 11040 1294 11054 1346
rect 11106 1294 11120 1346
rect 11040 1186 11120 1294
rect 11040 1134 11054 1186
rect 11106 1134 11120 1186
rect 11040 1026 11120 1134
rect 11040 974 11054 1026
rect 11106 974 11120 1026
rect 11040 857 11120 974
rect 11040 823 11063 857
rect 11097 823 11120 857
rect 11040 697 11120 823
rect 11040 663 11063 697
rect 11097 663 11120 697
rect 11040 546 11120 663
rect 11040 494 11054 546
rect 11106 494 11120 546
rect 11040 386 11120 494
rect 11040 334 11054 386
rect 11106 334 11120 386
rect 11040 226 11120 334
rect 11040 174 11054 226
rect 11106 174 11120 226
rect 11040 66 11120 174
rect 11040 14 11054 66
rect 11106 14 11120 66
rect 11040 0 11120 14
rect 11200 31417 11280 31440
rect 11200 31383 11223 31417
rect 11257 31383 11280 31417
rect 11200 31257 11280 31383
rect 11200 31223 11223 31257
rect 11257 31223 11280 31257
rect 11200 31097 11280 31223
rect 11200 31063 11223 31097
rect 11257 31063 11280 31097
rect 11200 30937 11280 31063
rect 11200 30903 11223 30937
rect 11257 30903 11280 30937
rect 11200 30777 11280 30903
rect 11200 30743 11223 30777
rect 11257 30743 11280 30777
rect 11200 30617 11280 30743
rect 11200 30583 11223 30617
rect 11257 30583 11280 30617
rect 11200 30457 11280 30583
rect 11200 30423 11223 30457
rect 11257 30423 11280 30457
rect 11200 30297 11280 30423
rect 11200 30263 11223 30297
rect 11257 30263 11280 30297
rect 11200 30137 11280 30263
rect 11200 30103 11223 30137
rect 11257 30103 11280 30137
rect 11200 29977 11280 30103
rect 11200 29943 11223 29977
rect 11257 29943 11280 29977
rect 11200 29817 11280 29943
rect 11200 29783 11223 29817
rect 11257 29783 11280 29817
rect 11200 29657 11280 29783
rect 11200 29623 11223 29657
rect 11257 29623 11280 29657
rect 11200 29497 11280 29623
rect 11200 29463 11223 29497
rect 11257 29463 11280 29497
rect 11200 29337 11280 29463
rect 11200 29303 11223 29337
rect 11257 29303 11280 29337
rect 11200 29177 11280 29303
rect 11200 29143 11223 29177
rect 11257 29143 11280 29177
rect 11200 29017 11280 29143
rect 11200 28983 11223 29017
rect 11257 28983 11280 29017
rect 11200 28857 11280 28983
rect 11200 28823 11223 28857
rect 11257 28823 11280 28857
rect 11200 28697 11280 28823
rect 11200 28663 11223 28697
rect 11257 28663 11280 28697
rect 11200 28537 11280 28663
rect 11200 28503 11223 28537
rect 11257 28503 11280 28537
rect 11200 28377 11280 28503
rect 11200 28343 11223 28377
rect 11257 28343 11280 28377
rect 11200 28217 11280 28343
rect 11200 28183 11223 28217
rect 11257 28183 11280 28217
rect 11200 28057 11280 28183
rect 11200 28023 11223 28057
rect 11257 28023 11280 28057
rect 11200 27897 11280 28023
rect 11200 27863 11223 27897
rect 11257 27863 11280 27897
rect 11200 27737 11280 27863
rect 11200 27703 11223 27737
rect 11257 27703 11280 27737
rect 11200 27577 11280 27703
rect 11200 27543 11223 27577
rect 11257 27543 11280 27577
rect 11200 27417 11280 27543
rect 11200 27383 11223 27417
rect 11257 27383 11280 27417
rect 11200 27257 11280 27383
rect 11200 27223 11223 27257
rect 11257 27223 11280 27257
rect 11200 27097 11280 27223
rect 11200 27063 11223 27097
rect 11257 27063 11280 27097
rect 11200 26937 11280 27063
rect 11200 26903 11223 26937
rect 11257 26903 11280 26937
rect 11200 26777 11280 26903
rect 11200 26743 11223 26777
rect 11257 26743 11280 26777
rect 11200 26617 11280 26743
rect 11200 26583 11223 26617
rect 11257 26583 11280 26617
rect 11200 26457 11280 26583
rect 11200 26423 11223 26457
rect 11257 26423 11280 26457
rect 11200 26297 11280 26423
rect 11200 26263 11223 26297
rect 11257 26263 11280 26297
rect 11200 26137 11280 26263
rect 11200 26103 11223 26137
rect 11257 26103 11280 26137
rect 11200 25977 11280 26103
rect 11200 25943 11223 25977
rect 11257 25943 11280 25977
rect 11200 25817 11280 25943
rect 11200 25783 11223 25817
rect 11257 25783 11280 25817
rect 11200 25657 11280 25783
rect 11200 25623 11223 25657
rect 11257 25623 11280 25657
rect 11200 25497 11280 25623
rect 11200 25463 11223 25497
rect 11257 25463 11280 25497
rect 11200 25337 11280 25463
rect 11200 25303 11223 25337
rect 11257 25303 11280 25337
rect 11200 25177 11280 25303
rect 11200 25143 11223 25177
rect 11257 25143 11280 25177
rect 11200 25017 11280 25143
rect 11200 24983 11223 25017
rect 11257 24983 11280 25017
rect 11200 24857 11280 24983
rect 11200 24823 11223 24857
rect 11257 24823 11280 24857
rect 11200 24697 11280 24823
rect 11200 24663 11223 24697
rect 11257 24663 11280 24697
rect 11200 24537 11280 24663
rect 11200 24503 11223 24537
rect 11257 24503 11280 24537
rect 11200 24377 11280 24503
rect 11200 24343 11223 24377
rect 11257 24343 11280 24377
rect 11200 24217 11280 24343
rect 11200 24183 11223 24217
rect 11257 24183 11280 24217
rect 11200 24057 11280 24183
rect 11200 24023 11223 24057
rect 11257 24023 11280 24057
rect 11200 23897 11280 24023
rect 11200 23863 11223 23897
rect 11257 23863 11280 23897
rect 11200 23737 11280 23863
rect 11200 23703 11223 23737
rect 11257 23703 11280 23737
rect 11200 23577 11280 23703
rect 11200 23543 11223 23577
rect 11257 23543 11280 23577
rect 11200 23417 11280 23543
rect 11200 23383 11223 23417
rect 11257 23383 11280 23417
rect 11200 23257 11280 23383
rect 11200 23223 11223 23257
rect 11257 23223 11280 23257
rect 11200 23097 11280 23223
rect 11200 23063 11223 23097
rect 11257 23063 11280 23097
rect 11200 22937 11280 23063
rect 11200 22903 11223 22937
rect 11257 22903 11280 22937
rect 11200 22777 11280 22903
rect 11200 22743 11223 22777
rect 11257 22743 11280 22777
rect 11200 22617 11280 22743
rect 11200 22583 11223 22617
rect 11257 22583 11280 22617
rect 11200 22457 11280 22583
rect 11200 22423 11223 22457
rect 11257 22423 11280 22457
rect 11200 22297 11280 22423
rect 11200 22263 11223 22297
rect 11257 22263 11280 22297
rect 11200 22137 11280 22263
rect 11200 22103 11223 22137
rect 11257 22103 11280 22137
rect 11200 21977 11280 22103
rect 11200 21943 11223 21977
rect 11257 21943 11280 21977
rect 11200 21817 11280 21943
rect 11200 21783 11223 21817
rect 11257 21783 11280 21817
rect 11200 21657 11280 21783
rect 11200 21623 11223 21657
rect 11257 21623 11280 21657
rect 11200 21497 11280 21623
rect 11200 21463 11223 21497
rect 11257 21463 11280 21497
rect 11200 21337 11280 21463
rect 11200 21303 11223 21337
rect 11257 21303 11280 21337
rect 11200 21177 11280 21303
rect 11200 21143 11223 21177
rect 11257 21143 11280 21177
rect 11200 21017 11280 21143
rect 11200 20983 11223 21017
rect 11257 20983 11280 21017
rect 11200 20857 11280 20983
rect 11200 20823 11223 20857
rect 11257 20823 11280 20857
rect 11200 20697 11280 20823
rect 11200 20663 11223 20697
rect 11257 20663 11280 20697
rect 11200 20537 11280 20663
rect 11200 20503 11223 20537
rect 11257 20503 11280 20537
rect 11200 20377 11280 20503
rect 11200 20343 11223 20377
rect 11257 20343 11280 20377
rect 11200 20217 11280 20343
rect 11200 20183 11223 20217
rect 11257 20183 11280 20217
rect 11200 20057 11280 20183
rect 11200 20023 11223 20057
rect 11257 20023 11280 20057
rect 11200 19897 11280 20023
rect 11200 19863 11223 19897
rect 11257 19863 11280 19897
rect 11200 19737 11280 19863
rect 11200 19703 11223 19737
rect 11257 19703 11280 19737
rect 11200 19577 11280 19703
rect 11200 19543 11223 19577
rect 11257 19543 11280 19577
rect 11200 19417 11280 19543
rect 11200 19383 11223 19417
rect 11257 19383 11280 19417
rect 11200 19257 11280 19383
rect 11200 19223 11223 19257
rect 11257 19223 11280 19257
rect 11200 19097 11280 19223
rect 11200 19063 11223 19097
rect 11257 19063 11280 19097
rect 11200 18937 11280 19063
rect 11200 18903 11223 18937
rect 11257 18903 11280 18937
rect 11200 18777 11280 18903
rect 11200 18743 11223 18777
rect 11257 18743 11280 18777
rect 11200 18617 11280 18743
rect 11200 18583 11223 18617
rect 11257 18583 11280 18617
rect 11200 18457 11280 18583
rect 11200 18423 11223 18457
rect 11257 18423 11280 18457
rect 11200 18297 11280 18423
rect 11200 18263 11223 18297
rect 11257 18263 11280 18297
rect 11200 18137 11280 18263
rect 11200 18103 11223 18137
rect 11257 18103 11280 18137
rect 11200 17977 11280 18103
rect 11200 17943 11223 17977
rect 11257 17943 11280 17977
rect 11200 17817 11280 17943
rect 11200 17783 11223 17817
rect 11257 17783 11280 17817
rect 11200 17657 11280 17783
rect 11200 17623 11223 17657
rect 11257 17623 11280 17657
rect 11200 17497 11280 17623
rect 11200 17463 11223 17497
rect 11257 17463 11280 17497
rect 11200 17337 11280 17463
rect 11200 17303 11223 17337
rect 11257 17303 11280 17337
rect 11200 17177 11280 17303
rect 11200 17143 11223 17177
rect 11257 17143 11280 17177
rect 11200 17017 11280 17143
rect 11200 16983 11223 17017
rect 11257 16983 11280 17017
rect 11200 16857 11280 16983
rect 11200 16823 11223 16857
rect 11257 16823 11280 16857
rect 11200 16697 11280 16823
rect 11200 16663 11223 16697
rect 11257 16663 11280 16697
rect 11200 16537 11280 16663
rect 11200 16503 11223 16537
rect 11257 16503 11280 16537
rect 11200 16377 11280 16503
rect 11200 16343 11223 16377
rect 11257 16343 11280 16377
rect 11200 16217 11280 16343
rect 11200 16183 11223 16217
rect 11257 16183 11280 16217
rect 11200 16057 11280 16183
rect 11200 16023 11223 16057
rect 11257 16023 11280 16057
rect 11200 15897 11280 16023
rect 11200 15863 11223 15897
rect 11257 15863 11280 15897
rect 11200 15737 11280 15863
rect 11200 15703 11223 15737
rect 11257 15703 11280 15737
rect 11200 15577 11280 15703
rect 11200 15543 11223 15577
rect 11257 15543 11280 15577
rect 11200 15417 11280 15543
rect 11200 15383 11223 15417
rect 11257 15383 11280 15417
rect 11200 15257 11280 15383
rect 11200 15223 11223 15257
rect 11257 15223 11280 15257
rect 11200 15097 11280 15223
rect 11200 15063 11223 15097
rect 11257 15063 11280 15097
rect 11200 14937 11280 15063
rect 11200 14903 11223 14937
rect 11257 14903 11280 14937
rect 11200 14777 11280 14903
rect 11200 14743 11223 14777
rect 11257 14743 11280 14777
rect 11200 14617 11280 14743
rect 11200 14583 11223 14617
rect 11257 14583 11280 14617
rect 11200 14457 11280 14583
rect 11200 14423 11223 14457
rect 11257 14423 11280 14457
rect 11200 14297 11280 14423
rect 11200 14263 11223 14297
rect 11257 14263 11280 14297
rect 11200 14137 11280 14263
rect 11200 14103 11223 14137
rect 11257 14103 11280 14137
rect 11200 13977 11280 14103
rect 11200 13943 11223 13977
rect 11257 13943 11280 13977
rect 11200 13817 11280 13943
rect 11200 13783 11223 13817
rect 11257 13783 11280 13817
rect 11200 13657 11280 13783
rect 11200 13623 11223 13657
rect 11257 13623 11280 13657
rect 11200 13497 11280 13623
rect 11200 13463 11223 13497
rect 11257 13463 11280 13497
rect 11200 13337 11280 13463
rect 11200 13303 11223 13337
rect 11257 13303 11280 13337
rect 11200 13177 11280 13303
rect 11200 13143 11223 13177
rect 11257 13143 11280 13177
rect 11200 13017 11280 13143
rect 11200 12983 11223 13017
rect 11257 12983 11280 13017
rect 11200 12857 11280 12983
rect 11200 12823 11223 12857
rect 11257 12823 11280 12857
rect 11200 12697 11280 12823
rect 11200 12663 11223 12697
rect 11257 12663 11280 12697
rect 11200 12537 11280 12663
rect 11200 12503 11223 12537
rect 11257 12503 11280 12537
rect 11200 12377 11280 12503
rect 11200 12343 11223 12377
rect 11257 12343 11280 12377
rect 11200 12217 11280 12343
rect 11200 12183 11223 12217
rect 11257 12183 11280 12217
rect 11200 12057 11280 12183
rect 11200 12023 11223 12057
rect 11257 12023 11280 12057
rect 11200 11897 11280 12023
rect 11200 11863 11223 11897
rect 11257 11863 11280 11897
rect 11200 11737 11280 11863
rect 11200 11703 11223 11737
rect 11257 11703 11280 11737
rect 11200 11577 11280 11703
rect 11200 11543 11223 11577
rect 11257 11543 11280 11577
rect 11200 11417 11280 11543
rect 11200 11383 11223 11417
rect 11257 11383 11280 11417
rect 11200 11257 11280 11383
rect 11200 11223 11223 11257
rect 11257 11223 11280 11257
rect 11200 11097 11280 11223
rect 11200 11063 11223 11097
rect 11257 11063 11280 11097
rect 11200 10937 11280 11063
rect 11200 10903 11223 10937
rect 11257 10903 11280 10937
rect 11200 10777 11280 10903
rect 11200 10743 11223 10777
rect 11257 10743 11280 10777
rect 11200 10617 11280 10743
rect 11200 10583 11223 10617
rect 11257 10583 11280 10617
rect 11200 10457 11280 10583
rect 11200 10423 11223 10457
rect 11257 10423 11280 10457
rect 11200 10297 11280 10423
rect 11200 10263 11223 10297
rect 11257 10263 11280 10297
rect 11200 10137 11280 10263
rect 11200 10103 11223 10137
rect 11257 10103 11280 10137
rect 11200 9977 11280 10103
rect 11200 9943 11223 9977
rect 11257 9943 11280 9977
rect 11200 9817 11280 9943
rect 11200 9783 11223 9817
rect 11257 9783 11280 9817
rect 11200 9657 11280 9783
rect 11200 9623 11223 9657
rect 11257 9623 11280 9657
rect 11200 9497 11280 9623
rect 11200 9463 11223 9497
rect 11257 9463 11280 9497
rect 11200 9337 11280 9463
rect 11200 9303 11223 9337
rect 11257 9303 11280 9337
rect 11200 9177 11280 9303
rect 11200 9143 11223 9177
rect 11257 9143 11280 9177
rect 11200 9017 11280 9143
rect 11200 8983 11223 9017
rect 11257 8983 11280 9017
rect 11200 8857 11280 8983
rect 11200 8823 11223 8857
rect 11257 8823 11280 8857
rect 11200 8697 11280 8823
rect 11200 8663 11223 8697
rect 11257 8663 11280 8697
rect 11200 8537 11280 8663
rect 11200 8503 11223 8537
rect 11257 8503 11280 8537
rect 11200 8377 11280 8503
rect 11200 8343 11223 8377
rect 11257 8343 11280 8377
rect 11200 8217 11280 8343
rect 11200 8183 11223 8217
rect 11257 8183 11280 8217
rect 11200 8057 11280 8183
rect 11200 8023 11223 8057
rect 11257 8023 11280 8057
rect 11200 7897 11280 8023
rect 11200 7863 11223 7897
rect 11257 7863 11280 7897
rect 11200 7737 11280 7863
rect 11200 7703 11223 7737
rect 11257 7703 11280 7737
rect 11200 7577 11280 7703
rect 11200 7543 11223 7577
rect 11257 7543 11280 7577
rect 11200 7417 11280 7543
rect 11200 7383 11223 7417
rect 11257 7383 11280 7417
rect 11200 7257 11280 7383
rect 11200 7223 11223 7257
rect 11257 7223 11280 7257
rect 11200 7097 11280 7223
rect 11200 7063 11223 7097
rect 11257 7063 11280 7097
rect 11200 6937 11280 7063
rect 11200 6903 11223 6937
rect 11257 6903 11280 6937
rect 11200 6777 11280 6903
rect 11200 6743 11223 6777
rect 11257 6743 11280 6777
rect 11200 6617 11280 6743
rect 11200 6583 11223 6617
rect 11257 6583 11280 6617
rect 11200 6457 11280 6583
rect 11200 6423 11223 6457
rect 11257 6423 11280 6457
rect 11200 6297 11280 6423
rect 11200 6263 11223 6297
rect 11257 6263 11280 6297
rect 11200 6137 11280 6263
rect 11200 6103 11223 6137
rect 11257 6103 11280 6137
rect 11200 5977 11280 6103
rect 11200 5943 11223 5977
rect 11257 5943 11280 5977
rect 11200 5817 11280 5943
rect 11200 5783 11223 5817
rect 11257 5783 11280 5817
rect 11200 5657 11280 5783
rect 11200 5623 11223 5657
rect 11257 5623 11280 5657
rect 11200 5497 11280 5623
rect 11200 5463 11223 5497
rect 11257 5463 11280 5497
rect 11200 5337 11280 5463
rect 11200 5303 11223 5337
rect 11257 5303 11280 5337
rect 11200 5177 11280 5303
rect 11200 5143 11223 5177
rect 11257 5143 11280 5177
rect 11200 5017 11280 5143
rect 11200 4983 11223 5017
rect 11257 4983 11280 5017
rect 11200 4857 11280 4983
rect 11200 4823 11223 4857
rect 11257 4823 11280 4857
rect 11200 4697 11280 4823
rect 11200 4663 11223 4697
rect 11257 4663 11280 4697
rect 11200 4537 11280 4663
rect 11200 4503 11223 4537
rect 11257 4503 11280 4537
rect 11200 4377 11280 4503
rect 11200 4343 11223 4377
rect 11257 4343 11280 4377
rect 11200 4217 11280 4343
rect 11200 4183 11223 4217
rect 11257 4183 11280 4217
rect 11200 4057 11280 4183
rect 11200 4023 11223 4057
rect 11257 4023 11280 4057
rect 11200 3897 11280 4023
rect 11200 3863 11223 3897
rect 11257 3863 11280 3897
rect 11200 3737 11280 3863
rect 11200 3703 11223 3737
rect 11257 3703 11280 3737
rect 11200 3577 11280 3703
rect 11200 3543 11223 3577
rect 11257 3543 11280 3577
rect 11200 3417 11280 3543
rect 11200 3383 11223 3417
rect 11257 3383 11280 3417
rect 11200 3257 11280 3383
rect 11200 3223 11223 3257
rect 11257 3223 11280 3257
rect 11200 3097 11280 3223
rect 11200 3063 11223 3097
rect 11257 3063 11280 3097
rect 11200 2937 11280 3063
rect 11200 2903 11223 2937
rect 11257 2903 11280 2937
rect 11200 2777 11280 2903
rect 11200 2743 11223 2777
rect 11257 2743 11280 2777
rect 11200 2617 11280 2743
rect 11200 2583 11223 2617
rect 11257 2583 11280 2617
rect 11200 2457 11280 2583
rect 11200 2423 11223 2457
rect 11257 2423 11280 2457
rect 11200 2297 11280 2423
rect 11200 2263 11223 2297
rect 11257 2263 11280 2297
rect 11200 2137 11280 2263
rect 11200 2103 11223 2137
rect 11257 2103 11280 2137
rect 11200 1977 11280 2103
rect 11200 1943 11223 1977
rect 11257 1943 11280 1977
rect 11200 1817 11280 1943
rect 11200 1783 11223 1817
rect 11257 1783 11280 1817
rect 11200 1657 11280 1783
rect 11200 1623 11223 1657
rect 11257 1623 11280 1657
rect 11200 1497 11280 1623
rect 11200 1463 11223 1497
rect 11257 1463 11280 1497
rect 11200 1337 11280 1463
rect 11200 1303 11223 1337
rect 11257 1303 11280 1337
rect 11200 1177 11280 1303
rect 11200 1143 11223 1177
rect 11257 1143 11280 1177
rect 11200 1017 11280 1143
rect 11200 983 11223 1017
rect 11257 983 11280 1017
rect 11200 857 11280 983
rect 11200 823 11223 857
rect 11257 823 11280 857
rect 11200 697 11280 823
rect 11200 663 11223 697
rect 11257 663 11280 697
rect 11200 537 11280 663
rect 11200 503 11223 537
rect 11257 503 11280 537
rect 11200 377 11280 503
rect 11200 343 11223 377
rect 11257 343 11280 377
rect 11200 217 11280 343
rect 11200 183 11223 217
rect 11257 183 11280 217
rect 11200 57 11280 183
rect 11200 23 11223 57
rect 11257 23 11280 57
rect 11200 0 11280 23
rect 11360 31426 11440 31440
rect 11360 31374 11374 31426
rect 11426 31374 11440 31426
rect 11360 31266 11440 31374
rect 11360 31214 11374 31266
rect 11426 31214 11440 31266
rect 11360 31106 11440 31214
rect 11360 31054 11374 31106
rect 11426 31054 11440 31106
rect 11360 30946 11440 31054
rect 11360 30894 11374 30946
rect 11426 30894 11440 30946
rect 11360 30786 11440 30894
rect 11360 30734 11374 30786
rect 11426 30734 11440 30786
rect 11360 30626 11440 30734
rect 11360 30574 11374 30626
rect 11426 30574 11440 30626
rect 11360 30466 11440 30574
rect 11360 30414 11374 30466
rect 11426 30414 11440 30466
rect 11360 30306 11440 30414
rect 11360 30254 11374 30306
rect 11426 30254 11440 30306
rect 11360 30137 11440 30254
rect 11360 30103 11383 30137
rect 11417 30103 11440 30137
rect 11360 29986 11440 30103
rect 11360 29934 11374 29986
rect 11426 29934 11440 29986
rect 11360 29826 11440 29934
rect 11360 29774 11374 29826
rect 11426 29774 11440 29826
rect 11360 29666 11440 29774
rect 11360 29614 11374 29666
rect 11426 29614 11440 29666
rect 11360 29506 11440 29614
rect 11360 29454 11374 29506
rect 11426 29454 11440 29506
rect 11360 29346 11440 29454
rect 11360 29294 11374 29346
rect 11426 29294 11440 29346
rect 11360 29186 11440 29294
rect 11360 29134 11374 29186
rect 11426 29134 11440 29186
rect 11360 29026 11440 29134
rect 11360 28974 11374 29026
rect 11426 28974 11440 29026
rect 11360 28866 11440 28974
rect 11360 28814 11374 28866
rect 11426 28814 11440 28866
rect 11360 28697 11440 28814
rect 11360 28663 11383 28697
rect 11417 28663 11440 28697
rect 11360 28537 11440 28663
rect 11360 28503 11383 28537
rect 11417 28503 11440 28537
rect 11360 28377 11440 28503
rect 11360 28343 11383 28377
rect 11417 28343 11440 28377
rect 11360 28217 11440 28343
rect 11360 28183 11383 28217
rect 11417 28183 11440 28217
rect 11360 28066 11440 28183
rect 11360 28014 11374 28066
rect 11426 28014 11440 28066
rect 11360 27906 11440 28014
rect 11360 27854 11374 27906
rect 11426 27854 11440 27906
rect 11360 27746 11440 27854
rect 11360 27694 11374 27746
rect 11426 27694 11440 27746
rect 11360 27586 11440 27694
rect 11360 27534 11374 27586
rect 11426 27534 11440 27586
rect 11360 27426 11440 27534
rect 11360 27374 11374 27426
rect 11426 27374 11440 27426
rect 11360 27266 11440 27374
rect 11360 27214 11374 27266
rect 11426 27214 11440 27266
rect 11360 27106 11440 27214
rect 11360 27054 11374 27106
rect 11426 27054 11440 27106
rect 11360 26946 11440 27054
rect 11360 26894 11374 26946
rect 11426 26894 11440 26946
rect 11360 26777 11440 26894
rect 11360 26743 11383 26777
rect 11417 26743 11440 26777
rect 11360 26617 11440 26743
rect 11360 26583 11383 26617
rect 11417 26583 11440 26617
rect 11360 26457 11440 26583
rect 11360 26423 11383 26457
rect 11417 26423 11440 26457
rect 11360 26297 11440 26423
rect 11360 26263 11383 26297
rect 11417 26263 11440 26297
rect 11360 26146 11440 26263
rect 11360 26094 11374 26146
rect 11426 26094 11440 26146
rect 11360 25986 11440 26094
rect 11360 25934 11374 25986
rect 11426 25934 11440 25986
rect 11360 25826 11440 25934
rect 11360 25774 11374 25826
rect 11426 25774 11440 25826
rect 11360 25666 11440 25774
rect 11360 25614 11374 25666
rect 11426 25614 11440 25666
rect 11360 25506 11440 25614
rect 11360 25454 11374 25506
rect 11426 25454 11440 25506
rect 11360 25346 11440 25454
rect 11360 25294 11374 25346
rect 11426 25294 11440 25346
rect 11360 25186 11440 25294
rect 11360 25134 11374 25186
rect 11426 25134 11440 25186
rect 11360 25026 11440 25134
rect 11360 24974 11374 25026
rect 11426 24974 11440 25026
rect 11360 24857 11440 24974
rect 11360 24823 11383 24857
rect 11417 24823 11440 24857
rect 11360 24706 11440 24823
rect 11360 24654 11374 24706
rect 11426 24654 11440 24706
rect 11360 24546 11440 24654
rect 11360 24494 11374 24546
rect 11426 24494 11440 24546
rect 11360 24386 11440 24494
rect 11360 24334 11374 24386
rect 11426 24334 11440 24386
rect 11360 24226 11440 24334
rect 11360 24174 11374 24226
rect 11426 24174 11440 24226
rect 11360 24066 11440 24174
rect 11360 24014 11374 24066
rect 11426 24014 11440 24066
rect 11360 23906 11440 24014
rect 11360 23854 11374 23906
rect 11426 23854 11440 23906
rect 11360 23746 11440 23854
rect 11360 23694 11374 23746
rect 11426 23694 11440 23746
rect 11360 23586 11440 23694
rect 11360 23534 11374 23586
rect 11426 23534 11440 23586
rect 11360 23426 11440 23534
rect 11360 23374 11374 23426
rect 11426 23374 11440 23426
rect 11360 23266 11440 23374
rect 11360 23214 11374 23266
rect 11426 23214 11440 23266
rect 11360 23106 11440 23214
rect 11360 23054 11374 23106
rect 11426 23054 11440 23106
rect 11360 22946 11440 23054
rect 11360 22894 11374 22946
rect 11426 22894 11440 22946
rect 11360 22786 11440 22894
rect 11360 22734 11374 22786
rect 11426 22734 11440 22786
rect 11360 22626 11440 22734
rect 11360 22574 11374 22626
rect 11426 22574 11440 22626
rect 11360 22466 11440 22574
rect 11360 22414 11374 22466
rect 11426 22414 11440 22466
rect 11360 22306 11440 22414
rect 11360 22254 11374 22306
rect 11426 22254 11440 22306
rect 11360 22146 11440 22254
rect 11360 22094 11374 22146
rect 11426 22094 11440 22146
rect 11360 21977 11440 22094
rect 11360 21943 11383 21977
rect 11417 21943 11440 21977
rect 11360 21826 11440 21943
rect 11360 21774 11374 21826
rect 11426 21774 11440 21826
rect 11360 21666 11440 21774
rect 11360 21614 11374 21666
rect 11426 21614 11440 21666
rect 11360 21506 11440 21614
rect 11360 21454 11374 21506
rect 11426 21454 11440 21506
rect 11360 21346 11440 21454
rect 11360 21294 11374 21346
rect 11426 21294 11440 21346
rect 11360 21186 11440 21294
rect 11360 21134 11374 21186
rect 11426 21134 11440 21186
rect 11360 21026 11440 21134
rect 11360 20974 11374 21026
rect 11426 20974 11440 21026
rect 11360 20866 11440 20974
rect 11360 20814 11374 20866
rect 11426 20814 11440 20866
rect 11360 20706 11440 20814
rect 11360 20654 11374 20706
rect 11426 20654 11440 20706
rect 11360 20537 11440 20654
rect 11360 20503 11383 20537
rect 11417 20503 11440 20537
rect 11360 20377 11440 20503
rect 11360 20343 11383 20377
rect 11417 20343 11440 20377
rect 11360 20217 11440 20343
rect 11360 20183 11383 20217
rect 11417 20183 11440 20217
rect 11360 20057 11440 20183
rect 11360 20023 11383 20057
rect 11417 20023 11440 20057
rect 11360 19906 11440 20023
rect 11360 19854 11374 19906
rect 11426 19854 11440 19906
rect 11360 19746 11440 19854
rect 11360 19694 11374 19746
rect 11426 19694 11440 19746
rect 11360 19586 11440 19694
rect 11360 19534 11374 19586
rect 11426 19534 11440 19586
rect 11360 19426 11440 19534
rect 11360 19374 11374 19426
rect 11426 19374 11440 19426
rect 11360 19266 11440 19374
rect 11360 19214 11374 19266
rect 11426 19214 11440 19266
rect 11360 19106 11440 19214
rect 11360 19054 11374 19106
rect 11426 19054 11440 19106
rect 11360 18946 11440 19054
rect 11360 18894 11374 18946
rect 11426 18894 11440 18946
rect 11360 18786 11440 18894
rect 11360 18734 11374 18786
rect 11426 18734 11440 18786
rect 11360 18617 11440 18734
rect 11360 18583 11383 18617
rect 11417 18583 11440 18617
rect 11360 18457 11440 18583
rect 11360 18423 11383 18457
rect 11417 18423 11440 18457
rect 11360 18297 11440 18423
rect 11360 18263 11383 18297
rect 11417 18263 11440 18297
rect 11360 18137 11440 18263
rect 11360 18103 11383 18137
rect 11417 18103 11440 18137
rect 11360 17986 11440 18103
rect 11360 17934 11374 17986
rect 11426 17934 11440 17986
rect 11360 17826 11440 17934
rect 11360 17774 11374 17826
rect 11426 17774 11440 17826
rect 11360 17666 11440 17774
rect 11360 17614 11374 17666
rect 11426 17614 11440 17666
rect 11360 17506 11440 17614
rect 11360 17454 11374 17506
rect 11426 17454 11440 17506
rect 11360 17346 11440 17454
rect 11360 17294 11374 17346
rect 11426 17294 11440 17346
rect 11360 17186 11440 17294
rect 11360 17134 11374 17186
rect 11426 17134 11440 17186
rect 11360 17026 11440 17134
rect 11360 16974 11374 17026
rect 11426 16974 11440 17026
rect 11360 16866 11440 16974
rect 11360 16814 11374 16866
rect 11426 16814 11440 16866
rect 11360 16697 11440 16814
rect 11360 16663 11383 16697
rect 11417 16663 11440 16697
rect 11360 16546 11440 16663
rect 11360 16494 11374 16546
rect 11426 16494 11440 16546
rect 11360 16386 11440 16494
rect 11360 16334 11374 16386
rect 11426 16334 11440 16386
rect 11360 16226 11440 16334
rect 11360 16174 11374 16226
rect 11426 16174 11440 16226
rect 11360 16066 11440 16174
rect 11360 16014 11374 16066
rect 11426 16014 11440 16066
rect 11360 15906 11440 16014
rect 11360 15854 11374 15906
rect 11426 15854 11440 15906
rect 11360 15746 11440 15854
rect 11360 15694 11374 15746
rect 11426 15694 11440 15746
rect 11360 15586 11440 15694
rect 11360 15534 11374 15586
rect 11426 15534 11440 15586
rect 11360 15426 11440 15534
rect 11360 15374 11374 15426
rect 11426 15374 11440 15426
rect 11360 15266 11440 15374
rect 11360 15214 11374 15266
rect 11426 15214 11440 15266
rect 11360 15106 11440 15214
rect 11360 15054 11374 15106
rect 11426 15054 11440 15106
rect 11360 14946 11440 15054
rect 11360 14894 11374 14946
rect 11426 14894 11440 14946
rect 11360 14786 11440 14894
rect 11360 14734 11374 14786
rect 11426 14734 11440 14786
rect 11360 14626 11440 14734
rect 11360 14574 11374 14626
rect 11426 14574 11440 14626
rect 11360 14466 11440 14574
rect 11360 14414 11374 14466
rect 11426 14414 11440 14466
rect 11360 14306 11440 14414
rect 11360 14254 11374 14306
rect 11426 14254 11440 14306
rect 11360 14146 11440 14254
rect 11360 14094 11374 14146
rect 11426 14094 11440 14146
rect 11360 13986 11440 14094
rect 11360 13934 11374 13986
rect 11426 13934 11440 13986
rect 11360 13817 11440 13934
rect 11360 13783 11383 13817
rect 11417 13783 11440 13817
rect 11360 13666 11440 13783
rect 11360 13614 11374 13666
rect 11426 13614 11440 13666
rect 11360 13506 11440 13614
rect 11360 13454 11374 13506
rect 11426 13454 11440 13506
rect 11360 13346 11440 13454
rect 11360 13294 11374 13346
rect 11426 13294 11440 13346
rect 11360 13186 11440 13294
rect 11360 13134 11374 13186
rect 11426 13134 11440 13186
rect 11360 13026 11440 13134
rect 11360 12974 11374 13026
rect 11426 12974 11440 13026
rect 11360 12866 11440 12974
rect 11360 12814 11374 12866
rect 11426 12814 11440 12866
rect 11360 12706 11440 12814
rect 11360 12654 11374 12706
rect 11426 12654 11440 12706
rect 11360 12546 11440 12654
rect 11360 12494 11374 12546
rect 11426 12494 11440 12546
rect 11360 12377 11440 12494
rect 11360 12343 11383 12377
rect 11417 12343 11440 12377
rect 11360 12217 11440 12343
rect 11360 12183 11383 12217
rect 11417 12183 11440 12217
rect 11360 12057 11440 12183
rect 11360 12023 11383 12057
rect 11417 12023 11440 12057
rect 11360 11897 11440 12023
rect 11360 11863 11383 11897
rect 11417 11863 11440 11897
rect 11360 11746 11440 11863
rect 11360 11694 11374 11746
rect 11426 11694 11440 11746
rect 11360 11586 11440 11694
rect 11360 11534 11374 11586
rect 11426 11534 11440 11586
rect 11360 11426 11440 11534
rect 11360 11374 11374 11426
rect 11426 11374 11440 11426
rect 11360 11266 11440 11374
rect 11360 11214 11374 11266
rect 11426 11214 11440 11266
rect 11360 11106 11440 11214
rect 11360 11054 11374 11106
rect 11426 11054 11440 11106
rect 11360 10946 11440 11054
rect 11360 10894 11374 10946
rect 11426 10894 11440 10946
rect 11360 10786 11440 10894
rect 11360 10734 11374 10786
rect 11426 10734 11440 10786
rect 11360 10626 11440 10734
rect 11360 10574 11374 10626
rect 11426 10574 11440 10626
rect 11360 10466 11440 10574
rect 11360 10414 11374 10466
rect 11426 10414 11440 10466
rect 11360 10306 11440 10414
rect 11360 10254 11374 10306
rect 11426 10254 11440 10306
rect 11360 10146 11440 10254
rect 11360 10094 11374 10146
rect 11426 10094 11440 10146
rect 11360 9986 11440 10094
rect 11360 9934 11374 9986
rect 11426 9934 11440 9986
rect 11360 9826 11440 9934
rect 11360 9774 11374 9826
rect 11426 9774 11440 9826
rect 11360 9657 11440 9774
rect 11360 9623 11383 9657
rect 11417 9623 11440 9657
rect 11360 9506 11440 9623
rect 11360 9454 11374 9506
rect 11426 9454 11440 9506
rect 11360 9346 11440 9454
rect 11360 9294 11374 9346
rect 11426 9294 11440 9346
rect 11360 9177 11440 9294
rect 11360 9143 11383 9177
rect 11417 9143 11440 9177
rect 11360 9026 11440 9143
rect 11360 8974 11374 9026
rect 11426 8974 11440 9026
rect 11360 8866 11440 8974
rect 11360 8814 11374 8866
rect 11426 8814 11440 8866
rect 11360 8706 11440 8814
rect 11360 8654 11374 8706
rect 11426 8654 11440 8706
rect 11360 8546 11440 8654
rect 11360 8494 11374 8546
rect 11426 8494 11440 8546
rect 11360 8386 11440 8494
rect 11360 8334 11374 8386
rect 11426 8334 11440 8386
rect 11360 8226 11440 8334
rect 11360 8174 11374 8226
rect 11426 8174 11440 8226
rect 11360 8066 11440 8174
rect 11360 8014 11374 8066
rect 11426 8014 11440 8066
rect 11360 7906 11440 8014
rect 11360 7854 11374 7906
rect 11426 7854 11440 7906
rect 11360 7746 11440 7854
rect 11360 7694 11374 7746
rect 11426 7694 11440 7746
rect 11360 7577 11440 7694
rect 11360 7543 11383 7577
rect 11417 7543 11440 7577
rect 11360 7426 11440 7543
rect 11360 7374 11374 7426
rect 11426 7374 11440 7426
rect 11360 7266 11440 7374
rect 11360 7214 11374 7266
rect 11426 7214 11440 7266
rect 11360 7097 11440 7214
rect 11360 7063 11383 7097
rect 11417 7063 11440 7097
rect 11360 6946 11440 7063
rect 11360 6894 11374 6946
rect 11426 6894 11440 6946
rect 11360 6786 11440 6894
rect 11360 6734 11374 6786
rect 11426 6734 11440 6786
rect 11360 6617 11440 6734
rect 11360 6583 11383 6617
rect 11417 6583 11440 6617
rect 11360 6466 11440 6583
rect 11360 6414 11374 6466
rect 11426 6414 11440 6466
rect 11360 6306 11440 6414
rect 11360 6254 11374 6306
rect 11426 6254 11440 6306
rect 11360 6146 11440 6254
rect 11360 6094 11374 6146
rect 11426 6094 11440 6146
rect 11360 5986 11440 6094
rect 11360 5934 11374 5986
rect 11426 5934 11440 5986
rect 11360 5826 11440 5934
rect 11360 5774 11374 5826
rect 11426 5774 11440 5826
rect 11360 5666 11440 5774
rect 11360 5614 11374 5666
rect 11426 5614 11440 5666
rect 11360 5506 11440 5614
rect 11360 5454 11374 5506
rect 11426 5454 11440 5506
rect 11360 5346 11440 5454
rect 11360 5294 11374 5346
rect 11426 5294 11440 5346
rect 11360 5186 11440 5294
rect 11360 5134 11374 5186
rect 11426 5134 11440 5186
rect 11360 5026 11440 5134
rect 11360 4974 11374 5026
rect 11426 4974 11440 5026
rect 11360 4866 11440 4974
rect 11360 4814 11374 4866
rect 11426 4814 11440 4866
rect 11360 4706 11440 4814
rect 11360 4654 11374 4706
rect 11426 4654 11440 4706
rect 11360 4546 11440 4654
rect 11360 4494 11374 4546
rect 11426 4494 11440 4546
rect 11360 4386 11440 4494
rect 11360 4334 11374 4386
rect 11426 4334 11440 4386
rect 11360 4226 11440 4334
rect 11360 4174 11374 4226
rect 11426 4174 11440 4226
rect 11360 4066 11440 4174
rect 11360 4014 11374 4066
rect 11426 4014 11440 4066
rect 11360 3906 11440 4014
rect 11360 3854 11374 3906
rect 11426 3854 11440 3906
rect 11360 3737 11440 3854
rect 11360 3703 11383 3737
rect 11417 3703 11440 3737
rect 11360 3577 11440 3703
rect 11360 3543 11383 3577
rect 11417 3543 11440 3577
rect 11360 3426 11440 3543
rect 11360 3374 11374 3426
rect 11426 3374 11440 3426
rect 11360 3266 11440 3374
rect 11360 3214 11374 3266
rect 11426 3214 11440 3266
rect 11360 3106 11440 3214
rect 11360 3054 11374 3106
rect 11426 3054 11440 3106
rect 11360 2946 11440 3054
rect 11360 2894 11374 2946
rect 11426 2894 11440 2946
rect 11360 2786 11440 2894
rect 11360 2734 11374 2786
rect 11426 2734 11440 2786
rect 11360 2626 11440 2734
rect 11360 2574 11374 2626
rect 11426 2574 11440 2626
rect 11360 2466 11440 2574
rect 11360 2414 11374 2466
rect 11426 2414 11440 2466
rect 11360 2306 11440 2414
rect 11360 2254 11374 2306
rect 11426 2254 11440 2306
rect 11360 2146 11440 2254
rect 11360 2094 11374 2146
rect 11426 2094 11440 2146
rect 11360 1986 11440 2094
rect 11360 1934 11374 1986
rect 11426 1934 11440 1986
rect 11360 1817 11440 1934
rect 11360 1783 11383 1817
rect 11417 1783 11440 1817
rect 11360 1666 11440 1783
rect 11360 1614 11374 1666
rect 11426 1614 11440 1666
rect 11360 1506 11440 1614
rect 11360 1454 11374 1506
rect 11426 1454 11440 1506
rect 11360 1346 11440 1454
rect 11360 1294 11374 1346
rect 11426 1294 11440 1346
rect 11360 1186 11440 1294
rect 11360 1134 11374 1186
rect 11426 1134 11440 1186
rect 11360 1026 11440 1134
rect 11360 974 11374 1026
rect 11426 974 11440 1026
rect 11360 857 11440 974
rect 11360 823 11383 857
rect 11417 823 11440 857
rect 11360 697 11440 823
rect 11360 663 11383 697
rect 11417 663 11440 697
rect 11360 546 11440 663
rect 11360 494 11374 546
rect 11426 494 11440 546
rect 11360 386 11440 494
rect 11360 334 11374 386
rect 11426 334 11440 386
rect 11360 226 11440 334
rect 11360 174 11374 226
rect 11426 174 11440 226
rect 11360 66 11440 174
rect 11360 14 11374 66
rect 11426 14 11440 66
rect 11360 0 11440 14
rect 11520 31426 11600 31440
rect 11520 31374 11534 31426
rect 11586 31374 11600 31426
rect 11520 31266 11600 31374
rect 11520 31214 11534 31266
rect 11586 31214 11600 31266
rect 11520 31106 11600 31214
rect 11520 31054 11534 31106
rect 11586 31054 11600 31106
rect 11520 30946 11600 31054
rect 11520 30894 11534 30946
rect 11586 30894 11600 30946
rect 11520 30786 11600 30894
rect 11520 30734 11534 30786
rect 11586 30734 11600 30786
rect 11520 30626 11600 30734
rect 11520 30574 11534 30626
rect 11586 30574 11600 30626
rect 11520 30466 11600 30574
rect 11520 30414 11534 30466
rect 11586 30414 11600 30466
rect 11520 30306 11600 30414
rect 11520 30254 11534 30306
rect 11586 30254 11600 30306
rect 11520 30137 11600 30254
rect 11520 30103 11543 30137
rect 11577 30103 11600 30137
rect 11520 29986 11600 30103
rect 11520 29934 11534 29986
rect 11586 29934 11600 29986
rect 11520 29826 11600 29934
rect 11520 29774 11534 29826
rect 11586 29774 11600 29826
rect 11520 29666 11600 29774
rect 11520 29614 11534 29666
rect 11586 29614 11600 29666
rect 11520 29506 11600 29614
rect 11520 29454 11534 29506
rect 11586 29454 11600 29506
rect 11520 29346 11600 29454
rect 11520 29294 11534 29346
rect 11586 29294 11600 29346
rect 11520 29186 11600 29294
rect 11520 29134 11534 29186
rect 11586 29134 11600 29186
rect 11520 29026 11600 29134
rect 11520 28974 11534 29026
rect 11586 28974 11600 29026
rect 11520 28866 11600 28974
rect 11520 28814 11534 28866
rect 11586 28814 11600 28866
rect 11520 28697 11600 28814
rect 11520 28663 11543 28697
rect 11577 28663 11600 28697
rect 11520 28537 11600 28663
rect 11520 28503 11543 28537
rect 11577 28503 11600 28537
rect 11520 28377 11600 28503
rect 11520 28343 11543 28377
rect 11577 28343 11600 28377
rect 11520 28217 11600 28343
rect 11520 28183 11543 28217
rect 11577 28183 11600 28217
rect 11520 28066 11600 28183
rect 11520 28014 11534 28066
rect 11586 28014 11600 28066
rect 11520 27906 11600 28014
rect 11520 27854 11534 27906
rect 11586 27854 11600 27906
rect 11520 27746 11600 27854
rect 11520 27694 11534 27746
rect 11586 27694 11600 27746
rect 11520 27586 11600 27694
rect 11520 27534 11534 27586
rect 11586 27534 11600 27586
rect 11520 27426 11600 27534
rect 11520 27374 11534 27426
rect 11586 27374 11600 27426
rect 11520 27266 11600 27374
rect 11520 27214 11534 27266
rect 11586 27214 11600 27266
rect 11520 27106 11600 27214
rect 11520 27054 11534 27106
rect 11586 27054 11600 27106
rect 11520 26946 11600 27054
rect 11520 26894 11534 26946
rect 11586 26894 11600 26946
rect 11520 26777 11600 26894
rect 11520 26743 11543 26777
rect 11577 26743 11600 26777
rect 11520 26617 11600 26743
rect 11520 26583 11543 26617
rect 11577 26583 11600 26617
rect 11520 26457 11600 26583
rect 11520 26423 11543 26457
rect 11577 26423 11600 26457
rect 11520 26297 11600 26423
rect 11520 26263 11543 26297
rect 11577 26263 11600 26297
rect 11520 26146 11600 26263
rect 11520 26094 11534 26146
rect 11586 26094 11600 26146
rect 11520 25986 11600 26094
rect 11520 25934 11534 25986
rect 11586 25934 11600 25986
rect 11520 25826 11600 25934
rect 11520 25774 11534 25826
rect 11586 25774 11600 25826
rect 11520 25666 11600 25774
rect 11520 25614 11534 25666
rect 11586 25614 11600 25666
rect 11520 25506 11600 25614
rect 11520 25454 11534 25506
rect 11586 25454 11600 25506
rect 11520 25346 11600 25454
rect 11520 25294 11534 25346
rect 11586 25294 11600 25346
rect 11520 25186 11600 25294
rect 11520 25134 11534 25186
rect 11586 25134 11600 25186
rect 11520 25026 11600 25134
rect 11520 24974 11534 25026
rect 11586 24974 11600 25026
rect 11520 24857 11600 24974
rect 11520 24823 11543 24857
rect 11577 24823 11600 24857
rect 11520 24706 11600 24823
rect 11520 24654 11534 24706
rect 11586 24654 11600 24706
rect 11520 24546 11600 24654
rect 11520 24494 11534 24546
rect 11586 24494 11600 24546
rect 11520 24386 11600 24494
rect 11520 24334 11534 24386
rect 11586 24334 11600 24386
rect 11520 24226 11600 24334
rect 11520 24174 11534 24226
rect 11586 24174 11600 24226
rect 11520 24066 11600 24174
rect 11520 24014 11534 24066
rect 11586 24014 11600 24066
rect 11520 23906 11600 24014
rect 11520 23854 11534 23906
rect 11586 23854 11600 23906
rect 11520 23746 11600 23854
rect 11520 23694 11534 23746
rect 11586 23694 11600 23746
rect 11520 23586 11600 23694
rect 11520 23534 11534 23586
rect 11586 23534 11600 23586
rect 11520 23426 11600 23534
rect 11520 23374 11534 23426
rect 11586 23374 11600 23426
rect 11520 23266 11600 23374
rect 11520 23214 11534 23266
rect 11586 23214 11600 23266
rect 11520 23106 11600 23214
rect 11520 23054 11534 23106
rect 11586 23054 11600 23106
rect 11520 22946 11600 23054
rect 11520 22894 11534 22946
rect 11586 22894 11600 22946
rect 11520 22786 11600 22894
rect 11520 22734 11534 22786
rect 11586 22734 11600 22786
rect 11520 22626 11600 22734
rect 11520 22574 11534 22626
rect 11586 22574 11600 22626
rect 11520 22466 11600 22574
rect 11520 22414 11534 22466
rect 11586 22414 11600 22466
rect 11520 22306 11600 22414
rect 11520 22254 11534 22306
rect 11586 22254 11600 22306
rect 11520 22146 11600 22254
rect 11520 22094 11534 22146
rect 11586 22094 11600 22146
rect 11520 21977 11600 22094
rect 11520 21943 11543 21977
rect 11577 21943 11600 21977
rect 11520 21826 11600 21943
rect 11520 21774 11534 21826
rect 11586 21774 11600 21826
rect 11520 21666 11600 21774
rect 11520 21614 11534 21666
rect 11586 21614 11600 21666
rect 11520 21506 11600 21614
rect 11520 21454 11534 21506
rect 11586 21454 11600 21506
rect 11520 21346 11600 21454
rect 11520 21294 11534 21346
rect 11586 21294 11600 21346
rect 11520 21186 11600 21294
rect 11520 21134 11534 21186
rect 11586 21134 11600 21186
rect 11520 21026 11600 21134
rect 11520 20974 11534 21026
rect 11586 20974 11600 21026
rect 11520 20866 11600 20974
rect 11520 20814 11534 20866
rect 11586 20814 11600 20866
rect 11520 20706 11600 20814
rect 11520 20654 11534 20706
rect 11586 20654 11600 20706
rect 11520 20537 11600 20654
rect 11520 20503 11543 20537
rect 11577 20503 11600 20537
rect 11520 20377 11600 20503
rect 11520 20343 11543 20377
rect 11577 20343 11600 20377
rect 11520 20217 11600 20343
rect 11520 20183 11543 20217
rect 11577 20183 11600 20217
rect 11520 20057 11600 20183
rect 11520 20023 11543 20057
rect 11577 20023 11600 20057
rect 11520 19906 11600 20023
rect 11520 19854 11534 19906
rect 11586 19854 11600 19906
rect 11520 19746 11600 19854
rect 11520 19694 11534 19746
rect 11586 19694 11600 19746
rect 11520 19586 11600 19694
rect 11520 19534 11534 19586
rect 11586 19534 11600 19586
rect 11520 19426 11600 19534
rect 11520 19374 11534 19426
rect 11586 19374 11600 19426
rect 11520 19266 11600 19374
rect 11520 19214 11534 19266
rect 11586 19214 11600 19266
rect 11520 19106 11600 19214
rect 11520 19054 11534 19106
rect 11586 19054 11600 19106
rect 11520 18946 11600 19054
rect 11520 18894 11534 18946
rect 11586 18894 11600 18946
rect 11520 18786 11600 18894
rect 11520 18734 11534 18786
rect 11586 18734 11600 18786
rect 11520 18617 11600 18734
rect 11520 18583 11543 18617
rect 11577 18583 11600 18617
rect 11520 18457 11600 18583
rect 11520 18423 11543 18457
rect 11577 18423 11600 18457
rect 11520 18297 11600 18423
rect 11520 18263 11543 18297
rect 11577 18263 11600 18297
rect 11520 18137 11600 18263
rect 11520 18103 11543 18137
rect 11577 18103 11600 18137
rect 11520 17986 11600 18103
rect 11520 17934 11534 17986
rect 11586 17934 11600 17986
rect 11520 17826 11600 17934
rect 11520 17774 11534 17826
rect 11586 17774 11600 17826
rect 11520 17666 11600 17774
rect 11520 17614 11534 17666
rect 11586 17614 11600 17666
rect 11520 17506 11600 17614
rect 11520 17454 11534 17506
rect 11586 17454 11600 17506
rect 11520 17346 11600 17454
rect 11520 17294 11534 17346
rect 11586 17294 11600 17346
rect 11520 17186 11600 17294
rect 11520 17134 11534 17186
rect 11586 17134 11600 17186
rect 11520 17026 11600 17134
rect 11520 16974 11534 17026
rect 11586 16974 11600 17026
rect 11520 16866 11600 16974
rect 11520 16814 11534 16866
rect 11586 16814 11600 16866
rect 11520 16697 11600 16814
rect 11520 16663 11543 16697
rect 11577 16663 11600 16697
rect 11520 16546 11600 16663
rect 11520 16494 11534 16546
rect 11586 16494 11600 16546
rect 11520 16386 11600 16494
rect 11520 16334 11534 16386
rect 11586 16334 11600 16386
rect 11520 16226 11600 16334
rect 11520 16174 11534 16226
rect 11586 16174 11600 16226
rect 11520 16066 11600 16174
rect 11520 16014 11534 16066
rect 11586 16014 11600 16066
rect 11520 15906 11600 16014
rect 11520 15854 11534 15906
rect 11586 15854 11600 15906
rect 11520 15746 11600 15854
rect 11520 15694 11534 15746
rect 11586 15694 11600 15746
rect 11520 15586 11600 15694
rect 11520 15534 11534 15586
rect 11586 15534 11600 15586
rect 11520 15426 11600 15534
rect 11520 15374 11534 15426
rect 11586 15374 11600 15426
rect 11520 15266 11600 15374
rect 11520 15214 11534 15266
rect 11586 15214 11600 15266
rect 11520 15106 11600 15214
rect 11520 15054 11534 15106
rect 11586 15054 11600 15106
rect 11520 14946 11600 15054
rect 11520 14894 11534 14946
rect 11586 14894 11600 14946
rect 11520 14786 11600 14894
rect 11520 14734 11534 14786
rect 11586 14734 11600 14786
rect 11520 14626 11600 14734
rect 11520 14574 11534 14626
rect 11586 14574 11600 14626
rect 11520 14466 11600 14574
rect 11520 14414 11534 14466
rect 11586 14414 11600 14466
rect 11520 14306 11600 14414
rect 11520 14254 11534 14306
rect 11586 14254 11600 14306
rect 11520 14146 11600 14254
rect 11520 14094 11534 14146
rect 11586 14094 11600 14146
rect 11520 13986 11600 14094
rect 11520 13934 11534 13986
rect 11586 13934 11600 13986
rect 11520 13817 11600 13934
rect 11520 13783 11543 13817
rect 11577 13783 11600 13817
rect 11520 13666 11600 13783
rect 11520 13614 11534 13666
rect 11586 13614 11600 13666
rect 11520 13506 11600 13614
rect 11520 13454 11534 13506
rect 11586 13454 11600 13506
rect 11520 13346 11600 13454
rect 11520 13294 11534 13346
rect 11586 13294 11600 13346
rect 11520 13186 11600 13294
rect 11520 13134 11534 13186
rect 11586 13134 11600 13186
rect 11520 13026 11600 13134
rect 11520 12974 11534 13026
rect 11586 12974 11600 13026
rect 11520 12866 11600 12974
rect 11520 12814 11534 12866
rect 11586 12814 11600 12866
rect 11520 12706 11600 12814
rect 11520 12654 11534 12706
rect 11586 12654 11600 12706
rect 11520 12546 11600 12654
rect 11520 12494 11534 12546
rect 11586 12494 11600 12546
rect 11520 12377 11600 12494
rect 11520 12343 11543 12377
rect 11577 12343 11600 12377
rect 11520 12217 11600 12343
rect 11520 12183 11543 12217
rect 11577 12183 11600 12217
rect 11520 12057 11600 12183
rect 11520 12023 11543 12057
rect 11577 12023 11600 12057
rect 11520 11897 11600 12023
rect 11520 11863 11543 11897
rect 11577 11863 11600 11897
rect 11520 11746 11600 11863
rect 11520 11694 11534 11746
rect 11586 11694 11600 11746
rect 11520 11586 11600 11694
rect 11520 11534 11534 11586
rect 11586 11534 11600 11586
rect 11520 11426 11600 11534
rect 11520 11374 11534 11426
rect 11586 11374 11600 11426
rect 11520 11266 11600 11374
rect 11520 11214 11534 11266
rect 11586 11214 11600 11266
rect 11520 11106 11600 11214
rect 11520 11054 11534 11106
rect 11586 11054 11600 11106
rect 11520 10946 11600 11054
rect 11520 10894 11534 10946
rect 11586 10894 11600 10946
rect 11520 10786 11600 10894
rect 11520 10734 11534 10786
rect 11586 10734 11600 10786
rect 11520 10626 11600 10734
rect 11520 10574 11534 10626
rect 11586 10574 11600 10626
rect 11520 10466 11600 10574
rect 11520 10414 11534 10466
rect 11586 10414 11600 10466
rect 11520 10306 11600 10414
rect 11520 10254 11534 10306
rect 11586 10254 11600 10306
rect 11520 10146 11600 10254
rect 11520 10094 11534 10146
rect 11586 10094 11600 10146
rect 11520 9986 11600 10094
rect 11520 9934 11534 9986
rect 11586 9934 11600 9986
rect 11520 9826 11600 9934
rect 11520 9774 11534 9826
rect 11586 9774 11600 9826
rect 11520 9657 11600 9774
rect 11520 9623 11543 9657
rect 11577 9623 11600 9657
rect 11520 9506 11600 9623
rect 11520 9454 11534 9506
rect 11586 9454 11600 9506
rect 11520 9346 11600 9454
rect 11520 9294 11534 9346
rect 11586 9294 11600 9346
rect 11520 9177 11600 9294
rect 11520 9143 11543 9177
rect 11577 9143 11600 9177
rect 11520 9026 11600 9143
rect 11520 8974 11534 9026
rect 11586 8974 11600 9026
rect 11520 8866 11600 8974
rect 11520 8814 11534 8866
rect 11586 8814 11600 8866
rect 11520 8706 11600 8814
rect 11520 8654 11534 8706
rect 11586 8654 11600 8706
rect 11520 8546 11600 8654
rect 11520 8494 11534 8546
rect 11586 8494 11600 8546
rect 11520 8386 11600 8494
rect 11520 8334 11534 8386
rect 11586 8334 11600 8386
rect 11520 8226 11600 8334
rect 11520 8174 11534 8226
rect 11586 8174 11600 8226
rect 11520 8066 11600 8174
rect 11520 8014 11534 8066
rect 11586 8014 11600 8066
rect 11520 7906 11600 8014
rect 11520 7854 11534 7906
rect 11586 7854 11600 7906
rect 11520 7746 11600 7854
rect 11520 7694 11534 7746
rect 11586 7694 11600 7746
rect 11520 7577 11600 7694
rect 11520 7543 11543 7577
rect 11577 7543 11600 7577
rect 11520 7426 11600 7543
rect 11520 7374 11534 7426
rect 11586 7374 11600 7426
rect 11520 7266 11600 7374
rect 11520 7214 11534 7266
rect 11586 7214 11600 7266
rect 11520 7097 11600 7214
rect 11520 7063 11543 7097
rect 11577 7063 11600 7097
rect 11520 6946 11600 7063
rect 11520 6894 11534 6946
rect 11586 6894 11600 6946
rect 11520 6786 11600 6894
rect 11520 6734 11534 6786
rect 11586 6734 11600 6786
rect 11520 6617 11600 6734
rect 11520 6583 11543 6617
rect 11577 6583 11600 6617
rect 11520 6466 11600 6583
rect 11520 6414 11534 6466
rect 11586 6414 11600 6466
rect 11520 6306 11600 6414
rect 11520 6254 11534 6306
rect 11586 6254 11600 6306
rect 11520 6146 11600 6254
rect 11520 6094 11534 6146
rect 11586 6094 11600 6146
rect 11520 5986 11600 6094
rect 11520 5934 11534 5986
rect 11586 5934 11600 5986
rect 11520 5826 11600 5934
rect 11520 5774 11534 5826
rect 11586 5774 11600 5826
rect 11520 5666 11600 5774
rect 11520 5614 11534 5666
rect 11586 5614 11600 5666
rect 11520 5506 11600 5614
rect 11520 5454 11534 5506
rect 11586 5454 11600 5506
rect 11520 5346 11600 5454
rect 11520 5294 11534 5346
rect 11586 5294 11600 5346
rect 11520 5186 11600 5294
rect 11520 5134 11534 5186
rect 11586 5134 11600 5186
rect 11520 5026 11600 5134
rect 11520 4974 11534 5026
rect 11586 4974 11600 5026
rect 11520 4866 11600 4974
rect 11520 4814 11534 4866
rect 11586 4814 11600 4866
rect 11520 4706 11600 4814
rect 11520 4654 11534 4706
rect 11586 4654 11600 4706
rect 11520 4546 11600 4654
rect 11520 4494 11534 4546
rect 11586 4494 11600 4546
rect 11520 4386 11600 4494
rect 11520 4334 11534 4386
rect 11586 4334 11600 4386
rect 11520 4226 11600 4334
rect 11520 4174 11534 4226
rect 11586 4174 11600 4226
rect 11520 4066 11600 4174
rect 11520 4014 11534 4066
rect 11586 4014 11600 4066
rect 11520 3906 11600 4014
rect 11520 3854 11534 3906
rect 11586 3854 11600 3906
rect 11520 3737 11600 3854
rect 11520 3703 11543 3737
rect 11577 3703 11600 3737
rect 11520 3577 11600 3703
rect 11520 3543 11543 3577
rect 11577 3543 11600 3577
rect 11520 3426 11600 3543
rect 11520 3374 11534 3426
rect 11586 3374 11600 3426
rect 11520 3266 11600 3374
rect 11520 3214 11534 3266
rect 11586 3214 11600 3266
rect 11520 3106 11600 3214
rect 11520 3054 11534 3106
rect 11586 3054 11600 3106
rect 11520 2946 11600 3054
rect 11520 2894 11534 2946
rect 11586 2894 11600 2946
rect 11520 2786 11600 2894
rect 11520 2734 11534 2786
rect 11586 2734 11600 2786
rect 11520 2626 11600 2734
rect 11520 2574 11534 2626
rect 11586 2574 11600 2626
rect 11520 2466 11600 2574
rect 11520 2414 11534 2466
rect 11586 2414 11600 2466
rect 11520 2306 11600 2414
rect 11520 2254 11534 2306
rect 11586 2254 11600 2306
rect 11520 2146 11600 2254
rect 11520 2094 11534 2146
rect 11586 2094 11600 2146
rect 11520 1986 11600 2094
rect 11520 1934 11534 1986
rect 11586 1934 11600 1986
rect 11520 1817 11600 1934
rect 11520 1783 11543 1817
rect 11577 1783 11600 1817
rect 11520 1666 11600 1783
rect 11520 1614 11534 1666
rect 11586 1614 11600 1666
rect 11520 1506 11600 1614
rect 11520 1454 11534 1506
rect 11586 1454 11600 1506
rect 11520 1346 11600 1454
rect 11520 1294 11534 1346
rect 11586 1294 11600 1346
rect 11520 1186 11600 1294
rect 11520 1134 11534 1186
rect 11586 1134 11600 1186
rect 11520 1026 11600 1134
rect 11520 974 11534 1026
rect 11586 974 11600 1026
rect 11520 857 11600 974
rect 11520 823 11543 857
rect 11577 823 11600 857
rect 11520 697 11600 823
rect 11520 663 11543 697
rect 11577 663 11600 697
rect 11520 546 11600 663
rect 11520 494 11534 546
rect 11586 494 11600 546
rect 11520 386 11600 494
rect 11520 334 11534 386
rect 11586 334 11600 386
rect 11520 226 11600 334
rect 11520 174 11534 226
rect 11586 174 11600 226
rect 11520 66 11600 174
rect 11520 14 11534 66
rect 11586 14 11600 66
rect 11520 0 11600 14
rect 11680 31417 11760 31440
rect 11680 31383 11703 31417
rect 11737 31383 11760 31417
rect 11680 31257 11760 31383
rect 11680 31223 11703 31257
rect 11737 31223 11760 31257
rect 11680 31097 11760 31223
rect 11680 31063 11703 31097
rect 11737 31063 11760 31097
rect 11680 30937 11760 31063
rect 11680 30903 11703 30937
rect 11737 30903 11760 30937
rect 11680 30777 11760 30903
rect 11680 30743 11703 30777
rect 11737 30743 11760 30777
rect 11680 30617 11760 30743
rect 11680 30583 11703 30617
rect 11737 30583 11760 30617
rect 11680 30457 11760 30583
rect 11680 30423 11703 30457
rect 11737 30423 11760 30457
rect 11680 30297 11760 30423
rect 11680 30263 11703 30297
rect 11737 30263 11760 30297
rect 11680 30137 11760 30263
rect 11680 30103 11703 30137
rect 11737 30103 11760 30137
rect 11680 29977 11760 30103
rect 11680 29943 11703 29977
rect 11737 29943 11760 29977
rect 11680 29817 11760 29943
rect 11680 29783 11703 29817
rect 11737 29783 11760 29817
rect 11680 29657 11760 29783
rect 11680 29623 11703 29657
rect 11737 29623 11760 29657
rect 11680 29497 11760 29623
rect 11680 29463 11703 29497
rect 11737 29463 11760 29497
rect 11680 29337 11760 29463
rect 11680 29303 11703 29337
rect 11737 29303 11760 29337
rect 11680 29177 11760 29303
rect 11680 29143 11703 29177
rect 11737 29143 11760 29177
rect 11680 29017 11760 29143
rect 11680 28983 11703 29017
rect 11737 28983 11760 29017
rect 11680 28857 11760 28983
rect 11680 28823 11703 28857
rect 11737 28823 11760 28857
rect 11680 28697 11760 28823
rect 11680 28663 11703 28697
rect 11737 28663 11760 28697
rect 11680 28537 11760 28663
rect 11680 28503 11703 28537
rect 11737 28503 11760 28537
rect 11680 28377 11760 28503
rect 11680 28343 11703 28377
rect 11737 28343 11760 28377
rect 11680 28217 11760 28343
rect 11680 28183 11703 28217
rect 11737 28183 11760 28217
rect 11680 28057 11760 28183
rect 11680 28023 11703 28057
rect 11737 28023 11760 28057
rect 11680 27897 11760 28023
rect 11680 27863 11703 27897
rect 11737 27863 11760 27897
rect 11680 27737 11760 27863
rect 11680 27703 11703 27737
rect 11737 27703 11760 27737
rect 11680 27577 11760 27703
rect 11680 27543 11703 27577
rect 11737 27543 11760 27577
rect 11680 27417 11760 27543
rect 11680 27383 11703 27417
rect 11737 27383 11760 27417
rect 11680 27257 11760 27383
rect 11680 27223 11703 27257
rect 11737 27223 11760 27257
rect 11680 27097 11760 27223
rect 11680 27063 11703 27097
rect 11737 27063 11760 27097
rect 11680 26937 11760 27063
rect 11680 26903 11703 26937
rect 11737 26903 11760 26937
rect 11680 26777 11760 26903
rect 11680 26743 11703 26777
rect 11737 26743 11760 26777
rect 11680 26617 11760 26743
rect 11680 26583 11703 26617
rect 11737 26583 11760 26617
rect 11680 26457 11760 26583
rect 11680 26423 11703 26457
rect 11737 26423 11760 26457
rect 11680 26297 11760 26423
rect 11680 26263 11703 26297
rect 11737 26263 11760 26297
rect 11680 26137 11760 26263
rect 11680 26103 11703 26137
rect 11737 26103 11760 26137
rect 11680 25977 11760 26103
rect 11680 25943 11703 25977
rect 11737 25943 11760 25977
rect 11680 25817 11760 25943
rect 11680 25783 11703 25817
rect 11737 25783 11760 25817
rect 11680 25657 11760 25783
rect 11680 25623 11703 25657
rect 11737 25623 11760 25657
rect 11680 25497 11760 25623
rect 11680 25463 11703 25497
rect 11737 25463 11760 25497
rect 11680 25337 11760 25463
rect 11680 25303 11703 25337
rect 11737 25303 11760 25337
rect 11680 25177 11760 25303
rect 11680 25143 11703 25177
rect 11737 25143 11760 25177
rect 11680 25017 11760 25143
rect 11680 24983 11703 25017
rect 11737 24983 11760 25017
rect 11680 24857 11760 24983
rect 11680 24823 11703 24857
rect 11737 24823 11760 24857
rect 11680 24697 11760 24823
rect 11680 24663 11703 24697
rect 11737 24663 11760 24697
rect 11680 24537 11760 24663
rect 11680 24503 11703 24537
rect 11737 24503 11760 24537
rect 11680 24377 11760 24503
rect 11680 24343 11703 24377
rect 11737 24343 11760 24377
rect 11680 24217 11760 24343
rect 11680 24183 11703 24217
rect 11737 24183 11760 24217
rect 11680 24057 11760 24183
rect 11680 24023 11703 24057
rect 11737 24023 11760 24057
rect 11680 23897 11760 24023
rect 11680 23863 11703 23897
rect 11737 23863 11760 23897
rect 11680 23737 11760 23863
rect 11680 23703 11703 23737
rect 11737 23703 11760 23737
rect 11680 23577 11760 23703
rect 11680 23543 11703 23577
rect 11737 23543 11760 23577
rect 11680 23417 11760 23543
rect 11680 23383 11703 23417
rect 11737 23383 11760 23417
rect 11680 23257 11760 23383
rect 11680 23223 11703 23257
rect 11737 23223 11760 23257
rect 11680 23097 11760 23223
rect 11680 23063 11703 23097
rect 11737 23063 11760 23097
rect 11680 22937 11760 23063
rect 11680 22903 11703 22937
rect 11737 22903 11760 22937
rect 11680 22777 11760 22903
rect 11680 22743 11703 22777
rect 11737 22743 11760 22777
rect 11680 22617 11760 22743
rect 11680 22583 11703 22617
rect 11737 22583 11760 22617
rect 11680 22457 11760 22583
rect 11680 22423 11703 22457
rect 11737 22423 11760 22457
rect 11680 22297 11760 22423
rect 11680 22263 11703 22297
rect 11737 22263 11760 22297
rect 11680 22137 11760 22263
rect 11680 22103 11703 22137
rect 11737 22103 11760 22137
rect 11680 21977 11760 22103
rect 11680 21943 11703 21977
rect 11737 21943 11760 21977
rect 11680 21817 11760 21943
rect 11680 21783 11703 21817
rect 11737 21783 11760 21817
rect 11680 21657 11760 21783
rect 11680 21623 11703 21657
rect 11737 21623 11760 21657
rect 11680 21497 11760 21623
rect 11680 21463 11703 21497
rect 11737 21463 11760 21497
rect 11680 21337 11760 21463
rect 11680 21303 11703 21337
rect 11737 21303 11760 21337
rect 11680 21177 11760 21303
rect 11680 21143 11703 21177
rect 11737 21143 11760 21177
rect 11680 21017 11760 21143
rect 11680 20983 11703 21017
rect 11737 20983 11760 21017
rect 11680 20857 11760 20983
rect 11680 20823 11703 20857
rect 11737 20823 11760 20857
rect 11680 20697 11760 20823
rect 11680 20663 11703 20697
rect 11737 20663 11760 20697
rect 11680 20537 11760 20663
rect 11680 20503 11703 20537
rect 11737 20503 11760 20537
rect 11680 20377 11760 20503
rect 11680 20343 11703 20377
rect 11737 20343 11760 20377
rect 11680 20217 11760 20343
rect 11680 20183 11703 20217
rect 11737 20183 11760 20217
rect 11680 20057 11760 20183
rect 11680 20023 11703 20057
rect 11737 20023 11760 20057
rect 11680 19897 11760 20023
rect 11680 19863 11703 19897
rect 11737 19863 11760 19897
rect 11680 19737 11760 19863
rect 11680 19703 11703 19737
rect 11737 19703 11760 19737
rect 11680 19577 11760 19703
rect 11680 19543 11703 19577
rect 11737 19543 11760 19577
rect 11680 19417 11760 19543
rect 11680 19383 11703 19417
rect 11737 19383 11760 19417
rect 11680 19257 11760 19383
rect 11680 19223 11703 19257
rect 11737 19223 11760 19257
rect 11680 19097 11760 19223
rect 11680 19063 11703 19097
rect 11737 19063 11760 19097
rect 11680 18937 11760 19063
rect 11680 18903 11703 18937
rect 11737 18903 11760 18937
rect 11680 18777 11760 18903
rect 11680 18743 11703 18777
rect 11737 18743 11760 18777
rect 11680 18617 11760 18743
rect 11680 18583 11703 18617
rect 11737 18583 11760 18617
rect 11680 18457 11760 18583
rect 11680 18423 11703 18457
rect 11737 18423 11760 18457
rect 11680 18297 11760 18423
rect 11680 18263 11703 18297
rect 11737 18263 11760 18297
rect 11680 18137 11760 18263
rect 11680 18103 11703 18137
rect 11737 18103 11760 18137
rect 11680 17977 11760 18103
rect 11680 17943 11703 17977
rect 11737 17943 11760 17977
rect 11680 17817 11760 17943
rect 11680 17783 11703 17817
rect 11737 17783 11760 17817
rect 11680 17657 11760 17783
rect 11680 17623 11703 17657
rect 11737 17623 11760 17657
rect 11680 17497 11760 17623
rect 11680 17463 11703 17497
rect 11737 17463 11760 17497
rect 11680 17337 11760 17463
rect 11680 17303 11703 17337
rect 11737 17303 11760 17337
rect 11680 17177 11760 17303
rect 11680 17143 11703 17177
rect 11737 17143 11760 17177
rect 11680 17017 11760 17143
rect 11680 16983 11703 17017
rect 11737 16983 11760 17017
rect 11680 16857 11760 16983
rect 11680 16823 11703 16857
rect 11737 16823 11760 16857
rect 11680 16697 11760 16823
rect 11680 16663 11703 16697
rect 11737 16663 11760 16697
rect 11680 16537 11760 16663
rect 11680 16503 11703 16537
rect 11737 16503 11760 16537
rect 11680 16377 11760 16503
rect 11680 16343 11703 16377
rect 11737 16343 11760 16377
rect 11680 16217 11760 16343
rect 11680 16183 11703 16217
rect 11737 16183 11760 16217
rect 11680 16057 11760 16183
rect 11680 16023 11703 16057
rect 11737 16023 11760 16057
rect 11680 15897 11760 16023
rect 11680 15863 11703 15897
rect 11737 15863 11760 15897
rect 11680 15737 11760 15863
rect 11680 15703 11703 15737
rect 11737 15703 11760 15737
rect 11680 15577 11760 15703
rect 11680 15543 11703 15577
rect 11737 15543 11760 15577
rect 11680 15417 11760 15543
rect 11680 15383 11703 15417
rect 11737 15383 11760 15417
rect 11680 15257 11760 15383
rect 11680 15223 11703 15257
rect 11737 15223 11760 15257
rect 11680 15097 11760 15223
rect 11680 15063 11703 15097
rect 11737 15063 11760 15097
rect 11680 14937 11760 15063
rect 11680 14903 11703 14937
rect 11737 14903 11760 14937
rect 11680 14777 11760 14903
rect 11680 14743 11703 14777
rect 11737 14743 11760 14777
rect 11680 14617 11760 14743
rect 11680 14583 11703 14617
rect 11737 14583 11760 14617
rect 11680 14457 11760 14583
rect 11680 14423 11703 14457
rect 11737 14423 11760 14457
rect 11680 14297 11760 14423
rect 11680 14263 11703 14297
rect 11737 14263 11760 14297
rect 11680 14137 11760 14263
rect 11680 14103 11703 14137
rect 11737 14103 11760 14137
rect 11680 13977 11760 14103
rect 11680 13943 11703 13977
rect 11737 13943 11760 13977
rect 11680 13817 11760 13943
rect 11680 13783 11703 13817
rect 11737 13783 11760 13817
rect 11680 13657 11760 13783
rect 11680 13623 11703 13657
rect 11737 13623 11760 13657
rect 11680 13497 11760 13623
rect 11680 13463 11703 13497
rect 11737 13463 11760 13497
rect 11680 13337 11760 13463
rect 11680 13303 11703 13337
rect 11737 13303 11760 13337
rect 11680 13177 11760 13303
rect 11680 13143 11703 13177
rect 11737 13143 11760 13177
rect 11680 13017 11760 13143
rect 11680 12983 11703 13017
rect 11737 12983 11760 13017
rect 11680 12857 11760 12983
rect 11680 12823 11703 12857
rect 11737 12823 11760 12857
rect 11680 12697 11760 12823
rect 11680 12663 11703 12697
rect 11737 12663 11760 12697
rect 11680 12537 11760 12663
rect 11680 12503 11703 12537
rect 11737 12503 11760 12537
rect 11680 12377 11760 12503
rect 11680 12343 11703 12377
rect 11737 12343 11760 12377
rect 11680 12217 11760 12343
rect 11680 12183 11703 12217
rect 11737 12183 11760 12217
rect 11680 12057 11760 12183
rect 11680 12023 11703 12057
rect 11737 12023 11760 12057
rect 11680 11897 11760 12023
rect 11680 11863 11703 11897
rect 11737 11863 11760 11897
rect 11680 11737 11760 11863
rect 11680 11703 11703 11737
rect 11737 11703 11760 11737
rect 11680 11577 11760 11703
rect 11680 11543 11703 11577
rect 11737 11543 11760 11577
rect 11680 11417 11760 11543
rect 11680 11383 11703 11417
rect 11737 11383 11760 11417
rect 11680 11257 11760 11383
rect 11680 11223 11703 11257
rect 11737 11223 11760 11257
rect 11680 11097 11760 11223
rect 11680 11063 11703 11097
rect 11737 11063 11760 11097
rect 11680 10937 11760 11063
rect 11680 10903 11703 10937
rect 11737 10903 11760 10937
rect 11680 10777 11760 10903
rect 11680 10743 11703 10777
rect 11737 10743 11760 10777
rect 11680 10617 11760 10743
rect 11680 10583 11703 10617
rect 11737 10583 11760 10617
rect 11680 10457 11760 10583
rect 11680 10423 11703 10457
rect 11737 10423 11760 10457
rect 11680 10297 11760 10423
rect 11680 10263 11703 10297
rect 11737 10263 11760 10297
rect 11680 10137 11760 10263
rect 11680 10103 11703 10137
rect 11737 10103 11760 10137
rect 11680 9977 11760 10103
rect 11680 9943 11703 9977
rect 11737 9943 11760 9977
rect 11680 9817 11760 9943
rect 11680 9783 11703 9817
rect 11737 9783 11760 9817
rect 11680 9657 11760 9783
rect 11680 9623 11703 9657
rect 11737 9623 11760 9657
rect 11680 9497 11760 9623
rect 11680 9463 11703 9497
rect 11737 9463 11760 9497
rect 11680 9337 11760 9463
rect 11680 9303 11703 9337
rect 11737 9303 11760 9337
rect 11680 9177 11760 9303
rect 11680 9143 11703 9177
rect 11737 9143 11760 9177
rect 11680 9017 11760 9143
rect 11680 8983 11703 9017
rect 11737 8983 11760 9017
rect 11680 8857 11760 8983
rect 11680 8823 11703 8857
rect 11737 8823 11760 8857
rect 11680 8697 11760 8823
rect 11680 8663 11703 8697
rect 11737 8663 11760 8697
rect 11680 8537 11760 8663
rect 11680 8503 11703 8537
rect 11737 8503 11760 8537
rect 11680 8377 11760 8503
rect 11680 8343 11703 8377
rect 11737 8343 11760 8377
rect 11680 8217 11760 8343
rect 11680 8183 11703 8217
rect 11737 8183 11760 8217
rect 11680 8057 11760 8183
rect 11680 8023 11703 8057
rect 11737 8023 11760 8057
rect 11680 7897 11760 8023
rect 11680 7863 11703 7897
rect 11737 7863 11760 7897
rect 11680 7737 11760 7863
rect 11680 7703 11703 7737
rect 11737 7703 11760 7737
rect 11680 7577 11760 7703
rect 11680 7543 11703 7577
rect 11737 7543 11760 7577
rect 11680 7417 11760 7543
rect 11680 7383 11703 7417
rect 11737 7383 11760 7417
rect 11680 7257 11760 7383
rect 11680 7223 11703 7257
rect 11737 7223 11760 7257
rect 11680 7097 11760 7223
rect 11680 7063 11703 7097
rect 11737 7063 11760 7097
rect 11680 6937 11760 7063
rect 11680 6903 11703 6937
rect 11737 6903 11760 6937
rect 11680 6777 11760 6903
rect 11680 6743 11703 6777
rect 11737 6743 11760 6777
rect 11680 6617 11760 6743
rect 11680 6583 11703 6617
rect 11737 6583 11760 6617
rect 11680 6457 11760 6583
rect 11680 6423 11703 6457
rect 11737 6423 11760 6457
rect 11680 6297 11760 6423
rect 11680 6263 11703 6297
rect 11737 6263 11760 6297
rect 11680 6137 11760 6263
rect 11680 6103 11703 6137
rect 11737 6103 11760 6137
rect 11680 5977 11760 6103
rect 11680 5943 11703 5977
rect 11737 5943 11760 5977
rect 11680 5817 11760 5943
rect 11680 5783 11703 5817
rect 11737 5783 11760 5817
rect 11680 5657 11760 5783
rect 11680 5623 11703 5657
rect 11737 5623 11760 5657
rect 11680 5497 11760 5623
rect 11680 5463 11703 5497
rect 11737 5463 11760 5497
rect 11680 5337 11760 5463
rect 11680 5303 11703 5337
rect 11737 5303 11760 5337
rect 11680 5177 11760 5303
rect 11680 5143 11703 5177
rect 11737 5143 11760 5177
rect 11680 5017 11760 5143
rect 11680 4983 11703 5017
rect 11737 4983 11760 5017
rect 11680 4857 11760 4983
rect 11680 4823 11703 4857
rect 11737 4823 11760 4857
rect 11680 4697 11760 4823
rect 11680 4663 11703 4697
rect 11737 4663 11760 4697
rect 11680 4537 11760 4663
rect 11680 4503 11703 4537
rect 11737 4503 11760 4537
rect 11680 4377 11760 4503
rect 11680 4343 11703 4377
rect 11737 4343 11760 4377
rect 11680 4217 11760 4343
rect 11680 4183 11703 4217
rect 11737 4183 11760 4217
rect 11680 4057 11760 4183
rect 11680 4023 11703 4057
rect 11737 4023 11760 4057
rect 11680 3897 11760 4023
rect 11680 3863 11703 3897
rect 11737 3863 11760 3897
rect 11680 3737 11760 3863
rect 11680 3703 11703 3737
rect 11737 3703 11760 3737
rect 11680 3577 11760 3703
rect 11680 3543 11703 3577
rect 11737 3543 11760 3577
rect 11680 3417 11760 3543
rect 11680 3383 11703 3417
rect 11737 3383 11760 3417
rect 11680 3257 11760 3383
rect 11680 3223 11703 3257
rect 11737 3223 11760 3257
rect 11680 3097 11760 3223
rect 11680 3063 11703 3097
rect 11737 3063 11760 3097
rect 11680 2937 11760 3063
rect 11680 2903 11703 2937
rect 11737 2903 11760 2937
rect 11680 2777 11760 2903
rect 11680 2743 11703 2777
rect 11737 2743 11760 2777
rect 11680 2617 11760 2743
rect 11680 2583 11703 2617
rect 11737 2583 11760 2617
rect 11680 2457 11760 2583
rect 11680 2423 11703 2457
rect 11737 2423 11760 2457
rect 11680 2297 11760 2423
rect 11680 2263 11703 2297
rect 11737 2263 11760 2297
rect 11680 2137 11760 2263
rect 11680 2103 11703 2137
rect 11737 2103 11760 2137
rect 11680 1977 11760 2103
rect 11680 1943 11703 1977
rect 11737 1943 11760 1977
rect 11680 1817 11760 1943
rect 11680 1783 11703 1817
rect 11737 1783 11760 1817
rect 11680 1657 11760 1783
rect 11680 1623 11703 1657
rect 11737 1623 11760 1657
rect 11680 1497 11760 1623
rect 11680 1463 11703 1497
rect 11737 1463 11760 1497
rect 11680 1337 11760 1463
rect 11680 1303 11703 1337
rect 11737 1303 11760 1337
rect 11680 1177 11760 1303
rect 11680 1143 11703 1177
rect 11737 1143 11760 1177
rect 11680 1017 11760 1143
rect 11680 983 11703 1017
rect 11737 983 11760 1017
rect 11680 857 11760 983
rect 11680 823 11703 857
rect 11737 823 11760 857
rect 11680 697 11760 823
rect 11680 663 11703 697
rect 11737 663 11760 697
rect 11680 537 11760 663
rect 11680 503 11703 537
rect 11737 503 11760 537
rect 11680 377 11760 503
rect 11680 343 11703 377
rect 11737 343 11760 377
rect 11680 217 11760 343
rect 11680 183 11703 217
rect 11737 183 11760 217
rect 11680 57 11760 183
rect 11680 23 11703 57
rect 11737 23 11760 57
rect 11680 0 11760 23
rect 11840 31426 11920 31440
rect 11840 31374 11854 31426
rect 11906 31374 11920 31426
rect 11840 31266 11920 31374
rect 11840 31214 11854 31266
rect 11906 31214 11920 31266
rect 11840 31106 11920 31214
rect 11840 31054 11854 31106
rect 11906 31054 11920 31106
rect 11840 30946 11920 31054
rect 11840 30894 11854 30946
rect 11906 30894 11920 30946
rect 11840 30786 11920 30894
rect 11840 30734 11854 30786
rect 11906 30734 11920 30786
rect 11840 30626 11920 30734
rect 11840 30574 11854 30626
rect 11906 30574 11920 30626
rect 11840 30466 11920 30574
rect 11840 30414 11854 30466
rect 11906 30414 11920 30466
rect 11840 30306 11920 30414
rect 11840 30254 11854 30306
rect 11906 30254 11920 30306
rect 11840 30137 11920 30254
rect 11840 30103 11863 30137
rect 11897 30103 11920 30137
rect 11840 29986 11920 30103
rect 11840 29934 11854 29986
rect 11906 29934 11920 29986
rect 11840 29826 11920 29934
rect 11840 29774 11854 29826
rect 11906 29774 11920 29826
rect 11840 29666 11920 29774
rect 11840 29614 11854 29666
rect 11906 29614 11920 29666
rect 11840 29506 11920 29614
rect 11840 29454 11854 29506
rect 11906 29454 11920 29506
rect 11840 29346 11920 29454
rect 11840 29294 11854 29346
rect 11906 29294 11920 29346
rect 11840 29186 11920 29294
rect 11840 29134 11854 29186
rect 11906 29134 11920 29186
rect 11840 29026 11920 29134
rect 11840 28974 11854 29026
rect 11906 28974 11920 29026
rect 11840 28866 11920 28974
rect 11840 28814 11854 28866
rect 11906 28814 11920 28866
rect 11840 28697 11920 28814
rect 11840 28663 11863 28697
rect 11897 28663 11920 28697
rect 11840 28537 11920 28663
rect 11840 28503 11863 28537
rect 11897 28503 11920 28537
rect 11840 28377 11920 28503
rect 11840 28343 11863 28377
rect 11897 28343 11920 28377
rect 11840 28217 11920 28343
rect 11840 28183 11863 28217
rect 11897 28183 11920 28217
rect 11840 28066 11920 28183
rect 11840 28014 11854 28066
rect 11906 28014 11920 28066
rect 11840 27906 11920 28014
rect 11840 27854 11854 27906
rect 11906 27854 11920 27906
rect 11840 27746 11920 27854
rect 11840 27694 11854 27746
rect 11906 27694 11920 27746
rect 11840 27586 11920 27694
rect 11840 27534 11854 27586
rect 11906 27534 11920 27586
rect 11840 27426 11920 27534
rect 11840 27374 11854 27426
rect 11906 27374 11920 27426
rect 11840 27266 11920 27374
rect 11840 27214 11854 27266
rect 11906 27214 11920 27266
rect 11840 27106 11920 27214
rect 11840 27054 11854 27106
rect 11906 27054 11920 27106
rect 11840 26946 11920 27054
rect 11840 26894 11854 26946
rect 11906 26894 11920 26946
rect 11840 26777 11920 26894
rect 11840 26743 11863 26777
rect 11897 26743 11920 26777
rect 11840 26617 11920 26743
rect 11840 26583 11863 26617
rect 11897 26583 11920 26617
rect 11840 26457 11920 26583
rect 11840 26423 11863 26457
rect 11897 26423 11920 26457
rect 11840 26297 11920 26423
rect 11840 26263 11863 26297
rect 11897 26263 11920 26297
rect 11840 26146 11920 26263
rect 11840 26094 11854 26146
rect 11906 26094 11920 26146
rect 11840 25986 11920 26094
rect 11840 25934 11854 25986
rect 11906 25934 11920 25986
rect 11840 25826 11920 25934
rect 11840 25774 11854 25826
rect 11906 25774 11920 25826
rect 11840 25666 11920 25774
rect 11840 25614 11854 25666
rect 11906 25614 11920 25666
rect 11840 25506 11920 25614
rect 11840 25454 11854 25506
rect 11906 25454 11920 25506
rect 11840 25346 11920 25454
rect 11840 25294 11854 25346
rect 11906 25294 11920 25346
rect 11840 25186 11920 25294
rect 11840 25134 11854 25186
rect 11906 25134 11920 25186
rect 11840 25026 11920 25134
rect 11840 24974 11854 25026
rect 11906 24974 11920 25026
rect 11840 24857 11920 24974
rect 11840 24823 11863 24857
rect 11897 24823 11920 24857
rect 11840 24706 11920 24823
rect 11840 24654 11854 24706
rect 11906 24654 11920 24706
rect 11840 24546 11920 24654
rect 11840 24494 11854 24546
rect 11906 24494 11920 24546
rect 11840 24386 11920 24494
rect 11840 24334 11854 24386
rect 11906 24334 11920 24386
rect 11840 24226 11920 24334
rect 11840 24174 11854 24226
rect 11906 24174 11920 24226
rect 11840 24066 11920 24174
rect 11840 24014 11854 24066
rect 11906 24014 11920 24066
rect 11840 23906 11920 24014
rect 11840 23854 11854 23906
rect 11906 23854 11920 23906
rect 11840 23746 11920 23854
rect 11840 23694 11854 23746
rect 11906 23694 11920 23746
rect 11840 23586 11920 23694
rect 11840 23534 11854 23586
rect 11906 23534 11920 23586
rect 11840 23426 11920 23534
rect 11840 23374 11854 23426
rect 11906 23374 11920 23426
rect 11840 23266 11920 23374
rect 11840 23214 11854 23266
rect 11906 23214 11920 23266
rect 11840 23106 11920 23214
rect 11840 23054 11854 23106
rect 11906 23054 11920 23106
rect 11840 22946 11920 23054
rect 11840 22894 11854 22946
rect 11906 22894 11920 22946
rect 11840 22786 11920 22894
rect 11840 22734 11854 22786
rect 11906 22734 11920 22786
rect 11840 22626 11920 22734
rect 11840 22574 11854 22626
rect 11906 22574 11920 22626
rect 11840 22466 11920 22574
rect 11840 22414 11854 22466
rect 11906 22414 11920 22466
rect 11840 22306 11920 22414
rect 11840 22254 11854 22306
rect 11906 22254 11920 22306
rect 11840 22146 11920 22254
rect 11840 22094 11854 22146
rect 11906 22094 11920 22146
rect 11840 21977 11920 22094
rect 11840 21943 11863 21977
rect 11897 21943 11920 21977
rect 11840 21826 11920 21943
rect 11840 21774 11854 21826
rect 11906 21774 11920 21826
rect 11840 21666 11920 21774
rect 11840 21614 11854 21666
rect 11906 21614 11920 21666
rect 11840 21506 11920 21614
rect 11840 21454 11854 21506
rect 11906 21454 11920 21506
rect 11840 21346 11920 21454
rect 11840 21294 11854 21346
rect 11906 21294 11920 21346
rect 11840 21186 11920 21294
rect 11840 21134 11854 21186
rect 11906 21134 11920 21186
rect 11840 21026 11920 21134
rect 11840 20974 11854 21026
rect 11906 20974 11920 21026
rect 11840 20866 11920 20974
rect 11840 20814 11854 20866
rect 11906 20814 11920 20866
rect 11840 20706 11920 20814
rect 11840 20654 11854 20706
rect 11906 20654 11920 20706
rect 11840 20537 11920 20654
rect 11840 20503 11863 20537
rect 11897 20503 11920 20537
rect 11840 20377 11920 20503
rect 11840 20343 11863 20377
rect 11897 20343 11920 20377
rect 11840 20217 11920 20343
rect 11840 20183 11863 20217
rect 11897 20183 11920 20217
rect 11840 20057 11920 20183
rect 11840 20023 11863 20057
rect 11897 20023 11920 20057
rect 11840 19906 11920 20023
rect 11840 19854 11854 19906
rect 11906 19854 11920 19906
rect 11840 19746 11920 19854
rect 11840 19694 11854 19746
rect 11906 19694 11920 19746
rect 11840 19586 11920 19694
rect 11840 19534 11854 19586
rect 11906 19534 11920 19586
rect 11840 19426 11920 19534
rect 11840 19374 11854 19426
rect 11906 19374 11920 19426
rect 11840 19266 11920 19374
rect 11840 19214 11854 19266
rect 11906 19214 11920 19266
rect 11840 19106 11920 19214
rect 11840 19054 11854 19106
rect 11906 19054 11920 19106
rect 11840 18946 11920 19054
rect 11840 18894 11854 18946
rect 11906 18894 11920 18946
rect 11840 18786 11920 18894
rect 11840 18734 11854 18786
rect 11906 18734 11920 18786
rect 11840 18617 11920 18734
rect 11840 18583 11863 18617
rect 11897 18583 11920 18617
rect 11840 18457 11920 18583
rect 11840 18423 11863 18457
rect 11897 18423 11920 18457
rect 11840 18297 11920 18423
rect 11840 18263 11863 18297
rect 11897 18263 11920 18297
rect 11840 18137 11920 18263
rect 11840 18103 11863 18137
rect 11897 18103 11920 18137
rect 11840 17986 11920 18103
rect 11840 17934 11854 17986
rect 11906 17934 11920 17986
rect 11840 17826 11920 17934
rect 11840 17774 11854 17826
rect 11906 17774 11920 17826
rect 11840 17666 11920 17774
rect 11840 17614 11854 17666
rect 11906 17614 11920 17666
rect 11840 17506 11920 17614
rect 11840 17454 11854 17506
rect 11906 17454 11920 17506
rect 11840 17346 11920 17454
rect 11840 17294 11854 17346
rect 11906 17294 11920 17346
rect 11840 17186 11920 17294
rect 11840 17134 11854 17186
rect 11906 17134 11920 17186
rect 11840 17026 11920 17134
rect 11840 16974 11854 17026
rect 11906 16974 11920 17026
rect 11840 16866 11920 16974
rect 11840 16814 11854 16866
rect 11906 16814 11920 16866
rect 11840 16697 11920 16814
rect 11840 16663 11863 16697
rect 11897 16663 11920 16697
rect 11840 16546 11920 16663
rect 11840 16494 11854 16546
rect 11906 16494 11920 16546
rect 11840 16386 11920 16494
rect 11840 16334 11854 16386
rect 11906 16334 11920 16386
rect 11840 16226 11920 16334
rect 11840 16174 11854 16226
rect 11906 16174 11920 16226
rect 11840 16066 11920 16174
rect 11840 16014 11854 16066
rect 11906 16014 11920 16066
rect 11840 15906 11920 16014
rect 11840 15854 11854 15906
rect 11906 15854 11920 15906
rect 11840 15746 11920 15854
rect 11840 15694 11854 15746
rect 11906 15694 11920 15746
rect 11840 15586 11920 15694
rect 11840 15534 11854 15586
rect 11906 15534 11920 15586
rect 11840 15426 11920 15534
rect 11840 15374 11854 15426
rect 11906 15374 11920 15426
rect 11840 15266 11920 15374
rect 11840 15214 11854 15266
rect 11906 15214 11920 15266
rect 11840 15106 11920 15214
rect 11840 15054 11854 15106
rect 11906 15054 11920 15106
rect 11840 14946 11920 15054
rect 11840 14894 11854 14946
rect 11906 14894 11920 14946
rect 11840 14786 11920 14894
rect 11840 14734 11854 14786
rect 11906 14734 11920 14786
rect 11840 14626 11920 14734
rect 11840 14574 11854 14626
rect 11906 14574 11920 14626
rect 11840 14466 11920 14574
rect 11840 14414 11854 14466
rect 11906 14414 11920 14466
rect 11840 14306 11920 14414
rect 11840 14254 11854 14306
rect 11906 14254 11920 14306
rect 11840 14146 11920 14254
rect 11840 14094 11854 14146
rect 11906 14094 11920 14146
rect 11840 13986 11920 14094
rect 11840 13934 11854 13986
rect 11906 13934 11920 13986
rect 11840 13817 11920 13934
rect 11840 13783 11863 13817
rect 11897 13783 11920 13817
rect 11840 13666 11920 13783
rect 11840 13614 11854 13666
rect 11906 13614 11920 13666
rect 11840 13506 11920 13614
rect 11840 13454 11854 13506
rect 11906 13454 11920 13506
rect 11840 13346 11920 13454
rect 11840 13294 11854 13346
rect 11906 13294 11920 13346
rect 11840 13186 11920 13294
rect 11840 13134 11854 13186
rect 11906 13134 11920 13186
rect 11840 13026 11920 13134
rect 11840 12974 11854 13026
rect 11906 12974 11920 13026
rect 11840 12866 11920 12974
rect 11840 12814 11854 12866
rect 11906 12814 11920 12866
rect 11840 12706 11920 12814
rect 11840 12654 11854 12706
rect 11906 12654 11920 12706
rect 11840 12546 11920 12654
rect 11840 12494 11854 12546
rect 11906 12494 11920 12546
rect 11840 12377 11920 12494
rect 11840 12343 11863 12377
rect 11897 12343 11920 12377
rect 11840 12217 11920 12343
rect 11840 12183 11863 12217
rect 11897 12183 11920 12217
rect 11840 12057 11920 12183
rect 11840 12023 11863 12057
rect 11897 12023 11920 12057
rect 11840 11897 11920 12023
rect 11840 11863 11863 11897
rect 11897 11863 11920 11897
rect 11840 11746 11920 11863
rect 11840 11694 11854 11746
rect 11906 11694 11920 11746
rect 11840 11586 11920 11694
rect 11840 11534 11854 11586
rect 11906 11534 11920 11586
rect 11840 11426 11920 11534
rect 11840 11374 11854 11426
rect 11906 11374 11920 11426
rect 11840 11266 11920 11374
rect 11840 11214 11854 11266
rect 11906 11214 11920 11266
rect 11840 11106 11920 11214
rect 11840 11054 11854 11106
rect 11906 11054 11920 11106
rect 11840 10946 11920 11054
rect 11840 10894 11854 10946
rect 11906 10894 11920 10946
rect 11840 10786 11920 10894
rect 11840 10734 11854 10786
rect 11906 10734 11920 10786
rect 11840 10626 11920 10734
rect 11840 10574 11854 10626
rect 11906 10574 11920 10626
rect 11840 10466 11920 10574
rect 11840 10414 11854 10466
rect 11906 10414 11920 10466
rect 11840 10306 11920 10414
rect 11840 10254 11854 10306
rect 11906 10254 11920 10306
rect 11840 10146 11920 10254
rect 11840 10094 11854 10146
rect 11906 10094 11920 10146
rect 11840 9986 11920 10094
rect 11840 9934 11854 9986
rect 11906 9934 11920 9986
rect 11840 9826 11920 9934
rect 11840 9774 11854 9826
rect 11906 9774 11920 9826
rect 11840 9657 11920 9774
rect 11840 9623 11863 9657
rect 11897 9623 11920 9657
rect 11840 9506 11920 9623
rect 11840 9454 11854 9506
rect 11906 9454 11920 9506
rect 11840 9346 11920 9454
rect 11840 9294 11854 9346
rect 11906 9294 11920 9346
rect 11840 9177 11920 9294
rect 11840 9143 11863 9177
rect 11897 9143 11920 9177
rect 11840 9026 11920 9143
rect 11840 8974 11854 9026
rect 11906 8974 11920 9026
rect 11840 8866 11920 8974
rect 11840 8814 11854 8866
rect 11906 8814 11920 8866
rect 11840 8706 11920 8814
rect 11840 8654 11854 8706
rect 11906 8654 11920 8706
rect 11840 8546 11920 8654
rect 11840 8494 11854 8546
rect 11906 8494 11920 8546
rect 11840 8386 11920 8494
rect 11840 8334 11854 8386
rect 11906 8334 11920 8386
rect 11840 8226 11920 8334
rect 11840 8174 11854 8226
rect 11906 8174 11920 8226
rect 11840 8066 11920 8174
rect 11840 8014 11854 8066
rect 11906 8014 11920 8066
rect 11840 7906 11920 8014
rect 11840 7854 11854 7906
rect 11906 7854 11920 7906
rect 11840 7746 11920 7854
rect 11840 7694 11854 7746
rect 11906 7694 11920 7746
rect 11840 7577 11920 7694
rect 11840 7543 11863 7577
rect 11897 7543 11920 7577
rect 11840 7426 11920 7543
rect 11840 7374 11854 7426
rect 11906 7374 11920 7426
rect 11840 7266 11920 7374
rect 11840 7214 11854 7266
rect 11906 7214 11920 7266
rect 11840 7097 11920 7214
rect 11840 7063 11863 7097
rect 11897 7063 11920 7097
rect 11840 6946 11920 7063
rect 11840 6894 11854 6946
rect 11906 6894 11920 6946
rect 11840 6786 11920 6894
rect 11840 6734 11854 6786
rect 11906 6734 11920 6786
rect 11840 6617 11920 6734
rect 11840 6583 11863 6617
rect 11897 6583 11920 6617
rect 11840 6466 11920 6583
rect 11840 6414 11854 6466
rect 11906 6414 11920 6466
rect 11840 6306 11920 6414
rect 11840 6254 11854 6306
rect 11906 6254 11920 6306
rect 11840 6146 11920 6254
rect 11840 6094 11854 6146
rect 11906 6094 11920 6146
rect 11840 5986 11920 6094
rect 11840 5934 11854 5986
rect 11906 5934 11920 5986
rect 11840 5826 11920 5934
rect 11840 5774 11854 5826
rect 11906 5774 11920 5826
rect 11840 5666 11920 5774
rect 11840 5614 11854 5666
rect 11906 5614 11920 5666
rect 11840 5506 11920 5614
rect 11840 5454 11854 5506
rect 11906 5454 11920 5506
rect 11840 5346 11920 5454
rect 11840 5294 11854 5346
rect 11906 5294 11920 5346
rect 11840 5186 11920 5294
rect 11840 5134 11854 5186
rect 11906 5134 11920 5186
rect 11840 5026 11920 5134
rect 11840 4974 11854 5026
rect 11906 4974 11920 5026
rect 11840 4866 11920 4974
rect 11840 4814 11854 4866
rect 11906 4814 11920 4866
rect 11840 4706 11920 4814
rect 11840 4654 11854 4706
rect 11906 4654 11920 4706
rect 11840 4546 11920 4654
rect 11840 4494 11854 4546
rect 11906 4494 11920 4546
rect 11840 4386 11920 4494
rect 11840 4334 11854 4386
rect 11906 4334 11920 4386
rect 11840 4226 11920 4334
rect 11840 4174 11854 4226
rect 11906 4174 11920 4226
rect 11840 4066 11920 4174
rect 11840 4014 11854 4066
rect 11906 4014 11920 4066
rect 11840 3906 11920 4014
rect 11840 3854 11854 3906
rect 11906 3854 11920 3906
rect 11840 3737 11920 3854
rect 11840 3703 11863 3737
rect 11897 3703 11920 3737
rect 11840 3577 11920 3703
rect 11840 3543 11863 3577
rect 11897 3543 11920 3577
rect 11840 3426 11920 3543
rect 11840 3374 11854 3426
rect 11906 3374 11920 3426
rect 11840 3266 11920 3374
rect 11840 3214 11854 3266
rect 11906 3214 11920 3266
rect 11840 3106 11920 3214
rect 11840 3054 11854 3106
rect 11906 3054 11920 3106
rect 11840 2946 11920 3054
rect 11840 2894 11854 2946
rect 11906 2894 11920 2946
rect 11840 2786 11920 2894
rect 11840 2734 11854 2786
rect 11906 2734 11920 2786
rect 11840 2626 11920 2734
rect 11840 2574 11854 2626
rect 11906 2574 11920 2626
rect 11840 2466 11920 2574
rect 11840 2414 11854 2466
rect 11906 2414 11920 2466
rect 11840 2306 11920 2414
rect 11840 2254 11854 2306
rect 11906 2254 11920 2306
rect 11840 2146 11920 2254
rect 11840 2094 11854 2146
rect 11906 2094 11920 2146
rect 11840 1986 11920 2094
rect 11840 1934 11854 1986
rect 11906 1934 11920 1986
rect 11840 1817 11920 1934
rect 11840 1783 11863 1817
rect 11897 1783 11920 1817
rect 11840 1666 11920 1783
rect 11840 1614 11854 1666
rect 11906 1614 11920 1666
rect 11840 1506 11920 1614
rect 11840 1454 11854 1506
rect 11906 1454 11920 1506
rect 11840 1346 11920 1454
rect 11840 1294 11854 1346
rect 11906 1294 11920 1346
rect 11840 1186 11920 1294
rect 11840 1134 11854 1186
rect 11906 1134 11920 1186
rect 11840 1026 11920 1134
rect 11840 974 11854 1026
rect 11906 974 11920 1026
rect 11840 857 11920 974
rect 11840 823 11863 857
rect 11897 823 11920 857
rect 11840 697 11920 823
rect 11840 663 11863 697
rect 11897 663 11920 697
rect 11840 546 11920 663
rect 11840 494 11854 546
rect 11906 494 11920 546
rect 11840 386 11920 494
rect 11840 334 11854 386
rect 11906 334 11920 386
rect 11840 226 11920 334
rect 11840 174 11854 226
rect 11906 174 11920 226
rect 11840 66 11920 174
rect 11840 14 11854 66
rect 11906 14 11920 66
rect 11840 0 11920 14
rect 12000 31426 12080 31440
rect 12000 31374 12014 31426
rect 12066 31374 12080 31426
rect 12000 31266 12080 31374
rect 12000 31214 12014 31266
rect 12066 31214 12080 31266
rect 12000 31106 12080 31214
rect 12000 31054 12014 31106
rect 12066 31054 12080 31106
rect 12000 30946 12080 31054
rect 12000 30894 12014 30946
rect 12066 30894 12080 30946
rect 12000 30786 12080 30894
rect 12000 30734 12014 30786
rect 12066 30734 12080 30786
rect 12000 30626 12080 30734
rect 12000 30574 12014 30626
rect 12066 30574 12080 30626
rect 12000 30466 12080 30574
rect 12000 30414 12014 30466
rect 12066 30414 12080 30466
rect 12000 30306 12080 30414
rect 12000 30254 12014 30306
rect 12066 30254 12080 30306
rect 12000 30137 12080 30254
rect 12000 30103 12023 30137
rect 12057 30103 12080 30137
rect 12000 29986 12080 30103
rect 12000 29934 12014 29986
rect 12066 29934 12080 29986
rect 12000 29826 12080 29934
rect 12000 29774 12014 29826
rect 12066 29774 12080 29826
rect 12000 29666 12080 29774
rect 12000 29614 12014 29666
rect 12066 29614 12080 29666
rect 12000 29506 12080 29614
rect 12000 29454 12014 29506
rect 12066 29454 12080 29506
rect 12000 29346 12080 29454
rect 12000 29294 12014 29346
rect 12066 29294 12080 29346
rect 12000 29186 12080 29294
rect 12000 29134 12014 29186
rect 12066 29134 12080 29186
rect 12000 29026 12080 29134
rect 12000 28974 12014 29026
rect 12066 28974 12080 29026
rect 12000 28866 12080 28974
rect 12000 28814 12014 28866
rect 12066 28814 12080 28866
rect 12000 28697 12080 28814
rect 12000 28663 12023 28697
rect 12057 28663 12080 28697
rect 12000 28537 12080 28663
rect 12000 28503 12023 28537
rect 12057 28503 12080 28537
rect 12000 28377 12080 28503
rect 12000 28343 12023 28377
rect 12057 28343 12080 28377
rect 12000 28217 12080 28343
rect 12000 28183 12023 28217
rect 12057 28183 12080 28217
rect 12000 28066 12080 28183
rect 12000 28014 12014 28066
rect 12066 28014 12080 28066
rect 12000 27906 12080 28014
rect 12000 27854 12014 27906
rect 12066 27854 12080 27906
rect 12000 27746 12080 27854
rect 12000 27694 12014 27746
rect 12066 27694 12080 27746
rect 12000 27586 12080 27694
rect 12000 27534 12014 27586
rect 12066 27534 12080 27586
rect 12000 27426 12080 27534
rect 12000 27374 12014 27426
rect 12066 27374 12080 27426
rect 12000 27266 12080 27374
rect 12000 27214 12014 27266
rect 12066 27214 12080 27266
rect 12000 27106 12080 27214
rect 12000 27054 12014 27106
rect 12066 27054 12080 27106
rect 12000 26946 12080 27054
rect 12000 26894 12014 26946
rect 12066 26894 12080 26946
rect 12000 26777 12080 26894
rect 12000 26743 12023 26777
rect 12057 26743 12080 26777
rect 12000 26617 12080 26743
rect 12000 26583 12023 26617
rect 12057 26583 12080 26617
rect 12000 26457 12080 26583
rect 12000 26423 12023 26457
rect 12057 26423 12080 26457
rect 12000 26297 12080 26423
rect 12000 26263 12023 26297
rect 12057 26263 12080 26297
rect 12000 26146 12080 26263
rect 12000 26094 12014 26146
rect 12066 26094 12080 26146
rect 12000 25986 12080 26094
rect 12000 25934 12014 25986
rect 12066 25934 12080 25986
rect 12000 25826 12080 25934
rect 12000 25774 12014 25826
rect 12066 25774 12080 25826
rect 12000 25666 12080 25774
rect 12000 25614 12014 25666
rect 12066 25614 12080 25666
rect 12000 25506 12080 25614
rect 12000 25454 12014 25506
rect 12066 25454 12080 25506
rect 12000 25346 12080 25454
rect 12000 25294 12014 25346
rect 12066 25294 12080 25346
rect 12000 25186 12080 25294
rect 12000 25134 12014 25186
rect 12066 25134 12080 25186
rect 12000 25026 12080 25134
rect 12000 24974 12014 25026
rect 12066 24974 12080 25026
rect 12000 24857 12080 24974
rect 12000 24823 12023 24857
rect 12057 24823 12080 24857
rect 12000 24706 12080 24823
rect 12000 24654 12014 24706
rect 12066 24654 12080 24706
rect 12000 24546 12080 24654
rect 12000 24494 12014 24546
rect 12066 24494 12080 24546
rect 12000 24386 12080 24494
rect 12000 24334 12014 24386
rect 12066 24334 12080 24386
rect 12000 24226 12080 24334
rect 12000 24174 12014 24226
rect 12066 24174 12080 24226
rect 12000 24066 12080 24174
rect 12000 24014 12014 24066
rect 12066 24014 12080 24066
rect 12000 23906 12080 24014
rect 12000 23854 12014 23906
rect 12066 23854 12080 23906
rect 12000 23746 12080 23854
rect 12000 23694 12014 23746
rect 12066 23694 12080 23746
rect 12000 23586 12080 23694
rect 12000 23534 12014 23586
rect 12066 23534 12080 23586
rect 12000 23426 12080 23534
rect 12000 23374 12014 23426
rect 12066 23374 12080 23426
rect 12000 23266 12080 23374
rect 12000 23214 12014 23266
rect 12066 23214 12080 23266
rect 12000 23106 12080 23214
rect 12000 23054 12014 23106
rect 12066 23054 12080 23106
rect 12000 22946 12080 23054
rect 12000 22894 12014 22946
rect 12066 22894 12080 22946
rect 12000 22786 12080 22894
rect 12000 22734 12014 22786
rect 12066 22734 12080 22786
rect 12000 22626 12080 22734
rect 12000 22574 12014 22626
rect 12066 22574 12080 22626
rect 12000 22466 12080 22574
rect 12000 22414 12014 22466
rect 12066 22414 12080 22466
rect 12000 22306 12080 22414
rect 12000 22254 12014 22306
rect 12066 22254 12080 22306
rect 12000 22146 12080 22254
rect 12000 22094 12014 22146
rect 12066 22094 12080 22146
rect 12000 21977 12080 22094
rect 12000 21943 12023 21977
rect 12057 21943 12080 21977
rect 12000 21826 12080 21943
rect 12000 21774 12014 21826
rect 12066 21774 12080 21826
rect 12000 21666 12080 21774
rect 12000 21614 12014 21666
rect 12066 21614 12080 21666
rect 12000 21506 12080 21614
rect 12000 21454 12014 21506
rect 12066 21454 12080 21506
rect 12000 21346 12080 21454
rect 12000 21294 12014 21346
rect 12066 21294 12080 21346
rect 12000 21186 12080 21294
rect 12000 21134 12014 21186
rect 12066 21134 12080 21186
rect 12000 21026 12080 21134
rect 12000 20974 12014 21026
rect 12066 20974 12080 21026
rect 12000 20866 12080 20974
rect 12000 20814 12014 20866
rect 12066 20814 12080 20866
rect 12000 20706 12080 20814
rect 12000 20654 12014 20706
rect 12066 20654 12080 20706
rect 12000 20537 12080 20654
rect 12000 20503 12023 20537
rect 12057 20503 12080 20537
rect 12000 20377 12080 20503
rect 12000 20343 12023 20377
rect 12057 20343 12080 20377
rect 12000 20217 12080 20343
rect 12000 20183 12023 20217
rect 12057 20183 12080 20217
rect 12000 20057 12080 20183
rect 12000 20023 12023 20057
rect 12057 20023 12080 20057
rect 12000 19906 12080 20023
rect 12000 19854 12014 19906
rect 12066 19854 12080 19906
rect 12000 19746 12080 19854
rect 12000 19694 12014 19746
rect 12066 19694 12080 19746
rect 12000 19586 12080 19694
rect 12000 19534 12014 19586
rect 12066 19534 12080 19586
rect 12000 19426 12080 19534
rect 12000 19374 12014 19426
rect 12066 19374 12080 19426
rect 12000 19266 12080 19374
rect 12000 19214 12014 19266
rect 12066 19214 12080 19266
rect 12000 19106 12080 19214
rect 12000 19054 12014 19106
rect 12066 19054 12080 19106
rect 12000 18946 12080 19054
rect 12000 18894 12014 18946
rect 12066 18894 12080 18946
rect 12000 18786 12080 18894
rect 12000 18734 12014 18786
rect 12066 18734 12080 18786
rect 12000 18617 12080 18734
rect 12000 18583 12023 18617
rect 12057 18583 12080 18617
rect 12000 18457 12080 18583
rect 12000 18423 12023 18457
rect 12057 18423 12080 18457
rect 12000 18297 12080 18423
rect 12000 18263 12023 18297
rect 12057 18263 12080 18297
rect 12000 18137 12080 18263
rect 12000 18103 12023 18137
rect 12057 18103 12080 18137
rect 12000 17986 12080 18103
rect 12000 17934 12014 17986
rect 12066 17934 12080 17986
rect 12000 17826 12080 17934
rect 12000 17774 12014 17826
rect 12066 17774 12080 17826
rect 12000 17666 12080 17774
rect 12000 17614 12014 17666
rect 12066 17614 12080 17666
rect 12000 17506 12080 17614
rect 12000 17454 12014 17506
rect 12066 17454 12080 17506
rect 12000 17346 12080 17454
rect 12000 17294 12014 17346
rect 12066 17294 12080 17346
rect 12000 17186 12080 17294
rect 12000 17134 12014 17186
rect 12066 17134 12080 17186
rect 12000 17026 12080 17134
rect 12000 16974 12014 17026
rect 12066 16974 12080 17026
rect 12000 16866 12080 16974
rect 12000 16814 12014 16866
rect 12066 16814 12080 16866
rect 12000 16697 12080 16814
rect 12000 16663 12023 16697
rect 12057 16663 12080 16697
rect 12000 16546 12080 16663
rect 12000 16494 12014 16546
rect 12066 16494 12080 16546
rect 12000 16386 12080 16494
rect 12000 16334 12014 16386
rect 12066 16334 12080 16386
rect 12000 16226 12080 16334
rect 12000 16174 12014 16226
rect 12066 16174 12080 16226
rect 12000 16066 12080 16174
rect 12000 16014 12014 16066
rect 12066 16014 12080 16066
rect 12000 15906 12080 16014
rect 12000 15854 12014 15906
rect 12066 15854 12080 15906
rect 12000 15746 12080 15854
rect 12000 15694 12014 15746
rect 12066 15694 12080 15746
rect 12000 15586 12080 15694
rect 12000 15534 12014 15586
rect 12066 15534 12080 15586
rect 12000 15426 12080 15534
rect 12000 15374 12014 15426
rect 12066 15374 12080 15426
rect 12000 15266 12080 15374
rect 12000 15214 12014 15266
rect 12066 15214 12080 15266
rect 12000 15106 12080 15214
rect 12000 15054 12014 15106
rect 12066 15054 12080 15106
rect 12000 14946 12080 15054
rect 12000 14894 12014 14946
rect 12066 14894 12080 14946
rect 12000 14786 12080 14894
rect 12000 14734 12014 14786
rect 12066 14734 12080 14786
rect 12000 14626 12080 14734
rect 12000 14574 12014 14626
rect 12066 14574 12080 14626
rect 12000 14466 12080 14574
rect 12000 14414 12014 14466
rect 12066 14414 12080 14466
rect 12000 14306 12080 14414
rect 12000 14254 12014 14306
rect 12066 14254 12080 14306
rect 12000 14146 12080 14254
rect 12000 14094 12014 14146
rect 12066 14094 12080 14146
rect 12000 13986 12080 14094
rect 12000 13934 12014 13986
rect 12066 13934 12080 13986
rect 12000 13817 12080 13934
rect 12000 13783 12023 13817
rect 12057 13783 12080 13817
rect 12000 13666 12080 13783
rect 12000 13614 12014 13666
rect 12066 13614 12080 13666
rect 12000 13506 12080 13614
rect 12000 13454 12014 13506
rect 12066 13454 12080 13506
rect 12000 13346 12080 13454
rect 12000 13294 12014 13346
rect 12066 13294 12080 13346
rect 12000 13186 12080 13294
rect 12000 13134 12014 13186
rect 12066 13134 12080 13186
rect 12000 13026 12080 13134
rect 12000 12974 12014 13026
rect 12066 12974 12080 13026
rect 12000 12866 12080 12974
rect 12000 12814 12014 12866
rect 12066 12814 12080 12866
rect 12000 12706 12080 12814
rect 12000 12654 12014 12706
rect 12066 12654 12080 12706
rect 12000 12546 12080 12654
rect 12000 12494 12014 12546
rect 12066 12494 12080 12546
rect 12000 12377 12080 12494
rect 12000 12343 12023 12377
rect 12057 12343 12080 12377
rect 12000 12217 12080 12343
rect 12000 12183 12023 12217
rect 12057 12183 12080 12217
rect 12000 12057 12080 12183
rect 12000 12023 12023 12057
rect 12057 12023 12080 12057
rect 12000 11897 12080 12023
rect 12000 11863 12023 11897
rect 12057 11863 12080 11897
rect 12000 11746 12080 11863
rect 12000 11694 12014 11746
rect 12066 11694 12080 11746
rect 12000 11586 12080 11694
rect 12000 11534 12014 11586
rect 12066 11534 12080 11586
rect 12000 11426 12080 11534
rect 12000 11374 12014 11426
rect 12066 11374 12080 11426
rect 12000 11266 12080 11374
rect 12000 11214 12014 11266
rect 12066 11214 12080 11266
rect 12000 11106 12080 11214
rect 12000 11054 12014 11106
rect 12066 11054 12080 11106
rect 12000 10946 12080 11054
rect 12000 10894 12014 10946
rect 12066 10894 12080 10946
rect 12000 10786 12080 10894
rect 12000 10734 12014 10786
rect 12066 10734 12080 10786
rect 12000 10626 12080 10734
rect 12000 10574 12014 10626
rect 12066 10574 12080 10626
rect 12000 10466 12080 10574
rect 12000 10414 12014 10466
rect 12066 10414 12080 10466
rect 12000 10306 12080 10414
rect 12000 10254 12014 10306
rect 12066 10254 12080 10306
rect 12000 10146 12080 10254
rect 12000 10094 12014 10146
rect 12066 10094 12080 10146
rect 12000 9986 12080 10094
rect 12000 9934 12014 9986
rect 12066 9934 12080 9986
rect 12000 9826 12080 9934
rect 12000 9774 12014 9826
rect 12066 9774 12080 9826
rect 12000 9657 12080 9774
rect 12000 9623 12023 9657
rect 12057 9623 12080 9657
rect 12000 9506 12080 9623
rect 12000 9454 12014 9506
rect 12066 9454 12080 9506
rect 12000 9346 12080 9454
rect 12000 9294 12014 9346
rect 12066 9294 12080 9346
rect 12000 9177 12080 9294
rect 12000 9143 12023 9177
rect 12057 9143 12080 9177
rect 12000 9026 12080 9143
rect 12000 8974 12014 9026
rect 12066 8974 12080 9026
rect 12000 8866 12080 8974
rect 12000 8814 12014 8866
rect 12066 8814 12080 8866
rect 12000 8706 12080 8814
rect 12000 8654 12014 8706
rect 12066 8654 12080 8706
rect 12000 8546 12080 8654
rect 12000 8494 12014 8546
rect 12066 8494 12080 8546
rect 12000 8386 12080 8494
rect 12000 8334 12014 8386
rect 12066 8334 12080 8386
rect 12000 8226 12080 8334
rect 12000 8174 12014 8226
rect 12066 8174 12080 8226
rect 12000 8066 12080 8174
rect 12000 8014 12014 8066
rect 12066 8014 12080 8066
rect 12000 7906 12080 8014
rect 12000 7854 12014 7906
rect 12066 7854 12080 7906
rect 12000 7746 12080 7854
rect 12000 7694 12014 7746
rect 12066 7694 12080 7746
rect 12000 7577 12080 7694
rect 12000 7543 12023 7577
rect 12057 7543 12080 7577
rect 12000 7426 12080 7543
rect 12000 7374 12014 7426
rect 12066 7374 12080 7426
rect 12000 7266 12080 7374
rect 12000 7214 12014 7266
rect 12066 7214 12080 7266
rect 12000 7097 12080 7214
rect 12000 7063 12023 7097
rect 12057 7063 12080 7097
rect 12000 6946 12080 7063
rect 12000 6894 12014 6946
rect 12066 6894 12080 6946
rect 12000 6786 12080 6894
rect 12000 6734 12014 6786
rect 12066 6734 12080 6786
rect 12000 6617 12080 6734
rect 12000 6583 12023 6617
rect 12057 6583 12080 6617
rect 12000 6466 12080 6583
rect 12000 6414 12014 6466
rect 12066 6414 12080 6466
rect 12000 6306 12080 6414
rect 12000 6254 12014 6306
rect 12066 6254 12080 6306
rect 12000 6146 12080 6254
rect 12000 6094 12014 6146
rect 12066 6094 12080 6146
rect 12000 5986 12080 6094
rect 12000 5934 12014 5986
rect 12066 5934 12080 5986
rect 12000 5826 12080 5934
rect 12000 5774 12014 5826
rect 12066 5774 12080 5826
rect 12000 5666 12080 5774
rect 12000 5614 12014 5666
rect 12066 5614 12080 5666
rect 12000 5506 12080 5614
rect 12000 5454 12014 5506
rect 12066 5454 12080 5506
rect 12000 5346 12080 5454
rect 12000 5294 12014 5346
rect 12066 5294 12080 5346
rect 12000 5186 12080 5294
rect 12000 5134 12014 5186
rect 12066 5134 12080 5186
rect 12000 5026 12080 5134
rect 12000 4974 12014 5026
rect 12066 4974 12080 5026
rect 12000 4866 12080 4974
rect 12000 4814 12014 4866
rect 12066 4814 12080 4866
rect 12000 4706 12080 4814
rect 12000 4654 12014 4706
rect 12066 4654 12080 4706
rect 12000 4546 12080 4654
rect 12000 4494 12014 4546
rect 12066 4494 12080 4546
rect 12000 4386 12080 4494
rect 12000 4334 12014 4386
rect 12066 4334 12080 4386
rect 12000 4226 12080 4334
rect 12000 4174 12014 4226
rect 12066 4174 12080 4226
rect 12000 4066 12080 4174
rect 12000 4014 12014 4066
rect 12066 4014 12080 4066
rect 12000 3906 12080 4014
rect 12000 3854 12014 3906
rect 12066 3854 12080 3906
rect 12000 3737 12080 3854
rect 12000 3703 12023 3737
rect 12057 3703 12080 3737
rect 12000 3577 12080 3703
rect 12000 3543 12023 3577
rect 12057 3543 12080 3577
rect 12000 3426 12080 3543
rect 12000 3374 12014 3426
rect 12066 3374 12080 3426
rect 12000 3266 12080 3374
rect 12000 3214 12014 3266
rect 12066 3214 12080 3266
rect 12000 3106 12080 3214
rect 12000 3054 12014 3106
rect 12066 3054 12080 3106
rect 12000 2946 12080 3054
rect 12000 2894 12014 2946
rect 12066 2894 12080 2946
rect 12000 2786 12080 2894
rect 12000 2734 12014 2786
rect 12066 2734 12080 2786
rect 12000 2626 12080 2734
rect 12000 2574 12014 2626
rect 12066 2574 12080 2626
rect 12000 2466 12080 2574
rect 12000 2414 12014 2466
rect 12066 2414 12080 2466
rect 12000 2306 12080 2414
rect 12000 2254 12014 2306
rect 12066 2254 12080 2306
rect 12000 2146 12080 2254
rect 12000 2094 12014 2146
rect 12066 2094 12080 2146
rect 12000 1986 12080 2094
rect 12000 1934 12014 1986
rect 12066 1934 12080 1986
rect 12000 1817 12080 1934
rect 12000 1783 12023 1817
rect 12057 1783 12080 1817
rect 12000 1666 12080 1783
rect 12000 1614 12014 1666
rect 12066 1614 12080 1666
rect 12000 1506 12080 1614
rect 12000 1454 12014 1506
rect 12066 1454 12080 1506
rect 12000 1346 12080 1454
rect 12000 1294 12014 1346
rect 12066 1294 12080 1346
rect 12000 1186 12080 1294
rect 12000 1134 12014 1186
rect 12066 1134 12080 1186
rect 12000 1026 12080 1134
rect 12000 974 12014 1026
rect 12066 974 12080 1026
rect 12000 857 12080 974
rect 12000 823 12023 857
rect 12057 823 12080 857
rect 12000 697 12080 823
rect 12000 663 12023 697
rect 12057 663 12080 697
rect 12000 546 12080 663
rect 12000 494 12014 546
rect 12066 494 12080 546
rect 12000 386 12080 494
rect 12000 334 12014 386
rect 12066 334 12080 386
rect 12000 226 12080 334
rect 12000 174 12014 226
rect 12066 174 12080 226
rect 12000 66 12080 174
rect 12000 14 12014 66
rect 12066 14 12080 66
rect 12000 0 12080 14
rect 12160 31417 12240 31440
rect 12160 31383 12183 31417
rect 12217 31383 12240 31417
rect 12160 31257 12240 31383
rect 12160 31223 12183 31257
rect 12217 31223 12240 31257
rect 12160 31097 12240 31223
rect 12160 31063 12183 31097
rect 12217 31063 12240 31097
rect 12160 30937 12240 31063
rect 12160 30903 12183 30937
rect 12217 30903 12240 30937
rect 12160 30777 12240 30903
rect 12160 30743 12183 30777
rect 12217 30743 12240 30777
rect 12160 30617 12240 30743
rect 12160 30583 12183 30617
rect 12217 30583 12240 30617
rect 12160 30457 12240 30583
rect 12160 30423 12183 30457
rect 12217 30423 12240 30457
rect 12160 30297 12240 30423
rect 12160 30263 12183 30297
rect 12217 30263 12240 30297
rect 12160 30137 12240 30263
rect 12160 30103 12183 30137
rect 12217 30103 12240 30137
rect 12160 29977 12240 30103
rect 12160 29943 12183 29977
rect 12217 29943 12240 29977
rect 12160 29817 12240 29943
rect 12160 29783 12183 29817
rect 12217 29783 12240 29817
rect 12160 29657 12240 29783
rect 12160 29623 12183 29657
rect 12217 29623 12240 29657
rect 12160 29497 12240 29623
rect 12160 29463 12183 29497
rect 12217 29463 12240 29497
rect 12160 29337 12240 29463
rect 12160 29303 12183 29337
rect 12217 29303 12240 29337
rect 12160 29177 12240 29303
rect 12160 29143 12183 29177
rect 12217 29143 12240 29177
rect 12160 29017 12240 29143
rect 12160 28983 12183 29017
rect 12217 28983 12240 29017
rect 12160 28857 12240 28983
rect 12160 28823 12183 28857
rect 12217 28823 12240 28857
rect 12160 28697 12240 28823
rect 12160 28663 12183 28697
rect 12217 28663 12240 28697
rect 12160 28537 12240 28663
rect 12160 28503 12183 28537
rect 12217 28503 12240 28537
rect 12160 28377 12240 28503
rect 12160 28343 12183 28377
rect 12217 28343 12240 28377
rect 12160 28217 12240 28343
rect 12160 28183 12183 28217
rect 12217 28183 12240 28217
rect 12160 28057 12240 28183
rect 12160 28023 12183 28057
rect 12217 28023 12240 28057
rect 12160 27897 12240 28023
rect 12160 27863 12183 27897
rect 12217 27863 12240 27897
rect 12160 27737 12240 27863
rect 12160 27703 12183 27737
rect 12217 27703 12240 27737
rect 12160 27577 12240 27703
rect 12160 27543 12183 27577
rect 12217 27543 12240 27577
rect 12160 27417 12240 27543
rect 12160 27383 12183 27417
rect 12217 27383 12240 27417
rect 12160 27257 12240 27383
rect 12160 27223 12183 27257
rect 12217 27223 12240 27257
rect 12160 27097 12240 27223
rect 12160 27063 12183 27097
rect 12217 27063 12240 27097
rect 12160 26937 12240 27063
rect 12160 26903 12183 26937
rect 12217 26903 12240 26937
rect 12160 26777 12240 26903
rect 12160 26743 12183 26777
rect 12217 26743 12240 26777
rect 12160 26617 12240 26743
rect 12160 26583 12183 26617
rect 12217 26583 12240 26617
rect 12160 26457 12240 26583
rect 12160 26423 12183 26457
rect 12217 26423 12240 26457
rect 12160 26297 12240 26423
rect 12160 26263 12183 26297
rect 12217 26263 12240 26297
rect 12160 26137 12240 26263
rect 12160 26103 12183 26137
rect 12217 26103 12240 26137
rect 12160 25977 12240 26103
rect 12160 25943 12183 25977
rect 12217 25943 12240 25977
rect 12160 25817 12240 25943
rect 12160 25783 12183 25817
rect 12217 25783 12240 25817
rect 12160 25657 12240 25783
rect 12160 25623 12183 25657
rect 12217 25623 12240 25657
rect 12160 25497 12240 25623
rect 12160 25463 12183 25497
rect 12217 25463 12240 25497
rect 12160 25337 12240 25463
rect 12160 25303 12183 25337
rect 12217 25303 12240 25337
rect 12160 25177 12240 25303
rect 12160 25143 12183 25177
rect 12217 25143 12240 25177
rect 12160 25017 12240 25143
rect 12160 24983 12183 25017
rect 12217 24983 12240 25017
rect 12160 24857 12240 24983
rect 12160 24823 12183 24857
rect 12217 24823 12240 24857
rect 12160 24697 12240 24823
rect 12160 24663 12183 24697
rect 12217 24663 12240 24697
rect 12160 24537 12240 24663
rect 12160 24503 12183 24537
rect 12217 24503 12240 24537
rect 12160 24377 12240 24503
rect 12160 24343 12183 24377
rect 12217 24343 12240 24377
rect 12160 24217 12240 24343
rect 12160 24183 12183 24217
rect 12217 24183 12240 24217
rect 12160 24057 12240 24183
rect 12160 24023 12183 24057
rect 12217 24023 12240 24057
rect 12160 23897 12240 24023
rect 12160 23863 12183 23897
rect 12217 23863 12240 23897
rect 12160 23737 12240 23863
rect 12160 23703 12183 23737
rect 12217 23703 12240 23737
rect 12160 23577 12240 23703
rect 12160 23543 12183 23577
rect 12217 23543 12240 23577
rect 12160 23417 12240 23543
rect 12160 23383 12183 23417
rect 12217 23383 12240 23417
rect 12160 23257 12240 23383
rect 12160 23223 12183 23257
rect 12217 23223 12240 23257
rect 12160 23097 12240 23223
rect 12160 23063 12183 23097
rect 12217 23063 12240 23097
rect 12160 22937 12240 23063
rect 12160 22903 12183 22937
rect 12217 22903 12240 22937
rect 12160 22777 12240 22903
rect 12160 22743 12183 22777
rect 12217 22743 12240 22777
rect 12160 22617 12240 22743
rect 12160 22583 12183 22617
rect 12217 22583 12240 22617
rect 12160 22457 12240 22583
rect 12160 22423 12183 22457
rect 12217 22423 12240 22457
rect 12160 22297 12240 22423
rect 12160 22263 12183 22297
rect 12217 22263 12240 22297
rect 12160 22137 12240 22263
rect 12160 22103 12183 22137
rect 12217 22103 12240 22137
rect 12160 21977 12240 22103
rect 12160 21943 12183 21977
rect 12217 21943 12240 21977
rect 12160 21817 12240 21943
rect 12160 21783 12183 21817
rect 12217 21783 12240 21817
rect 12160 21657 12240 21783
rect 12160 21623 12183 21657
rect 12217 21623 12240 21657
rect 12160 21497 12240 21623
rect 12160 21463 12183 21497
rect 12217 21463 12240 21497
rect 12160 21337 12240 21463
rect 12160 21303 12183 21337
rect 12217 21303 12240 21337
rect 12160 21177 12240 21303
rect 12160 21143 12183 21177
rect 12217 21143 12240 21177
rect 12160 21017 12240 21143
rect 12160 20983 12183 21017
rect 12217 20983 12240 21017
rect 12160 20857 12240 20983
rect 12160 20823 12183 20857
rect 12217 20823 12240 20857
rect 12160 20697 12240 20823
rect 12160 20663 12183 20697
rect 12217 20663 12240 20697
rect 12160 20537 12240 20663
rect 12160 20503 12183 20537
rect 12217 20503 12240 20537
rect 12160 20377 12240 20503
rect 12160 20343 12183 20377
rect 12217 20343 12240 20377
rect 12160 20217 12240 20343
rect 12160 20183 12183 20217
rect 12217 20183 12240 20217
rect 12160 20057 12240 20183
rect 12160 20023 12183 20057
rect 12217 20023 12240 20057
rect 12160 19897 12240 20023
rect 12160 19863 12183 19897
rect 12217 19863 12240 19897
rect 12160 19737 12240 19863
rect 12160 19703 12183 19737
rect 12217 19703 12240 19737
rect 12160 19577 12240 19703
rect 12160 19543 12183 19577
rect 12217 19543 12240 19577
rect 12160 19417 12240 19543
rect 12160 19383 12183 19417
rect 12217 19383 12240 19417
rect 12160 19257 12240 19383
rect 12160 19223 12183 19257
rect 12217 19223 12240 19257
rect 12160 19097 12240 19223
rect 12160 19063 12183 19097
rect 12217 19063 12240 19097
rect 12160 18937 12240 19063
rect 12160 18903 12183 18937
rect 12217 18903 12240 18937
rect 12160 18777 12240 18903
rect 12160 18743 12183 18777
rect 12217 18743 12240 18777
rect 12160 18617 12240 18743
rect 12160 18583 12183 18617
rect 12217 18583 12240 18617
rect 12160 18457 12240 18583
rect 12160 18423 12183 18457
rect 12217 18423 12240 18457
rect 12160 18297 12240 18423
rect 12160 18263 12183 18297
rect 12217 18263 12240 18297
rect 12160 18137 12240 18263
rect 12160 18103 12183 18137
rect 12217 18103 12240 18137
rect 12160 17977 12240 18103
rect 12160 17943 12183 17977
rect 12217 17943 12240 17977
rect 12160 17817 12240 17943
rect 12160 17783 12183 17817
rect 12217 17783 12240 17817
rect 12160 17657 12240 17783
rect 12160 17623 12183 17657
rect 12217 17623 12240 17657
rect 12160 17497 12240 17623
rect 12160 17463 12183 17497
rect 12217 17463 12240 17497
rect 12160 17337 12240 17463
rect 12160 17303 12183 17337
rect 12217 17303 12240 17337
rect 12160 17177 12240 17303
rect 12160 17143 12183 17177
rect 12217 17143 12240 17177
rect 12160 17017 12240 17143
rect 12160 16983 12183 17017
rect 12217 16983 12240 17017
rect 12160 16857 12240 16983
rect 12160 16823 12183 16857
rect 12217 16823 12240 16857
rect 12160 16697 12240 16823
rect 12160 16663 12183 16697
rect 12217 16663 12240 16697
rect 12160 16537 12240 16663
rect 12160 16503 12183 16537
rect 12217 16503 12240 16537
rect 12160 16377 12240 16503
rect 12160 16343 12183 16377
rect 12217 16343 12240 16377
rect 12160 16217 12240 16343
rect 12160 16183 12183 16217
rect 12217 16183 12240 16217
rect 12160 16057 12240 16183
rect 12160 16023 12183 16057
rect 12217 16023 12240 16057
rect 12160 15897 12240 16023
rect 12160 15863 12183 15897
rect 12217 15863 12240 15897
rect 12160 15737 12240 15863
rect 12160 15703 12183 15737
rect 12217 15703 12240 15737
rect 12160 15577 12240 15703
rect 12160 15543 12183 15577
rect 12217 15543 12240 15577
rect 12160 15417 12240 15543
rect 12160 15383 12183 15417
rect 12217 15383 12240 15417
rect 12160 15257 12240 15383
rect 12160 15223 12183 15257
rect 12217 15223 12240 15257
rect 12160 15097 12240 15223
rect 12160 15063 12183 15097
rect 12217 15063 12240 15097
rect 12160 14937 12240 15063
rect 12160 14903 12183 14937
rect 12217 14903 12240 14937
rect 12160 14777 12240 14903
rect 12160 14743 12183 14777
rect 12217 14743 12240 14777
rect 12160 14617 12240 14743
rect 12160 14583 12183 14617
rect 12217 14583 12240 14617
rect 12160 14457 12240 14583
rect 12160 14423 12183 14457
rect 12217 14423 12240 14457
rect 12160 14297 12240 14423
rect 12160 14263 12183 14297
rect 12217 14263 12240 14297
rect 12160 14137 12240 14263
rect 12160 14103 12183 14137
rect 12217 14103 12240 14137
rect 12160 13977 12240 14103
rect 12160 13943 12183 13977
rect 12217 13943 12240 13977
rect 12160 13817 12240 13943
rect 12160 13783 12183 13817
rect 12217 13783 12240 13817
rect 12160 13657 12240 13783
rect 12160 13623 12183 13657
rect 12217 13623 12240 13657
rect 12160 13497 12240 13623
rect 12160 13463 12183 13497
rect 12217 13463 12240 13497
rect 12160 13337 12240 13463
rect 12160 13303 12183 13337
rect 12217 13303 12240 13337
rect 12160 13177 12240 13303
rect 12160 13143 12183 13177
rect 12217 13143 12240 13177
rect 12160 13017 12240 13143
rect 12160 12983 12183 13017
rect 12217 12983 12240 13017
rect 12160 12857 12240 12983
rect 12160 12823 12183 12857
rect 12217 12823 12240 12857
rect 12160 12697 12240 12823
rect 12160 12663 12183 12697
rect 12217 12663 12240 12697
rect 12160 12537 12240 12663
rect 12160 12503 12183 12537
rect 12217 12503 12240 12537
rect 12160 12377 12240 12503
rect 12160 12343 12183 12377
rect 12217 12343 12240 12377
rect 12160 12217 12240 12343
rect 12160 12183 12183 12217
rect 12217 12183 12240 12217
rect 12160 12057 12240 12183
rect 12160 12023 12183 12057
rect 12217 12023 12240 12057
rect 12160 11897 12240 12023
rect 12160 11863 12183 11897
rect 12217 11863 12240 11897
rect 12160 11737 12240 11863
rect 12160 11703 12183 11737
rect 12217 11703 12240 11737
rect 12160 11577 12240 11703
rect 12160 11543 12183 11577
rect 12217 11543 12240 11577
rect 12160 11417 12240 11543
rect 12160 11383 12183 11417
rect 12217 11383 12240 11417
rect 12160 11257 12240 11383
rect 12160 11223 12183 11257
rect 12217 11223 12240 11257
rect 12160 11097 12240 11223
rect 12160 11063 12183 11097
rect 12217 11063 12240 11097
rect 12160 10937 12240 11063
rect 12160 10903 12183 10937
rect 12217 10903 12240 10937
rect 12160 10777 12240 10903
rect 12160 10743 12183 10777
rect 12217 10743 12240 10777
rect 12160 10617 12240 10743
rect 12160 10583 12183 10617
rect 12217 10583 12240 10617
rect 12160 10457 12240 10583
rect 12160 10423 12183 10457
rect 12217 10423 12240 10457
rect 12160 10297 12240 10423
rect 12160 10263 12183 10297
rect 12217 10263 12240 10297
rect 12160 10137 12240 10263
rect 12160 10103 12183 10137
rect 12217 10103 12240 10137
rect 12160 9977 12240 10103
rect 12160 9943 12183 9977
rect 12217 9943 12240 9977
rect 12160 9817 12240 9943
rect 12160 9783 12183 9817
rect 12217 9783 12240 9817
rect 12160 9657 12240 9783
rect 12160 9623 12183 9657
rect 12217 9623 12240 9657
rect 12160 9497 12240 9623
rect 12160 9463 12183 9497
rect 12217 9463 12240 9497
rect 12160 9337 12240 9463
rect 12160 9303 12183 9337
rect 12217 9303 12240 9337
rect 12160 9177 12240 9303
rect 12160 9143 12183 9177
rect 12217 9143 12240 9177
rect 12160 9017 12240 9143
rect 12160 8983 12183 9017
rect 12217 8983 12240 9017
rect 12160 8857 12240 8983
rect 12160 8823 12183 8857
rect 12217 8823 12240 8857
rect 12160 8697 12240 8823
rect 12160 8663 12183 8697
rect 12217 8663 12240 8697
rect 12160 8537 12240 8663
rect 12160 8503 12183 8537
rect 12217 8503 12240 8537
rect 12160 8377 12240 8503
rect 12160 8343 12183 8377
rect 12217 8343 12240 8377
rect 12160 8217 12240 8343
rect 12160 8183 12183 8217
rect 12217 8183 12240 8217
rect 12160 8057 12240 8183
rect 12160 8023 12183 8057
rect 12217 8023 12240 8057
rect 12160 7897 12240 8023
rect 12160 7863 12183 7897
rect 12217 7863 12240 7897
rect 12160 7737 12240 7863
rect 12160 7703 12183 7737
rect 12217 7703 12240 7737
rect 12160 7577 12240 7703
rect 12160 7543 12183 7577
rect 12217 7543 12240 7577
rect 12160 7417 12240 7543
rect 12160 7383 12183 7417
rect 12217 7383 12240 7417
rect 12160 7257 12240 7383
rect 12160 7223 12183 7257
rect 12217 7223 12240 7257
rect 12160 7097 12240 7223
rect 12160 7063 12183 7097
rect 12217 7063 12240 7097
rect 12160 6937 12240 7063
rect 12160 6903 12183 6937
rect 12217 6903 12240 6937
rect 12160 6777 12240 6903
rect 12160 6743 12183 6777
rect 12217 6743 12240 6777
rect 12160 6617 12240 6743
rect 12160 6583 12183 6617
rect 12217 6583 12240 6617
rect 12160 6457 12240 6583
rect 12160 6423 12183 6457
rect 12217 6423 12240 6457
rect 12160 6297 12240 6423
rect 12160 6263 12183 6297
rect 12217 6263 12240 6297
rect 12160 6137 12240 6263
rect 12160 6103 12183 6137
rect 12217 6103 12240 6137
rect 12160 5977 12240 6103
rect 12160 5943 12183 5977
rect 12217 5943 12240 5977
rect 12160 5817 12240 5943
rect 12160 5783 12183 5817
rect 12217 5783 12240 5817
rect 12160 5657 12240 5783
rect 12160 5623 12183 5657
rect 12217 5623 12240 5657
rect 12160 5497 12240 5623
rect 12160 5463 12183 5497
rect 12217 5463 12240 5497
rect 12160 5337 12240 5463
rect 12160 5303 12183 5337
rect 12217 5303 12240 5337
rect 12160 5177 12240 5303
rect 12160 5143 12183 5177
rect 12217 5143 12240 5177
rect 12160 5017 12240 5143
rect 12160 4983 12183 5017
rect 12217 4983 12240 5017
rect 12160 4857 12240 4983
rect 12160 4823 12183 4857
rect 12217 4823 12240 4857
rect 12160 4697 12240 4823
rect 12160 4663 12183 4697
rect 12217 4663 12240 4697
rect 12160 4537 12240 4663
rect 12160 4503 12183 4537
rect 12217 4503 12240 4537
rect 12160 4377 12240 4503
rect 12160 4343 12183 4377
rect 12217 4343 12240 4377
rect 12160 4217 12240 4343
rect 12160 4183 12183 4217
rect 12217 4183 12240 4217
rect 12160 4057 12240 4183
rect 12160 4023 12183 4057
rect 12217 4023 12240 4057
rect 12160 3897 12240 4023
rect 12160 3863 12183 3897
rect 12217 3863 12240 3897
rect 12160 3737 12240 3863
rect 12160 3703 12183 3737
rect 12217 3703 12240 3737
rect 12160 3577 12240 3703
rect 12160 3543 12183 3577
rect 12217 3543 12240 3577
rect 12160 3417 12240 3543
rect 12160 3383 12183 3417
rect 12217 3383 12240 3417
rect 12160 3257 12240 3383
rect 12160 3223 12183 3257
rect 12217 3223 12240 3257
rect 12160 3097 12240 3223
rect 12160 3063 12183 3097
rect 12217 3063 12240 3097
rect 12160 2937 12240 3063
rect 12160 2903 12183 2937
rect 12217 2903 12240 2937
rect 12160 2777 12240 2903
rect 12160 2743 12183 2777
rect 12217 2743 12240 2777
rect 12160 2617 12240 2743
rect 12160 2583 12183 2617
rect 12217 2583 12240 2617
rect 12160 2457 12240 2583
rect 12160 2423 12183 2457
rect 12217 2423 12240 2457
rect 12160 2297 12240 2423
rect 12160 2263 12183 2297
rect 12217 2263 12240 2297
rect 12160 2137 12240 2263
rect 12160 2103 12183 2137
rect 12217 2103 12240 2137
rect 12160 1977 12240 2103
rect 12160 1943 12183 1977
rect 12217 1943 12240 1977
rect 12160 1817 12240 1943
rect 12160 1783 12183 1817
rect 12217 1783 12240 1817
rect 12160 1657 12240 1783
rect 12160 1623 12183 1657
rect 12217 1623 12240 1657
rect 12160 1497 12240 1623
rect 12160 1463 12183 1497
rect 12217 1463 12240 1497
rect 12160 1337 12240 1463
rect 12160 1303 12183 1337
rect 12217 1303 12240 1337
rect 12160 1177 12240 1303
rect 12160 1143 12183 1177
rect 12217 1143 12240 1177
rect 12160 1017 12240 1143
rect 12160 983 12183 1017
rect 12217 983 12240 1017
rect 12160 857 12240 983
rect 12160 823 12183 857
rect 12217 823 12240 857
rect 12160 697 12240 823
rect 12160 663 12183 697
rect 12217 663 12240 697
rect 12160 537 12240 663
rect 12160 503 12183 537
rect 12217 503 12240 537
rect 12160 377 12240 503
rect 12160 343 12183 377
rect 12217 343 12240 377
rect 12160 217 12240 343
rect 12160 183 12183 217
rect 12217 183 12240 217
rect 12160 57 12240 183
rect 12160 23 12183 57
rect 12217 23 12240 57
rect 12160 0 12240 23
rect 12320 31426 12400 31440
rect 12320 31374 12334 31426
rect 12386 31374 12400 31426
rect 12320 31266 12400 31374
rect 12320 31214 12334 31266
rect 12386 31214 12400 31266
rect 12320 31106 12400 31214
rect 12320 31054 12334 31106
rect 12386 31054 12400 31106
rect 12320 30946 12400 31054
rect 12320 30894 12334 30946
rect 12386 30894 12400 30946
rect 12320 30786 12400 30894
rect 12320 30734 12334 30786
rect 12386 30734 12400 30786
rect 12320 30626 12400 30734
rect 12320 30574 12334 30626
rect 12386 30574 12400 30626
rect 12320 30466 12400 30574
rect 12320 30414 12334 30466
rect 12386 30414 12400 30466
rect 12320 30306 12400 30414
rect 12320 30254 12334 30306
rect 12386 30254 12400 30306
rect 12320 30137 12400 30254
rect 12320 30103 12343 30137
rect 12377 30103 12400 30137
rect 12320 29986 12400 30103
rect 12320 29934 12334 29986
rect 12386 29934 12400 29986
rect 12320 29826 12400 29934
rect 12320 29774 12334 29826
rect 12386 29774 12400 29826
rect 12320 29666 12400 29774
rect 12320 29614 12334 29666
rect 12386 29614 12400 29666
rect 12320 29506 12400 29614
rect 12320 29454 12334 29506
rect 12386 29454 12400 29506
rect 12320 29346 12400 29454
rect 12320 29294 12334 29346
rect 12386 29294 12400 29346
rect 12320 29186 12400 29294
rect 12320 29134 12334 29186
rect 12386 29134 12400 29186
rect 12320 29026 12400 29134
rect 12320 28974 12334 29026
rect 12386 28974 12400 29026
rect 12320 28866 12400 28974
rect 12320 28814 12334 28866
rect 12386 28814 12400 28866
rect 12320 28697 12400 28814
rect 12320 28663 12343 28697
rect 12377 28663 12400 28697
rect 12320 28537 12400 28663
rect 12320 28503 12343 28537
rect 12377 28503 12400 28537
rect 12320 28377 12400 28503
rect 12320 28343 12343 28377
rect 12377 28343 12400 28377
rect 12320 28217 12400 28343
rect 12320 28183 12343 28217
rect 12377 28183 12400 28217
rect 12320 28066 12400 28183
rect 12320 28014 12334 28066
rect 12386 28014 12400 28066
rect 12320 27906 12400 28014
rect 12320 27854 12334 27906
rect 12386 27854 12400 27906
rect 12320 27746 12400 27854
rect 12320 27694 12334 27746
rect 12386 27694 12400 27746
rect 12320 27586 12400 27694
rect 12320 27534 12334 27586
rect 12386 27534 12400 27586
rect 12320 27426 12400 27534
rect 12320 27374 12334 27426
rect 12386 27374 12400 27426
rect 12320 27266 12400 27374
rect 12320 27214 12334 27266
rect 12386 27214 12400 27266
rect 12320 27106 12400 27214
rect 12320 27054 12334 27106
rect 12386 27054 12400 27106
rect 12320 26946 12400 27054
rect 12320 26894 12334 26946
rect 12386 26894 12400 26946
rect 12320 26777 12400 26894
rect 12320 26743 12343 26777
rect 12377 26743 12400 26777
rect 12320 26617 12400 26743
rect 12320 26583 12343 26617
rect 12377 26583 12400 26617
rect 12320 26457 12400 26583
rect 12320 26423 12343 26457
rect 12377 26423 12400 26457
rect 12320 26297 12400 26423
rect 12320 26263 12343 26297
rect 12377 26263 12400 26297
rect 12320 26146 12400 26263
rect 12320 26094 12334 26146
rect 12386 26094 12400 26146
rect 12320 25986 12400 26094
rect 12320 25934 12334 25986
rect 12386 25934 12400 25986
rect 12320 25826 12400 25934
rect 12320 25774 12334 25826
rect 12386 25774 12400 25826
rect 12320 25666 12400 25774
rect 12320 25614 12334 25666
rect 12386 25614 12400 25666
rect 12320 25506 12400 25614
rect 12320 25454 12334 25506
rect 12386 25454 12400 25506
rect 12320 25346 12400 25454
rect 12320 25294 12334 25346
rect 12386 25294 12400 25346
rect 12320 25186 12400 25294
rect 12320 25134 12334 25186
rect 12386 25134 12400 25186
rect 12320 25026 12400 25134
rect 12320 24974 12334 25026
rect 12386 24974 12400 25026
rect 12320 24857 12400 24974
rect 12320 24823 12343 24857
rect 12377 24823 12400 24857
rect 12320 24706 12400 24823
rect 12320 24654 12334 24706
rect 12386 24654 12400 24706
rect 12320 24546 12400 24654
rect 12320 24494 12334 24546
rect 12386 24494 12400 24546
rect 12320 24386 12400 24494
rect 12320 24334 12334 24386
rect 12386 24334 12400 24386
rect 12320 24226 12400 24334
rect 12320 24174 12334 24226
rect 12386 24174 12400 24226
rect 12320 24066 12400 24174
rect 12320 24014 12334 24066
rect 12386 24014 12400 24066
rect 12320 23906 12400 24014
rect 12320 23854 12334 23906
rect 12386 23854 12400 23906
rect 12320 23746 12400 23854
rect 12320 23694 12334 23746
rect 12386 23694 12400 23746
rect 12320 23586 12400 23694
rect 12320 23534 12334 23586
rect 12386 23534 12400 23586
rect 12320 23426 12400 23534
rect 12320 23374 12334 23426
rect 12386 23374 12400 23426
rect 12320 23266 12400 23374
rect 12320 23214 12334 23266
rect 12386 23214 12400 23266
rect 12320 23106 12400 23214
rect 12320 23054 12334 23106
rect 12386 23054 12400 23106
rect 12320 22946 12400 23054
rect 12320 22894 12334 22946
rect 12386 22894 12400 22946
rect 12320 22786 12400 22894
rect 12320 22734 12334 22786
rect 12386 22734 12400 22786
rect 12320 22626 12400 22734
rect 12320 22574 12334 22626
rect 12386 22574 12400 22626
rect 12320 22466 12400 22574
rect 12320 22414 12334 22466
rect 12386 22414 12400 22466
rect 12320 22306 12400 22414
rect 12320 22254 12334 22306
rect 12386 22254 12400 22306
rect 12320 22146 12400 22254
rect 12320 22094 12334 22146
rect 12386 22094 12400 22146
rect 12320 21977 12400 22094
rect 12320 21943 12343 21977
rect 12377 21943 12400 21977
rect 12320 21826 12400 21943
rect 12320 21774 12334 21826
rect 12386 21774 12400 21826
rect 12320 21666 12400 21774
rect 12320 21614 12334 21666
rect 12386 21614 12400 21666
rect 12320 21506 12400 21614
rect 12320 21454 12334 21506
rect 12386 21454 12400 21506
rect 12320 21346 12400 21454
rect 12320 21294 12334 21346
rect 12386 21294 12400 21346
rect 12320 21186 12400 21294
rect 12320 21134 12334 21186
rect 12386 21134 12400 21186
rect 12320 21026 12400 21134
rect 12320 20974 12334 21026
rect 12386 20974 12400 21026
rect 12320 20866 12400 20974
rect 12320 20814 12334 20866
rect 12386 20814 12400 20866
rect 12320 20706 12400 20814
rect 12320 20654 12334 20706
rect 12386 20654 12400 20706
rect 12320 20537 12400 20654
rect 12320 20503 12343 20537
rect 12377 20503 12400 20537
rect 12320 20377 12400 20503
rect 12320 20343 12343 20377
rect 12377 20343 12400 20377
rect 12320 20217 12400 20343
rect 12320 20183 12343 20217
rect 12377 20183 12400 20217
rect 12320 20057 12400 20183
rect 12320 20023 12343 20057
rect 12377 20023 12400 20057
rect 12320 19906 12400 20023
rect 12320 19854 12334 19906
rect 12386 19854 12400 19906
rect 12320 19746 12400 19854
rect 12320 19694 12334 19746
rect 12386 19694 12400 19746
rect 12320 19586 12400 19694
rect 12320 19534 12334 19586
rect 12386 19534 12400 19586
rect 12320 19426 12400 19534
rect 12320 19374 12334 19426
rect 12386 19374 12400 19426
rect 12320 19266 12400 19374
rect 12320 19214 12334 19266
rect 12386 19214 12400 19266
rect 12320 19106 12400 19214
rect 12320 19054 12334 19106
rect 12386 19054 12400 19106
rect 12320 18946 12400 19054
rect 12320 18894 12334 18946
rect 12386 18894 12400 18946
rect 12320 18786 12400 18894
rect 12320 18734 12334 18786
rect 12386 18734 12400 18786
rect 12320 18617 12400 18734
rect 12320 18583 12343 18617
rect 12377 18583 12400 18617
rect 12320 18457 12400 18583
rect 12320 18423 12343 18457
rect 12377 18423 12400 18457
rect 12320 18297 12400 18423
rect 12320 18263 12343 18297
rect 12377 18263 12400 18297
rect 12320 18137 12400 18263
rect 12320 18103 12343 18137
rect 12377 18103 12400 18137
rect 12320 17986 12400 18103
rect 12320 17934 12334 17986
rect 12386 17934 12400 17986
rect 12320 17826 12400 17934
rect 12320 17774 12334 17826
rect 12386 17774 12400 17826
rect 12320 17666 12400 17774
rect 12320 17614 12334 17666
rect 12386 17614 12400 17666
rect 12320 17506 12400 17614
rect 12320 17454 12334 17506
rect 12386 17454 12400 17506
rect 12320 17346 12400 17454
rect 12320 17294 12334 17346
rect 12386 17294 12400 17346
rect 12320 17186 12400 17294
rect 12320 17134 12334 17186
rect 12386 17134 12400 17186
rect 12320 17026 12400 17134
rect 12320 16974 12334 17026
rect 12386 16974 12400 17026
rect 12320 16866 12400 16974
rect 12320 16814 12334 16866
rect 12386 16814 12400 16866
rect 12320 16697 12400 16814
rect 12320 16663 12343 16697
rect 12377 16663 12400 16697
rect 12320 16546 12400 16663
rect 12320 16494 12334 16546
rect 12386 16494 12400 16546
rect 12320 16386 12400 16494
rect 12320 16334 12334 16386
rect 12386 16334 12400 16386
rect 12320 16226 12400 16334
rect 12320 16174 12334 16226
rect 12386 16174 12400 16226
rect 12320 16066 12400 16174
rect 12320 16014 12334 16066
rect 12386 16014 12400 16066
rect 12320 15906 12400 16014
rect 12320 15854 12334 15906
rect 12386 15854 12400 15906
rect 12320 15746 12400 15854
rect 12320 15694 12334 15746
rect 12386 15694 12400 15746
rect 12320 15586 12400 15694
rect 12320 15534 12334 15586
rect 12386 15534 12400 15586
rect 12320 15426 12400 15534
rect 12320 15374 12334 15426
rect 12386 15374 12400 15426
rect 12320 15266 12400 15374
rect 12320 15214 12334 15266
rect 12386 15214 12400 15266
rect 12320 15106 12400 15214
rect 12320 15054 12334 15106
rect 12386 15054 12400 15106
rect 12320 14946 12400 15054
rect 12320 14894 12334 14946
rect 12386 14894 12400 14946
rect 12320 14786 12400 14894
rect 12320 14734 12334 14786
rect 12386 14734 12400 14786
rect 12320 14626 12400 14734
rect 12320 14574 12334 14626
rect 12386 14574 12400 14626
rect 12320 14466 12400 14574
rect 12320 14414 12334 14466
rect 12386 14414 12400 14466
rect 12320 14306 12400 14414
rect 12320 14254 12334 14306
rect 12386 14254 12400 14306
rect 12320 14146 12400 14254
rect 12320 14094 12334 14146
rect 12386 14094 12400 14146
rect 12320 13986 12400 14094
rect 12320 13934 12334 13986
rect 12386 13934 12400 13986
rect 12320 13817 12400 13934
rect 12320 13783 12343 13817
rect 12377 13783 12400 13817
rect 12320 13666 12400 13783
rect 12320 13614 12334 13666
rect 12386 13614 12400 13666
rect 12320 13506 12400 13614
rect 12320 13454 12334 13506
rect 12386 13454 12400 13506
rect 12320 13346 12400 13454
rect 12320 13294 12334 13346
rect 12386 13294 12400 13346
rect 12320 13186 12400 13294
rect 12320 13134 12334 13186
rect 12386 13134 12400 13186
rect 12320 13026 12400 13134
rect 12320 12974 12334 13026
rect 12386 12974 12400 13026
rect 12320 12866 12400 12974
rect 12320 12814 12334 12866
rect 12386 12814 12400 12866
rect 12320 12706 12400 12814
rect 12320 12654 12334 12706
rect 12386 12654 12400 12706
rect 12320 12546 12400 12654
rect 12320 12494 12334 12546
rect 12386 12494 12400 12546
rect 12320 12377 12400 12494
rect 12320 12343 12343 12377
rect 12377 12343 12400 12377
rect 12320 12217 12400 12343
rect 12320 12183 12343 12217
rect 12377 12183 12400 12217
rect 12320 12057 12400 12183
rect 12320 12023 12343 12057
rect 12377 12023 12400 12057
rect 12320 11897 12400 12023
rect 12320 11863 12343 11897
rect 12377 11863 12400 11897
rect 12320 11746 12400 11863
rect 12320 11694 12334 11746
rect 12386 11694 12400 11746
rect 12320 11586 12400 11694
rect 12320 11534 12334 11586
rect 12386 11534 12400 11586
rect 12320 11426 12400 11534
rect 12320 11374 12334 11426
rect 12386 11374 12400 11426
rect 12320 11266 12400 11374
rect 12320 11214 12334 11266
rect 12386 11214 12400 11266
rect 12320 11106 12400 11214
rect 12320 11054 12334 11106
rect 12386 11054 12400 11106
rect 12320 10946 12400 11054
rect 12320 10894 12334 10946
rect 12386 10894 12400 10946
rect 12320 10786 12400 10894
rect 12320 10734 12334 10786
rect 12386 10734 12400 10786
rect 12320 10626 12400 10734
rect 12320 10574 12334 10626
rect 12386 10574 12400 10626
rect 12320 10466 12400 10574
rect 12320 10414 12334 10466
rect 12386 10414 12400 10466
rect 12320 10306 12400 10414
rect 12320 10254 12334 10306
rect 12386 10254 12400 10306
rect 12320 10146 12400 10254
rect 12320 10094 12334 10146
rect 12386 10094 12400 10146
rect 12320 9986 12400 10094
rect 12320 9934 12334 9986
rect 12386 9934 12400 9986
rect 12320 9826 12400 9934
rect 12320 9774 12334 9826
rect 12386 9774 12400 9826
rect 12320 9657 12400 9774
rect 12320 9623 12343 9657
rect 12377 9623 12400 9657
rect 12320 9506 12400 9623
rect 12320 9454 12334 9506
rect 12386 9454 12400 9506
rect 12320 9346 12400 9454
rect 12320 9294 12334 9346
rect 12386 9294 12400 9346
rect 12320 9177 12400 9294
rect 12320 9143 12343 9177
rect 12377 9143 12400 9177
rect 12320 9026 12400 9143
rect 12320 8974 12334 9026
rect 12386 8974 12400 9026
rect 12320 8866 12400 8974
rect 12320 8814 12334 8866
rect 12386 8814 12400 8866
rect 12320 8706 12400 8814
rect 12320 8654 12334 8706
rect 12386 8654 12400 8706
rect 12320 8546 12400 8654
rect 12320 8494 12334 8546
rect 12386 8494 12400 8546
rect 12320 8386 12400 8494
rect 12320 8334 12334 8386
rect 12386 8334 12400 8386
rect 12320 8226 12400 8334
rect 12320 8174 12334 8226
rect 12386 8174 12400 8226
rect 12320 8066 12400 8174
rect 12320 8014 12334 8066
rect 12386 8014 12400 8066
rect 12320 7906 12400 8014
rect 12320 7854 12334 7906
rect 12386 7854 12400 7906
rect 12320 7746 12400 7854
rect 12320 7694 12334 7746
rect 12386 7694 12400 7746
rect 12320 7577 12400 7694
rect 12320 7543 12343 7577
rect 12377 7543 12400 7577
rect 12320 7426 12400 7543
rect 12320 7374 12334 7426
rect 12386 7374 12400 7426
rect 12320 7266 12400 7374
rect 12320 7214 12334 7266
rect 12386 7214 12400 7266
rect 12320 7097 12400 7214
rect 12320 7063 12343 7097
rect 12377 7063 12400 7097
rect 12320 6946 12400 7063
rect 12320 6894 12334 6946
rect 12386 6894 12400 6946
rect 12320 6786 12400 6894
rect 12320 6734 12334 6786
rect 12386 6734 12400 6786
rect 12320 6617 12400 6734
rect 12320 6583 12343 6617
rect 12377 6583 12400 6617
rect 12320 6466 12400 6583
rect 12320 6414 12334 6466
rect 12386 6414 12400 6466
rect 12320 6306 12400 6414
rect 12320 6254 12334 6306
rect 12386 6254 12400 6306
rect 12320 6146 12400 6254
rect 12320 6094 12334 6146
rect 12386 6094 12400 6146
rect 12320 5986 12400 6094
rect 12320 5934 12334 5986
rect 12386 5934 12400 5986
rect 12320 5826 12400 5934
rect 12320 5774 12334 5826
rect 12386 5774 12400 5826
rect 12320 5666 12400 5774
rect 12320 5614 12334 5666
rect 12386 5614 12400 5666
rect 12320 5506 12400 5614
rect 12320 5454 12334 5506
rect 12386 5454 12400 5506
rect 12320 5346 12400 5454
rect 12320 5294 12334 5346
rect 12386 5294 12400 5346
rect 12320 5186 12400 5294
rect 12320 5134 12334 5186
rect 12386 5134 12400 5186
rect 12320 5026 12400 5134
rect 12320 4974 12334 5026
rect 12386 4974 12400 5026
rect 12320 4866 12400 4974
rect 12320 4814 12334 4866
rect 12386 4814 12400 4866
rect 12320 4706 12400 4814
rect 12320 4654 12334 4706
rect 12386 4654 12400 4706
rect 12320 4546 12400 4654
rect 12320 4494 12334 4546
rect 12386 4494 12400 4546
rect 12320 4386 12400 4494
rect 12320 4334 12334 4386
rect 12386 4334 12400 4386
rect 12320 4226 12400 4334
rect 12320 4174 12334 4226
rect 12386 4174 12400 4226
rect 12320 4066 12400 4174
rect 12320 4014 12334 4066
rect 12386 4014 12400 4066
rect 12320 3906 12400 4014
rect 12320 3854 12334 3906
rect 12386 3854 12400 3906
rect 12320 3737 12400 3854
rect 12320 3703 12343 3737
rect 12377 3703 12400 3737
rect 12320 3577 12400 3703
rect 12320 3543 12343 3577
rect 12377 3543 12400 3577
rect 12320 3426 12400 3543
rect 12320 3374 12334 3426
rect 12386 3374 12400 3426
rect 12320 3266 12400 3374
rect 12320 3214 12334 3266
rect 12386 3214 12400 3266
rect 12320 3106 12400 3214
rect 12320 3054 12334 3106
rect 12386 3054 12400 3106
rect 12320 2946 12400 3054
rect 12320 2894 12334 2946
rect 12386 2894 12400 2946
rect 12320 2786 12400 2894
rect 12320 2734 12334 2786
rect 12386 2734 12400 2786
rect 12320 2626 12400 2734
rect 12320 2574 12334 2626
rect 12386 2574 12400 2626
rect 12320 2466 12400 2574
rect 12320 2414 12334 2466
rect 12386 2414 12400 2466
rect 12320 2306 12400 2414
rect 12320 2254 12334 2306
rect 12386 2254 12400 2306
rect 12320 2146 12400 2254
rect 12320 2094 12334 2146
rect 12386 2094 12400 2146
rect 12320 1986 12400 2094
rect 12320 1934 12334 1986
rect 12386 1934 12400 1986
rect 12320 1817 12400 1934
rect 12320 1783 12343 1817
rect 12377 1783 12400 1817
rect 12320 1666 12400 1783
rect 12320 1614 12334 1666
rect 12386 1614 12400 1666
rect 12320 1506 12400 1614
rect 12320 1454 12334 1506
rect 12386 1454 12400 1506
rect 12320 1346 12400 1454
rect 12320 1294 12334 1346
rect 12386 1294 12400 1346
rect 12320 1186 12400 1294
rect 12320 1134 12334 1186
rect 12386 1134 12400 1186
rect 12320 1026 12400 1134
rect 12320 974 12334 1026
rect 12386 974 12400 1026
rect 12320 857 12400 974
rect 12320 823 12343 857
rect 12377 823 12400 857
rect 12320 697 12400 823
rect 12320 663 12343 697
rect 12377 663 12400 697
rect 12320 546 12400 663
rect 12320 494 12334 546
rect 12386 494 12400 546
rect 12320 386 12400 494
rect 12320 334 12334 386
rect 12386 334 12400 386
rect 12320 226 12400 334
rect 12320 174 12334 226
rect 12386 174 12400 226
rect 12320 66 12400 174
rect 12320 14 12334 66
rect 12386 14 12400 66
rect 12320 0 12400 14
<< via1 >>
rect 8494 31417 8546 31426
rect 8494 31383 8503 31417
rect 8503 31383 8537 31417
rect 8537 31383 8546 31417
rect 8494 31374 8546 31383
rect 8494 31257 8546 31266
rect 8494 31223 8503 31257
rect 8503 31223 8537 31257
rect 8537 31223 8546 31257
rect 8494 31214 8546 31223
rect 8494 31097 8546 31106
rect 8494 31063 8503 31097
rect 8503 31063 8537 31097
rect 8537 31063 8546 31097
rect 8494 31054 8546 31063
rect 8494 30937 8546 30946
rect 8494 30903 8503 30937
rect 8503 30903 8537 30937
rect 8537 30903 8546 30937
rect 8494 30894 8546 30903
rect 8494 30777 8546 30786
rect 8494 30743 8503 30777
rect 8503 30743 8537 30777
rect 8537 30743 8546 30777
rect 8494 30734 8546 30743
rect 8494 30617 8546 30626
rect 8494 30583 8503 30617
rect 8503 30583 8537 30617
rect 8537 30583 8546 30617
rect 8494 30574 8546 30583
rect 8494 30457 8546 30466
rect 8494 30423 8503 30457
rect 8503 30423 8537 30457
rect 8537 30423 8546 30457
rect 8494 30414 8546 30423
rect 8494 30297 8546 30306
rect 8494 30263 8503 30297
rect 8503 30263 8537 30297
rect 8537 30263 8546 30297
rect 8494 30254 8546 30263
rect 8494 29977 8546 29986
rect 8494 29943 8503 29977
rect 8503 29943 8537 29977
rect 8537 29943 8546 29977
rect 8494 29934 8546 29943
rect 8494 29817 8546 29826
rect 8494 29783 8503 29817
rect 8503 29783 8537 29817
rect 8537 29783 8546 29817
rect 8494 29774 8546 29783
rect 8494 29657 8546 29666
rect 8494 29623 8503 29657
rect 8503 29623 8537 29657
rect 8537 29623 8546 29657
rect 8494 29614 8546 29623
rect 8494 29497 8546 29506
rect 8494 29463 8503 29497
rect 8503 29463 8537 29497
rect 8537 29463 8546 29497
rect 8494 29454 8546 29463
rect 8494 29337 8546 29346
rect 8494 29303 8503 29337
rect 8503 29303 8537 29337
rect 8537 29303 8546 29337
rect 8494 29294 8546 29303
rect 8494 29177 8546 29186
rect 8494 29143 8503 29177
rect 8503 29143 8537 29177
rect 8537 29143 8546 29177
rect 8494 29134 8546 29143
rect 8494 29017 8546 29026
rect 8494 28983 8503 29017
rect 8503 28983 8537 29017
rect 8537 28983 8546 29017
rect 8494 28974 8546 28983
rect 8494 28857 8546 28866
rect 8494 28823 8503 28857
rect 8503 28823 8537 28857
rect 8537 28823 8546 28857
rect 8494 28814 8546 28823
rect 8494 28057 8546 28066
rect 8494 28023 8503 28057
rect 8503 28023 8537 28057
rect 8537 28023 8546 28057
rect 8494 28014 8546 28023
rect 8494 27897 8546 27906
rect 8494 27863 8503 27897
rect 8503 27863 8537 27897
rect 8537 27863 8546 27897
rect 8494 27854 8546 27863
rect 8494 27737 8546 27746
rect 8494 27703 8503 27737
rect 8503 27703 8537 27737
rect 8537 27703 8546 27737
rect 8494 27694 8546 27703
rect 8494 27577 8546 27586
rect 8494 27543 8503 27577
rect 8503 27543 8537 27577
rect 8537 27543 8546 27577
rect 8494 27534 8546 27543
rect 8494 27417 8546 27426
rect 8494 27383 8503 27417
rect 8503 27383 8537 27417
rect 8537 27383 8546 27417
rect 8494 27374 8546 27383
rect 8494 27257 8546 27266
rect 8494 27223 8503 27257
rect 8503 27223 8537 27257
rect 8537 27223 8546 27257
rect 8494 27214 8546 27223
rect 8494 27097 8546 27106
rect 8494 27063 8503 27097
rect 8503 27063 8537 27097
rect 8537 27063 8546 27097
rect 8494 27054 8546 27063
rect 8494 26937 8546 26946
rect 8494 26903 8503 26937
rect 8503 26903 8537 26937
rect 8537 26903 8546 26937
rect 8494 26894 8546 26903
rect 8494 26137 8546 26146
rect 8494 26103 8503 26137
rect 8503 26103 8537 26137
rect 8537 26103 8546 26137
rect 8494 26094 8546 26103
rect 8494 25977 8546 25986
rect 8494 25943 8503 25977
rect 8503 25943 8537 25977
rect 8537 25943 8546 25977
rect 8494 25934 8546 25943
rect 8494 25817 8546 25826
rect 8494 25783 8503 25817
rect 8503 25783 8537 25817
rect 8537 25783 8546 25817
rect 8494 25774 8546 25783
rect 8494 25657 8546 25666
rect 8494 25623 8503 25657
rect 8503 25623 8537 25657
rect 8537 25623 8546 25657
rect 8494 25614 8546 25623
rect 8494 25497 8546 25506
rect 8494 25463 8503 25497
rect 8503 25463 8537 25497
rect 8537 25463 8546 25497
rect 8494 25454 8546 25463
rect 8494 25337 8546 25346
rect 8494 25303 8503 25337
rect 8503 25303 8537 25337
rect 8537 25303 8546 25337
rect 8494 25294 8546 25303
rect 8494 25177 8546 25186
rect 8494 25143 8503 25177
rect 8503 25143 8537 25177
rect 8537 25143 8546 25177
rect 8494 25134 8546 25143
rect 8494 25017 8546 25026
rect 8494 24983 8503 25017
rect 8503 24983 8537 25017
rect 8537 24983 8546 25017
rect 8494 24974 8546 24983
rect 8494 24697 8546 24706
rect 8494 24663 8503 24697
rect 8503 24663 8537 24697
rect 8537 24663 8546 24697
rect 8494 24654 8546 24663
rect 8494 24537 8546 24546
rect 8494 24503 8503 24537
rect 8503 24503 8537 24537
rect 8537 24503 8546 24537
rect 8494 24494 8546 24503
rect 8494 24377 8546 24386
rect 8494 24343 8503 24377
rect 8503 24343 8537 24377
rect 8537 24343 8546 24377
rect 8494 24334 8546 24343
rect 8494 24217 8546 24226
rect 8494 24183 8503 24217
rect 8503 24183 8537 24217
rect 8537 24183 8546 24217
rect 8494 24174 8546 24183
rect 8494 24057 8546 24066
rect 8494 24023 8503 24057
rect 8503 24023 8537 24057
rect 8537 24023 8546 24057
rect 8494 24014 8546 24023
rect 8494 23897 8546 23906
rect 8494 23863 8503 23897
rect 8503 23863 8537 23897
rect 8537 23863 8546 23897
rect 8494 23854 8546 23863
rect 8494 23737 8546 23746
rect 8494 23703 8503 23737
rect 8503 23703 8537 23737
rect 8537 23703 8546 23737
rect 8494 23694 8546 23703
rect 8494 23577 8546 23586
rect 8494 23543 8503 23577
rect 8503 23543 8537 23577
rect 8537 23543 8546 23577
rect 8494 23534 8546 23543
rect 8494 23417 8546 23426
rect 8494 23383 8503 23417
rect 8503 23383 8537 23417
rect 8537 23383 8546 23417
rect 8494 23374 8546 23383
rect 8494 23257 8546 23266
rect 8494 23223 8503 23257
rect 8503 23223 8537 23257
rect 8537 23223 8546 23257
rect 8494 23214 8546 23223
rect 8494 23097 8546 23106
rect 8494 23063 8503 23097
rect 8503 23063 8537 23097
rect 8537 23063 8546 23097
rect 8494 23054 8546 23063
rect 8494 22937 8546 22946
rect 8494 22903 8503 22937
rect 8503 22903 8537 22937
rect 8537 22903 8546 22937
rect 8494 22894 8546 22903
rect 8494 22777 8546 22786
rect 8494 22743 8503 22777
rect 8503 22743 8537 22777
rect 8537 22743 8546 22777
rect 8494 22734 8546 22743
rect 8494 22617 8546 22626
rect 8494 22583 8503 22617
rect 8503 22583 8537 22617
rect 8537 22583 8546 22617
rect 8494 22574 8546 22583
rect 8494 22457 8546 22466
rect 8494 22423 8503 22457
rect 8503 22423 8537 22457
rect 8537 22423 8546 22457
rect 8494 22414 8546 22423
rect 8494 22297 8546 22306
rect 8494 22263 8503 22297
rect 8503 22263 8537 22297
rect 8537 22263 8546 22297
rect 8494 22254 8546 22263
rect 8494 22137 8546 22146
rect 8494 22103 8503 22137
rect 8503 22103 8537 22137
rect 8537 22103 8546 22137
rect 8494 22094 8546 22103
rect 8494 21817 8546 21826
rect 8494 21783 8503 21817
rect 8503 21783 8537 21817
rect 8537 21783 8546 21817
rect 8494 21774 8546 21783
rect 8494 21657 8546 21666
rect 8494 21623 8503 21657
rect 8503 21623 8537 21657
rect 8537 21623 8546 21657
rect 8494 21614 8546 21623
rect 8494 21497 8546 21506
rect 8494 21463 8503 21497
rect 8503 21463 8537 21497
rect 8537 21463 8546 21497
rect 8494 21454 8546 21463
rect 8494 21337 8546 21346
rect 8494 21303 8503 21337
rect 8503 21303 8537 21337
rect 8537 21303 8546 21337
rect 8494 21294 8546 21303
rect 8494 21177 8546 21186
rect 8494 21143 8503 21177
rect 8503 21143 8537 21177
rect 8537 21143 8546 21177
rect 8494 21134 8546 21143
rect 8494 21017 8546 21026
rect 8494 20983 8503 21017
rect 8503 20983 8537 21017
rect 8537 20983 8546 21017
rect 8494 20974 8546 20983
rect 8494 20857 8546 20866
rect 8494 20823 8503 20857
rect 8503 20823 8537 20857
rect 8537 20823 8546 20857
rect 8494 20814 8546 20823
rect 8494 20697 8546 20706
rect 8494 20663 8503 20697
rect 8503 20663 8537 20697
rect 8537 20663 8546 20697
rect 8494 20654 8546 20663
rect 8494 19897 8546 19906
rect 8494 19863 8503 19897
rect 8503 19863 8537 19897
rect 8537 19863 8546 19897
rect 8494 19854 8546 19863
rect 8494 19737 8546 19746
rect 8494 19703 8503 19737
rect 8503 19703 8537 19737
rect 8537 19703 8546 19737
rect 8494 19694 8546 19703
rect 8494 19577 8546 19586
rect 8494 19543 8503 19577
rect 8503 19543 8537 19577
rect 8537 19543 8546 19577
rect 8494 19534 8546 19543
rect 8494 19417 8546 19426
rect 8494 19383 8503 19417
rect 8503 19383 8537 19417
rect 8537 19383 8546 19417
rect 8494 19374 8546 19383
rect 8494 19257 8546 19266
rect 8494 19223 8503 19257
rect 8503 19223 8537 19257
rect 8537 19223 8546 19257
rect 8494 19214 8546 19223
rect 8494 19097 8546 19106
rect 8494 19063 8503 19097
rect 8503 19063 8537 19097
rect 8537 19063 8546 19097
rect 8494 19054 8546 19063
rect 8494 18937 8546 18946
rect 8494 18903 8503 18937
rect 8503 18903 8537 18937
rect 8537 18903 8546 18937
rect 8494 18894 8546 18903
rect 8494 18777 8546 18786
rect 8494 18743 8503 18777
rect 8503 18743 8537 18777
rect 8537 18743 8546 18777
rect 8494 18734 8546 18743
rect 8494 17977 8546 17986
rect 8494 17943 8503 17977
rect 8503 17943 8537 17977
rect 8537 17943 8546 17977
rect 8494 17934 8546 17943
rect 8494 17817 8546 17826
rect 8494 17783 8503 17817
rect 8503 17783 8537 17817
rect 8537 17783 8546 17817
rect 8494 17774 8546 17783
rect 8494 17657 8546 17666
rect 8494 17623 8503 17657
rect 8503 17623 8537 17657
rect 8537 17623 8546 17657
rect 8494 17614 8546 17623
rect 8494 17497 8546 17506
rect 8494 17463 8503 17497
rect 8503 17463 8537 17497
rect 8537 17463 8546 17497
rect 8494 17454 8546 17463
rect 8494 17337 8546 17346
rect 8494 17303 8503 17337
rect 8503 17303 8537 17337
rect 8537 17303 8546 17337
rect 8494 17294 8546 17303
rect 8494 17177 8546 17186
rect 8494 17143 8503 17177
rect 8503 17143 8537 17177
rect 8537 17143 8546 17177
rect 8494 17134 8546 17143
rect 8494 17017 8546 17026
rect 8494 16983 8503 17017
rect 8503 16983 8537 17017
rect 8537 16983 8546 17017
rect 8494 16974 8546 16983
rect 8494 16857 8546 16866
rect 8494 16823 8503 16857
rect 8503 16823 8537 16857
rect 8537 16823 8546 16857
rect 8494 16814 8546 16823
rect 8494 16537 8546 16546
rect 8494 16503 8503 16537
rect 8503 16503 8537 16537
rect 8537 16503 8546 16537
rect 8494 16494 8546 16503
rect 8494 16377 8546 16386
rect 8494 16343 8503 16377
rect 8503 16343 8537 16377
rect 8537 16343 8546 16377
rect 8494 16334 8546 16343
rect 8494 16217 8546 16226
rect 8494 16183 8503 16217
rect 8503 16183 8537 16217
rect 8537 16183 8546 16217
rect 8494 16174 8546 16183
rect 8494 16057 8546 16066
rect 8494 16023 8503 16057
rect 8503 16023 8537 16057
rect 8537 16023 8546 16057
rect 8494 16014 8546 16023
rect 8494 15897 8546 15906
rect 8494 15863 8503 15897
rect 8503 15863 8537 15897
rect 8537 15863 8546 15897
rect 8494 15854 8546 15863
rect 8494 15737 8546 15746
rect 8494 15703 8503 15737
rect 8503 15703 8537 15737
rect 8537 15703 8546 15737
rect 8494 15694 8546 15703
rect 8494 15577 8546 15586
rect 8494 15543 8503 15577
rect 8503 15543 8537 15577
rect 8537 15543 8546 15577
rect 8494 15534 8546 15543
rect 8494 15417 8546 15426
rect 8494 15383 8503 15417
rect 8503 15383 8537 15417
rect 8537 15383 8546 15417
rect 8494 15374 8546 15383
rect 8494 15257 8546 15266
rect 8494 15223 8503 15257
rect 8503 15223 8537 15257
rect 8537 15223 8546 15257
rect 8494 15214 8546 15223
rect 8494 15097 8546 15106
rect 8494 15063 8503 15097
rect 8503 15063 8537 15097
rect 8537 15063 8546 15097
rect 8494 15054 8546 15063
rect 8494 14937 8546 14946
rect 8494 14903 8503 14937
rect 8503 14903 8537 14937
rect 8537 14903 8546 14937
rect 8494 14894 8546 14903
rect 8494 14777 8546 14786
rect 8494 14743 8503 14777
rect 8503 14743 8537 14777
rect 8537 14743 8546 14777
rect 8494 14734 8546 14743
rect 8494 14617 8546 14626
rect 8494 14583 8503 14617
rect 8503 14583 8537 14617
rect 8537 14583 8546 14617
rect 8494 14574 8546 14583
rect 8494 14457 8546 14466
rect 8494 14423 8503 14457
rect 8503 14423 8537 14457
rect 8537 14423 8546 14457
rect 8494 14414 8546 14423
rect 8494 14297 8546 14306
rect 8494 14263 8503 14297
rect 8503 14263 8537 14297
rect 8537 14263 8546 14297
rect 8494 14254 8546 14263
rect 8494 14137 8546 14146
rect 8494 14103 8503 14137
rect 8503 14103 8537 14137
rect 8537 14103 8546 14137
rect 8494 14094 8546 14103
rect 8494 13977 8546 13986
rect 8494 13943 8503 13977
rect 8503 13943 8537 13977
rect 8537 13943 8546 13977
rect 8494 13934 8546 13943
rect 8494 13657 8546 13666
rect 8494 13623 8503 13657
rect 8503 13623 8537 13657
rect 8537 13623 8546 13657
rect 8494 13614 8546 13623
rect 8494 13497 8546 13506
rect 8494 13463 8503 13497
rect 8503 13463 8537 13497
rect 8537 13463 8546 13497
rect 8494 13454 8546 13463
rect 8494 13337 8546 13346
rect 8494 13303 8503 13337
rect 8503 13303 8537 13337
rect 8537 13303 8546 13337
rect 8494 13294 8546 13303
rect 8494 13177 8546 13186
rect 8494 13143 8503 13177
rect 8503 13143 8537 13177
rect 8537 13143 8546 13177
rect 8494 13134 8546 13143
rect 8494 13017 8546 13026
rect 8494 12983 8503 13017
rect 8503 12983 8537 13017
rect 8537 12983 8546 13017
rect 8494 12974 8546 12983
rect 8494 12857 8546 12866
rect 8494 12823 8503 12857
rect 8503 12823 8537 12857
rect 8537 12823 8546 12857
rect 8494 12814 8546 12823
rect 8494 12697 8546 12706
rect 8494 12663 8503 12697
rect 8503 12663 8537 12697
rect 8537 12663 8546 12697
rect 8494 12654 8546 12663
rect 8494 12537 8546 12546
rect 8494 12503 8503 12537
rect 8503 12503 8537 12537
rect 8537 12503 8546 12537
rect 8494 12494 8546 12503
rect 8494 11737 8546 11746
rect 8494 11703 8503 11737
rect 8503 11703 8537 11737
rect 8537 11703 8546 11737
rect 8494 11694 8546 11703
rect 8494 11577 8546 11586
rect 8494 11543 8503 11577
rect 8503 11543 8537 11577
rect 8537 11543 8546 11577
rect 8494 11534 8546 11543
rect 8494 11417 8546 11426
rect 8494 11383 8503 11417
rect 8503 11383 8537 11417
rect 8537 11383 8546 11417
rect 8494 11374 8546 11383
rect 8494 11257 8546 11266
rect 8494 11223 8503 11257
rect 8503 11223 8537 11257
rect 8537 11223 8546 11257
rect 8494 11214 8546 11223
rect 8494 11097 8546 11106
rect 8494 11063 8503 11097
rect 8503 11063 8537 11097
rect 8537 11063 8546 11097
rect 8494 11054 8546 11063
rect 8494 10937 8546 10946
rect 8494 10903 8503 10937
rect 8503 10903 8537 10937
rect 8537 10903 8546 10937
rect 8494 10894 8546 10903
rect 8494 10777 8546 10786
rect 8494 10743 8503 10777
rect 8503 10743 8537 10777
rect 8537 10743 8546 10777
rect 8494 10734 8546 10743
rect 8494 10617 8546 10626
rect 8494 10583 8503 10617
rect 8503 10583 8537 10617
rect 8537 10583 8546 10617
rect 8494 10574 8546 10583
rect 8494 10457 8546 10466
rect 8494 10423 8503 10457
rect 8503 10423 8537 10457
rect 8537 10423 8546 10457
rect 8494 10414 8546 10423
rect 8494 10297 8546 10306
rect 8494 10263 8503 10297
rect 8503 10263 8537 10297
rect 8537 10263 8546 10297
rect 8494 10254 8546 10263
rect 8494 10137 8546 10146
rect 8494 10103 8503 10137
rect 8503 10103 8537 10137
rect 8537 10103 8546 10137
rect 8494 10094 8546 10103
rect 8494 9977 8546 9986
rect 8494 9943 8503 9977
rect 8503 9943 8537 9977
rect 8537 9943 8546 9977
rect 8494 9934 8546 9943
rect 8494 9817 8546 9826
rect 8494 9783 8503 9817
rect 8503 9783 8537 9817
rect 8537 9783 8546 9817
rect 8494 9774 8546 9783
rect 8494 9497 8546 9506
rect 8494 9463 8503 9497
rect 8503 9463 8537 9497
rect 8537 9463 8546 9497
rect 8494 9454 8546 9463
rect 8494 9337 8546 9346
rect 8494 9303 8503 9337
rect 8503 9303 8537 9337
rect 8537 9303 8546 9337
rect 8494 9294 8546 9303
rect 8494 9017 8546 9026
rect 8494 8983 8503 9017
rect 8503 8983 8537 9017
rect 8537 8983 8546 9017
rect 8494 8974 8546 8983
rect 8494 8857 8546 8866
rect 8494 8823 8503 8857
rect 8503 8823 8537 8857
rect 8537 8823 8546 8857
rect 8494 8814 8546 8823
rect 8494 8697 8546 8706
rect 8494 8663 8503 8697
rect 8503 8663 8537 8697
rect 8537 8663 8546 8697
rect 8494 8654 8546 8663
rect 8494 8537 8546 8546
rect 8494 8503 8503 8537
rect 8503 8503 8537 8537
rect 8537 8503 8546 8537
rect 8494 8494 8546 8503
rect 8494 8377 8546 8386
rect 8494 8343 8503 8377
rect 8503 8343 8537 8377
rect 8537 8343 8546 8377
rect 8494 8334 8546 8343
rect 8494 8217 8546 8226
rect 8494 8183 8503 8217
rect 8503 8183 8537 8217
rect 8537 8183 8546 8217
rect 8494 8174 8546 8183
rect 8494 8057 8546 8066
rect 8494 8023 8503 8057
rect 8503 8023 8537 8057
rect 8537 8023 8546 8057
rect 8494 8014 8546 8023
rect 8494 7897 8546 7906
rect 8494 7863 8503 7897
rect 8503 7863 8537 7897
rect 8537 7863 8546 7897
rect 8494 7854 8546 7863
rect 8494 7737 8546 7746
rect 8494 7703 8503 7737
rect 8503 7703 8537 7737
rect 8537 7703 8546 7737
rect 8494 7694 8546 7703
rect 8494 7417 8546 7426
rect 8494 7383 8503 7417
rect 8503 7383 8537 7417
rect 8537 7383 8546 7417
rect 8494 7374 8546 7383
rect 8494 7257 8546 7266
rect 8494 7223 8503 7257
rect 8503 7223 8537 7257
rect 8537 7223 8546 7257
rect 8494 7214 8546 7223
rect 8494 6937 8546 6946
rect 8494 6903 8503 6937
rect 8503 6903 8537 6937
rect 8537 6903 8546 6937
rect 8494 6894 8546 6903
rect 8494 6777 8546 6786
rect 8494 6743 8503 6777
rect 8503 6743 8537 6777
rect 8537 6743 8546 6777
rect 8494 6734 8546 6743
rect 8494 6457 8546 6466
rect 8494 6423 8503 6457
rect 8503 6423 8537 6457
rect 8537 6423 8546 6457
rect 8494 6414 8546 6423
rect 8494 6297 8546 6306
rect 8494 6263 8503 6297
rect 8503 6263 8537 6297
rect 8537 6263 8546 6297
rect 8494 6254 8546 6263
rect 8494 6137 8546 6146
rect 8494 6103 8503 6137
rect 8503 6103 8537 6137
rect 8537 6103 8546 6137
rect 8494 6094 8546 6103
rect 8494 5977 8546 5986
rect 8494 5943 8503 5977
rect 8503 5943 8537 5977
rect 8537 5943 8546 5977
rect 8494 5934 8546 5943
rect 8494 5817 8546 5826
rect 8494 5783 8503 5817
rect 8503 5783 8537 5817
rect 8537 5783 8546 5817
rect 8494 5774 8546 5783
rect 8494 5657 8546 5666
rect 8494 5623 8503 5657
rect 8503 5623 8537 5657
rect 8537 5623 8546 5657
rect 8494 5614 8546 5623
rect 8494 5497 8546 5506
rect 8494 5463 8503 5497
rect 8503 5463 8537 5497
rect 8537 5463 8546 5497
rect 8494 5454 8546 5463
rect 8494 5337 8546 5346
rect 8494 5303 8503 5337
rect 8503 5303 8537 5337
rect 8537 5303 8546 5337
rect 8494 5294 8546 5303
rect 8494 5177 8546 5186
rect 8494 5143 8503 5177
rect 8503 5143 8537 5177
rect 8537 5143 8546 5177
rect 8494 5134 8546 5143
rect 8494 5017 8546 5026
rect 8494 4983 8503 5017
rect 8503 4983 8537 5017
rect 8537 4983 8546 5017
rect 8494 4974 8546 4983
rect 8494 4857 8546 4866
rect 8494 4823 8503 4857
rect 8503 4823 8537 4857
rect 8537 4823 8546 4857
rect 8494 4814 8546 4823
rect 8494 4697 8546 4706
rect 8494 4663 8503 4697
rect 8503 4663 8537 4697
rect 8537 4663 8546 4697
rect 8494 4654 8546 4663
rect 8494 4537 8546 4546
rect 8494 4503 8503 4537
rect 8503 4503 8537 4537
rect 8537 4503 8546 4537
rect 8494 4494 8546 4503
rect 8494 4377 8546 4386
rect 8494 4343 8503 4377
rect 8503 4343 8537 4377
rect 8537 4343 8546 4377
rect 8494 4334 8546 4343
rect 8494 4217 8546 4226
rect 8494 4183 8503 4217
rect 8503 4183 8537 4217
rect 8537 4183 8546 4217
rect 8494 4174 8546 4183
rect 8494 4057 8546 4066
rect 8494 4023 8503 4057
rect 8503 4023 8537 4057
rect 8537 4023 8546 4057
rect 8494 4014 8546 4023
rect 8494 3897 8546 3906
rect 8494 3863 8503 3897
rect 8503 3863 8537 3897
rect 8537 3863 8546 3897
rect 8494 3854 8546 3863
rect 8494 3417 8546 3426
rect 8494 3383 8503 3417
rect 8503 3383 8537 3417
rect 8537 3383 8546 3417
rect 8494 3374 8546 3383
rect 8494 3257 8546 3266
rect 8494 3223 8503 3257
rect 8503 3223 8537 3257
rect 8537 3223 8546 3257
rect 8494 3214 8546 3223
rect 8494 3097 8546 3106
rect 8494 3063 8503 3097
rect 8503 3063 8537 3097
rect 8537 3063 8546 3097
rect 8494 3054 8546 3063
rect 8494 2937 8546 2946
rect 8494 2903 8503 2937
rect 8503 2903 8537 2937
rect 8537 2903 8546 2937
rect 8494 2894 8546 2903
rect 8494 2777 8546 2786
rect 8494 2743 8503 2777
rect 8503 2743 8537 2777
rect 8537 2743 8546 2777
rect 8494 2734 8546 2743
rect 8494 2617 8546 2626
rect 8494 2583 8503 2617
rect 8503 2583 8537 2617
rect 8537 2583 8546 2617
rect 8494 2574 8546 2583
rect 8494 2457 8546 2466
rect 8494 2423 8503 2457
rect 8503 2423 8537 2457
rect 8537 2423 8546 2457
rect 8494 2414 8546 2423
rect 8494 2297 8546 2306
rect 8494 2263 8503 2297
rect 8503 2263 8537 2297
rect 8537 2263 8546 2297
rect 8494 2254 8546 2263
rect 8494 2137 8546 2146
rect 8494 2103 8503 2137
rect 8503 2103 8537 2137
rect 8537 2103 8546 2137
rect 8494 2094 8546 2103
rect 8494 1977 8546 1986
rect 8494 1943 8503 1977
rect 8503 1943 8537 1977
rect 8537 1943 8546 1977
rect 8494 1934 8546 1943
rect 8494 1657 8546 1666
rect 8494 1623 8503 1657
rect 8503 1623 8537 1657
rect 8537 1623 8546 1657
rect 8494 1614 8546 1623
rect 8494 1497 8546 1506
rect 8494 1463 8503 1497
rect 8503 1463 8537 1497
rect 8537 1463 8546 1497
rect 8494 1454 8546 1463
rect 8494 1337 8546 1346
rect 8494 1303 8503 1337
rect 8503 1303 8537 1337
rect 8537 1303 8546 1337
rect 8494 1294 8546 1303
rect 8494 1177 8546 1186
rect 8494 1143 8503 1177
rect 8503 1143 8537 1177
rect 8537 1143 8546 1177
rect 8494 1134 8546 1143
rect 8494 1017 8546 1026
rect 8494 983 8503 1017
rect 8503 983 8537 1017
rect 8537 983 8546 1017
rect 8494 974 8546 983
rect 8494 537 8546 546
rect 8494 503 8503 537
rect 8503 503 8537 537
rect 8537 503 8546 537
rect 8494 494 8546 503
rect 8494 377 8546 386
rect 8494 343 8503 377
rect 8503 343 8537 377
rect 8537 343 8546 377
rect 8494 334 8546 343
rect 8494 217 8546 226
rect 8494 183 8503 217
rect 8503 183 8537 217
rect 8537 183 8546 217
rect 8494 174 8546 183
rect 8494 57 8546 66
rect 8494 23 8503 57
rect 8503 23 8537 57
rect 8537 23 8546 57
rect 8494 14 8546 23
rect 8814 31417 8866 31426
rect 8814 31383 8823 31417
rect 8823 31383 8857 31417
rect 8857 31383 8866 31417
rect 8814 31374 8866 31383
rect 8814 31257 8866 31266
rect 8814 31223 8823 31257
rect 8823 31223 8857 31257
rect 8857 31223 8866 31257
rect 8814 31214 8866 31223
rect 8814 31097 8866 31106
rect 8814 31063 8823 31097
rect 8823 31063 8857 31097
rect 8857 31063 8866 31097
rect 8814 31054 8866 31063
rect 8814 30937 8866 30946
rect 8814 30903 8823 30937
rect 8823 30903 8857 30937
rect 8857 30903 8866 30937
rect 8814 30894 8866 30903
rect 8814 30777 8866 30786
rect 8814 30743 8823 30777
rect 8823 30743 8857 30777
rect 8857 30743 8866 30777
rect 8814 30734 8866 30743
rect 8814 30617 8866 30626
rect 8814 30583 8823 30617
rect 8823 30583 8857 30617
rect 8857 30583 8866 30617
rect 8814 30574 8866 30583
rect 8814 30457 8866 30466
rect 8814 30423 8823 30457
rect 8823 30423 8857 30457
rect 8857 30423 8866 30457
rect 8814 30414 8866 30423
rect 8814 30297 8866 30306
rect 8814 30263 8823 30297
rect 8823 30263 8857 30297
rect 8857 30263 8866 30297
rect 8814 30254 8866 30263
rect 8814 29977 8866 29986
rect 8814 29943 8823 29977
rect 8823 29943 8857 29977
rect 8857 29943 8866 29977
rect 8814 29934 8866 29943
rect 8814 29817 8866 29826
rect 8814 29783 8823 29817
rect 8823 29783 8857 29817
rect 8857 29783 8866 29817
rect 8814 29774 8866 29783
rect 8814 29657 8866 29666
rect 8814 29623 8823 29657
rect 8823 29623 8857 29657
rect 8857 29623 8866 29657
rect 8814 29614 8866 29623
rect 8814 29497 8866 29506
rect 8814 29463 8823 29497
rect 8823 29463 8857 29497
rect 8857 29463 8866 29497
rect 8814 29454 8866 29463
rect 8814 29337 8866 29346
rect 8814 29303 8823 29337
rect 8823 29303 8857 29337
rect 8857 29303 8866 29337
rect 8814 29294 8866 29303
rect 8814 29177 8866 29186
rect 8814 29143 8823 29177
rect 8823 29143 8857 29177
rect 8857 29143 8866 29177
rect 8814 29134 8866 29143
rect 8814 29017 8866 29026
rect 8814 28983 8823 29017
rect 8823 28983 8857 29017
rect 8857 28983 8866 29017
rect 8814 28974 8866 28983
rect 8814 28857 8866 28866
rect 8814 28823 8823 28857
rect 8823 28823 8857 28857
rect 8857 28823 8866 28857
rect 8814 28814 8866 28823
rect 8814 28057 8866 28066
rect 8814 28023 8823 28057
rect 8823 28023 8857 28057
rect 8857 28023 8866 28057
rect 8814 28014 8866 28023
rect 8814 27897 8866 27906
rect 8814 27863 8823 27897
rect 8823 27863 8857 27897
rect 8857 27863 8866 27897
rect 8814 27854 8866 27863
rect 8814 27737 8866 27746
rect 8814 27703 8823 27737
rect 8823 27703 8857 27737
rect 8857 27703 8866 27737
rect 8814 27694 8866 27703
rect 8814 27577 8866 27586
rect 8814 27543 8823 27577
rect 8823 27543 8857 27577
rect 8857 27543 8866 27577
rect 8814 27534 8866 27543
rect 8814 27417 8866 27426
rect 8814 27383 8823 27417
rect 8823 27383 8857 27417
rect 8857 27383 8866 27417
rect 8814 27374 8866 27383
rect 8814 27257 8866 27266
rect 8814 27223 8823 27257
rect 8823 27223 8857 27257
rect 8857 27223 8866 27257
rect 8814 27214 8866 27223
rect 8814 27097 8866 27106
rect 8814 27063 8823 27097
rect 8823 27063 8857 27097
rect 8857 27063 8866 27097
rect 8814 27054 8866 27063
rect 8814 26937 8866 26946
rect 8814 26903 8823 26937
rect 8823 26903 8857 26937
rect 8857 26903 8866 26937
rect 8814 26894 8866 26903
rect 8814 26137 8866 26146
rect 8814 26103 8823 26137
rect 8823 26103 8857 26137
rect 8857 26103 8866 26137
rect 8814 26094 8866 26103
rect 8814 25977 8866 25986
rect 8814 25943 8823 25977
rect 8823 25943 8857 25977
rect 8857 25943 8866 25977
rect 8814 25934 8866 25943
rect 8814 25817 8866 25826
rect 8814 25783 8823 25817
rect 8823 25783 8857 25817
rect 8857 25783 8866 25817
rect 8814 25774 8866 25783
rect 8814 25657 8866 25666
rect 8814 25623 8823 25657
rect 8823 25623 8857 25657
rect 8857 25623 8866 25657
rect 8814 25614 8866 25623
rect 8814 25497 8866 25506
rect 8814 25463 8823 25497
rect 8823 25463 8857 25497
rect 8857 25463 8866 25497
rect 8814 25454 8866 25463
rect 8814 25337 8866 25346
rect 8814 25303 8823 25337
rect 8823 25303 8857 25337
rect 8857 25303 8866 25337
rect 8814 25294 8866 25303
rect 8814 25177 8866 25186
rect 8814 25143 8823 25177
rect 8823 25143 8857 25177
rect 8857 25143 8866 25177
rect 8814 25134 8866 25143
rect 8814 25017 8866 25026
rect 8814 24983 8823 25017
rect 8823 24983 8857 25017
rect 8857 24983 8866 25017
rect 8814 24974 8866 24983
rect 8814 24697 8866 24706
rect 8814 24663 8823 24697
rect 8823 24663 8857 24697
rect 8857 24663 8866 24697
rect 8814 24654 8866 24663
rect 8814 24537 8866 24546
rect 8814 24503 8823 24537
rect 8823 24503 8857 24537
rect 8857 24503 8866 24537
rect 8814 24494 8866 24503
rect 8814 24377 8866 24386
rect 8814 24343 8823 24377
rect 8823 24343 8857 24377
rect 8857 24343 8866 24377
rect 8814 24334 8866 24343
rect 8814 24217 8866 24226
rect 8814 24183 8823 24217
rect 8823 24183 8857 24217
rect 8857 24183 8866 24217
rect 8814 24174 8866 24183
rect 8814 24057 8866 24066
rect 8814 24023 8823 24057
rect 8823 24023 8857 24057
rect 8857 24023 8866 24057
rect 8814 24014 8866 24023
rect 8814 23897 8866 23906
rect 8814 23863 8823 23897
rect 8823 23863 8857 23897
rect 8857 23863 8866 23897
rect 8814 23854 8866 23863
rect 8814 23737 8866 23746
rect 8814 23703 8823 23737
rect 8823 23703 8857 23737
rect 8857 23703 8866 23737
rect 8814 23694 8866 23703
rect 8814 23577 8866 23586
rect 8814 23543 8823 23577
rect 8823 23543 8857 23577
rect 8857 23543 8866 23577
rect 8814 23534 8866 23543
rect 8814 23417 8866 23426
rect 8814 23383 8823 23417
rect 8823 23383 8857 23417
rect 8857 23383 8866 23417
rect 8814 23374 8866 23383
rect 8814 23257 8866 23266
rect 8814 23223 8823 23257
rect 8823 23223 8857 23257
rect 8857 23223 8866 23257
rect 8814 23214 8866 23223
rect 8814 23097 8866 23106
rect 8814 23063 8823 23097
rect 8823 23063 8857 23097
rect 8857 23063 8866 23097
rect 8814 23054 8866 23063
rect 8814 22937 8866 22946
rect 8814 22903 8823 22937
rect 8823 22903 8857 22937
rect 8857 22903 8866 22937
rect 8814 22894 8866 22903
rect 8814 22777 8866 22786
rect 8814 22743 8823 22777
rect 8823 22743 8857 22777
rect 8857 22743 8866 22777
rect 8814 22734 8866 22743
rect 8814 22617 8866 22626
rect 8814 22583 8823 22617
rect 8823 22583 8857 22617
rect 8857 22583 8866 22617
rect 8814 22574 8866 22583
rect 8814 22457 8866 22466
rect 8814 22423 8823 22457
rect 8823 22423 8857 22457
rect 8857 22423 8866 22457
rect 8814 22414 8866 22423
rect 8814 22297 8866 22306
rect 8814 22263 8823 22297
rect 8823 22263 8857 22297
rect 8857 22263 8866 22297
rect 8814 22254 8866 22263
rect 8814 22137 8866 22146
rect 8814 22103 8823 22137
rect 8823 22103 8857 22137
rect 8857 22103 8866 22137
rect 8814 22094 8866 22103
rect 8814 21817 8866 21826
rect 8814 21783 8823 21817
rect 8823 21783 8857 21817
rect 8857 21783 8866 21817
rect 8814 21774 8866 21783
rect 8814 21657 8866 21666
rect 8814 21623 8823 21657
rect 8823 21623 8857 21657
rect 8857 21623 8866 21657
rect 8814 21614 8866 21623
rect 8814 21497 8866 21506
rect 8814 21463 8823 21497
rect 8823 21463 8857 21497
rect 8857 21463 8866 21497
rect 8814 21454 8866 21463
rect 8814 21337 8866 21346
rect 8814 21303 8823 21337
rect 8823 21303 8857 21337
rect 8857 21303 8866 21337
rect 8814 21294 8866 21303
rect 8814 21177 8866 21186
rect 8814 21143 8823 21177
rect 8823 21143 8857 21177
rect 8857 21143 8866 21177
rect 8814 21134 8866 21143
rect 8814 21017 8866 21026
rect 8814 20983 8823 21017
rect 8823 20983 8857 21017
rect 8857 20983 8866 21017
rect 8814 20974 8866 20983
rect 8814 20857 8866 20866
rect 8814 20823 8823 20857
rect 8823 20823 8857 20857
rect 8857 20823 8866 20857
rect 8814 20814 8866 20823
rect 8814 20697 8866 20706
rect 8814 20663 8823 20697
rect 8823 20663 8857 20697
rect 8857 20663 8866 20697
rect 8814 20654 8866 20663
rect 8814 19897 8866 19906
rect 8814 19863 8823 19897
rect 8823 19863 8857 19897
rect 8857 19863 8866 19897
rect 8814 19854 8866 19863
rect 8814 19737 8866 19746
rect 8814 19703 8823 19737
rect 8823 19703 8857 19737
rect 8857 19703 8866 19737
rect 8814 19694 8866 19703
rect 8814 19577 8866 19586
rect 8814 19543 8823 19577
rect 8823 19543 8857 19577
rect 8857 19543 8866 19577
rect 8814 19534 8866 19543
rect 8814 19417 8866 19426
rect 8814 19383 8823 19417
rect 8823 19383 8857 19417
rect 8857 19383 8866 19417
rect 8814 19374 8866 19383
rect 8814 19257 8866 19266
rect 8814 19223 8823 19257
rect 8823 19223 8857 19257
rect 8857 19223 8866 19257
rect 8814 19214 8866 19223
rect 8814 19097 8866 19106
rect 8814 19063 8823 19097
rect 8823 19063 8857 19097
rect 8857 19063 8866 19097
rect 8814 19054 8866 19063
rect 8814 18937 8866 18946
rect 8814 18903 8823 18937
rect 8823 18903 8857 18937
rect 8857 18903 8866 18937
rect 8814 18894 8866 18903
rect 8814 18777 8866 18786
rect 8814 18743 8823 18777
rect 8823 18743 8857 18777
rect 8857 18743 8866 18777
rect 8814 18734 8866 18743
rect 8814 17977 8866 17986
rect 8814 17943 8823 17977
rect 8823 17943 8857 17977
rect 8857 17943 8866 17977
rect 8814 17934 8866 17943
rect 8814 17817 8866 17826
rect 8814 17783 8823 17817
rect 8823 17783 8857 17817
rect 8857 17783 8866 17817
rect 8814 17774 8866 17783
rect 8814 17657 8866 17666
rect 8814 17623 8823 17657
rect 8823 17623 8857 17657
rect 8857 17623 8866 17657
rect 8814 17614 8866 17623
rect 8814 17497 8866 17506
rect 8814 17463 8823 17497
rect 8823 17463 8857 17497
rect 8857 17463 8866 17497
rect 8814 17454 8866 17463
rect 8814 17337 8866 17346
rect 8814 17303 8823 17337
rect 8823 17303 8857 17337
rect 8857 17303 8866 17337
rect 8814 17294 8866 17303
rect 8814 17177 8866 17186
rect 8814 17143 8823 17177
rect 8823 17143 8857 17177
rect 8857 17143 8866 17177
rect 8814 17134 8866 17143
rect 8814 17017 8866 17026
rect 8814 16983 8823 17017
rect 8823 16983 8857 17017
rect 8857 16983 8866 17017
rect 8814 16974 8866 16983
rect 8814 16857 8866 16866
rect 8814 16823 8823 16857
rect 8823 16823 8857 16857
rect 8857 16823 8866 16857
rect 8814 16814 8866 16823
rect 8814 16537 8866 16546
rect 8814 16503 8823 16537
rect 8823 16503 8857 16537
rect 8857 16503 8866 16537
rect 8814 16494 8866 16503
rect 8814 16377 8866 16386
rect 8814 16343 8823 16377
rect 8823 16343 8857 16377
rect 8857 16343 8866 16377
rect 8814 16334 8866 16343
rect 8814 16217 8866 16226
rect 8814 16183 8823 16217
rect 8823 16183 8857 16217
rect 8857 16183 8866 16217
rect 8814 16174 8866 16183
rect 8814 16057 8866 16066
rect 8814 16023 8823 16057
rect 8823 16023 8857 16057
rect 8857 16023 8866 16057
rect 8814 16014 8866 16023
rect 8814 15897 8866 15906
rect 8814 15863 8823 15897
rect 8823 15863 8857 15897
rect 8857 15863 8866 15897
rect 8814 15854 8866 15863
rect 8814 15737 8866 15746
rect 8814 15703 8823 15737
rect 8823 15703 8857 15737
rect 8857 15703 8866 15737
rect 8814 15694 8866 15703
rect 8814 15577 8866 15586
rect 8814 15543 8823 15577
rect 8823 15543 8857 15577
rect 8857 15543 8866 15577
rect 8814 15534 8866 15543
rect 8814 15417 8866 15426
rect 8814 15383 8823 15417
rect 8823 15383 8857 15417
rect 8857 15383 8866 15417
rect 8814 15374 8866 15383
rect 8814 15257 8866 15266
rect 8814 15223 8823 15257
rect 8823 15223 8857 15257
rect 8857 15223 8866 15257
rect 8814 15214 8866 15223
rect 8814 15097 8866 15106
rect 8814 15063 8823 15097
rect 8823 15063 8857 15097
rect 8857 15063 8866 15097
rect 8814 15054 8866 15063
rect 8814 14937 8866 14946
rect 8814 14903 8823 14937
rect 8823 14903 8857 14937
rect 8857 14903 8866 14937
rect 8814 14894 8866 14903
rect 8814 14777 8866 14786
rect 8814 14743 8823 14777
rect 8823 14743 8857 14777
rect 8857 14743 8866 14777
rect 8814 14734 8866 14743
rect 8814 14617 8866 14626
rect 8814 14583 8823 14617
rect 8823 14583 8857 14617
rect 8857 14583 8866 14617
rect 8814 14574 8866 14583
rect 8814 14457 8866 14466
rect 8814 14423 8823 14457
rect 8823 14423 8857 14457
rect 8857 14423 8866 14457
rect 8814 14414 8866 14423
rect 8814 14297 8866 14306
rect 8814 14263 8823 14297
rect 8823 14263 8857 14297
rect 8857 14263 8866 14297
rect 8814 14254 8866 14263
rect 8814 14137 8866 14146
rect 8814 14103 8823 14137
rect 8823 14103 8857 14137
rect 8857 14103 8866 14137
rect 8814 14094 8866 14103
rect 8814 13977 8866 13986
rect 8814 13943 8823 13977
rect 8823 13943 8857 13977
rect 8857 13943 8866 13977
rect 8814 13934 8866 13943
rect 8814 13657 8866 13666
rect 8814 13623 8823 13657
rect 8823 13623 8857 13657
rect 8857 13623 8866 13657
rect 8814 13614 8866 13623
rect 8814 13497 8866 13506
rect 8814 13463 8823 13497
rect 8823 13463 8857 13497
rect 8857 13463 8866 13497
rect 8814 13454 8866 13463
rect 8814 13337 8866 13346
rect 8814 13303 8823 13337
rect 8823 13303 8857 13337
rect 8857 13303 8866 13337
rect 8814 13294 8866 13303
rect 8814 13177 8866 13186
rect 8814 13143 8823 13177
rect 8823 13143 8857 13177
rect 8857 13143 8866 13177
rect 8814 13134 8866 13143
rect 8814 13017 8866 13026
rect 8814 12983 8823 13017
rect 8823 12983 8857 13017
rect 8857 12983 8866 13017
rect 8814 12974 8866 12983
rect 8814 12857 8866 12866
rect 8814 12823 8823 12857
rect 8823 12823 8857 12857
rect 8857 12823 8866 12857
rect 8814 12814 8866 12823
rect 8814 12697 8866 12706
rect 8814 12663 8823 12697
rect 8823 12663 8857 12697
rect 8857 12663 8866 12697
rect 8814 12654 8866 12663
rect 8814 12537 8866 12546
rect 8814 12503 8823 12537
rect 8823 12503 8857 12537
rect 8857 12503 8866 12537
rect 8814 12494 8866 12503
rect 8814 11737 8866 11746
rect 8814 11703 8823 11737
rect 8823 11703 8857 11737
rect 8857 11703 8866 11737
rect 8814 11694 8866 11703
rect 8814 11577 8866 11586
rect 8814 11543 8823 11577
rect 8823 11543 8857 11577
rect 8857 11543 8866 11577
rect 8814 11534 8866 11543
rect 8814 11417 8866 11426
rect 8814 11383 8823 11417
rect 8823 11383 8857 11417
rect 8857 11383 8866 11417
rect 8814 11374 8866 11383
rect 8814 11257 8866 11266
rect 8814 11223 8823 11257
rect 8823 11223 8857 11257
rect 8857 11223 8866 11257
rect 8814 11214 8866 11223
rect 8814 11097 8866 11106
rect 8814 11063 8823 11097
rect 8823 11063 8857 11097
rect 8857 11063 8866 11097
rect 8814 11054 8866 11063
rect 8814 10937 8866 10946
rect 8814 10903 8823 10937
rect 8823 10903 8857 10937
rect 8857 10903 8866 10937
rect 8814 10894 8866 10903
rect 8814 10777 8866 10786
rect 8814 10743 8823 10777
rect 8823 10743 8857 10777
rect 8857 10743 8866 10777
rect 8814 10734 8866 10743
rect 8814 10617 8866 10626
rect 8814 10583 8823 10617
rect 8823 10583 8857 10617
rect 8857 10583 8866 10617
rect 8814 10574 8866 10583
rect 8814 10457 8866 10466
rect 8814 10423 8823 10457
rect 8823 10423 8857 10457
rect 8857 10423 8866 10457
rect 8814 10414 8866 10423
rect 8814 10297 8866 10306
rect 8814 10263 8823 10297
rect 8823 10263 8857 10297
rect 8857 10263 8866 10297
rect 8814 10254 8866 10263
rect 8814 10137 8866 10146
rect 8814 10103 8823 10137
rect 8823 10103 8857 10137
rect 8857 10103 8866 10137
rect 8814 10094 8866 10103
rect 8814 9977 8866 9986
rect 8814 9943 8823 9977
rect 8823 9943 8857 9977
rect 8857 9943 8866 9977
rect 8814 9934 8866 9943
rect 8814 9817 8866 9826
rect 8814 9783 8823 9817
rect 8823 9783 8857 9817
rect 8857 9783 8866 9817
rect 8814 9774 8866 9783
rect 8814 9497 8866 9506
rect 8814 9463 8823 9497
rect 8823 9463 8857 9497
rect 8857 9463 8866 9497
rect 8814 9454 8866 9463
rect 8814 9337 8866 9346
rect 8814 9303 8823 9337
rect 8823 9303 8857 9337
rect 8857 9303 8866 9337
rect 8814 9294 8866 9303
rect 8814 9017 8866 9026
rect 8814 8983 8823 9017
rect 8823 8983 8857 9017
rect 8857 8983 8866 9017
rect 8814 8974 8866 8983
rect 8814 8857 8866 8866
rect 8814 8823 8823 8857
rect 8823 8823 8857 8857
rect 8857 8823 8866 8857
rect 8814 8814 8866 8823
rect 8814 8697 8866 8706
rect 8814 8663 8823 8697
rect 8823 8663 8857 8697
rect 8857 8663 8866 8697
rect 8814 8654 8866 8663
rect 8814 8537 8866 8546
rect 8814 8503 8823 8537
rect 8823 8503 8857 8537
rect 8857 8503 8866 8537
rect 8814 8494 8866 8503
rect 8814 8377 8866 8386
rect 8814 8343 8823 8377
rect 8823 8343 8857 8377
rect 8857 8343 8866 8377
rect 8814 8334 8866 8343
rect 8814 8217 8866 8226
rect 8814 8183 8823 8217
rect 8823 8183 8857 8217
rect 8857 8183 8866 8217
rect 8814 8174 8866 8183
rect 8814 8057 8866 8066
rect 8814 8023 8823 8057
rect 8823 8023 8857 8057
rect 8857 8023 8866 8057
rect 8814 8014 8866 8023
rect 8814 7897 8866 7906
rect 8814 7863 8823 7897
rect 8823 7863 8857 7897
rect 8857 7863 8866 7897
rect 8814 7854 8866 7863
rect 8814 7737 8866 7746
rect 8814 7703 8823 7737
rect 8823 7703 8857 7737
rect 8857 7703 8866 7737
rect 8814 7694 8866 7703
rect 8814 7417 8866 7426
rect 8814 7383 8823 7417
rect 8823 7383 8857 7417
rect 8857 7383 8866 7417
rect 8814 7374 8866 7383
rect 8814 7257 8866 7266
rect 8814 7223 8823 7257
rect 8823 7223 8857 7257
rect 8857 7223 8866 7257
rect 8814 7214 8866 7223
rect 8814 6937 8866 6946
rect 8814 6903 8823 6937
rect 8823 6903 8857 6937
rect 8857 6903 8866 6937
rect 8814 6894 8866 6903
rect 8814 6777 8866 6786
rect 8814 6743 8823 6777
rect 8823 6743 8857 6777
rect 8857 6743 8866 6777
rect 8814 6734 8866 6743
rect 8814 6457 8866 6466
rect 8814 6423 8823 6457
rect 8823 6423 8857 6457
rect 8857 6423 8866 6457
rect 8814 6414 8866 6423
rect 8814 6297 8866 6306
rect 8814 6263 8823 6297
rect 8823 6263 8857 6297
rect 8857 6263 8866 6297
rect 8814 6254 8866 6263
rect 8814 6137 8866 6146
rect 8814 6103 8823 6137
rect 8823 6103 8857 6137
rect 8857 6103 8866 6137
rect 8814 6094 8866 6103
rect 8814 5977 8866 5986
rect 8814 5943 8823 5977
rect 8823 5943 8857 5977
rect 8857 5943 8866 5977
rect 8814 5934 8866 5943
rect 8814 5817 8866 5826
rect 8814 5783 8823 5817
rect 8823 5783 8857 5817
rect 8857 5783 8866 5817
rect 8814 5774 8866 5783
rect 8814 5657 8866 5666
rect 8814 5623 8823 5657
rect 8823 5623 8857 5657
rect 8857 5623 8866 5657
rect 8814 5614 8866 5623
rect 8814 5497 8866 5506
rect 8814 5463 8823 5497
rect 8823 5463 8857 5497
rect 8857 5463 8866 5497
rect 8814 5454 8866 5463
rect 8814 5337 8866 5346
rect 8814 5303 8823 5337
rect 8823 5303 8857 5337
rect 8857 5303 8866 5337
rect 8814 5294 8866 5303
rect 8814 5177 8866 5186
rect 8814 5143 8823 5177
rect 8823 5143 8857 5177
rect 8857 5143 8866 5177
rect 8814 5134 8866 5143
rect 8814 5017 8866 5026
rect 8814 4983 8823 5017
rect 8823 4983 8857 5017
rect 8857 4983 8866 5017
rect 8814 4974 8866 4983
rect 8814 4857 8866 4866
rect 8814 4823 8823 4857
rect 8823 4823 8857 4857
rect 8857 4823 8866 4857
rect 8814 4814 8866 4823
rect 8814 4697 8866 4706
rect 8814 4663 8823 4697
rect 8823 4663 8857 4697
rect 8857 4663 8866 4697
rect 8814 4654 8866 4663
rect 8814 4537 8866 4546
rect 8814 4503 8823 4537
rect 8823 4503 8857 4537
rect 8857 4503 8866 4537
rect 8814 4494 8866 4503
rect 8814 4377 8866 4386
rect 8814 4343 8823 4377
rect 8823 4343 8857 4377
rect 8857 4343 8866 4377
rect 8814 4334 8866 4343
rect 8814 4217 8866 4226
rect 8814 4183 8823 4217
rect 8823 4183 8857 4217
rect 8857 4183 8866 4217
rect 8814 4174 8866 4183
rect 8814 4057 8866 4066
rect 8814 4023 8823 4057
rect 8823 4023 8857 4057
rect 8857 4023 8866 4057
rect 8814 4014 8866 4023
rect 8814 3897 8866 3906
rect 8814 3863 8823 3897
rect 8823 3863 8857 3897
rect 8857 3863 8866 3897
rect 8814 3854 8866 3863
rect 8814 3417 8866 3426
rect 8814 3383 8823 3417
rect 8823 3383 8857 3417
rect 8857 3383 8866 3417
rect 8814 3374 8866 3383
rect 8814 3257 8866 3266
rect 8814 3223 8823 3257
rect 8823 3223 8857 3257
rect 8857 3223 8866 3257
rect 8814 3214 8866 3223
rect 8814 3097 8866 3106
rect 8814 3063 8823 3097
rect 8823 3063 8857 3097
rect 8857 3063 8866 3097
rect 8814 3054 8866 3063
rect 8814 2937 8866 2946
rect 8814 2903 8823 2937
rect 8823 2903 8857 2937
rect 8857 2903 8866 2937
rect 8814 2894 8866 2903
rect 8814 2777 8866 2786
rect 8814 2743 8823 2777
rect 8823 2743 8857 2777
rect 8857 2743 8866 2777
rect 8814 2734 8866 2743
rect 8814 2617 8866 2626
rect 8814 2583 8823 2617
rect 8823 2583 8857 2617
rect 8857 2583 8866 2617
rect 8814 2574 8866 2583
rect 8814 2457 8866 2466
rect 8814 2423 8823 2457
rect 8823 2423 8857 2457
rect 8857 2423 8866 2457
rect 8814 2414 8866 2423
rect 8814 2297 8866 2306
rect 8814 2263 8823 2297
rect 8823 2263 8857 2297
rect 8857 2263 8866 2297
rect 8814 2254 8866 2263
rect 8814 2137 8866 2146
rect 8814 2103 8823 2137
rect 8823 2103 8857 2137
rect 8857 2103 8866 2137
rect 8814 2094 8866 2103
rect 8814 1977 8866 1986
rect 8814 1943 8823 1977
rect 8823 1943 8857 1977
rect 8857 1943 8866 1977
rect 8814 1934 8866 1943
rect 8814 1657 8866 1666
rect 8814 1623 8823 1657
rect 8823 1623 8857 1657
rect 8857 1623 8866 1657
rect 8814 1614 8866 1623
rect 8814 1497 8866 1506
rect 8814 1463 8823 1497
rect 8823 1463 8857 1497
rect 8857 1463 8866 1497
rect 8814 1454 8866 1463
rect 8814 1337 8866 1346
rect 8814 1303 8823 1337
rect 8823 1303 8857 1337
rect 8857 1303 8866 1337
rect 8814 1294 8866 1303
rect 8814 1177 8866 1186
rect 8814 1143 8823 1177
rect 8823 1143 8857 1177
rect 8857 1143 8866 1177
rect 8814 1134 8866 1143
rect 8814 1017 8866 1026
rect 8814 983 8823 1017
rect 8823 983 8857 1017
rect 8857 983 8866 1017
rect 8814 974 8866 983
rect 8814 537 8866 546
rect 8814 503 8823 537
rect 8823 503 8857 537
rect 8857 503 8866 537
rect 8814 494 8866 503
rect 8814 377 8866 386
rect 8814 343 8823 377
rect 8823 343 8857 377
rect 8857 343 8866 377
rect 8814 334 8866 343
rect 8814 217 8866 226
rect 8814 183 8823 217
rect 8823 183 8857 217
rect 8857 183 8866 217
rect 8814 174 8866 183
rect 8814 57 8866 66
rect 8814 23 8823 57
rect 8823 23 8857 57
rect 8857 23 8866 57
rect 8814 14 8866 23
rect 8974 31417 9026 31426
rect 8974 31383 8983 31417
rect 8983 31383 9017 31417
rect 9017 31383 9026 31417
rect 8974 31374 9026 31383
rect 8974 31257 9026 31266
rect 8974 31223 8983 31257
rect 8983 31223 9017 31257
rect 9017 31223 9026 31257
rect 8974 31214 9026 31223
rect 8974 31097 9026 31106
rect 8974 31063 8983 31097
rect 8983 31063 9017 31097
rect 9017 31063 9026 31097
rect 8974 31054 9026 31063
rect 8974 30937 9026 30946
rect 8974 30903 8983 30937
rect 8983 30903 9017 30937
rect 9017 30903 9026 30937
rect 8974 30894 9026 30903
rect 8974 30777 9026 30786
rect 8974 30743 8983 30777
rect 8983 30743 9017 30777
rect 9017 30743 9026 30777
rect 8974 30734 9026 30743
rect 8974 30617 9026 30626
rect 8974 30583 8983 30617
rect 8983 30583 9017 30617
rect 9017 30583 9026 30617
rect 8974 30574 9026 30583
rect 8974 30457 9026 30466
rect 8974 30423 8983 30457
rect 8983 30423 9017 30457
rect 9017 30423 9026 30457
rect 8974 30414 9026 30423
rect 8974 30297 9026 30306
rect 8974 30263 8983 30297
rect 8983 30263 9017 30297
rect 9017 30263 9026 30297
rect 8974 30254 9026 30263
rect 8974 29977 9026 29986
rect 8974 29943 8983 29977
rect 8983 29943 9017 29977
rect 9017 29943 9026 29977
rect 8974 29934 9026 29943
rect 8974 29817 9026 29826
rect 8974 29783 8983 29817
rect 8983 29783 9017 29817
rect 9017 29783 9026 29817
rect 8974 29774 9026 29783
rect 8974 29657 9026 29666
rect 8974 29623 8983 29657
rect 8983 29623 9017 29657
rect 9017 29623 9026 29657
rect 8974 29614 9026 29623
rect 8974 29497 9026 29506
rect 8974 29463 8983 29497
rect 8983 29463 9017 29497
rect 9017 29463 9026 29497
rect 8974 29454 9026 29463
rect 8974 29337 9026 29346
rect 8974 29303 8983 29337
rect 8983 29303 9017 29337
rect 9017 29303 9026 29337
rect 8974 29294 9026 29303
rect 8974 29177 9026 29186
rect 8974 29143 8983 29177
rect 8983 29143 9017 29177
rect 9017 29143 9026 29177
rect 8974 29134 9026 29143
rect 8974 29017 9026 29026
rect 8974 28983 8983 29017
rect 8983 28983 9017 29017
rect 9017 28983 9026 29017
rect 8974 28974 9026 28983
rect 8974 28857 9026 28866
rect 8974 28823 8983 28857
rect 8983 28823 9017 28857
rect 9017 28823 9026 28857
rect 8974 28814 9026 28823
rect 8974 28057 9026 28066
rect 8974 28023 8983 28057
rect 8983 28023 9017 28057
rect 9017 28023 9026 28057
rect 8974 28014 9026 28023
rect 8974 27897 9026 27906
rect 8974 27863 8983 27897
rect 8983 27863 9017 27897
rect 9017 27863 9026 27897
rect 8974 27854 9026 27863
rect 8974 27737 9026 27746
rect 8974 27703 8983 27737
rect 8983 27703 9017 27737
rect 9017 27703 9026 27737
rect 8974 27694 9026 27703
rect 8974 27577 9026 27586
rect 8974 27543 8983 27577
rect 8983 27543 9017 27577
rect 9017 27543 9026 27577
rect 8974 27534 9026 27543
rect 8974 27417 9026 27426
rect 8974 27383 8983 27417
rect 8983 27383 9017 27417
rect 9017 27383 9026 27417
rect 8974 27374 9026 27383
rect 8974 27257 9026 27266
rect 8974 27223 8983 27257
rect 8983 27223 9017 27257
rect 9017 27223 9026 27257
rect 8974 27214 9026 27223
rect 8974 27097 9026 27106
rect 8974 27063 8983 27097
rect 8983 27063 9017 27097
rect 9017 27063 9026 27097
rect 8974 27054 9026 27063
rect 8974 26937 9026 26946
rect 8974 26903 8983 26937
rect 8983 26903 9017 26937
rect 9017 26903 9026 26937
rect 8974 26894 9026 26903
rect 8974 26137 9026 26146
rect 8974 26103 8983 26137
rect 8983 26103 9017 26137
rect 9017 26103 9026 26137
rect 8974 26094 9026 26103
rect 8974 25977 9026 25986
rect 8974 25943 8983 25977
rect 8983 25943 9017 25977
rect 9017 25943 9026 25977
rect 8974 25934 9026 25943
rect 8974 25817 9026 25826
rect 8974 25783 8983 25817
rect 8983 25783 9017 25817
rect 9017 25783 9026 25817
rect 8974 25774 9026 25783
rect 8974 25657 9026 25666
rect 8974 25623 8983 25657
rect 8983 25623 9017 25657
rect 9017 25623 9026 25657
rect 8974 25614 9026 25623
rect 8974 25497 9026 25506
rect 8974 25463 8983 25497
rect 8983 25463 9017 25497
rect 9017 25463 9026 25497
rect 8974 25454 9026 25463
rect 8974 25337 9026 25346
rect 8974 25303 8983 25337
rect 8983 25303 9017 25337
rect 9017 25303 9026 25337
rect 8974 25294 9026 25303
rect 8974 25177 9026 25186
rect 8974 25143 8983 25177
rect 8983 25143 9017 25177
rect 9017 25143 9026 25177
rect 8974 25134 9026 25143
rect 8974 25017 9026 25026
rect 8974 24983 8983 25017
rect 8983 24983 9017 25017
rect 9017 24983 9026 25017
rect 8974 24974 9026 24983
rect 8974 24697 9026 24706
rect 8974 24663 8983 24697
rect 8983 24663 9017 24697
rect 9017 24663 9026 24697
rect 8974 24654 9026 24663
rect 8974 24537 9026 24546
rect 8974 24503 8983 24537
rect 8983 24503 9017 24537
rect 9017 24503 9026 24537
rect 8974 24494 9026 24503
rect 8974 24377 9026 24386
rect 8974 24343 8983 24377
rect 8983 24343 9017 24377
rect 9017 24343 9026 24377
rect 8974 24334 9026 24343
rect 8974 24217 9026 24226
rect 8974 24183 8983 24217
rect 8983 24183 9017 24217
rect 9017 24183 9026 24217
rect 8974 24174 9026 24183
rect 8974 24057 9026 24066
rect 8974 24023 8983 24057
rect 8983 24023 9017 24057
rect 9017 24023 9026 24057
rect 8974 24014 9026 24023
rect 8974 23897 9026 23906
rect 8974 23863 8983 23897
rect 8983 23863 9017 23897
rect 9017 23863 9026 23897
rect 8974 23854 9026 23863
rect 8974 23737 9026 23746
rect 8974 23703 8983 23737
rect 8983 23703 9017 23737
rect 9017 23703 9026 23737
rect 8974 23694 9026 23703
rect 8974 23577 9026 23586
rect 8974 23543 8983 23577
rect 8983 23543 9017 23577
rect 9017 23543 9026 23577
rect 8974 23534 9026 23543
rect 8974 23417 9026 23426
rect 8974 23383 8983 23417
rect 8983 23383 9017 23417
rect 9017 23383 9026 23417
rect 8974 23374 9026 23383
rect 8974 23257 9026 23266
rect 8974 23223 8983 23257
rect 8983 23223 9017 23257
rect 9017 23223 9026 23257
rect 8974 23214 9026 23223
rect 8974 23097 9026 23106
rect 8974 23063 8983 23097
rect 8983 23063 9017 23097
rect 9017 23063 9026 23097
rect 8974 23054 9026 23063
rect 8974 22937 9026 22946
rect 8974 22903 8983 22937
rect 8983 22903 9017 22937
rect 9017 22903 9026 22937
rect 8974 22894 9026 22903
rect 8974 22777 9026 22786
rect 8974 22743 8983 22777
rect 8983 22743 9017 22777
rect 9017 22743 9026 22777
rect 8974 22734 9026 22743
rect 8974 22617 9026 22626
rect 8974 22583 8983 22617
rect 8983 22583 9017 22617
rect 9017 22583 9026 22617
rect 8974 22574 9026 22583
rect 8974 22457 9026 22466
rect 8974 22423 8983 22457
rect 8983 22423 9017 22457
rect 9017 22423 9026 22457
rect 8974 22414 9026 22423
rect 8974 22297 9026 22306
rect 8974 22263 8983 22297
rect 8983 22263 9017 22297
rect 9017 22263 9026 22297
rect 8974 22254 9026 22263
rect 8974 22137 9026 22146
rect 8974 22103 8983 22137
rect 8983 22103 9017 22137
rect 9017 22103 9026 22137
rect 8974 22094 9026 22103
rect 8974 21817 9026 21826
rect 8974 21783 8983 21817
rect 8983 21783 9017 21817
rect 9017 21783 9026 21817
rect 8974 21774 9026 21783
rect 8974 21657 9026 21666
rect 8974 21623 8983 21657
rect 8983 21623 9017 21657
rect 9017 21623 9026 21657
rect 8974 21614 9026 21623
rect 8974 21497 9026 21506
rect 8974 21463 8983 21497
rect 8983 21463 9017 21497
rect 9017 21463 9026 21497
rect 8974 21454 9026 21463
rect 8974 21337 9026 21346
rect 8974 21303 8983 21337
rect 8983 21303 9017 21337
rect 9017 21303 9026 21337
rect 8974 21294 9026 21303
rect 8974 21177 9026 21186
rect 8974 21143 8983 21177
rect 8983 21143 9017 21177
rect 9017 21143 9026 21177
rect 8974 21134 9026 21143
rect 8974 21017 9026 21026
rect 8974 20983 8983 21017
rect 8983 20983 9017 21017
rect 9017 20983 9026 21017
rect 8974 20974 9026 20983
rect 8974 20857 9026 20866
rect 8974 20823 8983 20857
rect 8983 20823 9017 20857
rect 9017 20823 9026 20857
rect 8974 20814 9026 20823
rect 8974 20697 9026 20706
rect 8974 20663 8983 20697
rect 8983 20663 9017 20697
rect 9017 20663 9026 20697
rect 8974 20654 9026 20663
rect 8974 19897 9026 19906
rect 8974 19863 8983 19897
rect 8983 19863 9017 19897
rect 9017 19863 9026 19897
rect 8974 19854 9026 19863
rect 8974 19737 9026 19746
rect 8974 19703 8983 19737
rect 8983 19703 9017 19737
rect 9017 19703 9026 19737
rect 8974 19694 9026 19703
rect 8974 19577 9026 19586
rect 8974 19543 8983 19577
rect 8983 19543 9017 19577
rect 9017 19543 9026 19577
rect 8974 19534 9026 19543
rect 8974 19417 9026 19426
rect 8974 19383 8983 19417
rect 8983 19383 9017 19417
rect 9017 19383 9026 19417
rect 8974 19374 9026 19383
rect 8974 19257 9026 19266
rect 8974 19223 8983 19257
rect 8983 19223 9017 19257
rect 9017 19223 9026 19257
rect 8974 19214 9026 19223
rect 8974 19097 9026 19106
rect 8974 19063 8983 19097
rect 8983 19063 9017 19097
rect 9017 19063 9026 19097
rect 8974 19054 9026 19063
rect 8974 18937 9026 18946
rect 8974 18903 8983 18937
rect 8983 18903 9017 18937
rect 9017 18903 9026 18937
rect 8974 18894 9026 18903
rect 8974 18777 9026 18786
rect 8974 18743 8983 18777
rect 8983 18743 9017 18777
rect 9017 18743 9026 18777
rect 8974 18734 9026 18743
rect 8974 17977 9026 17986
rect 8974 17943 8983 17977
rect 8983 17943 9017 17977
rect 9017 17943 9026 17977
rect 8974 17934 9026 17943
rect 8974 17817 9026 17826
rect 8974 17783 8983 17817
rect 8983 17783 9017 17817
rect 9017 17783 9026 17817
rect 8974 17774 9026 17783
rect 8974 17657 9026 17666
rect 8974 17623 8983 17657
rect 8983 17623 9017 17657
rect 9017 17623 9026 17657
rect 8974 17614 9026 17623
rect 8974 17497 9026 17506
rect 8974 17463 8983 17497
rect 8983 17463 9017 17497
rect 9017 17463 9026 17497
rect 8974 17454 9026 17463
rect 8974 17337 9026 17346
rect 8974 17303 8983 17337
rect 8983 17303 9017 17337
rect 9017 17303 9026 17337
rect 8974 17294 9026 17303
rect 8974 17177 9026 17186
rect 8974 17143 8983 17177
rect 8983 17143 9017 17177
rect 9017 17143 9026 17177
rect 8974 17134 9026 17143
rect 8974 17017 9026 17026
rect 8974 16983 8983 17017
rect 8983 16983 9017 17017
rect 9017 16983 9026 17017
rect 8974 16974 9026 16983
rect 8974 16857 9026 16866
rect 8974 16823 8983 16857
rect 8983 16823 9017 16857
rect 9017 16823 9026 16857
rect 8974 16814 9026 16823
rect 8974 16537 9026 16546
rect 8974 16503 8983 16537
rect 8983 16503 9017 16537
rect 9017 16503 9026 16537
rect 8974 16494 9026 16503
rect 8974 16377 9026 16386
rect 8974 16343 8983 16377
rect 8983 16343 9017 16377
rect 9017 16343 9026 16377
rect 8974 16334 9026 16343
rect 8974 16217 9026 16226
rect 8974 16183 8983 16217
rect 8983 16183 9017 16217
rect 9017 16183 9026 16217
rect 8974 16174 9026 16183
rect 8974 16057 9026 16066
rect 8974 16023 8983 16057
rect 8983 16023 9017 16057
rect 9017 16023 9026 16057
rect 8974 16014 9026 16023
rect 8974 15897 9026 15906
rect 8974 15863 8983 15897
rect 8983 15863 9017 15897
rect 9017 15863 9026 15897
rect 8974 15854 9026 15863
rect 8974 15737 9026 15746
rect 8974 15703 8983 15737
rect 8983 15703 9017 15737
rect 9017 15703 9026 15737
rect 8974 15694 9026 15703
rect 8974 15577 9026 15586
rect 8974 15543 8983 15577
rect 8983 15543 9017 15577
rect 9017 15543 9026 15577
rect 8974 15534 9026 15543
rect 8974 15417 9026 15426
rect 8974 15383 8983 15417
rect 8983 15383 9017 15417
rect 9017 15383 9026 15417
rect 8974 15374 9026 15383
rect 8974 15257 9026 15266
rect 8974 15223 8983 15257
rect 8983 15223 9017 15257
rect 9017 15223 9026 15257
rect 8974 15214 9026 15223
rect 8974 15097 9026 15106
rect 8974 15063 8983 15097
rect 8983 15063 9017 15097
rect 9017 15063 9026 15097
rect 8974 15054 9026 15063
rect 8974 14937 9026 14946
rect 8974 14903 8983 14937
rect 8983 14903 9017 14937
rect 9017 14903 9026 14937
rect 8974 14894 9026 14903
rect 8974 14777 9026 14786
rect 8974 14743 8983 14777
rect 8983 14743 9017 14777
rect 9017 14743 9026 14777
rect 8974 14734 9026 14743
rect 8974 14617 9026 14626
rect 8974 14583 8983 14617
rect 8983 14583 9017 14617
rect 9017 14583 9026 14617
rect 8974 14574 9026 14583
rect 8974 14457 9026 14466
rect 8974 14423 8983 14457
rect 8983 14423 9017 14457
rect 9017 14423 9026 14457
rect 8974 14414 9026 14423
rect 8974 14297 9026 14306
rect 8974 14263 8983 14297
rect 8983 14263 9017 14297
rect 9017 14263 9026 14297
rect 8974 14254 9026 14263
rect 8974 14137 9026 14146
rect 8974 14103 8983 14137
rect 8983 14103 9017 14137
rect 9017 14103 9026 14137
rect 8974 14094 9026 14103
rect 8974 13977 9026 13986
rect 8974 13943 8983 13977
rect 8983 13943 9017 13977
rect 9017 13943 9026 13977
rect 8974 13934 9026 13943
rect 8974 13657 9026 13666
rect 8974 13623 8983 13657
rect 8983 13623 9017 13657
rect 9017 13623 9026 13657
rect 8974 13614 9026 13623
rect 8974 13497 9026 13506
rect 8974 13463 8983 13497
rect 8983 13463 9017 13497
rect 9017 13463 9026 13497
rect 8974 13454 9026 13463
rect 8974 13337 9026 13346
rect 8974 13303 8983 13337
rect 8983 13303 9017 13337
rect 9017 13303 9026 13337
rect 8974 13294 9026 13303
rect 8974 13177 9026 13186
rect 8974 13143 8983 13177
rect 8983 13143 9017 13177
rect 9017 13143 9026 13177
rect 8974 13134 9026 13143
rect 8974 13017 9026 13026
rect 8974 12983 8983 13017
rect 8983 12983 9017 13017
rect 9017 12983 9026 13017
rect 8974 12974 9026 12983
rect 8974 12857 9026 12866
rect 8974 12823 8983 12857
rect 8983 12823 9017 12857
rect 9017 12823 9026 12857
rect 8974 12814 9026 12823
rect 8974 12697 9026 12706
rect 8974 12663 8983 12697
rect 8983 12663 9017 12697
rect 9017 12663 9026 12697
rect 8974 12654 9026 12663
rect 8974 12537 9026 12546
rect 8974 12503 8983 12537
rect 8983 12503 9017 12537
rect 9017 12503 9026 12537
rect 8974 12494 9026 12503
rect 8974 11737 9026 11746
rect 8974 11703 8983 11737
rect 8983 11703 9017 11737
rect 9017 11703 9026 11737
rect 8974 11694 9026 11703
rect 8974 11577 9026 11586
rect 8974 11543 8983 11577
rect 8983 11543 9017 11577
rect 9017 11543 9026 11577
rect 8974 11534 9026 11543
rect 8974 11417 9026 11426
rect 8974 11383 8983 11417
rect 8983 11383 9017 11417
rect 9017 11383 9026 11417
rect 8974 11374 9026 11383
rect 8974 11257 9026 11266
rect 8974 11223 8983 11257
rect 8983 11223 9017 11257
rect 9017 11223 9026 11257
rect 8974 11214 9026 11223
rect 8974 11097 9026 11106
rect 8974 11063 8983 11097
rect 8983 11063 9017 11097
rect 9017 11063 9026 11097
rect 8974 11054 9026 11063
rect 8974 10937 9026 10946
rect 8974 10903 8983 10937
rect 8983 10903 9017 10937
rect 9017 10903 9026 10937
rect 8974 10894 9026 10903
rect 8974 10777 9026 10786
rect 8974 10743 8983 10777
rect 8983 10743 9017 10777
rect 9017 10743 9026 10777
rect 8974 10734 9026 10743
rect 8974 10617 9026 10626
rect 8974 10583 8983 10617
rect 8983 10583 9017 10617
rect 9017 10583 9026 10617
rect 8974 10574 9026 10583
rect 8974 10457 9026 10466
rect 8974 10423 8983 10457
rect 8983 10423 9017 10457
rect 9017 10423 9026 10457
rect 8974 10414 9026 10423
rect 8974 10297 9026 10306
rect 8974 10263 8983 10297
rect 8983 10263 9017 10297
rect 9017 10263 9026 10297
rect 8974 10254 9026 10263
rect 8974 10137 9026 10146
rect 8974 10103 8983 10137
rect 8983 10103 9017 10137
rect 9017 10103 9026 10137
rect 8974 10094 9026 10103
rect 8974 9977 9026 9986
rect 8974 9943 8983 9977
rect 8983 9943 9017 9977
rect 9017 9943 9026 9977
rect 8974 9934 9026 9943
rect 8974 9817 9026 9826
rect 8974 9783 8983 9817
rect 8983 9783 9017 9817
rect 9017 9783 9026 9817
rect 8974 9774 9026 9783
rect 8974 9497 9026 9506
rect 8974 9463 8983 9497
rect 8983 9463 9017 9497
rect 9017 9463 9026 9497
rect 8974 9454 9026 9463
rect 8974 9337 9026 9346
rect 8974 9303 8983 9337
rect 8983 9303 9017 9337
rect 9017 9303 9026 9337
rect 8974 9294 9026 9303
rect 8974 9017 9026 9026
rect 8974 8983 8983 9017
rect 8983 8983 9017 9017
rect 9017 8983 9026 9017
rect 8974 8974 9026 8983
rect 8974 8857 9026 8866
rect 8974 8823 8983 8857
rect 8983 8823 9017 8857
rect 9017 8823 9026 8857
rect 8974 8814 9026 8823
rect 8974 8697 9026 8706
rect 8974 8663 8983 8697
rect 8983 8663 9017 8697
rect 9017 8663 9026 8697
rect 8974 8654 9026 8663
rect 8974 8537 9026 8546
rect 8974 8503 8983 8537
rect 8983 8503 9017 8537
rect 9017 8503 9026 8537
rect 8974 8494 9026 8503
rect 8974 8377 9026 8386
rect 8974 8343 8983 8377
rect 8983 8343 9017 8377
rect 9017 8343 9026 8377
rect 8974 8334 9026 8343
rect 8974 8217 9026 8226
rect 8974 8183 8983 8217
rect 8983 8183 9017 8217
rect 9017 8183 9026 8217
rect 8974 8174 9026 8183
rect 8974 8057 9026 8066
rect 8974 8023 8983 8057
rect 8983 8023 9017 8057
rect 9017 8023 9026 8057
rect 8974 8014 9026 8023
rect 8974 7897 9026 7906
rect 8974 7863 8983 7897
rect 8983 7863 9017 7897
rect 9017 7863 9026 7897
rect 8974 7854 9026 7863
rect 8974 7737 9026 7746
rect 8974 7703 8983 7737
rect 8983 7703 9017 7737
rect 9017 7703 9026 7737
rect 8974 7694 9026 7703
rect 8974 7417 9026 7426
rect 8974 7383 8983 7417
rect 8983 7383 9017 7417
rect 9017 7383 9026 7417
rect 8974 7374 9026 7383
rect 8974 7257 9026 7266
rect 8974 7223 8983 7257
rect 8983 7223 9017 7257
rect 9017 7223 9026 7257
rect 8974 7214 9026 7223
rect 8974 6937 9026 6946
rect 8974 6903 8983 6937
rect 8983 6903 9017 6937
rect 9017 6903 9026 6937
rect 8974 6894 9026 6903
rect 8974 6777 9026 6786
rect 8974 6743 8983 6777
rect 8983 6743 9017 6777
rect 9017 6743 9026 6777
rect 8974 6734 9026 6743
rect 8974 6457 9026 6466
rect 8974 6423 8983 6457
rect 8983 6423 9017 6457
rect 9017 6423 9026 6457
rect 8974 6414 9026 6423
rect 8974 6297 9026 6306
rect 8974 6263 8983 6297
rect 8983 6263 9017 6297
rect 9017 6263 9026 6297
rect 8974 6254 9026 6263
rect 8974 6137 9026 6146
rect 8974 6103 8983 6137
rect 8983 6103 9017 6137
rect 9017 6103 9026 6137
rect 8974 6094 9026 6103
rect 8974 5977 9026 5986
rect 8974 5943 8983 5977
rect 8983 5943 9017 5977
rect 9017 5943 9026 5977
rect 8974 5934 9026 5943
rect 8974 5817 9026 5826
rect 8974 5783 8983 5817
rect 8983 5783 9017 5817
rect 9017 5783 9026 5817
rect 8974 5774 9026 5783
rect 8974 5657 9026 5666
rect 8974 5623 8983 5657
rect 8983 5623 9017 5657
rect 9017 5623 9026 5657
rect 8974 5614 9026 5623
rect 8974 5497 9026 5506
rect 8974 5463 8983 5497
rect 8983 5463 9017 5497
rect 9017 5463 9026 5497
rect 8974 5454 9026 5463
rect 8974 5337 9026 5346
rect 8974 5303 8983 5337
rect 8983 5303 9017 5337
rect 9017 5303 9026 5337
rect 8974 5294 9026 5303
rect 8974 5177 9026 5186
rect 8974 5143 8983 5177
rect 8983 5143 9017 5177
rect 9017 5143 9026 5177
rect 8974 5134 9026 5143
rect 8974 5017 9026 5026
rect 8974 4983 8983 5017
rect 8983 4983 9017 5017
rect 9017 4983 9026 5017
rect 8974 4974 9026 4983
rect 8974 4857 9026 4866
rect 8974 4823 8983 4857
rect 8983 4823 9017 4857
rect 9017 4823 9026 4857
rect 8974 4814 9026 4823
rect 8974 4697 9026 4706
rect 8974 4663 8983 4697
rect 8983 4663 9017 4697
rect 9017 4663 9026 4697
rect 8974 4654 9026 4663
rect 8974 4537 9026 4546
rect 8974 4503 8983 4537
rect 8983 4503 9017 4537
rect 9017 4503 9026 4537
rect 8974 4494 9026 4503
rect 8974 4377 9026 4386
rect 8974 4343 8983 4377
rect 8983 4343 9017 4377
rect 9017 4343 9026 4377
rect 8974 4334 9026 4343
rect 8974 4217 9026 4226
rect 8974 4183 8983 4217
rect 8983 4183 9017 4217
rect 9017 4183 9026 4217
rect 8974 4174 9026 4183
rect 8974 4057 9026 4066
rect 8974 4023 8983 4057
rect 8983 4023 9017 4057
rect 9017 4023 9026 4057
rect 8974 4014 9026 4023
rect 8974 3897 9026 3906
rect 8974 3863 8983 3897
rect 8983 3863 9017 3897
rect 9017 3863 9026 3897
rect 8974 3854 9026 3863
rect 8974 3417 9026 3426
rect 8974 3383 8983 3417
rect 8983 3383 9017 3417
rect 9017 3383 9026 3417
rect 8974 3374 9026 3383
rect 8974 3257 9026 3266
rect 8974 3223 8983 3257
rect 8983 3223 9017 3257
rect 9017 3223 9026 3257
rect 8974 3214 9026 3223
rect 8974 3097 9026 3106
rect 8974 3063 8983 3097
rect 8983 3063 9017 3097
rect 9017 3063 9026 3097
rect 8974 3054 9026 3063
rect 8974 2937 9026 2946
rect 8974 2903 8983 2937
rect 8983 2903 9017 2937
rect 9017 2903 9026 2937
rect 8974 2894 9026 2903
rect 8974 2777 9026 2786
rect 8974 2743 8983 2777
rect 8983 2743 9017 2777
rect 9017 2743 9026 2777
rect 8974 2734 9026 2743
rect 8974 2617 9026 2626
rect 8974 2583 8983 2617
rect 8983 2583 9017 2617
rect 9017 2583 9026 2617
rect 8974 2574 9026 2583
rect 8974 2457 9026 2466
rect 8974 2423 8983 2457
rect 8983 2423 9017 2457
rect 9017 2423 9026 2457
rect 8974 2414 9026 2423
rect 8974 2297 9026 2306
rect 8974 2263 8983 2297
rect 8983 2263 9017 2297
rect 9017 2263 9026 2297
rect 8974 2254 9026 2263
rect 8974 2137 9026 2146
rect 8974 2103 8983 2137
rect 8983 2103 9017 2137
rect 9017 2103 9026 2137
rect 8974 2094 9026 2103
rect 8974 1977 9026 1986
rect 8974 1943 8983 1977
rect 8983 1943 9017 1977
rect 9017 1943 9026 1977
rect 8974 1934 9026 1943
rect 8974 1657 9026 1666
rect 8974 1623 8983 1657
rect 8983 1623 9017 1657
rect 9017 1623 9026 1657
rect 8974 1614 9026 1623
rect 8974 1497 9026 1506
rect 8974 1463 8983 1497
rect 8983 1463 9017 1497
rect 9017 1463 9026 1497
rect 8974 1454 9026 1463
rect 8974 1337 9026 1346
rect 8974 1303 8983 1337
rect 8983 1303 9017 1337
rect 9017 1303 9026 1337
rect 8974 1294 9026 1303
rect 8974 1177 9026 1186
rect 8974 1143 8983 1177
rect 8983 1143 9017 1177
rect 9017 1143 9026 1177
rect 8974 1134 9026 1143
rect 8974 1017 9026 1026
rect 8974 983 8983 1017
rect 8983 983 9017 1017
rect 9017 983 9026 1017
rect 8974 974 9026 983
rect 8974 537 9026 546
rect 8974 503 8983 537
rect 8983 503 9017 537
rect 9017 503 9026 537
rect 8974 494 9026 503
rect 8974 377 9026 386
rect 8974 343 8983 377
rect 8983 343 9017 377
rect 9017 343 9026 377
rect 8974 334 9026 343
rect 8974 217 9026 226
rect 8974 183 8983 217
rect 8983 183 9017 217
rect 9017 183 9026 217
rect 8974 174 9026 183
rect 8974 57 9026 66
rect 8974 23 8983 57
rect 8983 23 9017 57
rect 9017 23 9026 57
rect 8974 14 9026 23
rect 9294 31417 9346 31426
rect 9294 31383 9303 31417
rect 9303 31383 9337 31417
rect 9337 31383 9346 31417
rect 9294 31374 9346 31383
rect 9294 31257 9346 31266
rect 9294 31223 9303 31257
rect 9303 31223 9337 31257
rect 9337 31223 9346 31257
rect 9294 31214 9346 31223
rect 9294 31097 9346 31106
rect 9294 31063 9303 31097
rect 9303 31063 9337 31097
rect 9337 31063 9346 31097
rect 9294 31054 9346 31063
rect 9294 30937 9346 30946
rect 9294 30903 9303 30937
rect 9303 30903 9337 30937
rect 9337 30903 9346 30937
rect 9294 30894 9346 30903
rect 9294 30777 9346 30786
rect 9294 30743 9303 30777
rect 9303 30743 9337 30777
rect 9337 30743 9346 30777
rect 9294 30734 9346 30743
rect 9294 30617 9346 30626
rect 9294 30583 9303 30617
rect 9303 30583 9337 30617
rect 9337 30583 9346 30617
rect 9294 30574 9346 30583
rect 9294 30457 9346 30466
rect 9294 30423 9303 30457
rect 9303 30423 9337 30457
rect 9337 30423 9346 30457
rect 9294 30414 9346 30423
rect 9294 30297 9346 30306
rect 9294 30263 9303 30297
rect 9303 30263 9337 30297
rect 9337 30263 9346 30297
rect 9294 30254 9346 30263
rect 9294 29977 9346 29986
rect 9294 29943 9303 29977
rect 9303 29943 9337 29977
rect 9337 29943 9346 29977
rect 9294 29934 9346 29943
rect 9294 29817 9346 29826
rect 9294 29783 9303 29817
rect 9303 29783 9337 29817
rect 9337 29783 9346 29817
rect 9294 29774 9346 29783
rect 9294 29657 9346 29666
rect 9294 29623 9303 29657
rect 9303 29623 9337 29657
rect 9337 29623 9346 29657
rect 9294 29614 9346 29623
rect 9294 29497 9346 29506
rect 9294 29463 9303 29497
rect 9303 29463 9337 29497
rect 9337 29463 9346 29497
rect 9294 29454 9346 29463
rect 9294 29337 9346 29346
rect 9294 29303 9303 29337
rect 9303 29303 9337 29337
rect 9337 29303 9346 29337
rect 9294 29294 9346 29303
rect 9294 29177 9346 29186
rect 9294 29143 9303 29177
rect 9303 29143 9337 29177
rect 9337 29143 9346 29177
rect 9294 29134 9346 29143
rect 9294 29017 9346 29026
rect 9294 28983 9303 29017
rect 9303 28983 9337 29017
rect 9337 28983 9346 29017
rect 9294 28974 9346 28983
rect 9294 28857 9346 28866
rect 9294 28823 9303 28857
rect 9303 28823 9337 28857
rect 9337 28823 9346 28857
rect 9294 28814 9346 28823
rect 9294 28057 9346 28066
rect 9294 28023 9303 28057
rect 9303 28023 9337 28057
rect 9337 28023 9346 28057
rect 9294 28014 9346 28023
rect 9294 27897 9346 27906
rect 9294 27863 9303 27897
rect 9303 27863 9337 27897
rect 9337 27863 9346 27897
rect 9294 27854 9346 27863
rect 9294 27737 9346 27746
rect 9294 27703 9303 27737
rect 9303 27703 9337 27737
rect 9337 27703 9346 27737
rect 9294 27694 9346 27703
rect 9294 27577 9346 27586
rect 9294 27543 9303 27577
rect 9303 27543 9337 27577
rect 9337 27543 9346 27577
rect 9294 27534 9346 27543
rect 9294 27417 9346 27426
rect 9294 27383 9303 27417
rect 9303 27383 9337 27417
rect 9337 27383 9346 27417
rect 9294 27374 9346 27383
rect 9294 27257 9346 27266
rect 9294 27223 9303 27257
rect 9303 27223 9337 27257
rect 9337 27223 9346 27257
rect 9294 27214 9346 27223
rect 9294 27097 9346 27106
rect 9294 27063 9303 27097
rect 9303 27063 9337 27097
rect 9337 27063 9346 27097
rect 9294 27054 9346 27063
rect 9294 26937 9346 26946
rect 9294 26903 9303 26937
rect 9303 26903 9337 26937
rect 9337 26903 9346 26937
rect 9294 26894 9346 26903
rect 9294 26137 9346 26146
rect 9294 26103 9303 26137
rect 9303 26103 9337 26137
rect 9337 26103 9346 26137
rect 9294 26094 9346 26103
rect 9294 25977 9346 25986
rect 9294 25943 9303 25977
rect 9303 25943 9337 25977
rect 9337 25943 9346 25977
rect 9294 25934 9346 25943
rect 9294 25817 9346 25826
rect 9294 25783 9303 25817
rect 9303 25783 9337 25817
rect 9337 25783 9346 25817
rect 9294 25774 9346 25783
rect 9294 25657 9346 25666
rect 9294 25623 9303 25657
rect 9303 25623 9337 25657
rect 9337 25623 9346 25657
rect 9294 25614 9346 25623
rect 9294 25497 9346 25506
rect 9294 25463 9303 25497
rect 9303 25463 9337 25497
rect 9337 25463 9346 25497
rect 9294 25454 9346 25463
rect 9294 25337 9346 25346
rect 9294 25303 9303 25337
rect 9303 25303 9337 25337
rect 9337 25303 9346 25337
rect 9294 25294 9346 25303
rect 9294 25177 9346 25186
rect 9294 25143 9303 25177
rect 9303 25143 9337 25177
rect 9337 25143 9346 25177
rect 9294 25134 9346 25143
rect 9294 25017 9346 25026
rect 9294 24983 9303 25017
rect 9303 24983 9337 25017
rect 9337 24983 9346 25017
rect 9294 24974 9346 24983
rect 9294 24697 9346 24706
rect 9294 24663 9303 24697
rect 9303 24663 9337 24697
rect 9337 24663 9346 24697
rect 9294 24654 9346 24663
rect 9294 24537 9346 24546
rect 9294 24503 9303 24537
rect 9303 24503 9337 24537
rect 9337 24503 9346 24537
rect 9294 24494 9346 24503
rect 9294 24377 9346 24386
rect 9294 24343 9303 24377
rect 9303 24343 9337 24377
rect 9337 24343 9346 24377
rect 9294 24334 9346 24343
rect 9294 24217 9346 24226
rect 9294 24183 9303 24217
rect 9303 24183 9337 24217
rect 9337 24183 9346 24217
rect 9294 24174 9346 24183
rect 9294 24057 9346 24066
rect 9294 24023 9303 24057
rect 9303 24023 9337 24057
rect 9337 24023 9346 24057
rect 9294 24014 9346 24023
rect 9294 23897 9346 23906
rect 9294 23863 9303 23897
rect 9303 23863 9337 23897
rect 9337 23863 9346 23897
rect 9294 23854 9346 23863
rect 9294 23737 9346 23746
rect 9294 23703 9303 23737
rect 9303 23703 9337 23737
rect 9337 23703 9346 23737
rect 9294 23694 9346 23703
rect 9294 23577 9346 23586
rect 9294 23543 9303 23577
rect 9303 23543 9337 23577
rect 9337 23543 9346 23577
rect 9294 23534 9346 23543
rect 9294 23417 9346 23426
rect 9294 23383 9303 23417
rect 9303 23383 9337 23417
rect 9337 23383 9346 23417
rect 9294 23374 9346 23383
rect 9294 23257 9346 23266
rect 9294 23223 9303 23257
rect 9303 23223 9337 23257
rect 9337 23223 9346 23257
rect 9294 23214 9346 23223
rect 9294 23097 9346 23106
rect 9294 23063 9303 23097
rect 9303 23063 9337 23097
rect 9337 23063 9346 23097
rect 9294 23054 9346 23063
rect 9294 22937 9346 22946
rect 9294 22903 9303 22937
rect 9303 22903 9337 22937
rect 9337 22903 9346 22937
rect 9294 22894 9346 22903
rect 9294 22777 9346 22786
rect 9294 22743 9303 22777
rect 9303 22743 9337 22777
rect 9337 22743 9346 22777
rect 9294 22734 9346 22743
rect 9294 22617 9346 22626
rect 9294 22583 9303 22617
rect 9303 22583 9337 22617
rect 9337 22583 9346 22617
rect 9294 22574 9346 22583
rect 9294 22457 9346 22466
rect 9294 22423 9303 22457
rect 9303 22423 9337 22457
rect 9337 22423 9346 22457
rect 9294 22414 9346 22423
rect 9294 22297 9346 22306
rect 9294 22263 9303 22297
rect 9303 22263 9337 22297
rect 9337 22263 9346 22297
rect 9294 22254 9346 22263
rect 9294 22137 9346 22146
rect 9294 22103 9303 22137
rect 9303 22103 9337 22137
rect 9337 22103 9346 22137
rect 9294 22094 9346 22103
rect 9294 21817 9346 21826
rect 9294 21783 9303 21817
rect 9303 21783 9337 21817
rect 9337 21783 9346 21817
rect 9294 21774 9346 21783
rect 9294 21657 9346 21666
rect 9294 21623 9303 21657
rect 9303 21623 9337 21657
rect 9337 21623 9346 21657
rect 9294 21614 9346 21623
rect 9294 21497 9346 21506
rect 9294 21463 9303 21497
rect 9303 21463 9337 21497
rect 9337 21463 9346 21497
rect 9294 21454 9346 21463
rect 9294 21337 9346 21346
rect 9294 21303 9303 21337
rect 9303 21303 9337 21337
rect 9337 21303 9346 21337
rect 9294 21294 9346 21303
rect 9294 21177 9346 21186
rect 9294 21143 9303 21177
rect 9303 21143 9337 21177
rect 9337 21143 9346 21177
rect 9294 21134 9346 21143
rect 9294 21017 9346 21026
rect 9294 20983 9303 21017
rect 9303 20983 9337 21017
rect 9337 20983 9346 21017
rect 9294 20974 9346 20983
rect 9294 20857 9346 20866
rect 9294 20823 9303 20857
rect 9303 20823 9337 20857
rect 9337 20823 9346 20857
rect 9294 20814 9346 20823
rect 9294 20697 9346 20706
rect 9294 20663 9303 20697
rect 9303 20663 9337 20697
rect 9337 20663 9346 20697
rect 9294 20654 9346 20663
rect 9294 19897 9346 19906
rect 9294 19863 9303 19897
rect 9303 19863 9337 19897
rect 9337 19863 9346 19897
rect 9294 19854 9346 19863
rect 9294 19737 9346 19746
rect 9294 19703 9303 19737
rect 9303 19703 9337 19737
rect 9337 19703 9346 19737
rect 9294 19694 9346 19703
rect 9294 19577 9346 19586
rect 9294 19543 9303 19577
rect 9303 19543 9337 19577
rect 9337 19543 9346 19577
rect 9294 19534 9346 19543
rect 9294 19417 9346 19426
rect 9294 19383 9303 19417
rect 9303 19383 9337 19417
rect 9337 19383 9346 19417
rect 9294 19374 9346 19383
rect 9294 19257 9346 19266
rect 9294 19223 9303 19257
rect 9303 19223 9337 19257
rect 9337 19223 9346 19257
rect 9294 19214 9346 19223
rect 9294 19097 9346 19106
rect 9294 19063 9303 19097
rect 9303 19063 9337 19097
rect 9337 19063 9346 19097
rect 9294 19054 9346 19063
rect 9294 18937 9346 18946
rect 9294 18903 9303 18937
rect 9303 18903 9337 18937
rect 9337 18903 9346 18937
rect 9294 18894 9346 18903
rect 9294 18777 9346 18786
rect 9294 18743 9303 18777
rect 9303 18743 9337 18777
rect 9337 18743 9346 18777
rect 9294 18734 9346 18743
rect 9294 17977 9346 17986
rect 9294 17943 9303 17977
rect 9303 17943 9337 17977
rect 9337 17943 9346 17977
rect 9294 17934 9346 17943
rect 9294 17817 9346 17826
rect 9294 17783 9303 17817
rect 9303 17783 9337 17817
rect 9337 17783 9346 17817
rect 9294 17774 9346 17783
rect 9294 17657 9346 17666
rect 9294 17623 9303 17657
rect 9303 17623 9337 17657
rect 9337 17623 9346 17657
rect 9294 17614 9346 17623
rect 9294 17497 9346 17506
rect 9294 17463 9303 17497
rect 9303 17463 9337 17497
rect 9337 17463 9346 17497
rect 9294 17454 9346 17463
rect 9294 17337 9346 17346
rect 9294 17303 9303 17337
rect 9303 17303 9337 17337
rect 9337 17303 9346 17337
rect 9294 17294 9346 17303
rect 9294 17177 9346 17186
rect 9294 17143 9303 17177
rect 9303 17143 9337 17177
rect 9337 17143 9346 17177
rect 9294 17134 9346 17143
rect 9294 17017 9346 17026
rect 9294 16983 9303 17017
rect 9303 16983 9337 17017
rect 9337 16983 9346 17017
rect 9294 16974 9346 16983
rect 9294 16857 9346 16866
rect 9294 16823 9303 16857
rect 9303 16823 9337 16857
rect 9337 16823 9346 16857
rect 9294 16814 9346 16823
rect 9294 16537 9346 16546
rect 9294 16503 9303 16537
rect 9303 16503 9337 16537
rect 9337 16503 9346 16537
rect 9294 16494 9346 16503
rect 9294 16377 9346 16386
rect 9294 16343 9303 16377
rect 9303 16343 9337 16377
rect 9337 16343 9346 16377
rect 9294 16334 9346 16343
rect 9294 16217 9346 16226
rect 9294 16183 9303 16217
rect 9303 16183 9337 16217
rect 9337 16183 9346 16217
rect 9294 16174 9346 16183
rect 9294 16057 9346 16066
rect 9294 16023 9303 16057
rect 9303 16023 9337 16057
rect 9337 16023 9346 16057
rect 9294 16014 9346 16023
rect 9294 15897 9346 15906
rect 9294 15863 9303 15897
rect 9303 15863 9337 15897
rect 9337 15863 9346 15897
rect 9294 15854 9346 15863
rect 9294 15737 9346 15746
rect 9294 15703 9303 15737
rect 9303 15703 9337 15737
rect 9337 15703 9346 15737
rect 9294 15694 9346 15703
rect 9294 15577 9346 15586
rect 9294 15543 9303 15577
rect 9303 15543 9337 15577
rect 9337 15543 9346 15577
rect 9294 15534 9346 15543
rect 9294 15417 9346 15426
rect 9294 15383 9303 15417
rect 9303 15383 9337 15417
rect 9337 15383 9346 15417
rect 9294 15374 9346 15383
rect 9294 15257 9346 15266
rect 9294 15223 9303 15257
rect 9303 15223 9337 15257
rect 9337 15223 9346 15257
rect 9294 15214 9346 15223
rect 9294 15097 9346 15106
rect 9294 15063 9303 15097
rect 9303 15063 9337 15097
rect 9337 15063 9346 15097
rect 9294 15054 9346 15063
rect 9294 14937 9346 14946
rect 9294 14903 9303 14937
rect 9303 14903 9337 14937
rect 9337 14903 9346 14937
rect 9294 14894 9346 14903
rect 9294 14777 9346 14786
rect 9294 14743 9303 14777
rect 9303 14743 9337 14777
rect 9337 14743 9346 14777
rect 9294 14734 9346 14743
rect 9294 14617 9346 14626
rect 9294 14583 9303 14617
rect 9303 14583 9337 14617
rect 9337 14583 9346 14617
rect 9294 14574 9346 14583
rect 9294 14457 9346 14466
rect 9294 14423 9303 14457
rect 9303 14423 9337 14457
rect 9337 14423 9346 14457
rect 9294 14414 9346 14423
rect 9294 14297 9346 14306
rect 9294 14263 9303 14297
rect 9303 14263 9337 14297
rect 9337 14263 9346 14297
rect 9294 14254 9346 14263
rect 9294 14137 9346 14146
rect 9294 14103 9303 14137
rect 9303 14103 9337 14137
rect 9337 14103 9346 14137
rect 9294 14094 9346 14103
rect 9294 13977 9346 13986
rect 9294 13943 9303 13977
rect 9303 13943 9337 13977
rect 9337 13943 9346 13977
rect 9294 13934 9346 13943
rect 9294 13657 9346 13666
rect 9294 13623 9303 13657
rect 9303 13623 9337 13657
rect 9337 13623 9346 13657
rect 9294 13614 9346 13623
rect 9294 13497 9346 13506
rect 9294 13463 9303 13497
rect 9303 13463 9337 13497
rect 9337 13463 9346 13497
rect 9294 13454 9346 13463
rect 9294 13337 9346 13346
rect 9294 13303 9303 13337
rect 9303 13303 9337 13337
rect 9337 13303 9346 13337
rect 9294 13294 9346 13303
rect 9294 13177 9346 13186
rect 9294 13143 9303 13177
rect 9303 13143 9337 13177
rect 9337 13143 9346 13177
rect 9294 13134 9346 13143
rect 9294 13017 9346 13026
rect 9294 12983 9303 13017
rect 9303 12983 9337 13017
rect 9337 12983 9346 13017
rect 9294 12974 9346 12983
rect 9294 12857 9346 12866
rect 9294 12823 9303 12857
rect 9303 12823 9337 12857
rect 9337 12823 9346 12857
rect 9294 12814 9346 12823
rect 9294 12697 9346 12706
rect 9294 12663 9303 12697
rect 9303 12663 9337 12697
rect 9337 12663 9346 12697
rect 9294 12654 9346 12663
rect 9294 12537 9346 12546
rect 9294 12503 9303 12537
rect 9303 12503 9337 12537
rect 9337 12503 9346 12537
rect 9294 12494 9346 12503
rect 9294 11737 9346 11746
rect 9294 11703 9303 11737
rect 9303 11703 9337 11737
rect 9337 11703 9346 11737
rect 9294 11694 9346 11703
rect 9294 11577 9346 11586
rect 9294 11543 9303 11577
rect 9303 11543 9337 11577
rect 9337 11543 9346 11577
rect 9294 11534 9346 11543
rect 9294 11417 9346 11426
rect 9294 11383 9303 11417
rect 9303 11383 9337 11417
rect 9337 11383 9346 11417
rect 9294 11374 9346 11383
rect 9294 11257 9346 11266
rect 9294 11223 9303 11257
rect 9303 11223 9337 11257
rect 9337 11223 9346 11257
rect 9294 11214 9346 11223
rect 9294 11097 9346 11106
rect 9294 11063 9303 11097
rect 9303 11063 9337 11097
rect 9337 11063 9346 11097
rect 9294 11054 9346 11063
rect 9294 10937 9346 10946
rect 9294 10903 9303 10937
rect 9303 10903 9337 10937
rect 9337 10903 9346 10937
rect 9294 10894 9346 10903
rect 9294 10777 9346 10786
rect 9294 10743 9303 10777
rect 9303 10743 9337 10777
rect 9337 10743 9346 10777
rect 9294 10734 9346 10743
rect 9294 10617 9346 10626
rect 9294 10583 9303 10617
rect 9303 10583 9337 10617
rect 9337 10583 9346 10617
rect 9294 10574 9346 10583
rect 9294 10457 9346 10466
rect 9294 10423 9303 10457
rect 9303 10423 9337 10457
rect 9337 10423 9346 10457
rect 9294 10414 9346 10423
rect 9294 10297 9346 10306
rect 9294 10263 9303 10297
rect 9303 10263 9337 10297
rect 9337 10263 9346 10297
rect 9294 10254 9346 10263
rect 9294 10137 9346 10146
rect 9294 10103 9303 10137
rect 9303 10103 9337 10137
rect 9337 10103 9346 10137
rect 9294 10094 9346 10103
rect 9294 9977 9346 9986
rect 9294 9943 9303 9977
rect 9303 9943 9337 9977
rect 9337 9943 9346 9977
rect 9294 9934 9346 9943
rect 9294 9817 9346 9826
rect 9294 9783 9303 9817
rect 9303 9783 9337 9817
rect 9337 9783 9346 9817
rect 9294 9774 9346 9783
rect 9294 9497 9346 9506
rect 9294 9463 9303 9497
rect 9303 9463 9337 9497
rect 9337 9463 9346 9497
rect 9294 9454 9346 9463
rect 9294 9337 9346 9346
rect 9294 9303 9303 9337
rect 9303 9303 9337 9337
rect 9337 9303 9346 9337
rect 9294 9294 9346 9303
rect 9294 9017 9346 9026
rect 9294 8983 9303 9017
rect 9303 8983 9337 9017
rect 9337 8983 9346 9017
rect 9294 8974 9346 8983
rect 9294 8857 9346 8866
rect 9294 8823 9303 8857
rect 9303 8823 9337 8857
rect 9337 8823 9346 8857
rect 9294 8814 9346 8823
rect 9294 8697 9346 8706
rect 9294 8663 9303 8697
rect 9303 8663 9337 8697
rect 9337 8663 9346 8697
rect 9294 8654 9346 8663
rect 9294 8537 9346 8546
rect 9294 8503 9303 8537
rect 9303 8503 9337 8537
rect 9337 8503 9346 8537
rect 9294 8494 9346 8503
rect 9294 8377 9346 8386
rect 9294 8343 9303 8377
rect 9303 8343 9337 8377
rect 9337 8343 9346 8377
rect 9294 8334 9346 8343
rect 9294 8217 9346 8226
rect 9294 8183 9303 8217
rect 9303 8183 9337 8217
rect 9337 8183 9346 8217
rect 9294 8174 9346 8183
rect 9294 8057 9346 8066
rect 9294 8023 9303 8057
rect 9303 8023 9337 8057
rect 9337 8023 9346 8057
rect 9294 8014 9346 8023
rect 9294 7897 9346 7906
rect 9294 7863 9303 7897
rect 9303 7863 9337 7897
rect 9337 7863 9346 7897
rect 9294 7854 9346 7863
rect 9294 7737 9346 7746
rect 9294 7703 9303 7737
rect 9303 7703 9337 7737
rect 9337 7703 9346 7737
rect 9294 7694 9346 7703
rect 9294 7417 9346 7426
rect 9294 7383 9303 7417
rect 9303 7383 9337 7417
rect 9337 7383 9346 7417
rect 9294 7374 9346 7383
rect 9294 7257 9346 7266
rect 9294 7223 9303 7257
rect 9303 7223 9337 7257
rect 9337 7223 9346 7257
rect 9294 7214 9346 7223
rect 9294 6937 9346 6946
rect 9294 6903 9303 6937
rect 9303 6903 9337 6937
rect 9337 6903 9346 6937
rect 9294 6894 9346 6903
rect 9294 6777 9346 6786
rect 9294 6743 9303 6777
rect 9303 6743 9337 6777
rect 9337 6743 9346 6777
rect 9294 6734 9346 6743
rect 9294 6457 9346 6466
rect 9294 6423 9303 6457
rect 9303 6423 9337 6457
rect 9337 6423 9346 6457
rect 9294 6414 9346 6423
rect 9294 6297 9346 6306
rect 9294 6263 9303 6297
rect 9303 6263 9337 6297
rect 9337 6263 9346 6297
rect 9294 6254 9346 6263
rect 9294 6137 9346 6146
rect 9294 6103 9303 6137
rect 9303 6103 9337 6137
rect 9337 6103 9346 6137
rect 9294 6094 9346 6103
rect 9294 5977 9346 5986
rect 9294 5943 9303 5977
rect 9303 5943 9337 5977
rect 9337 5943 9346 5977
rect 9294 5934 9346 5943
rect 9294 5817 9346 5826
rect 9294 5783 9303 5817
rect 9303 5783 9337 5817
rect 9337 5783 9346 5817
rect 9294 5774 9346 5783
rect 9294 5657 9346 5666
rect 9294 5623 9303 5657
rect 9303 5623 9337 5657
rect 9337 5623 9346 5657
rect 9294 5614 9346 5623
rect 9294 5497 9346 5506
rect 9294 5463 9303 5497
rect 9303 5463 9337 5497
rect 9337 5463 9346 5497
rect 9294 5454 9346 5463
rect 9294 5337 9346 5346
rect 9294 5303 9303 5337
rect 9303 5303 9337 5337
rect 9337 5303 9346 5337
rect 9294 5294 9346 5303
rect 9294 5177 9346 5186
rect 9294 5143 9303 5177
rect 9303 5143 9337 5177
rect 9337 5143 9346 5177
rect 9294 5134 9346 5143
rect 9294 5017 9346 5026
rect 9294 4983 9303 5017
rect 9303 4983 9337 5017
rect 9337 4983 9346 5017
rect 9294 4974 9346 4983
rect 9294 4857 9346 4866
rect 9294 4823 9303 4857
rect 9303 4823 9337 4857
rect 9337 4823 9346 4857
rect 9294 4814 9346 4823
rect 9294 4697 9346 4706
rect 9294 4663 9303 4697
rect 9303 4663 9337 4697
rect 9337 4663 9346 4697
rect 9294 4654 9346 4663
rect 9294 4537 9346 4546
rect 9294 4503 9303 4537
rect 9303 4503 9337 4537
rect 9337 4503 9346 4537
rect 9294 4494 9346 4503
rect 9294 4377 9346 4386
rect 9294 4343 9303 4377
rect 9303 4343 9337 4377
rect 9337 4343 9346 4377
rect 9294 4334 9346 4343
rect 9294 4217 9346 4226
rect 9294 4183 9303 4217
rect 9303 4183 9337 4217
rect 9337 4183 9346 4217
rect 9294 4174 9346 4183
rect 9294 4057 9346 4066
rect 9294 4023 9303 4057
rect 9303 4023 9337 4057
rect 9337 4023 9346 4057
rect 9294 4014 9346 4023
rect 9294 3897 9346 3906
rect 9294 3863 9303 3897
rect 9303 3863 9337 3897
rect 9337 3863 9346 3897
rect 9294 3854 9346 3863
rect 9294 3417 9346 3426
rect 9294 3383 9303 3417
rect 9303 3383 9337 3417
rect 9337 3383 9346 3417
rect 9294 3374 9346 3383
rect 9294 3257 9346 3266
rect 9294 3223 9303 3257
rect 9303 3223 9337 3257
rect 9337 3223 9346 3257
rect 9294 3214 9346 3223
rect 9294 3097 9346 3106
rect 9294 3063 9303 3097
rect 9303 3063 9337 3097
rect 9337 3063 9346 3097
rect 9294 3054 9346 3063
rect 9294 2937 9346 2946
rect 9294 2903 9303 2937
rect 9303 2903 9337 2937
rect 9337 2903 9346 2937
rect 9294 2894 9346 2903
rect 9294 2777 9346 2786
rect 9294 2743 9303 2777
rect 9303 2743 9337 2777
rect 9337 2743 9346 2777
rect 9294 2734 9346 2743
rect 9294 2617 9346 2626
rect 9294 2583 9303 2617
rect 9303 2583 9337 2617
rect 9337 2583 9346 2617
rect 9294 2574 9346 2583
rect 9294 2457 9346 2466
rect 9294 2423 9303 2457
rect 9303 2423 9337 2457
rect 9337 2423 9346 2457
rect 9294 2414 9346 2423
rect 9294 2297 9346 2306
rect 9294 2263 9303 2297
rect 9303 2263 9337 2297
rect 9337 2263 9346 2297
rect 9294 2254 9346 2263
rect 9294 2137 9346 2146
rect 9294 2103 9303 2137
rect 9303 2103 9337 2137
rect 9337 2103 9346 2137
rect 9294 2094 9346 2103
rect 9294 1977 9346 1986
rect 9294 1943 9303 1977
rect 9303 1943 9337 1977
rect 9337 1943 9346 1977
rect 9294 1934 9346 1943
rect 9294 1657 9346 1666
rect 9294 1623 9303 1657
rect 9303 1623 9337 1657
rect 9337 1623 9346 1657
rect 9294 1614 9346 1623
rect 9294 1497 9346 1506
rect 9294 1463 9303 1497
rect 9303 1463 9337 1497
rect 9337 1463 9346 1497
rect 9294 1454 9346 1463
rect 9294 1337 9346 1346
rect 9294 1303 9303 1337
rect 9303 1303 9337 1337
rect 9337 1303 9346 1337
rect 9294 1294 9346 1303
rect 9294 1177 9346 1186
rect 9294 1143 9303 1177
rect 9303 1143 9337 1177
rect 9337 1143 9346 1177
rect 9294 1134 9346 1143
rect 9294 1017 9346 1026
rect 9294 983 9303 1017
rect 9303 983 9337 1017
rect 9337 983 9346 1017
rect 9294 974 9346 983
rect 9294 537 9346 546
rect 9294 503 9303 537
rect 9303 503 9337 537
rect 9337 503 9346 537
rect 9294 494 9346 503
rect 9294 377 9346 386
rect 9294 343 9303 377
rect 9303 343 9337 377
rect 9337 343 9346 377
rect 9294 334 9346 343
rect 9294 217 9346 226
rect 9294 183 9303 217
rect 9303 183 9337 217
rect 9337 183 9346 217
rect 9294 174 9346 183
rect 9294 57 9346 66
rect 9294 23 9303 57
rect 9303 23 9337 57
rect 9337 23 9346 57
rect 9294 14 9346 23
rect 9454 31417 9506 31426
rect 9454 31383 9463 31417
rect 9463 31383 9497 31417
rect 9497 31383 9506 31417
rect 9454 31374 9506 31383
rect 9454 31257 9506 31266
rect 9454 31223 9463 31257
rect 9463 31223 9497 31257
rect 9497 31223 9506 31257
rect 9454 31214 9506 31223
rect 9454 31097 9506 31106
rect 9454 31063 9463 31097
rect 9463 31063 9497 31097
rect 9497 31063 9506 31097
rect 9454 31054 9506 31063
rect 9454 30937 9506 30946
rect 9454 30903 9463 30937
rect 9463 30903 9497 30937
rect 9497 30903 9506 30937
rect 9454 30894 9506 30903
rect 9454 30777 9506 30786
rect 9454 30743 9463 30777
rect 9463 30743 9497 30777
rect 9497 30743 9506 30777
rect 9454 30734 9506 30743
rect 9454 30617 9506 30626
rect 9454 30583 9463 30617
rect 9463 30583 9497 30617
rect 9497 30583 9506 30617
rect 9454 30574 9506 30583
rect 9454 30457 9506 30466
rect 9454 30423 9463 30457
rect 9463 30423 9497 30457
rect 9497 30423 9506 30457
rect 9454 30414 9506 30423
rect 9454 30297 9506 30306
rect 9454 30263 9463 30297
rect 9463 30263 9497 30297
rect 9497 30263 9506 30297
rect 9454 30254 9506 30263
rect 9454 29977 9506 29986
rect 9454 29943 9463 29977
rect 9463 29943 9497 29977
rect 9497 29943 9506 29977
rect 9454 29934 9506 29943
rect 9454 29817 9506 29826
rect 9454 29783 9463 29817
rect 9463 29783 9497 29817
rect 9497 29783 9506 29817
rect 9454 29774 9506 29783
rect 9454 29657 9506 29666
rect 9454 29623 9463 29657
rect 9463 29623 9497 29657
rect 9497 29623 9506 29657
rect 9454 29614 9506 29623
rect 9454 29497 9506 29506
rect 9454 29463 9463 29497
rect 9463 29463 9497 29497
rect 9497 29463 9506 29497
rect 9454 29454 9506 29463
rect 9454 29337 9506 29346
rect 9454 29303 9463 29337
rect 9463 29303 9497 29337
rect 9497 29303 9506 29337
rect 9454 29294 9506 29303
rect 9454 29177 9506 29186
rect 9454 29143 9463 29177
rect 9463 29143 9497 29177
rect 9497 29143 9506 29177
rect 9454 29134 9506 29143
rect 9454 29017 9506 29026
rect 9454 28983 9463 29017
rect 9463 28983 9497 29017
rect 9497 28983 9506 29017
rect 9454 28974 9506 28983
rect 9454 28857 9506 28866
rect 9454 28823 9463 28857
rect 9463 28823 9497 28857
rect 9497 28823 9506 28857
rect 9454 28814 9506 28823
rect 9454 28057 9506 28066
rect 9454 28023 9463 28057
rect 9463 28023 9497 28057
rect 9497 28023 9506 28057
rect 9454 28014 9506 28023
rect 9454 27897 9506 27906
rect 9454 27863 9463 27897
rect 9463 27863 9497 27897
rect 9497 27863 9506 27897
rect 9454 27854 9506 27863
rect 9454 27737 9506 27746
rect 9454 27703 9463 27737
rect 9463 27703 9497 27737
rect 9497 27703 9506 27737
rect 9454 27694 9506 27703
rect 9454 27577 9506 27586
rect 9454 27543 9463 27577
rect 9463 27543 9497 27577
rect 9497 27543 9506 27577
rect 9454 27534 9506 27543
rect 9454 27417 9506 27426
rect 9454 27383 9463 27417
rect 9463 27383 9497 27417
rect 9497 27383 9506 27417
rect 9454 27374 9506 27383
rect 9454 27257 9506 27266
rect 9454 27223 9463 27257
rect 9463 27223 9497 27257
rect 9497 27223 9506 27257
rect 9454 27214 9506 27223
rect 9454 27097 9506 27106
rect 9454 27063 9463 27097
rect 9463 27063 9497 27097
rect 9497 27063 9506 27097
rect 9454 27054 9506 27063
rect 9454 26937 9506 26946
rect 9454 26903 9463 26937
rect 9463 26903 9497 26937
rect 9497 26903 9506 26937
rect 9454 26894 9506 26903
rect 9454 26137 9506 26146
rect 9454 26103 9463 26137
rect 9463 26103 9497 26137
rect 9497 26103 9506 26137
rect 9454 26094 9506 26103
rect 9454 25977 9506 25986
rect 9454 25943 9463 25977
rect 9463 25943 9497 25977
rect 9497 25943 9506 25977
rect 9454 25934 9506 25943
rect 9454 25817 9506 25826
rect 9454 25783 9463 25817
rect 9463 25783 9497 25817
rect 9497 25783 9506 25817
rect 9454 25774 9506 25783
rect 9454 25657 9506 25666
rect 9454 25623 9463 25657
rect 9463 25623 9497 25657
rect 9497 25623 9506 25657
rect 9454 25614 9506 25623
rect 9454 25497 9506 25506
rect 9454 25463 9463 25497
rect 9463 25463 9497 25497
rect 9497 25463 9506 25497
rect 9454 25454 9506 25463
rect 9454 25337 9506 25346
rect 9454 25303 9463 25337
rect 9463 25303 9497 25337
rect 9497 25303 9506 25337
rect 9454 25294 9506 25303
rect 9454 25177 9506 25186
rect 9454 25143 9463 25177
rect 9463 25143 9497 25177
rect 9497 25143 9506 25177
rect 9454 25134 9506 25143
rect 9454 25017 9506 25026
rect 9454 24983 9463 25017
rect 9463 24983 9497 25017
rect 9497 24983 9506 25017
rect 9454 24974 9506 24983
rect 9454 24697 9506 24706
rect 9454 24663 9463 24697
rect 9463 24663 9497 24697
rect 9497 24663 9506 24697
rect 9454 24654 9506 24663
rect 9454 24537 9506 24546
rect 9454 24503 9463 24537
rect 9463 24503 9497 24537
rect 9497 24503 9506 24537
rect 9454 24494 9506 24503
rect 9454 24377 9506 24386
rect 9454 24343 9463 24377
rect 9463 24343 9497 24377
rect 9497 24343 9506 24377
rect 9454 24334 9506 24343
rect 9454 24217 9506 24226
rect 9454 24183 9463 24217
rect 9463 24183 9497 24217
rect 9497 24183 9506 24217
rect 9454 24174 9506 24183
rect 9454 24057 9506 24066
rect 9454 24023 9463 24057
rect 9463 24023 9497 24057
rect 9497 24023 9506 24057
rect 9454 24014 9506 24023
rect 9454 23897 9506 23906
rect 9454 23863 9463 23897
rect 9463 23863 9497 23897
rect 9497 23863 9506 23897
rect 9454 23854 9506 23863
rect 9454 23737 9506 23746
rect 9454 23703 9463 23737
rect 9463 23703 9497 23737
rect 9497 23703 9506 23737
rect 9454 23694 9506 23703
rect 9454 23577 9506 23586
rect 9454 23543 9463 23577
rect 9463 23543 9497 23577
rect 9497 23543 9506 23577
rect 9454 23534 9506 23543
rect 9454 23417 9506 23426
rect 9454 23383 9463 23417
rect 9463 23383 9497 23417
rect 9497 23383 9506 23417
rect 9454 23374 9506 23383
rect 9454 23257 9506 23266
rect 9454 23223 9463 23257
rect 9463 23223 9497 23257
rect 9497 23223 9506 23257
rect 9454 23214 9506 23223
rect 9454 23097 9506 23106
rect 9454 23063 9463 23097
rect 9463 23063 9497 23097
rect 9497 23063 9506 23097
rect 9454 23054 9506 23063
rect 9454 22937 9506 22946
rect 9454 22903 9463 22937
rect 9463 22903 9497 22937
rect 9497 22903 9506 22937
rect 9454 22894 9506 22903
rect 9454 22777 9506 22786
rect 9454 22743 9463 22777
rect 9463 22743 9497 22777
rect 9497 22743 9506 22777
rect 9454 22734 9506 22743
rect 9454 22617 9506 22626
rect 9454 22583 9463 22617
rect 9463 22583 9497 22617
rect 9497 22583 9506 22617
rect 9454 22574 9506 22583
rect 9454 22457 9506 22466
rect 9454 22423 9463 22457
rect 9463 22423 9497 22457
rect 9497 22423 9506 22457
rect 9454 22414 9506 22423
rect 9454 22297 9506 22306
rect 9454 22263 9463 22297
rect 9463 22263 9497 22297
rect 9497 22263 9506 22297
rect 9454 22254 9506 22263
rect 9454 22137 9506 22146
rect 9454 22103 9463 22137
rect 9463 22103 9497 22137
rect 9497 22103 9506 22137
rect 9454 22094 9506 22103
rect 9454 21817 9506 21826
rect 9454 21783 9463 21817
rect 9463 21783 9497 21817
rect 9497 21783 9506 21817
rect 9454 21774 9506 21783
rect 9454 21657 9506 21666
rect 9454 21623 9463 21657
rect 9463 21623 9497 21657
rect 9497 21623 9506 21657
rect 9454 21614 9506 21623
rect 9454 21497 9506 21506
rect 9454 21463 9463 21497
rect 9463 21463 9497 21497
rect 9497 21463 9506 21497
rect 9454 21454 9506 21463
rect 9454 21337 9506 21346
rect 9454 21303 9463 21337
rect 9463 21303 9497 21337
rect 9497 21303 9506 21337
rect 9454 21294 9506 21303
rect 9454 21177 9506 21186
rect 9454 21143 9463 21177
rect 9463 21143 9497 21177
rect 9497 21143 9506 21177
rect 9454 21134 9506 21143
rect 9454 21017 9506 21026
rect 9454 20983 9463 21017
rect 9463 20983 9497 21017
rect 9497 20983 9506 21017
rect 9454 20974 9506 20983
rect 9454 20857 9506 20866
rect 9454 20823 9463 20857
rect 9463 20823 9497 20857
rect 9497 20823 9506 20857
rect 9454 20814 9506 20823
rect 9454 20697 9506 20706
rect 9454 20663 9463 20697
rect 9463 20663 9497 20697
rect 9497 20663 9506 20697
rect 9454 20654 9506 20663
rect 9454 19897 9506 19906
rect 9454 19863 9463 19897
rect 9463 19863 9497 19897
rect 9497 19863 9506 19897
rect 9454 19854 9506 19863
rect 9454 19737 9506 19746
rect 9454 19703 9463 19737
rect 9463 19703 9497 19737
rect 9497 19703 9506 19737
rect 9454 19694 9506 19703
rect 9454 19577 9506 19586
rect 9454 19543 9463 19577
rect 9463 19543 9497 19577
rect 9497 19543 9506 19577
rect 9454 19534 9506 19543
rect 9454 19417 9506 19426
rect 9454 19383 9463 19417
rect 9463 19383 9497 19417
rect 9497 19383 9506 19417
rect 9454 19374 9506 19383
rect 9454 19257 9506 19266
rect 9454 19223 9463 19257
rect 9463 19223 9497 19257
rect 9497 19223 9506 19257
rect 9454 19214 9506 19223
rect 9454 19097 9506 19106
rect 9454 19063 9463 19097
rect 9463 19063 9497 19097
rect 9497 19063 9506 19097
rect 9454 19054 9506 19063
rect 9454 18937 9506 18946
rect 9454 18903 9463 18937
rect 9463 18903 9497 18937
rect 9497 18903 9506 18937
rect 9454 18894 9506 18903
rect 9454 18777 9506 18786
rect 9454 18743 9463 18777
rect 9463 18743 9497 18777
rect 9497 18743 9506 18777
rect 9454 18734 9506 18743
rect 9454 17977 9506 17986
rect 9454 17943 9463 17977
rect 9463 17943 9497 17977
rect 9497 17943 9506 17977
rect 9454 17934 9506 17943
rect 9454 17817 9506 17826
rect 9454 17783 9463 17817
rect 9463 17783 9497 17817
rect 9497 17783 9506 17817
rect 9454 17774 9506 17783
rect 9454 17657 9506 17666
rect 9454 17623 9463 17657
rect 9463 17623 9497 17657
rect 9497 17623 9506 17657
rect 9454 17614 9506 17623
rect 9454 17497 9506 17506
rect 9454 17463 9463 17497
rect 9463 17463 9497 17497
rect 9497 17463 9506 17497
rect 9454 17454 9506 17463
rect 9454 17337 9506 17346
rect 9454 17303 9463 17337
rect 9463 17303 9497 17337
rect 9497 17303 9506 17337
rect 9454 17294 9506 17303
rect 9454 17177 9506 17186
rect 9454 17143 9463 17177
rect 9463 17143 9497 17177
rect 9497 17143 9506 17177
rect 9454 17134 9506 17143
rect 9454 17017 9506 17026
rect 9454 16983 9463 17017
rect 9463 16983 9497 17017
rect 9497 16983 9506 17017
rect 9454 16974 9506 16983
rect 9454 16857 9506 16866
rect 9454 16823 9463 16857
rect 9463 16823 9497 16857
rect 9497 16823 9506 16857
rect 9454 16814 9506 16823
rect 9454 16537 9506 16546
rect 9454 16503 9463 16537
rect 9463 16503 9497 16537
rect 9497 16503 9506 16537
rect 9454 16494 9506 16503
rect 9454 16377 9506 16386
rect 9454 16343 9463 16377
rect 9463 16343 9497 16377
rect 9497 16343 9506 16377
rect 9454 16334 9506 16343
rect 9454 16217 9506 16226
rect 9454 16183 9463 16217
rect 9463 16183 9497 16217
rect 9497 16183 9506 16217
rect 9454 16174 9506 16183
rect 9454 16057 9506 16066
rect 9454 16023 9463 16057
rect 9463 16023 9497 16057
rect 9497 16023 9506 16057
rect 9454 16014 9506 16023
rect 9454 15897 9506 15906
rect 9454 15863 9463 15897
rect 9463 15863 9497 15897
rect 9497 15863 9506 15897
rect 9454 15854 9506 15863
rect 9454 15737 9506 15746
rect 9454 15703 9463 15737
rect 9463 15703 9497 15737
rect 9497 15703 9506 15737
rect 9454 15694 9506 15703
rect 9454 15577 9506 15586
rect 9454 15543 9463 15577
rect 9463 15543 9497 15577
rect 9497 15543 9506 15577
rect 9454 15534 9506 15543
rect 9454 15417 9506 15426
rect 9454 15383 9463 15417
rect 9463 15383 9497 15417
rect 9497 15383 9506 15417
rect 9454 15374 9506 15383
rect 9454 15257 9506 15266
rect 9454 15223 9463 15257
rect 9463 15223 9497 15257
rect 9497 15223 9506 15257
rect 9454 15214 9506 15223
rect 9454 15097 9506 15106
rect 9454 15063 9463 15097
rect 9463 15063 9497 15097
rect 9497 15063 9506 15097
rect 9454 15054 9506 15063
rect 9454 14937 9506 14946
rect 9454 14903 9463 14937
rect 9463 14903 9497 14937
rect 9497 14903 9506 14937
rect 9454 14894 9506 14903
rect 9454 14777 9506 14786
rect 9454 14743 9463 14777
rect 9463 14743 9497 14777
rect 9497 14743 9506 14777
rect 9454 14734 9506 14743
rect 9454 14617 9506 14626
rect 9454 14583 9463 14617
rect 9463 14583 9497 14617
rect 9497 14583 9506 14617
rect 9454 14574 9506 14583
rect 9454 14457 9506 14466
rect 9454 14423 9463 14457
rect 9463 14423 9497 14457
rect 9497 14423 9506 14457
rect 9454 14414 9506 14423
rect 9454 14297 9506 14306
rect 9454 14263 9463 14297
rect 9463 14263 9497 14297
rect 9497 14263 9506 14297
rect 9454 14254 9506 14263
rect 9454 14137 9506 14146
rect 9454 14103 9463 14137
rect 9463 14103 9497 14137
rect 9497 14103 9506 14137
rect 9454 14094 9506 14103
rect 9454 13977 9506 13986
rect 9454 13943 9463 13977
rect 9463 13943 9497 13977
rect 9497 13943 9506 13977
rect 9454 13934 9506 13943
rect 9454 13657 9506 13666
rect 9454 13623 9463 13657
rect 9463 13623 9497 13657
rect 9497 13623 9506 13657
rect 9454 13614 9506 13623
rect 9454 13497 9506 13506
rect 9454 13463 9463 13497
rect 9463 13463 9497 13497
rect 9497 13463 9506 13497
rect 9454 13454 9506 13463
rect 9454 13337 9506 13346
rect 9454 13303 9463 13337
rect 9463 13303 9497 13337
rect 9497 13303 9506 13337
rect 9454 13294 9506 13303
rect 9454 13177 9506 13186
rect 9454 13143 9463 13177
rect 9463 13143 9497 13177
rect 9497 13143 9506 13177
rect 9454 13134 9506 13143
rect 9454 13017 9506 13026
rect 9454 12983 9463 13017
rect 9463 12983 9497 13017
rect 9497 12983 9506 13017
rect 9454 12974 9506 12983
rect 9454 12857 9506 12866
rect 9454 12823 9463 12857
rect 9463 12823 9497 12857
rect 9497 12823 9506 12857
rect 9454 12814 9506 12823
rect 9454 12697 9506 12706
rect 9454 12663 9463 12697
rect 9463 12663 9497 12697
rect 9497 12663 9506 12697
rect 9454 12654 9506 12663
rect 9454 12537 9506 12546
rect 9454 12503 9463 12537
rect 9463 12503 9497 12537
rect 9497 12503 9506 12537
rect 9454 12494 9506 12503
rect 9454 11737 9506 11746
rect 9454 11703 9463 11737
rect 9463 11703 9497 11737
rect 9497 11703 9506 11737
rect 9454 11694 9506 11703
rect 9454 11577 9506 11586
rect 9454 11543 9463 11577
rect 9463 11543 9497 11577
rect 9497 11543 9506 11577
rect 9454 11534 9506 11543
rect 9454 11417 9506 11426
rect 9454 11383 9463 11417
rect 9463 11383 9497 11417
rect 9497 11383 9506 11417
rect 9454 11374 9506 11383
rect 9454 11257 9506 11266
rect 9454 11223 9463 11257
rect 9463 11223 9497 11257
rect 9497 11223 9506 11257
rect 9454 11214 9506 11223
rect 9454 11097 9506 11106
rect 9454 11063 9463 11097
rect 9463 11063 9497 11097
rect 9497 11063 9506 11097
rect 9454 11054 9506 11063
rect 9454 10937 9506 10946
rect 9454 10903 9463 10937
rect 9463 10903 9497 10937
rect 9497 10903 9506 10937
rect 9454 10894 9506 10903
rect 9454 10777 9506 10786
rect 9454 10743 9463 10777
rect 9463 10743 9497 10777
rect 9497 10743 9506 10777
rect 9454 10734 9506 10743
rect 9454 10617 9506 10626
rect 9454 10583 9463 10617
rect 9463 10583 9497 10617
rect 9497 10583 9506 10617
rect 9454 10574 9506 10583
rect 9454 10457 9506 10466
rect 9454 10423 9463 10457
rect 9463 10423 9497 10457
rect 9497 10423 9506 10457
rect 9454 10414 9506 10423
rect 9454 10297 9506 10306
rect 9454 10263 9463 10297
rect 9463 10263 9497 10297
rect 9497 10263 9506 10297
rect 9454 10254 9506 10263
rect 9454 10137 9506 10146
rect 9454 10103 9463 10137
rect 9463 10103 9497 10137
rect 9497 10103 9506 10137
rect 9454 10094 9506 10103
rect 9454 9977 9506 9986
rect 9454 9943 9463 9977
rect 9463 9943 9497 9977
rect 9497 9943 9506 9977
rect 9454 9934 9506 9943
rect 9454 9817 9506 9826
rect 9454 9783 9463 9817
rect 9463 9783 9497 9817
rect 9497 9783 9506 9817
rect 9454 9774 9506 9783
rect 9454 9497 9506 9506
rect 9454 9463 9463 9497
rect 9463 9463 9497 9497
rect 9497 9463 9506 9497
rect 9454 9454 9506 9463
rect 9454 9337 9506 9346
rect 9454 9303 9463 9337
rect 9463 9303 9497 9337
rect 9497 9303 9506 9337
rect 9454 9294 9506 9303
rect 9454 9017 9506 9026
rect 9454 8983 9463 9017
rect 9463 8983 9497 9017
rect 9497 8983 9506 9017
rect 9454 8974 9506 8983
rect 9454 8857 9506 8866
rect 9454 8823 9463 8857
rect 9463 8823 9497 8857
rect 9497 8823 9506 8857
rect 9454 8814 9506 8823
rect 9454 8697 9506 8706
rect 9454 8663 9463 8697
rect 9463 8663 9497 8697
rect 9497 8663 9506 8697
rect 9454 8654 9506 8663
rect 9454 8537 9506 8546
rect 9454 8503 9463 8537
rect 9463 8503 9497 8537
rect 9497 8503 9506 8537
rect 9454 8494 9506 8503
rect 9454 8377 9506 8386
rect 9454 8343 9463 8377
rect 9463 8343 9497 8377
rect 9497 8343 9506 8377
rect 9454 8334 9506 8343
rect 9454 8217 9506 8226
rect 9454 8183 9463 8217
rect 9463 8183 9497 8217
rect 9497 8183 9506 8217
rect 9454 8174 9506 8183
rect 9454 8057 9506 8066
rect 9454 8023 9463 8057
rect 9463 8023 9497 8057
rect 9497 8023 9506 8057
rect 9454 8014 9506 8023
rect 9454 7897 9506 7906
rect 9454 7863 9463 7897
rect 9463 7863 9497 7897
rect 9497 7863 9506 7897
rect 9454 7854 9506 7863
rect 9454 7737 9506 7746
rect 9454 7703 9463 7737
rect 9463 7703 9497 7737
rect 9497 7703 9506 7737
rect 9454 7694 9506 7703
rect 9454 7417 9506 7426
rect 9454 7383 9463 7417
rect 9463 7383 9497 7417
rect 9497 7383 9506 7417
rect 9454 7374 9506 7383
rect 9454 7257 9506 7266
rect 9454 7223 9463 7257
rect 9463 7223 9497 7257
rect 9497 7223 9506 7257
rect 9454 7214 9506 7223
rect 9454 6937 9506 6946
rect 9454 6903 9463 6937
rect 9463 6903 9497 6937
rect 9497 6903 9506 6937
rect 9454 6894 9506 6903
rect 9454 6777 9506 6786
rect 9454 6743 9463 6777
rect 9463 6743 9497 6777
rect 9497 6743 9506 6777
rect 9454 6734 9506 6743
rect 9454 6457 9506 6466
rect 9454 6423 9463 6457
rect 9463 6423 9497 6457
rect 9497 6423 9506 6457
rect 9454 6414 9506 6423
rect 9454 6297 9506 6306
rect 9454 6263 9463 6297
rect 9463 6263 9497 6297
rect 9497 6263 9506 6297
rect 9454 6254 9506 6263
rect 9454 6137 9506 6146
rect 9454 6103 9463 6137
rect 9463 6103 9497 6137
rect 9497 6103 9506 6137
rect 9454 6094 9506 6103
rect 9454 5977 9506 5986
rect 9454 5943 9463 5977
rect 9463 5943 9497 5977
rect 9497 5943 9506 5977
rect 9454 5934 9506 5943
rect 9454 5817 9506 5826
rect 9454 5783 9463 5817
rect 9463 5783 9497 5817
rect 9497 5783 9506 5817
rect 9454 5774 9506 5783
rect 9454 5657 9506 5666
rect 9454 5623 9463 5657
rect 9463 5623 9497 5657
rect 9497 5623 9506 5657
rect 9454 5614 9506 5623
rect 9454 5497 9506 5506
rect 9454 5463 9463 5497
rect 9463 5463 9497 5497
rect 9497 5463 9506 5497
rect 9454 5454 9506 5463
rect 9454 5337 9506 5346
rect 9454 5303 9463 5337
rect 9463 5303 9497 5337
rect 9497 5303 9506 5337
rect 9454 5294 9506 5303
rect 9454 5177 9506 5186
rect 9454 5143 9463 5177
rect 9463 5143 9497 5177
rect 9497 5143 9506 5177
rect 9454 5134 9506 5143
rect 9454 5017 9506 5026
rect 9454 4983 9463 5017
rect 9463 4983 9497 5017
rect 9497 4983 9506 5017
rect 9454 4974 9506 4983
rect 9454 4857 9506 4866
rect 9454 4823 9463 4857
rect 9463 4823 9497 4857
rect 9497 4823 9506 4857
rect 9454 4814 9506 4823
rect 9454 4697 9506 4706
rect 9454 4663 9463 4697
rect 9463 4663 9497 4697
rect 9497 4663 9506 4697
rect 9454 4654 9506 4663
rect 9454 4537 9506 4546
rect 9454 4503 9463 4537
rect 9463 4503 9497 4537
rect 9497 4503 9506 4537
rect 9454 4494 9506 4503
rect 9454 4377 9506 4386
rect 9454 4343 9463 4377
rect 9463 4343 9497 4377
rect 9497 4343 9506 4377
rect 9454 4334 9506 4343
rect 9454 4217 9506 4226
rect 9454 4183 9463 4217
rect 9463 4183 9497 4217
rect 9497 4183 9506 4217
rect 9454 4174 9506 4183
rect 9454 4057 9506 4066
rect 9454 4023 9463 4057
rect 9463 4023 9497 4057
rect 9497 4023 9506 4057
rect 9454 4014 9506 4023
rect 9454 3897 9506 3906
rect 9454 3863 9463 3897
rect 9463 3863 9497 3897
rect 9497 3863 9506 3897
rect 9454 3854 9506 3863
rect 9454 3417 9506 3426
rect 9454 3383 9463 3417
rect 9463 3383 9497 3417
rect 9497 3383 9506 3417
rect 9454 3374 9506 3383
rect 9454 3257 9506 3266
rect 9454 3223 9463 3257
rect 9463 3223 9497 3257
rect 9497 3223 9506 3257
rect 9454 3214 9506 3223
rect 9454 3097 9506 3106
rect 9454 3063 9463 3097
rect 9463 3063 9497 3097
rect 9497 3063 9506 3097
rect 9454 3054 9506 3063
rect 9454 2937 9506 2946
rect 9454 2903 9463 2937
rect 9463 2903 9497 2937
rect 9497 2903 9506 2937
rect 9454 2894 9506 2903
rect 9454 2777 9506 2786
rect 9454 2743 9463 2777
rect 9463 2743 9497 2777
rect 9497 2743 9506 2777
rect 9454 2734 9506 2743
rect 9454 2617 9506 2626
rect 9454 2583 9463 2617
rect 9463 2583 9497 2617
rect 9497 2583 9506 2617
rect 9454 2574 9506 2583
rect 9454 2457 9506 2466
rect 9454 2423 9463 2457
rect 9463 2423 9497 2457
rect 9497 2423 9506 2457
rect 9454 2414 9506 2423
rect 9454 2297 9506 2306
rect 9454 2263 9463 2297
rect 9463 2263 9497 2297
rect 9497 2263 9506 2297
rect 9454 2254 9506 2263
rect 9454 2137 9506 2146
rect 9454 2103 9463 2137
rect 9463 2103 9497 2137
rect 9497 2103 9506 2137
rect 9454 2094 9506 2103
rect 9454 1977 9506 1986
rect 9454 1943 9463 1977
rect 9463 1943 9497 1977
rect 9497 1943 9506 1977
rect 9454 1934 9506 1943
rect 9454 1657 9506 1666
rect 9454 1623 9463 1657
rect 9463 1623 9497 1657
rect 9497 1623 9506 1657
rect 9454 1614 9506 1623
rect 9454 1497 9506 1506
rect 9454 1463 9463 1497
rect 9463 1463 9497 1497
rect 9497 1463 9506 1497
rect 9454 1454 9506 1463
rect 9454 1337 9506 1346
rect 9454 1303 9463 1337
rect 9463 1303 9497 1337
rect 9497 1303 9506 1337
rect 9454 1294 9506 1303
rect 9454 1177 9506 1186
rect 9454 1143 9463 1177
rect 9463 1143 9497 1177
rect 9497 1143 9506 1177
rect 9454 1134 9506 1143
rect 9454 1017 9506 1026
rect 9454 983 9463 1017
rect 9463 983 9497 1017
rect 9497 983 9506 1017
rect 9454 974 9506 983
rect 9454 537 9506 546
rect 9454 503 9463 537
rect 9463 503 9497 537
rect 9497 503 9506 537
rect 9454 494 9506 503
rect 9454 377 9506 386
rect 9454 343 9463 377
rect 9463 343 9497 377
rect 9497 343 9506 377
rect 9454 334 9506 343
rect 9454 217 9506 226
rect 9454 183 9463 217
rect 9463 183 9497 217
rect 9497 183 9506 217
rect 9454 174 9506 183
rect 9454 57 9506 66
rect 9454 23 9463 57
rect 9463 23 9497 57
rect 9497 23 9506 57
rect 9454 14 9506 23
rect 9774 31417 9826 31426
rect 9774 31383 9783 31417
rect 9783 31383 9817 31417
rect 9817 31383 9826 31417
rect 9774 31374 9826 31383
rect 9774 31257 9826 31266
rect 9774 31223 9783 31257
rect 9783 31223 9817 31257
rect 9817 31223 9826 31257
rect 9774 31214 9826 31223
rect 9774 31097 9826 31106
rect 9774 31063 9783 31097
rect 9783 31063 9817 31097
rect 9817 31063 9826 31097
rect 9774 31054 9826 31063
rect 9774 30937 9826 30946
rect 9774 30903 9783 30937
rect 9783 30903 9817 30937
rect 9817 30903 9826 30937
rect 9774 30894 9826 30903
rect 9774 30777 9826 30786
rect 9774 30743 9783 30777
rect 9783 30743 9817 30777
rect 9817 30743 9826 30777
rect 9774 30734 9826 30743
rect 9774 30617 9826 30626
rect 9774 30583 9783 30617
rect 9783 30583 9817 30617
rect 9817 30583 9826 30617
rect 9774 30574 9826 30583
rect 9774 30457 9826 30466
rect 9774 30423 9783 30457
rect 9783 30423 9817 30457
rect 9817 30423 9826 30457
rect 9774 30414 9826 30423
rect 9774 30297 9826 30306
rect 9774 30263 9783 30297
rect 9783 30263 9817 30297
rect 9817 30263 9826 30297
rect 9774 30254 9826 30263
rect 9774 29977 9826 29986
rect 9774 29943 9783 29977
rect 9783 29943 9817 29977
rect 9817 29943 9826 29977
rect 9774 29934 9826 29943
rect 9774 29817 9826 29826
rect 9774 29783 9783 29817
rect 9783 29783 9817 29817
rect 9817 29783 9826 29817
rect 9774 29774 9826 29783
rect 9774 29657 9826 29666
rect 9774 29623 9783 29657
rect 9783 29623 9817 29657
rect 9817 29623 9826 29657
rect 9774 29614 9826 29623
rect 9774 29497 9826 29506
rect 9774 29463 9783 29497
rect 9783 29463 9817 29497
rect 9817 29463 9826 29497
rect 9774 29454 9826 29463
rect 9774 29337 9826 29346
rect 9774 29303 9783 29337
rect 9783 29303 9817 29337
rect 9817 29303 9826 29337
rect 9774 29294 9826 29303
rect 9774 29177 9826 29186
rect 9774 29143 9783 29177
rect 9783 29143 9817 29177
rect 9817 29143 9826 29177
rect 9774 29134 9826 29143
rect 9774 29017 9826 29026
rect 9774 28983 9783 29017
rect 9783 28983 9817 29017
rect 9817 28983 9826 29017
rect 9774 28974 9826 28983
rect 9774 28857 9826 28866
rect 9774 28823 9783 28857
rect 9783 28823 9817 28857
rect 9817 28823 9826 28857
rect 9774 28814 9826 28823
rect 9774 28057 9826 28066
rect 9774 28023 9783 28057
rect 9783 28023 9817 28057
rect 9817 28023 9826 28057
rect 9774 28014 9826 28023
rect 9774 27897 9826 27906
rect 9774 27863 9783 27897
rect 9783 27863 9817 27897
rect 9817 27863 9826 27897
rect 9774 27854 9826 27863
rect 9774 27737 9826 27746
rect 9774 27703 9783 27737
rect 9783 27703 9817 27737
rect 9817 27703 9826 27737
rect 9774 27694 9826 27703
rect 9774 27577 9826 27586
rect 9774 27543 9783 27577
rect 9783 27543 9817 27577
rect 9817 27543 9826 27577
rect 9774 27534 9826 27543
rect 9774 27417 9826 27426
rect 9774 27383 9783 27417
rect 9783 27383 9817 27417
rect 9817 27383 9826 27417
rect 9774 27374 9826 27383
rect 9774 27257 9826 27266
rect 9774 27223 9783 27257
rect 9783 27223 9817 27257
rect 9817 27223 9826 27257
rect 9774 27214 9826 27223
rect 9774 27097 9826 27106
rect 9774 27063 9783 27097
rect 9783 27063 9817 27097
rect 9817 27063 9826 27097
rect 9774 27054 9826 27063
rect 9774 26937 9826 26946
rect 9774 26903 9783 26937
rect 9783 26903 9817 26937
rect 9817 26903 9826 26937
rect 9774 26894 9826 26903
rect 9774 26137 9826 26146
rect 9774 26103 9783 26137
rect 9783 26103 9817 26137
rect 9817 26103 9826 26137
rect 9774 26094 9826 26103
rect 9774 25977 9826 25986
rect 9774 25943 9783 25977
rect 9783 25943 9817 25977
rect 9817 25943 9826 25977
rect 9774 25934 9826 25943
rect 9774 25817 9826 25826
rect 9774 25783 9783 25817
rect 9783 25783 9817 25817
rect 9817 25783 9826 25817
rect 9774 25774 9826 25783
rect 9774 25657 9826 25666
rect 9774 25623 9783 25657
rect 9783 25623 9817 25657
rect 9817 25623 9826 25657
rect 9774 25614 9826 25623
rect 9774 25497 9826 25506
rect 9774 25463 9783 25497
rect 9783 25463 9817 25497
rect 9817 25463 9826 25497
rect 9774 25454 9826 25463
rect 9774 25337 9826 25346
rect 9774 25303 9783 25337
rect 9783 25303 9817 25337
rect 9817 25303 9826 25337
rect 9774 25294 9826 25303
rect 9774 25177 9826 25186
rect 9774 25143 9783 25177
rect 9783 25143 9817 25177
rect 9817 25143 9826 25177
rect 9774 25134 9826 25143
rect 9774 25017 9826 25026
rect 9774 24983 9783 25017
rect 9783 24983 9817 25017
rect 9817 24983 9826 25017
rect 9774 24974 9826 24983
rect 9774 24697 9826 24706
rect 9774 24663 9783 24697
rect 9783 24663 9817 24697
rect 9817 24663 9826 24697
rect 9774 24654 9826 24663
rect 9774 24537 9826 24546
rect 9774 24503 9783 24537
rect 9783 24503 9817 24537
rect 9817 24503 9826 24537
rect 9774 24494 9826 24503
rect 9774 24377 9826 24386
rect 9774 24343 9783 24377
rect 9783 24343 9817 24377
rect 9817 24343 9826 24377
rect 9774 24334 9826 24343
rect 9774 24217 9826 24226
rect 9774 24183 9783 24217
rect 9783 24183 9817 24217
rect 9817 24183 9826 24217
rect 9774 24174 9826 24183
rect 9774 24057 9826 24066
rect 9774 24023 9783 24057
rect 9783 24023 9817 24057
rect 9817 24023 9826 24057
rect 9774 24014 9826 24023
rect 9774 23897 9826 23906
rect 9774 23863 9783 23897
rect 9783 23863 9817 23897
rect 9817 23863 9826 23897
rect 9774 23854 9826 23863
rect 9774 23737 9826 23746
rect 9774 23703 9783 23737
rect 9783 23703 9817 23737
rect 9817 23703 9826 23737
rect 9774 23694 9826 23703
rect 9774 23577 9826 23586
rect 9774 23543 9783 23577
rect 9783 23543 9817 23577
rect 9817 23543 9826 23577
rect 9774 23534 9826 23543
rect 9774 23417 9826 23426
rect 9774 23383 9783 23417
rect 9783 23383 9817 23417
rect 9817 23383 9826 23417
rect 9774 23374 9826 23383
rect 9774 23257 9826 23266
rect 9774 23223 9783 23257
rect 9783 23223 9817 23257
rect 9817 23223 9826 23257
rect 9774 23214 9826 23223
rect 9774 23097 9826 23106
rect 9774 23063 9783 23097
rect 9783 23063 9817 23097
rect 9817 23063 9826 23097
rect 9774 23054 9826 23063
rect 9774 22937 9826 22946
rect 9774 22903 9783 22937
rect 9783 22903 9817 22937
rect 9817 22903 9826 22937
rect 9774 22894 9826 22903
rect 9774 22777 9826 22786
rect 9774 22743 9783 22777
rect 9783 22743 9817 22777
rect 9817 22743 9826 22777
rect 9774 22734 9826 22743
rect 9774 22617 9826 22626
rect 9774 22583 9783 22617
rect 9783 22583 9817 22617
rect 9817 22583 9826 22617
rect 9774 22574 9826 22583
rect 9774 22457 9826 22466
rect 9774 22423 9783 22457
rect 9783 22423 9817 22457
rect 9817 22423 9826 22457
rect 9774 22414 9826 22423
rect 9774 22297 9826 22306
rect 9774 22263 9783 22297
rect 9783 22263 9817 22297
rect 9817 22263 9826 22297
rect 9774 22254 9826 22263
rect 9774 22137 9826 22146
rect 9774 22103 9783 22137
rect 9783 22103 9817 22137
rect 9817 22103 9826 22137
rect 9774 22094 9826 22103
rect 9774 21817 9826 21826
rect 9774 21783 9783 21817
rect 9783 21783 9817 21817
rect 9817 21783 9826 21817
rect 9774 21774 9826 21783
rect 9774 21657 9826 21666
rect 9774 21623 9783 21657
rect 9783 21623 9817 21657
rect 9817 21623 9826 21657
rect 9774 21614 9826 21623
rect 9774 21497 9826 21506
rect 9774 21463 9783 21497
rect 9783 21463 9817 21497
rect 9817 21463 9826 21497
rect 9774 21454 9826 21463
rect 9774 21337 9826 21346
rect 9774 21303 9783 21337
rect 9783 21303 9817 21337
rect 9817 21303 9826 21337
rect 9774 21294 9826 21303
rect 9774 21177 9826 21186
rect 9774 21143 9783 21177
rect 9783 21143 9817 21177
rect 9817 21143 9826 21177
rect 9774 21134 9826 21143
rect 9774 21017 9826 21026
rect 9774 20983 9783 21017
rect 9783 20983 9817 21017
rect 9817 20983 9826 21017
rect 9774 20974 9826 20983
rect 9774 20857 9826 20866
rect 9774 20823 9783 20857
rect 9783 20823 9817 20857
rect 9817 20823 9826 20857
rect 9774 20814 9826 20823
rect 9774 20697 9826 20706
rect 9774 20663 9783 20697
rect 9783 20663 9817 20697
rect 9817 20663 9826 20697
rect 9774 20654 9826 20663
rect 9774 19897 9826 19906
rect 9774 19863 9783 19897
rect 9783 19863 9817 19897
rect 9817 19863 9826 19897
rect 9774 19854 9826 19863
rect 9774 19737 9826 19746
rect 9774 19703 9783 19737
rect 9783 19703 9817 19737
rect 9817 19703 9826 19737
rect 9774 19694 9826 19703
rect 9774 19577 9826 19586
rect 9774 19543 9783 19577
rect 9783 19543 9817 19577
rect 9817 19543 9826 19577
rect 9774 19534 9826 19543
rect 9774 19417 9826 19426
rect 9774 19383 9783 19417
rect 9783 19383 9817 19417
rect 9817 19383 9826 19417
rect 9774 19374 9826 19383
rect 9774 19257 9826 19266
rect 9774 19223 9783 19257
rect 9783 19223 9817 19257
rect 9817 19223 9826 19257
rect 9774 19214 9826 19223
rect 9774 19097 9826 19106
rect 9774 19063 9783 19097
rect 9783 19063 9817 19097
rect 9817 19063 9826 19097
rect 9774 19054 9826 19063
rect 9774 18937 9826 18946
rect 9774 18903 9783 18937
rect 9783 18903 9817 18937
rect 9817 18903 9826 18937
rect 9774 18894 9826 18903
rect 9774 18777 9826 18786
rect 9774 18743 9783 18777
rect 9783 18743 9817 18777
rect 9817 18743 9826 18777
rect 9774 18734 9826 18743
rect 9774 17977 9826 17986
rect 9774 17943 9783 17977
rect 9783 17943 9817 17977
rect 9817 17943 9826 17977
rect 9774 17934 9826 17943
rect 9774 17817 9826 17826
rect 9774 17783 9783 17817
rect 9783 17783 9817 17817
rect 9817 17783 9826 17817
rect 9774 17774 9826 17783
rect 9774 17657 9826 17666
rect 9774 17623 9783 17657
rect 9783 17623 9817 17657
rect 9817 17623 9826 17657
rect 9774 17614 9826 17623
rect 9774 17497 9826 17506
rect 9774 17463 9783 17497
rect 9783 17463 9817 17497
rect 9817 17463 9826 17497
rect 9774 17454 9826 17463
rect 9774 17337 9826 17346
rect 9774 17303 9783 17337
rect 9783 17303 9817 17337
rect 9817 17303 9826 17337
rect 9774 17294 9826 17303
rect 9774 17177 9826 17186
rect 9774 17143 9783 17177
rect 9783 17143 9817 17177
rect 9817 17143 9826 17177
rect 9774 17134 9826 17143
rect 9774 17017 9826 17026
rect 9774 16983 9783 17017
rect 9783 16983 9817 17017
rect 9817 16983 9826 17017
rect 9774 16974 9826 16983
rect 9774 16857 9826 16866
rect 9774 16823 9783 16857
rect 9783 16823 9817 16857
rect 9817 16823 9826 16857
rect 9774 16814 9826 16823
rect 9774 16537 9826 16546
rect 9774 16503 9783 16537
rect 9783 16503 9817 16537
rect 9817 16503 9826 16537
rect 9774 16494 9826 16503
rect 9774 16377 9826 16386
rect 9774 16343 9783 16377
rect 9783 16343 9817 16377
rect 9817 16343 9826 16377
rect 9774 16334 9826 16343
rect 9774 16217 9826 16226
rect 9774 16183 9783 16217
rect 9783 16183 9817 16217
rect 9817 16183 9826 16217
rect 9774 16174 9826 16183
rect 9774 16057 9826 16066
rect 9774 16023 9783 16057
rect 9783 16023 9817 16057
rect 9817 16023 9826 16057
rect 9774 16014 9826 16023
rect 9774 15897 9826 15906
rect 9774 15863 9783 15897
rect 9783 15863 9817 15897
rect 9817 15863 9826 15897
rect 9774 15854 9826 15863
rect 9774 15737 9826 15746
rect 9774 15703 9783 15737
rect 9783 15703 9817 15737
rect 9817 15703 9826 15737
rect 9774 15694 9826 15703
rect 9774 15577 9826 15586
rect 9774 15543 9783 15577
rect 9783 15543 9817 15577
rect 9817 15543 9826 15577
rect 9774 15534 9826 15543
rect 9774 15417 9826 15426
rect 9774 15383 9783 15417
rect 9783 15383 9817 15417
rect 9817 15383 9826 15417
rect 9774 15374 9826 15383
rect 9774 15257 9826 15266
rect 9774 15223 9783 15257
rect 9783 15223 9817 15257
rect 9817 15223 9826 15257
rect 9774 15214 9826 15223
rect 9774 15097 9826 15106
rect 9774 15063 9783 15097
rect 9783 15063 9817 15097
rect 9817 15063 9826 15097
rect 9774 15054 9826 15063
rect 9774 14937 9826 14946
rect 9774 14903 9783 14937
rect 9783 14903 9817 14937
rect 9817 14903 9826 14937
rect 9774 14894 9826 14903
rect 9774 14777 9826 14786
rect 9774 14743 9783 14777
rect 9783 14743 9817 14777
rect 9817 14743 9826 14777
rect 9774 14734 9826 14743
rect 9774 14617 9826 14626
rect 9774 14583 9783 14617
rect 9783 14583 9817 14617
rect 9817 14583 9826 14617
rect 9774 14574 9826 14583
rect 9774 14457 9826 14466
rect 9774 14423 9783 14457
rect 9783 14423 9817 14457
rect 9817 14423 9826 14457
rect 9774 14414 9826 14423
rect 9774 14297 9826 14306
rect 9774 14263 9783 14297
rect 9783 14263 9817 14297
rect 9817 14263 9826 14297
rect 9774 14254 9826 14263
rect 9774 14137 9826 14146
rect 9774 14103 9783 14137
rect 9783 14103 9817 14137
rect 9817 14103 9826 14137
rect 9774 14094 9826 14103
rect 9774 13977 9826 13986
rect 9774 13943 9783 13977
rect 9783 13943 9817 13977
rect 9817 13943 9826 13977
rect 9774 13934 9826 13943
rect 9774 13657 9826 13666
rect 9774 13623 9783 13657
rect 9783 13623 9817 13657
rect 9817 13623 9826 13657
rect 9774 13614 9826 13623
rect 9774 13497 9826 13506
rect 9774 13463 9783 13497
rect 9783 13463 9817 13497
rect 9817 13463 9826 13497
rect 9774 13454 9826 13463
rect 9774 13337 9826 13346
rect 9774 13303 9783 13337
rect 9783 13303 9817 13337
rect 9817 13303 9826 13337
rect 9774 13294 9826 13303
rect 9774 13177 9826 13186
rect 9774 13143 9783 13177
rect 9783 13143 9817 13177
rect 9817 13143 9826 13177
rect 9774 13134 9826 13143
rect 9774 13017 9826 13026
rect 9774 12983 9783 13017
rect 9783 12983 9817 13017
rect 9817 12983 9826 13017
rect 9774 12974 9826 12983
rect 9774 12857 9826 12866
rect 9774 12823 9783 12857
rect 9783 12823 9817 12857
rect 9817 12823 9826 12857
rect 9774 12814 9826 12823
rect 9774 12697 9826 12706
rect 9774 12663 9783 12697
rect 9783 12663 9817 12697
rect 9817 12663 9826 12697
rect 9774 12654 9826 12663
rect 9774 12537 9826 12546
rect 9774 12503 9783 12537
rect 9783 12503 9817 12537
rect 9817 12503 9826 12537
rect 9774 12494 9826 12503
rect 9774 11737 9826 11746
rect 9774 11703 9783 11737
rect 9783 11703 9817 11737
rect 9817 11703 9826 11737
rect 9774 11694 9826 11703
rect 9774 11577 9826 11586
rect 9774 11543 9783 11577
rect 9783 11543 9817 11577
rect 9817 11543 9826 11577
rect 9774 11534 9826 11543
rect 9774 11417 9826 11426
rect 9774 11383 9783 11417
rect 9783 11383 9817 11417
rect 9817 11383 9826 11417
rect 9774 11374 9826 11383
rect 9774 11257 9826 11266
rect 9774 11223 9783 11257
rect 9783 11223 9817 11257
rect 9817 11223 9826 11257
rect 9774 11214 9826 11223
rect 9774 11097 9826 11106
rect 9774 11063 9783 11097
rect 9783 11063 9817 11097
rect 9817 11063 9826 11097
rect 9774 11054 9826 11063
rect 9774 10937 9826 10946
rect 9774 10903 9783 10937
rect 9783 10903 9817 10937
rect 9817 10903 9826 10937
rect 9774 10894 9826 10903
rect 9774 10777 9826 10786
rect 9774 10743 9783 10777
rect 9783 10743 9817 10777
rect 9817 10743 9826 10777
rect 9774 10734 9826 10743
rect 9774 10617 9826 10626
rect 9774 10583 9783 10617
rect 9783 10583 9817 10617
rect 9817 10583 9826 10617
rect 9774 10574 9826 10583
rect 9774 10457 9826 10466
rect 9774 10423 9783 10457
rect 9783 10423 9817 10457
rect 9817 10423 9826 10457
rect 9774 10414 9826 10423
rect 9774 10297 9826 10306
rect 9774 10263 9783 10297
rect 9783 10263 9817 10297
rect 9817 10263 9826 10297
rect 9774 10254 9826 10263
rect 9774 10137 9826 10146
rect 9774 10103 9783 10137
rect 9783 10103 9817 10137
rect 9817 10103 9826 10137
rect 9774 10094 9826 10103
rect 9774 9977 9826 9986
rect 9774 9943 9783 9977
rect 9783 9943 9817 9977
rect 9817 9943 9826 9977
rect 9774 9934 9826 9943
rect 9774 9817 9826 9826
rect 9774 9783 9783 9817
rect 9783 9783 9817 9817
rect 9817 9783 9826 9817
rect 9774 9774 9826 9783
rect 9774 9497 9826 9506
rect 9774 9463 9783 9497
rect 9783 9463 9817 9497
rect 9817 9463 9826 9497
rect 9774 9454 9826 9463
rect 9774 9337 9826 9346
rect 9774 9303 9783 9337
rect 9783 9303 9817 9337
rect 9817 9303 9826 9337
rect 9774 9294 9826 9303
rect 9774 9017 9826 9026
rect 9774 8983 9783 9017
rect 9783 8983 9817 9017
rect 9817 8983 9826 9017
rect 9774 8974 9826 8983
rect 9774 8857 9826 8866
rect 9774 8823 9783 8857
rect 9783 8823 9817 8857
rect 9817 8823 9826 8857
rect 9774 8814 9826 8823
rect 9774 8697 9826 8706
rect 9774 8663 9783 8697
rect 9783 8663 9817 8697
rect 9817 8663 9826 8697
rect 9774 8654 9826 8663
rect 9774 8537 9826 8546
rect 9774 8503 9783 8537
rect 9783 8503 9817 8537
rect 9817 8503 9826 8537
rect 9774 8494 9826 8503
rect 9774 8377 9826 8386
rect 9774 8343 9783 8377
rect 9783 8343 9817 8377
rect 9817 8343 9826 8377
rect 9774 8334 9826 8343
rect 9774 8217 9826 8226
rect 9774 8183 9783 8217
rect 9783 8183 9817 8217
rect 9817 8183 9826 8217
rect 9774 8174 9826 8183
rect 9774 8057 9826 8066
rect 9774 8023 9783 8057
rect 9783 8023 9817 8057
rect 9817 8023 9826 8057
rect 9774 8014 9826 8023
rect 9774 7897 9826 7906
rect 9774 7863 9783 7897
rect 9783 7863 9817 7897
rect 9817 7863 9826 7897
rect 9774 7854 9826 7863
rect 9774 7737 9826 7746
rect 9774 7703 9783 7737
rect 9783 7703 9817 7737
rect 9817 7703 9826 7737
rect 9774 7694 9826 7703
rect 9774 7417 9826 7426
rect 9774 7383 9783 7417
rect 9783 7383 9817 7417
rect 9817 7383 9826 7417
rect 9774 7374 9826 7383
rect 9774 7257 9826 7266
rect 9774 7223 9783 7257
rect 9783 7223 9817 7257
rect 9817 7223 9826 7257
rect 9774 7214 9826 7223
rect 9774 6937 9826 6946
rect 9774 6903 9783 6937
rect 9783 6903 9817 6937
rect 9817 6903 9826 6937
rect 9774 6894 9826 6903
rect 9774 6777 9826 6786
rect 9774 6743 9783 6777
rect 9783 6743 9817 6777
rect 9817 6743 9826 6777
rect 9774 6734 9826 6743
rect 9774 6457 9826 6466
rect 9774 6423 9783 6457
rect 9783 6423 9817 6457
rect 9817 6423 9826 6457
rect 9774 6414 9826 6423
rect 9774 6297 9826 6306
rect 9774 6263 9783 6297
rect 9783 6263 9817 6297
rect 9817 6263 9826 6297
rect 9774 6254 9826 6263
rect 9774 6137 9826 6146
rect 9774 6103 9783 6137
rect 9783 6103 9817 6137
rect 9817 6103 9826 6137
rect 9774 6094 9826 6103
rect 9774 5977 9826 5986
rect 9774 5943 9783 5977
rect 9783 5943 9817 5977
rect 9817 5943 9826 5977
rect 9774 5934 9826 5943
rect 9774 5817 9826 5826
rect 9774 5783 9783 5817
rect 9783 5783 9817 5817
rect 9817 5783 9826 5817
rect 9774 5774 9826 5783
rect 9774 5657 9826 5666
rect 9774 5623 9783 5657
rect 9783 5623 9817 5657
rect 9817 5623 9826 5657
rect 9774 5614 9826 5623
rect 9774 5497 9826 5506
rect 9774 5463 9783 5497
rect 9783 5463 9817 5497
rect 9817 5463 9826 5497
rect 9774 5454 9826 5463
rect 9774 5337 9826 5346
rect 9774 5303 9783 5337
rect 9783 5303 9817 5337
rect 9817 5303 9826 5337
rect 9774 5294 9826 5303
rect 9774 5177 9826 5186
rect 9774 5143 9783 5177
rect 9783 5143 9817 5177
rect 9817 5143 9826 5177
rect 9774 5134 9826 5143
rect 9774 5017 9826 5026
rect 9774 4983 9783 5017
rect 9783 4983 9817 5017
rect 9817 4983 9826 5017
rect 9774 4974 9826 4983
rect 9774 4857 9826 4866
rect 9774 4823 9783 4857
rect 9783 4823 9817 4857
rect 9817 4823 9826 4857
rect 9774 4814 9826 4823
rect 9774 4697 9826 4706
rect 9774 4663 9783 4697
rect 9783 4663 9817 4697
rect 9817 4663 9826 4697
rect 9774 4654 9826 4663
rect 9774 4537 9826 4546
rect 9774 4503 9783 4537
rect 9783 4503 9817 4537
rect 9817 4503 9826 4537
rect 9774 4494 9826 4503
rect 9774 4377 9826 4386
rect 9774 4343 9783 4377
rect 9783 4343 9817 4377
rect 9817 4343 9826 4377
rect 9774 4334 9826 4343
rect 9774 4217 9826 4226
rect 9774 4183 9783 4217
rect 9783 4183 9817 4217
rect 9817 4183 9826 4217
rect 9774 4174 9826 4183
rect 9774 4057 9826 4066
rect 9774 4023 9783 4057
rect 9783 4023 9817 4057
rect 9817 4023 9826 4057
rect 9774 4014 9826 4023
rect 9774 3897 9826 3906
rect 9774 3863 9783 3897
rect 9783 3863 9817 3897
rect 9817 3863 9826 3897
rect 9774 3854 9826 3863
rect 9774 3417 9826 3426
rect 9774 3383 9783 3417
rect 9783 3383 9817 3417
rect 9817 3383 9826 3417
rect 9774 3374 9826 3383
rect 9774 3257 9826 3266
rect 9774 3223 9783 3257
rect 9783 3223 9817 3257
rect 9817 3223 9826 3257
rect 9774 3214 9826 3223
rect 9774 3097 9826 3106
rect 9774 3063 9783 3097
rect 9783 3063 9817 3097
rect 9817 3063 9826 3097
rect 9774 3054 9826 3063
rect 9774 2937 9826 2946
rect 9774 2903 9783 2937
rect 9783 2903 9817 2937
rect 9817 2903 9826 2937
rect 9774 2894 9826 2903
rect 9774 2777 9826 2786
rect 9774 2743 9783 2777
rect 9783 2743 9817 2777
rect 9817 2743 9826 2777
rect 9774 2734 9826 2743
rect 9774 2617 9826 2626
rect 9774 2583 9783 2617
rect 9783 2583 9817 2617
rect 9817 2583 9826 2617
rect 9774 2574 9826 2583
rect 9774 2457 9826 2466
rect 9774 2423 9783 2457
rect 9783 2423 9817 2457
rect 9817 2423 9826 2457
rect 9774 2414 9826 2423
rect 9774 2297 9826 2306
rect 9774 2263 9783 2297
rect 9783 2263 9817 2297
rect 9817 2263 9826 2297
rect 9774 2254 9826 2263
rect 9774 2137 9826 2146
rect 9774 2103 9783 2137
rect 9783 2103 9817 2137
rect 9817 2103 9826 2137
rect 9774 2094 9826 2103
rect 9774 1977 9826 1986
rect 9774 1943 9783 1977
rect 9783 1943 9817 1977
rect 9817 1943 9826 1977
rect 9774 1934 9826 1943
rect 9774 1657 9826 1666
rect 9774 1623 9783 1657
rect 9783 1623 9817 1657
rect 9817 1623 9826 1657
rect 9774 1614 9826 1623
rect 9774 1497 9826 1506
rect 9774 1463 9783 1497
rect 9783 1463 9817 1497
rect 9817 1463 9826 1497
rect 9774 1454 9826 1463
rect 9774 1337 9826 1346
rect 9774 1303 9783 1337
rect 9783 1303 9817 1337
rect 9817 1303 9826 1337
rect 9774 1294 9826 1303
rect 9774 1177 9826 1186
rect 9774 1143 9783 1177
rect 9783 1143 9817 1177
rect 9817 1143 9826 1177
rect 9774 1134 9826 1143
rect 9774 1017 9826 1026
rect 9774 983 9783 1017
rect 9783 983 9817 1017
rect 9817 983 9826 1017
rect 9774 974 9826 983
rect 9774 537 9826 546
rect 9774 503 9783 537
rect 9783 503 9817 537
rect 9817 503 9826 537
rect 9774 494 9826 503
rect 9774 377 9826 386
rect 9774 343 9783 377
rect 9783 343 9817 377
rect 9817 343 9826 377
rect 9774 334 9826 343
rect 9774 217 9826 226
rect 9774 183 9783 217
rect 9783 183 9817 217
rect 9817 183 9826 217
rect 9774 174 9826 183
rect 9774 57 9826 66
rect 9774 23 9783 57
rect 9783 23 9817 57
rect 9817 23 9826 57
rect 9774 14 9826 23
rect 10094 31417 10146 31426
rect 10094 31383 10103 31417
rect 10103 31383 10137 31417
rect 10137 31383 10146 31417
rect 10094 31374 10146 31383
rect 10094 31257 10146 31266
rect 10094 31223 10103 31257
rect 10103 31223 10137 31257
rect 10137 31223 10146 31257
rect 10094 31214 10146 31223
rect 10094 31097 10146 31106
rect 10094 31063 10103 31097
rect 10103 31063 10137 31097
rect 10137 31063 10146 31097
rect 10094 31054 10146 31063
rect 10094 30937 10146 30946
rect 10094 30903 10103 30937
rect 10103 30903 10137 30937
rect 10137 30903 10146 30937
rect 10094 30894 10146 30903
rect 10094 30777 10146 30786
rect 10094 30743 10103 30777
rect 10103 30743 10137 30777
rect 10137 30743 10146 30777
rect 10094 30734 10146 30743
rect 10094 30617 10146 30626
rect 10094 30583 10103 30617
rect 10103 30583 10137 30617
rect 10137 30583 10146 30617
rect 10094 30574 10146 30583
rect 10094 30457 10146 30466
rect 10094 30423 10103 30457
rect 10103 30423 10137 30457
rect 10137 30423 10146 30457
rect 10094 30414 10146 30423
rect 10094 30297 10146 30306
rect 10094 30263 10103 30297
rect 10103 30263 10137 30297
rect 10137 30263 10146 30297
rect 10094 30254 10146 30263
rect 10094 29977 10146 29986
rect 10094 29943 10103 29977
rect 10103 29943 10137 29977
rect 10137 29943 10146 29977
rect 10094 29934 10146 29943
rect 10094 29817 10146 29826
rect 10094 29783 10103 29817
rect 10103 29783 10137 29817
rect 10137 29783 10146 29817
rect 10094 29774 10146 29783
rect 10094 29657 10146 29666
rect 10094 29623 10103 29657
rect 10103 29623 10137 29657
rect 10137 29623 10146 29657
rect 10094 29614 10146 29623
rect 10094 29497 10146 29506
rect 10094 29463 10103 29497
rect 10103 29463 10137 29497
rect 10137 29463 10146 29497
rect 10094 29454 10146 29463
rect 10094 29337 10146 29346
rect 10094 29303 10103 29337
rect 10103 29303 10137 29337
rect 10137 29303 10146 29337
rect 10094 29294 10146 29303
rect 10094 29177 10146 29186
rect 10094 29143 10103 29177
rect 10103 29143 10137 29177
rect 10137 29143 10146 29177
rect 10094 29134 10146 29143
rect 10094 29017 10146 29026
rect 10094 28983 10103 29017
rect 10103 28983 10137 29017
rect 10137 28983 10146 29017
rect 10094 28974 10146 28983
rect 10094 28857 10146 28866
rect 10094 28823 10103 28857
rect 10103 28823 10137 28857
rect 10137 28823 10146 28857
rect 10094 28814 10146 28823
rect 10094 28057 10146 28066
rect 10094 28023 10103 28057
rect 10103 28023 10137 28057
rect 10137 28023 10146 28057
rect 10094 28014 10146 28023
rect 10094 27897 10146 27906
rect 10094 27863 10103 27897
rect 10103 27863 10137 27897
rect 10137 27863 10146 27897
rect 10094 27854 10146 27863
rect 10094 27737 10146 27746
rect 10094 27703 10103 27737
rect 10103 27703 10137 27737
rect 10137 27703 10146 27737
rect 10094 27694 10146 27703
rect 10094 27577 10146 27586
rect 10094 27543 10103 27577
rect 10103 27543 10137 27577
rect 10137 27543 10146 27577
rect 10094 27534 10146 27543
rect 10094 27417 10146 27426
rect 10094 27383 10103 27417
rect 10103 27383 10137 27417
rect 10137 27383 10146 27417
rect 10094 27374 10146 27383
rect 10094 27257 10146 27266
rect 10094 27223 10103 27257
rect 10103 27223 10137 27257
rect 10137 27223 10146 27257
rect 10094 27214 10146 27223
rect 10094 27097 10146 27106
rect 10094 27063 10103 27097
rect 10103 27063 10137 27097
rect 10137 27063 10146 27097
rect 10094 27054 10146 27063
rect 10094 26937 10146 26946
rect 10094 26903 10103 26937
rect 10103 26903 10137 26937
rect 10137 26903 10146 26937
rect 10094 26894 10146 26903
rect 10094 26137 10146 26146
rect 10094 26103 10103 26137
rect 10103 26103 10137 26137
rect 10137 26103 10146 26137
rect 10094 26094 10146 26103
rect 10094 25977 10146 25986
rect 10094 25943 10103 25977
rect 10103 25943 10137 25977
rect 10137 25943 10146 25977
rect 10094 25934 10146 25943
rect 10094 25817 10146 25826
rect 10094 25783 10103 25817
rect 10103 25783 10137 25817
rect 10137 25783 10146 25817
rect 10094 25774 10146 25783
rect 10094 25657 10146 25666
rect 10094 25623 10103 25657
rect 10103 25623 10137 25657
rect 10137 25623 10146 25657
rect 10094 25614 10146 25623
rect 10094 25497 10146 25506
rect 10094 25463 10103 25497
rect 10103 25463 10137 25497
rect 10137 25463 10146 25497
rect 10094 25454 10146 25463
rect 10094 25337 10146 25346
rect 10094 25303 10103 25337
rect 10103 25303 10137 25337
rect 10137 25303 10146 25337
rect 10094 25294 10146 25303
rect 10094 25177 10146 25186
rect 10094 25143 10103 25177
rect 10103 25143 10137 25177
rect 10137 25143 10146 25177
rect 10094 25134 10146 25143
rect 10094 25017 10146 25026
rect 10094 24983 10103 25017
rect 10103 24983 10137 25017
rect 10137 24983 10146 25017
rect 10094 24974 10146 24983
rect 10094 24697 10146 24706
rect 10094 24663 10103 24697
rect 10103 24663 10137 24697
rect 10137 24663 10146 24697
rect 10094 24654 10146 24663
rect 10094 24537 10146 24546
rect 10094 24503 10103 24537
rect 10103 24503 10137 24537
rect 10137 24503 10146 24537
rect 10094 24494 10146 24503
rect 10094 24377 10146 24386
rect 10094 24343 10103 24377
rect 10103 24343 10137 24377
rect 10137 24343 10146 24377
rect 10094 24334 10146 24343
rect 10094 24217 10146 24226
rect 10094 24183 10103 24217
rect 10103 24183 10137 24217
rect 10137 24183 10146 24217
rect 10094 24174 10146 24183
rect 10094 24057 10146 24066
rect 10094 24023 10103 24057
rect 10103 24023 10137 24057
rect 10137 24023 10146 24057
rect 10094 24014 10146 24023
rect 10094 23897 10146 23906
rect 10094 23863 10103 23897
rect 10103 23863 10137 23897
rect 10137 23863 10146 23897
rect 10094 23854 10146 23863
rect 10094 23737 10146 23746
rect 10094 23703 10103 23737
rect 10103 23703 10137 23737
rect 10137 23703 10146 23737
rect 10094 23694 10146 23703
rect 10094 23577 10146 23586
rect 10094 23543 10103 23577
rect 10103 23543 10137 23577
rect 10137 23543 10146 23577
rect 10094 23534 10146 23543
rect 10094 23417 10146 23426
rect 10094 23383 10103 23417
rect 10103 23383 10137 23417
rect 10137 23383 10146 23417
rect 10094 23374 10146 23383
rect 10094 23257 10146 23266
rect 10094 23223 10103 23257
rect 10103 23223 10137 23257
rect 10137 23223 10146 23257
rect 10094 23214 10146 23223
rect 10094 23097 10146 23106
rect 10094 23063 10103 23097
rect 10103 23063 10137 23097
rect 10137 23063 10146 23097
rect 10094 23054 10146 23063
rect 10094 22937 10146 22946
rect 10094 22903 10103 22937
rect 10103 22903 10137 22937
rect 10137 22903 10146 22937
rect 10094 22894 10146 22903
rect 10094 22777 10146 22786
rect 10094 22743 10103 22777
rect 10103 22743 10137 22777
rect 10137 22743 10146 22777
rect 10094 22734 10146 22743
rect 10094 22617 10146 22626
rect 10094 22583 10103 22617
rect 10103 22583 10137 22617
rect 10137 22583 10146 22617
rect 10094 22574 10146 22583
rect 10094 22457 10146 22466
rect 10094 22423 10103 22457
rect 10103 22423 10137 22457
rect 10137 22423 10146 22457
rect 10094 22414 10146 22423
rect 10094 22297 10146 22306
rect 10094 22263 10103 22297
rect 10103 22263 10137 22297
rect 10137 22263 10146 22297
rect 10094 22254 10146 22263
rect 10094 22137 10146 22146
rect 10094 22103 10103 22137
rect 10103 22103 10137 22137
rect 10137 22103 10146 22137
rect 10094 22094 10146 22103
rect 10094 21817 10146 21826
rect 10094 21783 10103 21817
rect 10103 21783 10137 21817
rect 10137 21783 10146 21817
rect 10094 21774 10146 21783
rect 10094 21657 10146 21666
rect 10094 21623 10103 21657
rect 10103 21623 10137 21657
rect 10137 21623 10146 21657
rect 10094 21614 10146 21623
rect 10094 21497 10146 21506
rect 10094 21463 10103 21497
rect 10103 21463 10137 21497
rect 10137 21463 10146 21497
rect 10094 21454 10146 21463
rect 10094 21337 10146 21346
rect 10094 21303 10103 21337
rect 10103 21303 10137 21337
rect 10137 21303 10146 21337
rect 10094 21294 10146 21303
rect 10094 21177 10146 21186
rect 10094 21143 10103 21177
rect 10103 21143 10137 21177
rect 10137 21143 10146 21177
rect 10094 21134 10146 21143
rect 10094 21017 10146 21026
rect 10094 20983 10103 21017
rect 10103 20983 10137 21017
rect 10137 20983 10146 21017
rect 10094 20974 10146 20983
rect 10094 20857 10146 20866
rect 10094 20823 10103 20857
rect 10103 20823 10137 20857
rect 10137 20823 10146 20857
rect 10094 20814 10146 20823
rect 10094 20697 10146 20706
rect 10094 20663 10103 20697
rect 10103 20663 10137 20697
rect 10137 20663 10146 20697
rect 10094 20654 10146 20663
rect 10094 19897 10146 19906
rect 10094 19863 10103 19897
rect 10103 19863 10137 19897
rect 10137 19863 10146 19897
rect 10094 19854 10146 19863
rect 10094 19737 10146 19746
rect 10094 19703 10103 19737
rect 10103 19703 10137 19737
rect 10137 19703 10146 19737
rect 10094 19694 10146 19703
rect 10094 19577 10146 19586
rect 10094 19543 10103 19577
rect 10103 19543 10137 19577
rect 10137 19543 10146 19577
rect 10094 19534 10146 19543
rect 10094 19417 10146 19426
rect 10094 19383 10103 19417
rect 10103 19383 10137 19417
rect 10137 19383 10146 19417
rect 10094 19374 10146 19383
rect 10094 19257 10146 19266
rect 10094 19223 10103 19257
rect 10103 19223 10137 19257
rect 10137 19223 10146 19257
rect 10094 19214 10146 19223
rect 10094 19097 10146 19106
rect 10094 19063 10103 19097
rect 10103 19063 10137 19097
rect 10137 19063 10146 19097
rect 10094 19054 10146 19063
rect 10094 18937 10146 18946
rect 10094 18903 10103 18937
rect 10103 18903 10137 18937
rect 10137 18903 10146 18937
rect 10094 18894 10146 18903
rect 10094 18777 10146 18786
rect 10094 18743 10103 18777
rect 10103 18743 10137 18777
rect 10137 18743 10146 18777
rect 10094 18734 10146 18743
rect 10094 17977 10146 17986
rect 10094 17943 10103 17977
rect 10103 17943 10137 17977
rect 10137 17943 10146 17977
rect 10094 17934 10146 17943
rect 10094 17817 10146 17826
rect 10094 17783 10103 17817
rect 10103 17783 10137 17817
rect 10137 17783 10146 17817
rect 10094 17774 10146 17783
rect 10094 17657 10146 17666
rect 10094 17623 10103 17657
rect 10103 17623 10137 17657
rect 10137 17623 10146 17657
rect 10094 17614 10146 17623
rect 10094 17497 10146 17506
rect 10094 17463 10103 17497
rect 10103 17463 10137 17497
rect 10137 17463 10146 17497
rect 10094 17454 10146 17463
rect 10094 17337 10146 17346
rect 10094 17303 10103 17337
rect 10103 17303 10137 17337
rect 10137 17303 10146 17337
rect 10094 17294 10146 17303
rect 10094 17177 10146 17186
rect 10094 17143 10103 17177
rect 10103 17143 10137 17177
rect 10137 17143 10146 17177
rect 10094 17134 10146 17143
rect 10094 17017 10146 17026
rect 10094 16983 10103 17017
rect 10103 16983 10137 17017
rect 10137 16983 10146 17017
rect 10094 16974 10146 16983
rect 10094 16857 10146 16866
rect 10094 16823 10103 16857
rect 10103 16823 10137 16857
rect 10137 16823 10146 16857
rect 10094 16814 10146 16823
rect 10094 16537 10146 16546
rect 10094 16503 10103 16537
rect 10103 16503 10137 16537
rect 10137 16503 10146 16537
rect 10094 16494 10146 16503
rect 10094 16377 10146 16386
rect 10094 16343 10103 16377
rect 10103 16343 10137 16377
rect 10137 16343 10146 16377
rect 10094 16334 10146 16343
rect 10094 16217 10146 16226
rect 10094 16183 10103 16217
rect 10103 16183 10137 16217
rect 10137 16183 10146 16217
rect 10094 16174 10146 16183
rect 10094 16057 10146 16066
rect 10094 16023 10103 16057
rect 10103 16023 10137 16057
rect 10137 16023 10146 16057
rect 10094 16014 10146 16023
rect 10094 15897 10146 15906
rect 10094 15863 10103 15897
rect 10103 15863 10137 15897
rect 10137 15863 10146 15897
rect 10094 15854 10146 15863
rect 10094 15737 10146 15746
rect 10094 15703 10103 15737
rect 10103 15703 10137 15737
rect 10137 15703 10146 15737
rect 10094 15694 10146 15703
rect 10094 15577 10146 15586
rect 10094 15543 10103 15577
rect 10103 15543 10137 15577
rect 10137 15543 10146 15577
rect 10094 15534 10146 15543
rect 10094 15417 10146 15426
rect 10094 15383 10103 15417
rect 10103 15383 10137 15417
rect 10137 15383 10146 15417
rect 10094 15374 10146 15383
rect 10094 15257 10146 15266
rect 10094 15223 10103 15257
rect 10103 15223 10137 15257
rect 10137 15223 10146 15257
rect 10094 15214 10146 15223
rect 10094 15097 10146 15106
rect 10094 15063 10103 15097
rect 10103 15063 10137 15097
rect 10137 15063 10146 15097
rect 10094 15054 10146 15063
rect 10094 14937 10146 14946
rect 10094 14903 10103 14937
rect 10103 14903 10137 14937
rect 10137 14903 10146 14937
rect 10094 14894 10146 14903
rect 10094 14777 10146 14786
rect 10094 14743 10103 14777
rect 10103 14743 10137 14777
rect 10137 14743 10146 14777
rect 10094 14734 10146 14743
rect 10094 14617 10146 14626
rect 10094 14583 10103 14617
rect 10103 14583 10137 14617
rect 10137 14583 10146 14617
rect 10094 14574 10146 14583
rect 10094 14457 10146 14466
rect 10094 14423 10103 14457
rect 10103 14423 10137 14457
rect 10137 14423 10146 14457
rect 10094 14414 10146 14423
rect 10094 14297 10146 14306
rect 10094 14263 10103 14297
rect 10103 14263 10137 14297
rect 10137 14263 10146 14297
rect 10094 14254 10146 14263
rect 10094 14137 10146 14146
rect 10094 14103 10103 14137
rect 10103 14103 10137 14137
rect 10137 14103 10146 14137
rect 10094 14094 10146 14103
rect 10094 13977 10146 13986
rect 10094 13943 10103 13977
rect 10103 13943 10137 13977
rect 10137 13943 10146 13977
rect 10094 13934 10146 13943
rect 10094 13657 10146 13666
rect 10094 13623 10103 13657
rect 10103 13623 10137 13657
rect 10137 13623 10146 13657
rect 10094 13614 10146 13623
rect 10094 13497 10146 13506
rect 10094 13463 10103 13497
rect 10103 13463 10137 13497
rect 10137 13463 10146 13497
rect 10094 13454 10146 13463
rect 10094 13337 10146 13346
rect 10094 13303 10103 13337
rect 10103 13303 10137 13337
rect 10137 13303 10146 13337
rect 10094 13294 10146 13303
rect 10094 13177 10146 13186
rect 10094 13143 10103 13177
rect 10103 13143 10137 13177
rect 10137 13143 10146 13177
rect 10094 13134 10146 13143
rect 10094 13017 10146 13026
rect 10094 12983 10103 13017
rect 10103 12983 10137 13017
rect 10137 12983 10146 13017
rect 10094 12974 10146 12983
rect 10094 12857 10146 12866
rect 10094 12823 10103 12857
rect 10103 12823 10137 12857
rect 10137 12823 10146 12857
rect 10094 12814 10146 12823
rect 10094 12697 10146 12706
rect 10094 12663 10103 12697
rect 10103 12663 10137 12697
rect 10137 12663 10146 12697
rect 10094 12654 10146 12663
rect 10094 12537 10146 12546
rect 10094 12503 10103 12537
rect 10103 12503 10137 12537
rect 10137 12503 10146 12537
rect 10094 12494 10146 12503
rect 10094 11737 10146 11746
rect 10094 11703 10103 11737
rect 10103 11703 10137 11737
rect 10137 11703 10146 11737
rect 10094 11694 10146 11703
rect 10094 11577 10146 11586
rect 10094 11543 10103 11577
rect 10103 11543 10137 11577
rect 10137 11543 10146 11577
rect 10094 11534 10146 11543
rect 10094 11417 10146 11426
rect 10094 11383 10103 11417
rect 10103 11383 10137 11417
rect 10137 11383 10146 11417
rect 10094 11374 10146 11383
rect 10094 11257 10146 11266
rect 10094 11223 10103 11257
rect 10103 11223 10137 11257
rect 10137 11223 10146 11257
rect 10094 11214 10146 11223
rect 10094 11097 10146 11106
rect 10094 11063 10103 11097
rect 10103 11063 10137 11097
rect 10137 11063 10146 11097
rect 10094 11054 10146 11063
rect 10094 10937 10146 10946
rect 10094 10903 10103 10937
rect 10103 10903 10137 10937
rect 10137 10903 10146 10937
rect 10094 10894 10146 10903
rect 10094 10777 10146 10786
rect 10094 10743 10103 10777
rect 10103 10743 10137 10777
rect 10137 10743 10146 10777
rect 10094 10734 10146 10743
rect 10094 10617 10146 10626
rect 10094 10583 10103 10617
rect 10103 10583 10137 10617
rect 10137 10583 10146 10617
rect 10094 10574 10146 10583
rect 10094 10457 10146 10466
rect 10094 10423 10103 10457
rect 10103 10423 10137 10457
rect 10137 10423 10146 10457
rect 10094 10414 10146 10423
rect 10094 10297 10146 10306
rect 10094 10263 10103 10297
rect 10103 10263 10137 10297
rect 10137 10263 10146 10297
rect 10094 10254 10146 10263
rect 10094 10137 10146 10146
rect 10094 10103 10103 10137
rect 10103 10103 10137 10137
rect 10137 10103 10146 10137
rect 10094 10094 10146 10103
rect 10094 9977 10146 9986
rect 10094 9943 10103 9977
rect 10103 9943 10137 9977
rect 10137 9943 10146 9977
rect 10094 9934 10146 9943
rect 10094 9817 10146 9826
rect 10094 9783 10103 9817
rect 10103 9783 10137 9817
rect 10137 9783 10146 9817
rect 10094 9774 10146 9783
rect 10094 9497 10146 9506
rect 10094 9463 10103 9497
rect 10103 9463 10137 9497
rect 10137 9463 10146 9497
rect 10094 9454 10146 9463
rect 10094 9337 10146 9346
rect 10094 9303 10103 9337
rect 10103 9303 10137 9337
rect 10137 9303 10146 9337
rect 10094 9294 10146 9303
rect 10094 9017 10146 9026
rect 10094 8983 10103 9017
rect 10103 8983 10137 9017
rect 10137 8983 10146 9017
rect 10094 8974 10146 8983
rect 10094 8857 10146 8866
rect 10094 8823 10103 8857
rect 10103 8823 10137 8857
rect 10137 8823 10146 8857
rect 10094 8814 10146 8823
rect 10094 8697 10146 8706
rect 10094 8663 10103 8697
rect 10103 8663 10137 8697
rect 10137 8663 10146 8697
rect 10094 8654 10146 8663
rect 10094 8537 10146 8546
rect 10094 8503 10103 8537
rect 10103 8503 10137 8537
rect 10137 8503 10146 8537
rect 10094 8494 10146 8503
rect 10094 8377 10146 8386
rect 10094 8343 10103 8377
rect 10103 8343 10137 8377
rect 10137 8343 10146 8377
rect 10094 8334 10146 8343
rect 10094 8217 10146 8226
rect 10094 8183 10103 8217
rect 10103 8183 10137 8217
rect 10137 8183 10146 8217
rect 10094 8174 10146 8183
rect 10094 8057 10146 8066
rect 10094 8023 10103 8057
rect 10103 8023 10137 8057
rect 10137 8023 10146 8057
rect 10094 8014 10146 8023
rect 10094 7897 10146 7906
rect 10094 7863 10103 7897
rect 10103 7863 10137 7897
rect 10137 7863 10146 7897
rect 10094 7854 10146 7863
rect 10094 7737 10146 7746
rect 10094 7703 10103 7737
rect 10103 7703 10137 7737
rect 10137 7703 10146 7737
rect 10094 7694 10146 7703
rect 10094 7417 10146 7426
rect 10094 7383 10103 7417
rect 10103 7383 10137 7417
rect 10137 7383 10146 7417
rect 10094 7374 10146 7383
rect 10094 7257 10146 7266
rect 10094 7223 10103 7257
rect 10103 7223 10137 7257
rect 10137 7223 10146 7257
rect 10094 7214 10146 7223
rect 10094 6937 10146 6946
rect 10094 6903 10103 6937
rect 10103 6903 10137 6937
rect 10137 6903 10146 6937
rect 10094 6894 10146 6903
rect 10094 6777 10146 6786
rect 10094 6743 10103 6777
rect 10103 6743 10137 6777
rect 10137 6743 10146 6777
rect 10094 6734 10146 6743
rect 10094 6457 10146 6466
rect 10094 6423 10103 6457
rect 10103 6423 10137 6457
rect 10137 6423 10146 6457
rect 10094 6414 10146 6423
rect 10094 6297 10146 6306
rect 10094 6263 10103 6297
rect 10103 6263 10137 6297
rect 10137 6263 10146 6297
rect 10094 6254 10146 6263
rect 10094 6137 10146 6146
rect 10094 6103 10103 6137
rect 10103 6103 10137 6137
rect 10137 6103 10146 6137
rect 10094 6094 10146 6103
rect 10094 5977 10146 5986
rect 10094 5943 10103 5977
rect 10103 5943 10137 5977
rect 10137 5943 10146 5977
rect 10094 5934 10146 5943
rect 10094 5817 10146 5826
rect 10094 5783 10103 5817
rect 10103 5783 10137 5817
rect 10137 5783 10146 5817
rect 10094 5774 10146 5783
rect 10094 5657 10146 5666
rect 10094 5623 10103 5657
rect 10103 5623 10137 5657
rect 10137 5623 10146 5657
rect 10094 5614 10146 5623
rect 10094 5497 10146 5506
rect 10094 5463 10103 5497
rect 10103 5463 10137 5497
rect 10137 5463 10146 5497
rect 10094 5454 10146 5463
rect 10094 5337 10146 5346
rect 10094 5303 10103 5337
rect 10103 5303 10137 5337
rect 10137 5303 10146 5337
rect 10094 5294 10146 5303
rect 10094 5177 10146 5186
rect 10094 5143 10103 5177
rect 10103 5143 10137 5177
rect 10137 5143 10146 5177
rect 10094 5134 10146 5143
rect 10094 5017 10146 5026
rect 10094 4983 10103 5017
rect 10103 4983 10137 5017
rect 10137 4983 10146 5017
rect 10094 4974 10146 4983
rect 10094 4857 10146 4866
rect 10094 4823 10103 4857
rect 10103 4823 10137 4857
rect 10137 4823 10146 4857
rect 10094 4814 10146 4823
rect 10094 4697 10146 4706
rect 10094 4663 10103 4697
rect 10103 4663 10137 4697
rect 10137 4663 10146 4697
rect 10094 4654 10146 4663
rect 10094 4537 10146 4546
rect 10094 4503 10103 4537
rect 10103 4503 10137 4537
rect 10137 4503 10146 4537
rect 10094 4494 10146 4503
rect 10094 4377 10146 4386
rect 10094 4343 10103 4377
rect 10103 4343 10137 4377
rect 10137 4343 10146 4377
rect 10094 4334 10146 4343
rect 10094 4217 10146 4226
rect 10094 4183 10103 4217
rect 10103 4183 10137 4217
rect 10137 4183 10146 4217
rect 10094 4174 10146 4183
rect 10094 4057 10146 4066
rect 10094 4023 10103 4057
rect 10103 4023 10137 4057
rect 10137 4023 10146 4057
rect 10094 4014 10146 4023
rect 10094 3897 10146 3906
rect 10094 3863 10103 3897
rect 10103 3863 10137 3897
rect 10137 3863 10146 3897
rect 10094 3854 10146 3863
rect 10094 3417 10146 3426
rect 10094 3383 10103 3417
rect 10103 3383 10137 3417
rect 10137 3383 10146 3417
rect 10094 3374 10146 3383
rect 10094 3257 10146 3266
rect 10094 3223 10103 3257
rect 10103 3223 10137 3257
rect 10137 3223 10146 3257
rect 10094 3214 10146 3223
rect 10094 3097 10146 3106
rect 10094 3063 10103 3097
rect 10103 3063 10137 3097
rect 10137 3063 10146 3097
rect 10094 3054 10146 3063
rect 10094 2937 10146 2946
rect 10094 2903 10103 2937
rect 10103 2903 10137 2937
rect 10137 2903 10146 2937
rect 10094 2894 10146 2903
rect 10094 2777 10146 2786
rect 10094 2743 10103 2777
rect 10103 2743 10137 2777
rect 10137 2743 10146 2777
rect 10094 2734 10146 2743
rect 10094 2617 10146 2626
rect 10094 2583 10103 2617
rect 10103 2583 10137 2617
rect 10137 2583 10146 2617
rect 10094 2574 10146 2583
rect 10094 2457 10146 2466
rect 10094 2423 10103 2457
rect 10103 2423 10137 2457
rect 10137 2423 10146 2457
rect 10094 2414 10146 2423
rect 10094 2297 10146 2306
rect 10094 2263 10103 2297
rect 10103 2263 10137 2297
rect 10137 2263 10146 2297
rect 10094 2254 10146 2263
rect 10094 2137 10146 2146
rect 10094 2103 10103 2137
rect 10103 2103 10137 2137
rect 10137 2103 10146 2137
rect 10094 2094 10146 2103
rect 10094 1977 10146 1986
rect 10094 1943 10103 1977
rect 10103 1943 10137 1977
rect 10137 1943 10146 1977
rect 10094 1934 10146 1943
rect 10094 1657 10146 1666
rect 10094 1623 10103 1657
rect 10103 1623 10137 1657
rect 10137 1623 10146 1657
rect 10094 1614 10146 1623
rect 10094 1497 10146 1506
rect 10094 1463 10103 1497
rect 10103 1463 10137 1497
rect 10137 1463 10146 1497
rect 10094 1454 10146 1463
rect 10094 1337 10146 1346
rect 10094 1303 10103 1337
rect 10103 1303 10137 1337
rect 10137 1303 10146 1337
rect 10094 1294 10146 1303
rect 10094 1177 10146 1186
rect 10094 1143 10103 1177
rect 10103 1143 10137 1177
rect 10137 1143 10146 1177
rect 10094 1134 10146 1143
rect 10094 1017 10146 1026
rect 10094 983 10103 1017
rect 10103 983 10137 1017
rect 10137 983 10146 1017
rect 10094 974 10146 983
rect 10094 537 10146 546
rect 10094 503 10103 537
rect 10103 503 10137 537
rect 10137 503 10146 537
rect 10094 494 10146 503
rect 10094 377 10146 386
rect 10094 343 10103 377
rect 10103 343 10137 377
rect 10137 343 10146 377
rect 10094 334 10146 343
rect 10094 217 10146 226
rect 10094 183 10103 217
rect 10103 183 10137 217
rect 10137 183 10146 217
rect 10094 174 10146 183
rect 10094 57 10146 66
rect 10094 23 10103 57
rect 10103 23 10137 57
rect 10137 23 10146 57
rect 10094 14 10146 23
rect 10414 31417 10466 31426
rect 10414 31383 10423 31417
rect 10423 31383 10457 31417
rect 10457 31383 10466 31417
rect 10414 31374 10466 31383
rect 10414 31257 10466 31266
rect 10414 31223 10423 31257
rect 10423 31223 10457 31257
rect 10457 31223 10466 31257
rect 10414 31214 10466 31223
rect 10414 31097 10466 31106
rect 10414 31063 10423 31097
rect 10423 31063 10457 31097
rect 10457 31063 10466 31097
rect 10414 31054 10466 31063
rect 10414 30937 10466 30946
rect 10414 30903 10423 30937
rect 10423 30903 10457 30937
rect 10457 30903 10466 30937
rect 10414 30894 10466 30903
rect 10414 30777 10466 30786
rect 10414 30743 10423 30777
rect 10423 30743 10457 30777
rect 10457 30743 10466 30777
rect 10414 30734 10466 30743
rect 10414 30617 10466 30626
rect 10414 30583 10423 30617
rect 10423 30583 10457 30617
rect 10457 30583 10466 30617
rect 10414 30574 10466 30583
rect 10414 30457 10466 30466
rect 10414 30423 10423 30457
rect 10423 30423 10457 30457
rect 10457 30423 10466 30457
rect 10414 30414 10466 30423
rect 10414 30297 10466 30306
rect 10414 30263 10423 30297
rect 10423 30263 10457 30297
rect 10457 30263 10466 30297
rect 10414 30254 10466 30263
rect 10414 29977 10466 29986
rect 10414 29943 10423 29977
rect 10423 29943 10457 29977
rect 10457 29943 10466 29977
rect 10414 29934 10466 29943
rect 10414 29817 10466 29826
rect 10414 29783 10423 29817
rect 10423 29783 10457 29817
rect 10457 29783 10466 29817
rect 10414 29774 10466 29783
rect 10414 29657 10466 29666
rect 10414 29623 10423 29657
rect 10423 29623 10457 29657
rect 10457 29623 10466 29657
rect 10414 29614 10466 29623
rect 10414 29497 10466 29506
rect 10414 29463 10423 29497
rect 10423 29463 10457 29497
rect 10457 29463 10466 29497
rect 10414 29454 10466 29463
rect 10414 29337 10466 29346
rect 10414 29303 10423 29337
rect 10423 29303 10457 29337
rect 10457 29303 10466 29337
rect 10414 29294 10466 29303
rect 10414 29177 10466 29186
rect 10414 29143 10423 29177
rect 10423 29143 10457 29177
rect 10457 29143 10466 29177
rect 10414 29134 10466 29143
rect 10414 29017 10466 29026
rect 10414 28983 10423 29017
rect 10423 28983 10457 29017
rect 10457 28983 10466 29017
rect 10414 28974 10466 28983
rect 10414 28857 10466 28866
rect 10414 28823 10423 28857
rect 10423 28823 10457 28857
rect 10457 28823 10466 28857
rect 10414 28814 10466 28823
rect 10414 28057 10466 28066
rect 10414 28023 10423 28057
rect 10423 28023 10457 28057
rect 10457 28023 10466 28057
rect 10414 28014 10466 28023
rect 10414 27897 10466 27906
rect 10414 27863 10423 27897
rect 10423 27863 10457 27897
rect 10457 27863 10466 27897
rect 10414 27854 10466 27863
rect 10414 27737 10466 27746
rect 10414 27703 10423 27737
rect 10423 27703 10457 27737
rect 10457 27703 10466 27737
rect 10414 27694 10466 27703
rect 10414 27577 10466 27586
rect 10414 27543 10423 27577
rect 10423 27543 10457 27577
rect 10457 27543 10466 27577
rect 10414 27534 10466 27543
rect 10414 27417 10466 27426
rect 10414 27383 10423 27417
rect 10423 27383 10457 27417
rect 10457 27383 10466 27417
rect 10414 27374 10466 27383
rect 10414 27257 10466 27266
rect 10414 27223 10423 27257
rect 10423 27223 10457 27257
rect 10457 27223 10466 27257
rect 10414 27214 10466 27223
rect 10414 27097 10466 27106
rect 10414 27063 10423 27097
rect 10423 27063 10457 27097
rect 10457 27063 10466 27097
rect 10414 27054 10466 27063
rect 10414 26937 10466 26946
rect 10414 26903 10423 26937
rect 10423 26903 10457 26937
rect 10457 26903 10466 26937
rect 10414 26894 10466 26903
rect 10414 26137 10466 26146
rect 10414 26103 10423 26137
rect 10423 26103 10457 26137
rect 10457 26103 10466 26137
rect 10414 26094 10466 26103
rect 10414 25977 10466 25986
rect 10414 25943 10423 25977
rect 10423 25943 10457 25977
rect 10457 25943 10466 25977
rect 10414 25934 10466 25943
rect 10414 25817 10466 25826
rect 10414 25783 10423 25817
rect 10423 25783 10457 25817
rect 10457 25783 10466 25817
rect 10414 25774 10466 25783
rect 10414 25657 10466 25666
rect 10414 25623 10423 25657
rect 10423 25623 10457 25657
rect 10457 25623 10466 25657
rect 10414 25614 10466 25623
rect 10414 25497 10466 25506
rect 10414 25463 10423 25497
rect 10423 25463 10457 25497
rect 10457 25463 10466 25497
rect 10414 25454 10466 25463
rect 10414 25337 10466 25346
rect 10414 25303 10423 25337
rect 10423 25303 10457 25337
rect 10457 25303 10466 25337
rect 10414 25294 10466 25303
rect 10414 25177 10466 25186
rect 10414 25143 10423 25177
rect 10423 25143 10457 25177
rect 10457 25143 10466 25177
rect 10414 25134 10466 25143
rect 10414 25017 10466 25026
rect 10414 24983 10423 25017
rect 10423 24983 10457 25017
rect 10457 24983 10466 25017
rect 10414 24974 10466 24983
rect 10414 24697 10466 24706
rect 10414 24663 10423 24697
rect 10423 24663 10457 24697
rect 10457 24663 10466 24697
rect 10414 24654 10466 24663
rect 10414 24537 10466 24546
rect 10414 24503 10423 24537
rect 10423 24503 10457 24537
rect 10457 24503 10466 24537
rect 10414 24494 10466 24503
rect 10414 24377 10466 24386
rect 10414 24343 10423 24377
rect 10423 24343 10457 24377
rect 10457 24343 10466 24377
rect 10414 24334 10466 24343
rect 10414 24217 10466 24226
rect 10414 24183 10423 24217
rect 10423 24183 10457 24217
rect 10457 24183 10466 24217
rect 10414 24174 10466 24183
rect 10414 24057 10466 24066
rect 10414 24023 10423 24057
rect 10423 24023 10457 24057
rect 10457 24023 10466 24057
rect 10414 24014 10466 24023
rect 10414 23897 10466 23906
rect 10414 23863 10423 23897
rect 10423 23863 10457 23897
rect 10457 23863 10466 23897
rect 10414 23854 10466 23863
rect 10414 23737 10466 23746
rect 10414 23703 10423 23737
rect 10423 23703 10457 23737
rect 10457 23703 10466 23737
rect 10414 23694 10466 23703
rect 10414 23577 10466 23586
rect 10414 23543 10423 23577
rect 10423 23543 10457 23577
rect 10457 23543 10466 23577
rect 10414 23534 10466 23543
rect 10414 23417 10466 23426
rect 10414 23383 10423 23417
rect 10423 23383 10457 23417
rect 10457 23383 10466 23417
rect 10414 23374 10466 23383
rect 10414 23257 10466 23266
rect 10414 23223 10423 23257
rect 10423 23223 10457 23257
rect 10457 23223 10466 23257
rect 10414 23214 10466 23223
rect 10414 23097 10466 23106
rect 10414 23063 10423 23097
rect 10423 23063 10457 23097
rect 10457 23063 10466 23097
rect 10414 23054 10466 23063
rect 10414 22937 10466 22946
rect 10414 22903 10423 22937
rect 10423 22903 10457 22937
rect 10457 22903 10466 22937
rect 10414 22894 10466 22903
rect 10414 22777 10466 22786
rect 10414 22743 10423 22777
rect 10423 22743 10457 22777
rect 10457 22743 10466 22777
rect 10414 22734 10466 22743
rect 10414 22617 10466 22626
rect 10414 22583 10423 22617
rect 10423 22583 10457 22617
rect 10457 22583 10466 22617
rect 10414 22574 10466 22583
rect 10414 22457 10466 22466
rect 10414 22423 10423 22457
rect 10423 22423 10457 22457
rect 10457 22423 10466 22457
rect 10414 22414 10466 22423
rect 10414 22297 10466 22306
rect 10414 22263 10423 22297
rect 10423 22263 10457 22297
rect 10457 22263 10466 22297
rect 10414 22254 10466 22263
rect 10414 22137 10466 22146
rect 10414 22103 10423 22137
rect 10423 22103 10457 22137
rect 10457 22103 10466 22137
rect 10414 22094 10466 22103
rect 10414 21817 10466 21826
rect 10414 21783 10423 21817
rect 10423 21783 10457 21817
rect 10457 21783 10466 21817
rect 10414 21774 10466 21783
rect 10414 21657 10466 21666
rect 10414 21623 10423 21657
rect 10423 21623 10457 21657
rect 10457 21623 10466 21657
rect 10414 21614 10466 21623
rect 10414 21497 10466 21506
rect 10414 21463 10423 21497
rect 10423 21463 10457 21497
rect 10457 21463 10466 21497
rect 10414 21454 10466 21463
rect 10414 21337 10466 21346
rect 10414 21303 10423 21337
rect 10423 21303 10457 21337
rect 10457 21303 10466 21337
rect 10414 21294 10466 21303
rect 10414 21177 10466 21186
rect 10414 21143 10423 21177
rect 10423 21143 10457 21177
rect 10457 21143 10466 21177
rect 10414 21134 10466 21143
rect 10414 21017 10466 21026
rect 10414 20983 10423 21017
rect 10423 20983 10457 21017
rect 10457 20983 10466 21017
rect 10414 20974 10466 20983
rect 10414 20857 10466 20866
rect 10414 20823 10423 20857
rect 10423 20823 10457 20857
rect 10457 20823 10466 20857
rect 10414 20814 10466 20823
rect 10414 20697 10466 20706
rect 10414 20663 10423 20697
rect 10423 20663 10457 20697
rect 10457 20663 10466 20697
rect 10414 20654 10466 20663
rect 10414 19897 10466 19906
rect 10414 19863 10423 19897
rect 10423 19863 10457 19897
rect 10457 19863 10466 19897
rect 10414 19854 10466 19863
rect 10414 19737 10466 19746
rect 10414 19703 10423 19737
rect 10423 19703 10457 19737
rect 10457 19703 10466 19737
rect 10414 19694 10466 19703
rect 10414 19577 10466 19586
rect 10414 19543 10423 19577
rect 10423 19543 10457 19577
rect 10457 19543 10466 19577
rect 10414 19534 10466 19543
rect 10414 19417 10466 19426
rect 10414 19383 10423 19417
rect 10423 19383 10457 19417
rect 10457 19383 10466 19417
rect 10414 19374 10466 19383
rect 10414 19257 10466 19266
rect 10414 19223 10423 19257
rect 10423 19223 10457 19257
rect 10457 19223 10466 19257
rect 10414 19214 10466 19223
rect 10414 19097 10466 19106
rect 10414 19063 10423 19097
rect 10423 19063 10457 19097
rect 10457 19063 10466 19097
rect 10414 19054 10466 19063
rect 10414 18937 10466 18946
rect 10414 18903 10423 18937
rect 10423 18903 10457 18937
rect 10457 18903 10466 18937
rect 10414 18894 10466 18903
rect 10414 18777 10466 18786
rect 10414 18743 10423 18777
rect 10423 18743 10457 18777
rect 10457 18743 10466 18777
rect 10414 18734 10466 18743
rect 10414 17977 10466 17986
rect 10414 17943 10423 17977
rect 10423 17943 10457 17977
rect 10457 17943 10466 17977
rect 10414 17934 10466 17943
rect 10414 17817 10466 17826
rect 10414 17783 10423 17817
rect 10423 17783 10457 17817
rect 10457 17783 10466 17817
rect 10414 17774 10466 17783
rect 10414 17657 10466 17666
rect 10414 17623 10423 17657
rect 10423 17623 10457 17657
rect 10457 17623 10466 17657
rect 10414 17614 10466 17623
rect 10414 17497 10466 17506
rect 10414 17463 10423 17497
rect 10423 17463 10457 17497
rect 10457 17463 10466 17497
rect 10414 17454 10466 17463
rect 10414 17337 10466 17346
rect 10414 17303 10423 17337
rect 10423 17303 10457 17337
rect 10457 17303 10466 17337
rect 10414 17294 10466 17303
rect 10414 17177 10466 17186
rect 10414 17143 10423 17177
rect 10423 17143 10457 17177
rect 10457 17143 10466 17177
rect 10414 17134 10466 17143
rect 10414 17017 10466 17026
rect 10414 16983 10423 17017
rect 10423 16983 10457 17017
rect 10457 16983 10466 17017
rect 10414 16974 10466 16983
rect 10414 16857 10466 16866
rect 10414 16823 10423 16857
rect 10423 16823 10457 16857
rect 10457 16823 10466 16857
rect 10414 16814 10466 16823
rect 10414 16537 10466 16546
rect 10414 16503 10423 16537
rect 10423 16503 10457 16537
rect 10457 16503 10466 16537
rect 10414 16494 10466 16503
rect 10414 16377 10466 16386
rect 10414 16343 10423 16377
rect 10423 16343 10457 16377
rect 10457 16343 10466 16377
rect 10414 16334 10466 16343
rect 10414 16217 10466 16226
rect 10414 16183 10423 16217
rect 10423 16183 10457 16217
rect 10457 16183 10466 16217
rect 10414 16174 10466 16183
rect 10414 16057 10466 16066
rect 10414 16023 10423 16057
rect 10423 16023 10457 16057
rect 10457 16023 10466 16057
rect 10414 16014 10466 16023
rect 10414 15897 10466 15906
rect 10414 15863 10423 15897
rect 10423 15863 10457 15897
rect 10457 15863 10466 15897
rect 10414 15854 10466 15863
rect 10414 15737 10466 15746
rect 10414 15703 10423 15737
rect 10423 15703 10457 15737
rect 10457 15703 10466 15737
rect 10414 15694 10466 15703
rect 10414 15577 10466 15586
rect 10414 15543 10423 15577
rect 10423 15543 10457 15577
rect 10457 15543 10466 15577
rect 10414 15534 10466 15543
rect 10414 15417 10466 15426
rect 10414 15383 10423 15417
rect 10423 15383 10457 15417
rect 10457 15383 10466 15417
rect 10414 15374 10466 15383
rect 10414 15257 10466 15266
rect 10414 15223 10423 15257
rect 10423 15223 10457 15257
rect 10457 15223 10466 15257
rect 10414 15214 10466 15223
rect 10414 15097 10466 15106
rect 10414 15063 10423 15097
rect 10423 15063 10457 15097
rect 10457 15063 10466 15097
rect 10414 15054 10466 15063
rect 10414 14937 10466 14946
rect 10414 14903 10423 14937
rect 10423 14903 10457 14937
rect 10457 14903 10466 14937
rect 10414 14894 10466 14903
rect 10414 14777 10466 14786
rect 10414 14743 10423 14777
rect 10423 14743 10457 14777
rect 10457 14743 10466 14777
rect 10414 14734 10466 14743
rect 10414 14617 10466 14626
rect 10414 14583 10423 14617
rect 10423 14583 10457 14617
rect 10457 14583 10466 14617
rect 10414 14574 10466 14583
rect 10414 14457 10466 14466
rect 10414 14423 10423 14457
rect 10423 14423 10457 14457
rect 10457 14423 10466 14457
rect 10414 14414 10466 14423
rect 10414 14297 10466 14306
rect 10414 14263 10423 14297
rect 10423 14263 10457 14297
rect 10457 14263 10466 14297
rect 10414 14254 10466 14263
rect 10414 14137 10466 14146
rect 10414 14103 10423 14137
rect 10423 14103 10457 14137
rect 10457 14103 10466 14137
rect 10414 14094 10466 14103
rect 10414 13977 10466 13986
rect 10414 13943 10423 13977
rect 10423 13943 10457 13977
rect 10457 13943 10466 13977
rect 10414 13934 10466 13943
rect 10414 13657 10466 13666
rect 10414 13623 10423 13657
rect 10423 13623 10457 13657
rect 10457 13623 10466 13657
rect 10414 13614 10466 13623
rect 10414 13497 10466 13506
rect 10414 13463 10423 13497
rect 10423 13463 10457 13497
rect 10457 13463 10466 13497
rect 10414 13454 10466 13463
rect 10414 13337 10466 13346
rect 10414 13303 10423 13337
rect 10423 13303 10457 13337
rect 10457 13303 10466 13337
rect 10414 13294 10466 13303
rect 10414 13177 10466 13186
rect 10414 13143 10423 13177
rect 10423 13143 10457 13177
rect 10457 13143 10466 13177
rect 10414 13134 10466 13143
rect 10414 13017 10466 13026
rect 10414 12983 10423 13017
rect 10423 12983 10457 13017
rect 10457 12983 10466 13017
rect 10414 12974 10466 12983
rect 10414 12857 10466 12866
rect 10414 12823 10423 12857
rect 10423 12823 10457 12857
rect 10457 12823 10466 12857
rect 10414 12814 10466 12823
rect 10414 12697 10466 12706
rect 10414 12663 10423 12697
rect 10423 12663 10457 12697
rect 10457 12663 10466 12697
rect 10414 12654 10466 12663
rect 10414 12537 10466 12546
rect 10414 12503 10423 12537
rect 10423 12503 10457 12537
rect 10457 12503 10466 12537
rect 10414 12494 10466 12503
rect 10414 11737 10466 11746
rect 10414 11703 10423 11737
rect 10423 11703 10457 11737
rect 10457 11703 10466 11737
rect 10414 11694 10466 11703
rect 10414 11577 10466 11586
rect 10414 11543 10423 11577
rect 10423 11543 10457 11577
rect 10457 11543 10466 11577
rect 10414 11534 10466 11543
rect 10414 11417 10466 11426
rect 10414 11383 10423 11417
rect 10423 11383 10457 11417
rect 10457 11383 10466 11417
rect 10414 11374 10466 11383
rect 10414 11257 10466 11266
rect 10414 11223 10423 11257
rect 10423 11223 10457 11257
rect 10457 11223 10466 11257
rect 10414 11214 10466 11223
rect 10414 11097 10466 11106
rect 10414 11063 10423 11097
rect 10423 11063 10457 11097
rect 10457 11063 10466 11097
rect 10414 11054 10466 11063
rect 10414 10937 10466 10946
rect 10414 10903 10423 10937
rect 10423 10903 10457 10937
rect 10457 10903 10466 10937
rect 10414 10894 10466 10903
rect 10414 10777 10466 10786
rect 10414 10743 10423 10777
rect 10423 10743 10457 10777
rect 10457 10743 10466 10777
rect 10414 10734 10466 10743
rect 10414 10617 10466 10626
rect 10414 10583 10423 10617
rect 10423 10583 10457 10617
rect 10457 10583 10466 10617
rect 10414 10574 10466 10583
rect 10414 10457 10466 10466
rect 10414 10423 10423 10457
rect 10423 10423 10457 10457
rect 10457 10423 10466 10457
rect 10414 10414 10466 10423
rect 10414 10297 10466 10306
rect 10414 10263 10423 10297
rect 10423 10263 10457 10297
rect 10457 10263 10466 10297
rect 10414 10254 10466 10263
rect 10414 10137 10466 10146
rect 10414 10103 10423 10137
rect 10423 10103 10457 10137
rect 10457 10103 10466 10137
rect 10414 10094 10466 10103
rect 10414 9977 10466 9986
rect 10414 9943 10423 9977
rect 10423 9943 10457 9977
rect 10457 9943 10466 9977
rect 10414 9934 10466 9943
rect 10414 9817 10466 9826
rect 10414 9783 10423 9817
rect 10423 9783 10457 9817
rect 10457 9783 10466 9817
rect 10414 9774 10466 9783
rect 10414 9497 10466 9506
rect 10414 9463 10423 9497
rect 10423 9463 10457 9497
rect 10457 9463 10466 9497
rect 10414 9454 10466 9463
rect 10414 9337 10466 9346
rect 10414 9303 10423 9337
rect 10423 9303 10457 9337
rect 10457 9303 10466 9337
rect 10414 9294 10466 9303
rect 10414 9017 10466 9026
rect 10414 8983 10423 9017
rect 10423 8983 10457 9017
rect 10457 8983 10466 9017
rect 10414 8974 10466 8983
rect 10414 8857 10466 8866
rect 10414 8823 10423 8857
rect 10423 8823 10457 8857
rect 10457 8823 10466 8857
rect 10414 8814 10466 8823
rect 10414 8697 10466 8706
rect 10414 8663 10423 8697
rect 10423 8663 10457 8697
rect 10457 8663 10466 8697
rect 10414 8654 10466 8663
rect 10414 8537 10466 8546
rect 10414 8503 10423 8537
rect 10423 8503 10457 8537
rect 10457 8503 10466 8537
rect 10414 8494 10466 8503
rect 10414 8377 10466 8386
rect 10414 8343 10423 8377
rect 10423 8343 10457 8377
rect 10457 8343 10466 8377
rect 10414 8334 10466 8343
rect 10414 8217 10466 8226
rect 10414 8183 10423 8217
rect 10423 8183 10457 8217
rect 10457 8183 10466 8217
rect 10414 8174 10466 8183
rect 10414 8057 10466 8066
rect 10414 8023 10423 8057
rect 10423 8023 10457 8057
rect 10457 8023 10466 8057
rect 10414 8014 10466 8023
rect 10414 7897 10466 7906
rect 10414 7863 10423 7897
rect 10423 7863 10457 7897
rect 10457 7863 10466 7897
rect 10414 7854 10466 7863
rect 10414 7737 10466 7746
rect 10414 7703 10423 7737
rect 10423 7703 10457 7737
rect 10457 7703 10466 7737
rect 10414 7694 10466 7703
rect 10414 7417 10466 7426
rect 10414 7383 10423 7417
rect 10423 7383 10457 7417
rect 10457 7383 10466 7417
rect 10414 7374 10466 7383
rect 10414 7257 10466 7266
rect 10414 7223 10423 7257
rect 10423 7223 10457 7257
rect 10457 7223 10466 7257
rect 10414 7214 10466 7223
rect 10414 6937 10466 6946
rect 10414 6903 10423 6937
rect 10423 6903 10457 6937
rect 10457 6903 10466 6937
rect 10414 6894 10466 6903
rect 10414 6777 10466 6786
rect 10414 6743 10423 6777
rect 10423 6743 10457 6777
rect 10457 6743 10466 6777
rect 10414 6734 10466 6743
rect 10414 6457 10466 6466
rect 10414 6423 10423 6457
rect 10423 6423 10457 6457
rect 10457 6423 10466 6457
rect 10414 6414 10466 6423
rect 10414 6297 10466 6306
rect 10414 6263 10423 6297
rect 10423 6263 10457 6297
rect 10457 6263 10466 6297
rect 10414 6254 10466 6263
rect 10414 6137 10466 6146
rect 10414 6103 10423 6137
rect 10423 6103 10457 6137
rect 10457 6103 10466 6137
rect 10414 6094 10466 6103
rect 10414 5977 10466 5986
rect 10414 5943 10423 5977
rect 10423 5943 10457 5977
rect 10457 5943 10466 5977
rect 10414 5934 10466 5943
rect 10414 5817 10466 5826
rect 10414 5783 10423 5817
rect 10423 5783 10457 5817
rect 10457 5783 10466 5817
rect 10414 5774 10466 5783
rect 10414 5657 10466 5666
rect 10414 5623 10423 5657
rect 10423 5623 10457 5657
rect 10457 5623 10466 5657
rect 10414 5614 10466 5623
rect 10414 5497 10466 5506
rect 10414 5463 10423 5497
rect 10423 5463 10457 5497
rect 10457 5463 10466 5497
rect 10414 5454 10466 5463
rect 10414 5337 10466 5346
rect 10414 5303 10423 5337
rect 10423 5303 10457 5337
rect 10457 5303 10466 5337
rect 10414 5294 10466 5303
rect 10414 5177 10466 5186
rect 10414 5143 10423 5177
rect 10423 5143 10457 5177
rect 10457 5143 10466 5177
rect 10414 5134 10466 5143
rect 10414 5017 10466 5026
rect 10414 4983 10423 5017
rect 10423 4983 10457 5017
rect 10457 4983 10466 5017
rect 10414 4974 10466 4983
rect 10414 4857 10466 4866
rect 10414 4823 10423 4857
rect 10423 4823 10457 4857
rect 10457 4823 10466 4857
rect 10414 4814 10466 4823
rect 10414 4697 10466 4706
rect 10414 4663 10423 4697
rect 10423 4663 10457 4697
rect 10457 4663 10466 4697
rect 10414 4654 10466 4663
rect 10414 4537 10466 4546
rect 10414 4503 10423 4537
rect 10423 4503 10457 4537
rect 10457 4503 10466 4537
rect 10414 4494 10466 4503
rect 10414 4377 10466 4386
rect 10414 4343 10423 4377
rect 10423 4343 10457 4377
rect 10457 4343 10466 4377
rect 10414 4334 10466 4343
rect 10414 4217 10466 4226
rect 10414 4183 10423 4217
rect 10423 4183 10457 4217
rect 10457 4183 10466 4217
rect 10414 4174 10466 4183
rect 10414 4057 10466 4066
rect 10414 4023 10423 4057
rect 10423 4023 10457 4057
rect 10457 4023 10466 4057
rect 10414 4014 10466 4023
rect 10414 3897 10466 3906
rect 10414 3863 10423 3897
rect 10423 3863 10457 3897
rect 10457 3863 10466 3897
rect 10414 3854 10466 3863
rect 10414 3417 10466 3426
rect 10414 3383 10423 3417
rect 10423 3383 10457 3417
rect 10457 3383 10466 3417
rect 10414 3374 10466 3383
rect 10414 3257 10466 3266
rect 10414 3223 10423 3257
rect 10423 3223 10457 3257
rect 10457 3223 10466 3257
rect 10414 3214 10466 3223
rect 10414 3097 10466 3106
rect 10414 3063 10423 3097
rect 10423 3063 10457 3097
rect 10457 3063 10466 3097
rect 10414 3054 10466 3063
rect 10414 2937 10466 2946
rect 10414 2903 10423 2937
rect 10423 2903 10457 2937
rect 10457 2903 10466 2937
rect 10414 2894 10466 2903
rect 10414 2777 10466 2786
rect 10414 2743 10423 2777
rect 10423 2743 10457 2777
rect 10457 2743 10466 2777
rect 10414 2734 10466 2743
rect 10414 2617 10466 2626
rect 10414 2583 10423 2617
rect 10423 2583 10457 2617
rect 10457 2583 10466 2617
rect 10414 2574 10466 2583
rect 10414 2457 10466 2466
rect 10414 2423 10423 2457
rect 10423 2423 10457 2457
rect 10457 2423 10466 2457
rect 10414 2414 10466 2423
rect 10414 2297 10466 2306
rect 10414 2263 10423 2297
rect 10423 2263 10457 2297
rect 10457 2263 10466 2297
rect 10414 2254 10466 2263
rect 10414 2137 10466 2146
rect 10414 2103 10423 2137
rect 10423 2103 10457 2137
rect 10457 2103 10466 2137
rect 10414 2094 10466 2103
rect 10414 1977 10466 1986
rect 10414 1943 10423 1977
rect 10423 1943 10457 1977
rect 10457 1943 10466 1977
rect 10414 1934 10466 1943
rect 10414 1657 10466 1666
rect 10414 1623 10423 1657
rect 10423 1623 10457 1657
rect 10457 1623 10466 1657
rect 10414 1614 10466 1623
rect 10414 1497 10466 1506
rect 10414 1463 10423 1497
rect 10423 1463 10457 1497
rect 10457 1463 10466 1497
rect 10414 1454 10466 1463
rect 10414 1337 10466 1346
rect 10414 1303 10423 1337
rect 10423 1303 10457 1337
rect 10457 1303 10466 1337
rect 10414 1294 10466 1303
rect 10414 1177 10466 1186
rect 10414 1143 10423 1177
rect 10423 1143 10457 1177
rect 10457 1143 10466 1177
rect 10414 1134 10466 1143
rect 10414 1017 10466 1026
rect 10414 983 10423 1017
rect 10423 983 10457 1017
rect 10457 983 10466 1017
rect 10414 974 10466 983
rect 10414 537 10466 546
rect 10414 503 10423 537
rect 10423 503 10457 537
rect 10457 503 10466 537
rect 10414 494 10466 503
rect 10414 377 10466 386
rect 10414 343 10423 377
rect 10423 343 10457 377
rect 10457 343 10466 377
rect 10414 334 10466 343
rect 10414 217 10466 226
rect 10414 183 10423 217
rect 10423 183 10457 217
rect 10457 183 10466 217
rect 10414 174 10466 183
rect 10414 57 10466 66
rect 10414 23 10423 57
rect 10423 23 10457 57
rect 10457 23 10466 57
rect 10414 14 10466 23
rect 10734 31417 10786 31426
rect 10734 31383 10743 31417
rect 10743 31383 10777 31417
rect 10777 31383 10786 31417
rect 10734 31374 10786 31383
rect 10734 31257 10786 31266
rect 10734 31223 10743 31257
rect 10743 31223 10777 31257
rect 10777 31223 10786 31257
rect 10734 31214 10786 31223
rect 10734 31097 10786 31106
rect 10734 31063 10743 31097
rect 10743 31063 10777 31097
rect 10777 31063 10786 31097
rect 10734 31054 10786 31063
rect 10734 30937 10786 30946
rect 10734 30903 10743 30937
rect 10743 30903 10777 30937
rect 10777 30903 10786 30937
rect 10734 30894 10786 30903
rect 10734 30777 10786 30786
rect 10734 30743 10743 30777
rect 10743 30743 10777 30777
rect 10777 30743 10786 30777
rect 10734 30734 10786 30743
rect 10734 30617 10786 30626
rect 10734 30583 10743 30617
rect 10743 30583 10777 30617
rect 10777 30583 10786 30617
rect 10734 30574 10786 30583
rect 10734 30457 10786 30466
rect 10734 30423 10743 30457
rect 10743 30423 10777 30457
rect 10777 30423 10786 30457
rect 10734 30414 10786 30423
rect 10734 30297 10786 30306
rect 10734 30263 10743 30297
rect 10743 30263 10777 30297
rect 10777 30263 10786 30297
rect 10734 30254 10786 30263
rect 10734 29977 10786 29986
rect 10734 29943 10743 29977
rect 10743 29943 10777 29977
rect 10777 29943 10786 29977
rect 10734 29934 10786 29943
rect 10734 29817 10786 29826
rect 10734 29783 10743 29817
rect 10743 29783 10777 29817
rect 10777 29783 10786 29817
rect 10734 29774 10786 29783
rect 10734 29657 10786 29666
rect 10734 29623 10743 29657
rect 10743 29623 10777 29657
rect 10777 29623 10786 29657
rect 10734 29614 10786 29623
rect 10734 29497 10786 29506
rect 10734 29463 10743 29497
rect 10743 29463 10777 29497
rect 10777 29463 10786 29497
rect 10734 29454 10786 29463
rect 10734 29337 10786 29346
rect 10734 29303 10743 29337
rect 10743 29303 10777 29337
rect 10777 29303 10786 29337
rect 10734 29294 10786 29303
rect 10734 29177 10786 29186
rect 10734 29143 10743 29177
rect 10743 29143 10777 29177
rect 10777 29143 10786 29177
rect 10734 29134 10786 29143
rect 10734 29017 10786 29026
rect 10734 28983 10743 29017
rect 10743 28983 10777 29017
rect 10777 28983 10786 29017
rect 10734 28974 10786 28983
rect 10734 28857 10786 28866
rect 10734 28823 10743 28857
rect 10743 28823 10777 28857
rect 10777 28823 10786 28857
rect 10734 28814 10786 28823
rect 10734 28057 10786 28066
rect 10734 28023 10743 28057
rect 10743 28023 10777 28057
rect 10777 28023 10786 28057
rect 10734 28014 10786 28023
rect 10734 27897 10786 27906
rect 10734 27863 10743 27897
rect 10743 27863 10777 27897
rect 10777 27863 10786 27897
rect 10734 27854 10786 27863
rect 10734 27737 10786 27746
rect 10734 27703 10743 27737
rect 10743 27703 10777 27737
rect 10777 27703 10786 27737
rect 10734 27694 10786 27703
rect 10734 27577 10786 27586
rect 10734 27543 10743 27577
rect 10743 27543 10777 27577
rect 10777 27543 10786 27577
rect 10734 27534 10786 27543
rect 10734 27417 10786 27426
rect 10734 27383 10743 27417
rect 10743 27383 10777 27417
rect 10777 27383 10786 27417
rect 10734 27374 10786 27383
rect 10734 27257 10786 27266
rect 10734 27223 10743 27257
rect 10743 27223 10777 27257
rect 10777 27223 10786 27257
rect 10734 27214 10786 27223
rect 10734 27097 10786 27106
rect 10734 27063 10743 27097
rect 10743 27063 10777 27097
rect 10777 27063 10786 27097
rect 10734 27054 10786 27063
rect 10734 26937 10786 26946
rect 10734 26903 10743 26937
rect 10743 26903 10777 26937
rect 10777 26903 10786 26937
rect 10734 26894 10786 26903
rect 10734 26137 10786 26146
rect 10734 26103 10743 26137
rect 10743 26103 10777 26137
rect 10777 26103 10786 26137
rect 10734 26094 10786 26103
rect 10734 25977 10786 25986
rect 10734 25943 10743 25977
rect 10743 25943 10777 25977
rect 10777 25943 10786 25977
rect 10734 25934 10786 25943
rect 10734 25817 10786 25826
rect 10734 25783 10743 25817
rect 10743 25783 10777 25817
rect 10777 25783 10786 25817
rect 10734 25774 10786 25783
rect 10734 25657 10786 25666
rect 10734 25623 10743 25657
rect 10743 25623 10777 25657
rect 10777 25623 10786 25657
rect 10734 25614 10786 25623
rect 10734 25497 10786 25506
rect 10734 25463 10743 25497
rect 10743 25463 10777 25497
rect 10777 25463 10786 25497
rect 10734 25454 10786 25463
rect 10734 25337 10786 25346
rect 10734 25303 10743 25337
rect 10743 25303 10777 25337
rect 10777 25303 10786 25337
rect 10734 25294 10786 25303
rect 10734 25177 10786 25186
rect 10734 25143 10743 25177
rect 10743 25143 10777 25177
rect 10777 25143 10786 25177
rect 10734 25134 10786 25143
rect 10734 25017 10786 25026
rect 10734 24983 10743 25017
rect 10743 24983 10777 25017
rect 10777 24983 10786 25017
rect 10734 24974 10786 24983
rect 10734 24697 10786 24706
rect 10734 24663 10743 24697
rect 10743 24663 10777 24697
rect 10777 24663 10786 24697
rect 10734 24654 10786 24663
rect 10734 24537 10786 24546
rect 10734 24503 10743 24537
rect 10743 24503 10777 24537
rect 10777 24503 10786 24537
rect 10734 24494 10786 24503
rect 10734 24377 10786 24386
rect 10734 24343 10743 24377
rect 10743 24343 10777 24377
rect 10777 24343 10786 24377
rect 10734 24334 10786 24343
rect 10734 24217 10786 24226
rect 10734 24183 10743 24217
rect 10743 24183 10777 24217
rect 10777 24183 10786 24217
rect 10734 24174 10786 24183
rect 10734 24057 10786 24066
rect 10734 24023 10743 24057
rect 10743 24023 10777 24057
rect 10777 24023 10786 24057
rect 10734 24014 10786 24023
rect 10734 23897 10786 23906
rect 10734 23863 10743 23897
rect 10743 23863 10777 23897
rect 10777 23863 10786 23897
rect 10734 23854 10786 23863
rect 10734 23737 10786 23746
rect 10734 23703 10743 23737
rect 10743 23703 10777 23737
rect 10777 23703 10786 23737
rect 10734 23694 10786 23703
rect 10734 23577 10786 23586
rect 10734 23543 10743 23577
rect 10743 23543 10777 23577
rect 10777 23543 10786 23577
rect 10734 23534 10786 23543
rect 10734 23417 10786 23426
rect 10734 23383 10743 23417
rect 10743 23383 10777 23417
rect 10777 23383 10786 23417
rect 10734 23374 10786 23383
rect 10734 23257 10786 23266
rect 10734 23223 10743 23257
rect 10743 23223 10777 23257
rect 10777 23223 10786 23257
rect 10734 23214 10786 23223
rect 10734 23097 10786 23106
rect 10734 23063 10743 23097
rect 10743 23063 10777 23097
rect 10777 23063 10786 23097
rect 10734 23054 10786 23063
rect 10734 22937 10786 22946
rect 10734 22903 10743 22937
rect 10743 22903 10777 22937
rect 10777 22903 10786 22937
rect 10734 22894 10786 22903
rect 10734 22777 10786 22786
rect 10734 22743 10743 22777
rect 10743 22743 10777 22777
rect 10777 22743 10786 22777
rect 10734 22734 10786 22743
rect 10734 22617 10786 22626
rect 10734 22583 10743 22617
rect 10743 22583 10777 22617
rect 10777 22583 10786 22617
rect 10734 22574 10786 22583
rect 10734 22457 10786 22466
rect 10734 22423 10743 22457
rect 10743 22423 10777 22457
rect 10777 22423 10786 22457
rect 10734 22414 10786 22423
rect 10734 22297 10786 22306
rect 10734 22263 10743 22297
rect 10743 22263 10777 22297
rect 10777 22263 10786 22297
rect 10734 22254 10786 22263
rect 10734 22137 10786 22146
rect 10734 22103 10743 22137
rect 10743 22103 10777 22137
rect 10777 22103 10786 22137
rect 10734 22094 10786 22103
rect 10734 21817 10786 21826
rect 10734 21783 10743 21817
rect 10743 21783 10777 21817
rect 10777 21783 10786 21817
rect 10734 21774 10786 21783
rect 10734 21657 10786 21666
rect 10734 21623 10743 21657
rect 10743 21623 10777 21657
rect 10777 21623 10786 21657
rect 10734 21614 10786 21623
rect 10734 21497 10786 21506
rect 10734 21463 10743 21497
rect 10743 21463 10777 21497
rect 10777 21463 10786 21497
rect 10734 21454 10786 21463
rect 10734 21337 10786 21346
rect 10734 21303 10743 21337
rect 10743 21303 10777 21337
rect 10777 21303 10786 21337
rect 10734 21294 10786 21303
rect 10734 21177 10786 21186
rect 10734 21143 10743 21177
rect 10743 21143 10777 21177
rect 10777 21143 10786 21177
rect 10734 21134 10786 21143
rect 10734 21017 10786 21026
rect 10734 20983 10743 21017
rect 10743 20983 10777 21017
rect 10777 20983 10786 21017
rect 10734 20974 10786 20983
rect 10734 20857 10786 20866
rect 10734 20823 10743 20857
rect 10743 20823 10777 20857
rect 10777 20823 10786 20857
rect 10734 20814 10786 20823
rect 10734 20697 10786 20706
rect 10734 20663 10743 20697
rect 10743 20663 10777 20697
rect 10777 20663 10786 20697
rect 10734 20654 10786 20663
rect 10734 19897 10786 19906
rect 10734 19863 10743 19897
rect 10743 19863 10777 19897
rect 10777 19863 10786 19897
rect 10734 19854 10786 19863
rect 10734 19737 10786 19746
rect 10734 19703 10743 19737
rect 10743 19703 10777 19737
rect 10777 19703 10786 19737
rect 10734 19694 10786 19703
rect 10734 19577 10786 19586
rect 10734 19543 10743 19577
rect 10743 19543 10777 19577
rect 10777 19543 10786 19577
rect 10734 19534 10786 19543
rect 10734 19417 10786 19426
rect 10734 19383 10743 19417
rect 10743 19383 10777 19417
rect 10777 19383 10786 19417
rect 10734 19374 10786 19383
rect 10734 19257 10786 19266
rect 10734 19223 10743 19257
rect 10743 19223 10777 19257
rect 10777 19223 10786 19257
rect 10734 19214 10786 19223
rect 10734 19097 10786 19106
rect 10734 19063 10743 19097
rect 10743 19063 10777 19097
rect 10777 19063 10786 19097
rect 10734 19054 10786 19063
rect 10734 18937 10786 18946
rect 10734 18903 10743 18937
rect 10743 18903 10777 18937
rect 10777 18903 10786 18937
rect 10734 18894 10786 18903
rect 10734 18777 10786 18786
rect 10734 18743 10743 18777
rect 10743 18743 10777 18777
rect 10777 18743 10786 18777
rect 10734 18734 10786 18743
rect 10734 17977 10786 17986
rect 10734 17943 10743 17977
rect 10743 17943 10777 17977
rect 10777 17943 10786 17977
rect 10734 17934 10786 17943
rect 10734 17817 10786 17826
rect 10734 17783 10743 17817
rect 10743 17783 10777 17817
rect 10777 17783 10786 17817
rect 10734 17774 10786 17783
rect 10734 17657 10786 17666
rect 10734 17623 10743 17657
rect 10743 17623 10777 17657
rect 10777 17623 10786 17657
rect 10734 17614 10786 17623
rect 10734 17497 10786 17506
rect 10734 17463 10743 17497
rect 10743 17463 10777 17497
rect 10777 17463 10786 17497
rect 10734 17454 10786 17463
rect 10734 17337 10786 17346
rect 10734 17303 10743 17337
rect 10743 17303 10777 17337
rect 10777 17303 10786 17337
rect 10734 17294 10786 17303
rect 10734 17177 10786 17186
rect 10734 17143 10743 17177
rect 10743 17143 10777 17177
rect 10777 17143 10786 17177
rect 10734 17134 10786 17143
rect 10734 17017 10786 17026
rect 10734 16983 10743 17017
rect 10743 16983 10777 17017
rect 10777 16983 10786 17017
rect 10734 16974 10786 16983
rect 10734 16857 10786 16866
rect 10734 16823 10743 16857
rect 10743 16823 10777 16857
rect 10777 16823 10786 16857
rect 10734 16814 10786 16823
rect 10734 16537 10786 16546
rect 10734 16503 10743 16537
rect 10743 16503 10777 16537
rect 10777 16503 10786 16537
rect 10734 16494 10786 16503
rect 10734 16377 10786 16386
rect 10734 16343 10743 16377
rect 10743 16343 10777 16377
rect 10777 16343 10786 16377
rect 10734 16334 10786 16343
rect 10734 16217 10786 16226
rect 10734 16183 10743 16217
rect 10743 16183 10777 16217
rect 10777 16183 10786 16217
rect 10734 16174 10786 16183
rect 10734 16057 10786 16066
rect 10734 16023 10743 16057
rect 10743 16023 10777 16057
rect 10777 16023 10786 16057
rect 10734 16014 10786 16023
rect 10734 15897 10786 15906
rect 10734 15863 10743 15897
rect 10743 15863 10777 15897
rect 10777 15863 10786 15897
rect 10734 15854 10786 15863
rect 10734 15737 10786 15746
rect 10734 15703 10743 15737
rect 10743 15703 10777 15737
rect 10777 15703 10786 15737
rect 10734 15694 10786 15703
rect 10734 15577 10786 15586
rect 10734 15543 10743 15577
rect 10743 15543 10777 15577
rect 10777 15543 10786 15577
rect 10734 15534 10786 15543
rect 10734 15417 10786 15426
rect 10734 15383 10743 15417
rect 10743 15383 10777 15417
rect 10777 15383 10786 15417
rect 10734 15374 10786 15383
rect 10734 15257 10786 15266
rect 10734 15223 10743 15257
rect 10743 15223 10777 15257
rect 10777 15223 10786 15257
rect 10734 15214 10786 15223
rect 10734 15097 10786 15106
rect 10734 15063 10743 15097
rect 10743 15063 10777 15097
rect 10777 15063 10786 15097
rect 10734 15054 10786 15063
rect 10734 14937 10786 14946
rect 10734 14903 10743 14937
rect 10743 14903 10777 14937
rect 10777 14903 10786 14937
rect 10734 14894 10786 14903
rect 10734 14777 10786 14786
rect 10734 14743 10743 14777
rect 10743 14743 10777 14777
rect 10777 14743 10786 14777
rect 10734 14734 10786 14743
rect 10734 14617 10786 14626
rect 10734 14583 10743 14617
rect 10743 14583 10777 14617
rect 10777 14583 10786 14617
rect 10734 14574 10786 14583
rect 10734 14457 10786 14466
rect 10734 14423 10743 14457
rect 10743 14423 10777 14457
rect 10777 14423 10786 14457
rect 10734 14414 10786 14423
rect 10734 14297 10786 14306
rect 10734 14263 10743 14297
rect 10743 14263 10777 14297
rect 10777 14263 10786 14297
rect 10734 14254 10786 14263
rect 10734 14137 10786 14146
rect 10734 14103 10743 14137
rect 10743 14103 10777 14137
rect 10777 14103 10786 14137
rect 10734 14094 10786 14103
rect 10734 13977 10786 13986
rect 10734 13943 10743 13977
rect 10743 13943 10777 13977
rect 10777 13943 10786 13977
rect 10734 13934 10786 13943
rect 10734 13657 10786 13666
rect 10734 13623 10743 13657
rect 10743 13623 10777 13657
rect 10777 13623 10786 13657
rect 10734 13614 10786 13623
rect 10734 13497 10786 13506
rect 10734 13463 10743 13497
rect 10743 13463 10777 13497
rect 10777 13463 10786 13497
rect 10734 13454 10786 13463
rect 10734 13337 10786 13346
rect 10734 13303 10743 13337
rect 10743 13303 10777 13337
rect 10777 13303 10786 13337
rect 10734 13294 10786 13303
rect 10734 13177 10786 13186
rect 10734 13143 10743 13177
rect 10743 13143 10777 13177
rect 10777 13143 10786 13177
rect 10734 13134 10786 13143
rect 10734 13017 10786 13026
rect 10734 12983 10743 13017
rect 10743 12983 10777 13017
rect 10777 12983 10786 13017
rect 10734 12974 10786 12983
rect 10734 12857 10786 12866
rect 10734 12823 10743 12857
rect 10743 12823 10777 12857
rect 10777 12823 10786 12857
rect 10734 12814 10786 12823
rect 10734 12697 10786 12706
rect 10734 12663 10743 12697
rect 10743 12663 10777 12697
rect 10777 12663 10786 12697
rect 10734 12654 10786 12663
rect 10734 12537 10786 12546
rect 10734 12503 10743 12537
rect 10743 12503 10777 12537
rect 10777 12503 10786 12537
rect 10734 12494 10786 12503
rect 10734 11737 10786 11746
rect 10734 11703 10743 11737
rect 10743 11703 10777 11737
rect 10777 11703 10786 11737
rect 10734 11694 10786 11703
rect 10734 11577 10786 11586
rect 10734 11543 10743 11577
rect 10743 11543 10777 11577
rect 10777 11543 10786 11577
rect 10734 11534 10786 11543
rect 10734 11417 10786 11426
rect 10734 11383 10743 11417
rect 10743 11383 10777 11417
rect 10777 11383 10786 11417
rect 10734 11374 10786 11383
rect 10734 11257 10786 11266
rect 10734 11223 10743 11257
rect 10743 11223 10777 11257
rect 10777 11223 10786 11257
rect 10734 11214 10786 11223
rect 10734 11097 10786 11106
rect 10734 11063 10743 11097
rect 10743 11063 10777 11097
rect 10777 11063 10786 11097
rect 10734 11054 10786 11063
rect 10734 10937 10786 10946
rect 10734 10903 10743 10937
rect 10743 10903 10777 10937
rect 10777 10903 10786 10937
rect 10734 10894 10786 10903
rect 10734 10777 10786 10786
rect 10734 10743 10743 10777
rect 10743 10743 10777 10777
rect 10777 10743 10786 10777
rect 10734 10734 10786 10743
rect 10734 10617 10786 10626
rect 10734 10583 10743 10617
rect 10743 10583 10777 10617
rect 10777 10583 10786 10617
rect 10734 10574 10786 10583
rect 10734 10457 10786 10466
rect 10734 10423 10743 10457
rect 10743 10423 10777 10457
rect 10777 10423 10786 10457
rect 10734 10414 10786 10423
rect 10734 10297 10786 10306
rect 10734 10263 10743 10297
rect 10743 10263 10777 10297
rect 10777 10263 10786 10297
rect 10734 10254 10786 10263
rect 10734 10137 10786 10146
rect 10734 10103 10743 10137
rect 10743 10103 10777 10137
rect 10777 10103 10786 10137
rect 10734 10094 10786 10103
rect 10734 9977 10786 9986
rect 10734 9943 10743 9977
rect 10743 9943 10777 9977
rect 10777 9943 10786 9977
rect 10734 9934 10786 9943
rect 10734 9817 10786 9826
rect 10734 9783 10743 9817
rect 10743 9783 10777 9817
rect 10777 9783 10786 9817
rect 10734 9774 10786 9783
rect 10734 9497 10786 9506
rect 10734 9463 10743 9497
rect 10743 9463 10777 9497
rect 10777 9463 10786 9497
rect 10734 9454 10786 9463
rect 10734 9337 10786 9346
rect 10734 9303 10743 9337
rect 10743 9303 10777 9337
rect 10777 9303 10786 9337
rect 10734 9294 10786 9303
rect 10734 9017 10786 9026
rect 10734 8983 10743 9017
rect 10743 8983 10777 9017
rect 10777 8983 10786 9017
rect 10734 8974 10786 8983
rect 10734 8857 10786 8866
rect 10734 8823 10743 8857
rect 10743 8823 10777 8857
rect 10777 8823 10786 8857
rect 10734 8814 10786 8823
rect 10734 8697 10786 8706
rect 10734 8663 10743 8697
rect 10743 8663 10777 8697
rect 10777 8663 10786 8697
rect 10734 8654 10786 8663
rect 10734 8537 10786 8546
rect 10734 8503 10743 8537
rect 10743 8503 10777 8537
rect 10777 8503 10786 8537
rect 10734 8494 10786 8503
rect 10734 8377 10786 8386
rect 10734 8343 10743 8377
rect 10743 8343 10777 8377
rect 10777 8343 10786 8377
rect 10734 8334 10786 8343
rect 10734 8217 10786 8226
rect 10734 8183 10743 8217
rect 10743 8183 10777 8217
rect 10777 8183 10786 8217
rect 10734 8174 10786 8183
rect 10734 8057 10786 8066
rect 10734 8023 10743 8057
rect 10743 8023 10777 8057
rect 10777 8023 10786 8057
rect 10734 8014 10786 8023
rect 10734 7897 10786 7906
rect 10734 7863 10743 7897
rect 10743 7863 10777 7897
rect 10777 7863 10786 7897
rect 10734 7854 10786 7863
rect 10734 7737 10786 7746
rect 10734 7703 10743 7737
rect 10743 7703 10777 7737
rect 10777 7703 10786 7737
rect 10734 7694 10786 7703
rect 10734 7417 10786 7426
rect 10734 7383 10743 7417
rect 10743 7383 10777 7417
rect 10777 7383 10786 7417
rect 10734 7374 10786 7383
rect 10734 7257 10786 7266
rect 10734 7223 10743 7257
rect 10743 7223 10777 7257
rect 10777 7223 10786 7257
rect 10734 7214 10786 7223
rect 10734 6937 10786 6946
rect 10734 6903 10743 6937
rect 10743 6903 10777 6937
rect 10777 6903 10786 6937
rect 10734 6894 10786 6903
rect 10734 6777 10786 6786
rect 10734 6743 10743 6777
rect 10743 6743 10777 6777
rect 10777 6743 10786 6777
rect 10734 6734 10786 6743
rect 10734 6457 10786 6466
rect 10734 6423 10743 6457
rect 10743 6423 10777 6457
rect 10777 6423 10786 6457
rect 10734 6414 10786 6423
rect 10734 6297 10786 6306
rect 10734 6263 10743 6297
rect 10743 6263 10777 6297
rect 10777 6263 10786 6297
rect 10734 6254 10786 6263
rect 10734 6137 10786 6146
rect 10734 6103 10743 6137
rect 10743 6103 10777 6137
rect 10777 6103 10786 6137
rect 10734 6094 10786 6103
rect 10734 5977 10786 5986
rect 10734 5943 10743 5977
rect 10743 5943 10777 5977
rect 10777 5943 10786 5977
rect 10734 5934 10786 5943
rect 10734 5817 10786 5826
rect 10734 5783 10743 5817
rect 10743 5783 10777 5817
rect 10777 5783 10786 5817
rect 10734 5774 10786 5783
rect 10734 5657 10786 5666
rect 10734 5623 10743 5657
rect 10743 5623 10777 5657
rect 10777 5623 10786 5657
rect 10734 5614 10786 5623
rect 10734 5497 10786 5506
rect 10734 5463 10743 5497
rect 10743 5463 10777 5497
rect 10777 5463 10786 5497
rect 10734 5454 10786 5463
rect 10734 5337 10786 5346
rect 10734 5303 10743 5337
rect 10743 5303 10777 5337
rect 10777 5303 10786 5337
rect 10734 5294 10786 5303
rect 10734 5177 10786 5186
rect 10734 5143 10743 5177
rect 10743 5143 10777 5177
rect 10777 5143 10786 5177
rect 10734 5134 10786 5143
rect 10734 5017 10786 5026
rect 10734 4983 10743 5017
rect 10743 4983 10777 5017
rect 10777 4983 10786 5017
rect 10734 4974 10786 4983
rect 10734 4857 10786 4866
rect 10734 4823 10743 4857
rect 10743 4823 10777 4857
rect 10777 4823 10786 4857
rect 10734 4814 10786 4823
rect 10734 4697 10786 4706
rect 10734 4663 10743 4697
rect 10743 4663 10777 4697
rect 10777 4663 10786 4697
rect 10734 4654 10786 4663
rect 10734 4537 10786 4546
rect 10734 4503 10743 4537
rect 10743 4503 10777 4537
rect 10777 4503 10786 4537
rect 10734 4494 10786 4503
rect 10734 4377 10786 4386
rect 10734 4343 10743 4377
rect 10743 4343 10777 4377
rect 10777 4343 10786 4377
rect 10734 4334 10786 4343
rect 10734 4217 10786 4226
rect 10734 4183 10743 4217
rect 10743 4183 10777 4217
rect 10777 4183 10786 4217
rect 10734 4174 10786 4183
rect 10734 4057 10786 4066
rect 10734 4023 10743 4057
rect 10743 4023 10777 4057
rect 10777 4023 10786 4057
rect 10734 4014 10786 4023
rect 10734 3897 10786 3906
rect 10734 3863 10743 3897
rect 10743 3863 10777 3897
rect 10777 3863 10786 3897
rect 10734 3854 10786 3863
rect 10734 3417 10786 3426
rect 10734 3383 10743 3417
rect 10743 3383 10777 3417
rect 10777 3383 10786 3417
rect 10734 3374 10786 3383
rect 10734 3257 10786 3266
rect 10734 3223 10743 3257
rect 10743 3223 10777 3257
rect 10777 3223 10786 3257
rect 10734 3214 10786 3223
rect 10734 3097 10786 3106
rect 10734 3063 10743 3097
rect 10743 3063 10777 3097
rect 10777 3063 10786 3097
rect 10734 3054 10786 3063
rect 10734 2937 10786 2946
rect 10734 2903 10743 2937
rect 10743 2903 10777 2937
rect 10777 2903 10786 2937
rect 10734 2894 10786 2903
rect 10734 2777 10786 2786
rect 10734 2743 10743 2777
rect 10743 2743 10777 2777
rect 10777 2743 10786 2777
rect 10734 2734 10786 2743
rect 10734 2617 10786 2626
rect 10734 2583 10743 2617
rect 10743 2583 10777 2617
rect 10777 2583 10786 2617
rect 10734 2574 10786 2583
rect 10734 2457 10786 2466
rect 10734 2423 10743 2457
rect 10743 2423 10777 2457
rect 10777 2423 10786 2457
rect 10734 2414 10786 2423
rect 10734 2297 10786 2306
rect 10734 2263 10743 2297
rect 10743 2263 10777 2297
rect 10777 2263 10786 2297
rect 10734 2254 10786 2263
rect 10734 2137 10786 2146
rect 10734 2103 10743 2137
rect 10743 2103 10777 2137
rect 10777 2103 10786 2137
rect 10734 2094 10786 2103
rect 10734 1977 10786 1986
rect 10734 1943 10743 1977
rect 10743 1943 10777 1977
rect 10777 1943 10786 1977
rect 10734 1934 10786 1943
rect 10734 1657 10786 1666
rect 10734 1623 10743 1657
rect 10743 1623 10777 1657
rect 10777 1623 10786 1657
rect 10734 1614 10786 1623
rect 10734 1497 10786 1506
rect 10734 1463 10743 1497
rect 10743 1463 10777 1497
rect 10777 1463 10786 1497
rect 10734 1454 10786 1463
rect 10734 1337 10786 1346
rect 10734 1303 10743 1337
rect 10743 1303 10777 1337
rect 10777 1303 10786 1337
rect 10734 1294 10786 1303
rect 10734 1177 10786 1186
rect 10734 1143 10743 1177
rect 10743 1143 10777 1177
rect 10777 1143 10786 1177
rect 10734 1134 10786 1143
rect 10734 1017 10786 1026
rect 10734 983 10743 1017
rect 10743 983 10777 1017
rect 10777 983 10786 1017
rect 10734 974 10786 983
rect 10734 537 10786 546
rect 10734 503 10743 537
rect 10743 503 10777 537
rect 10777 503 10786 537
rect 10734 494 10786 503
rect 10734 377 10786 386
rect 10734 343 10743 377
rect 10743 343 10777 377
rect 10777 343 10786 377
rect 10734 334 10786 343
rect 10734 217 10786 226
rect 10734 183 10743 217
rect 10743 183 10777 217
rect 10777 183 10786 217
rect 10734 174 10786 183
rect 10734 57 10786 66
rect 10734 23 10743 57
rect 10743 23 10777 57
rect 10777 23 10786 57
rect 10734 14 10786 23
rect 11054 31417 11106 31426
rect 11054 31383 11063 31417
rect 11063 31383 11097 31417
rect 11097 31383 11106 31417
rect 11054 31374 11106 31383
rect 11054 31257 11106 31266
rect 11054 31223 11063 31257
rect 11063 31223 11097 31257
rect 11097 31223 11106 31257
rect 11054 31214 11106 31223
rect 11054 31097 11106 31106
rect 11054 31063 11063 31097
rect 11063 31063 11097 31097
rect 11097 31063 11106 31097
rect 11054 31054 11106 31063
rect 11054 30937 11106 30946
rect 11054 30903 11063 30937
rect 11063 30903 11097 30937
rect 11097 30903 11106 30937
rect 11054 30894 11106 30903
rect 11054 30777 11106 30786
rect 11054 30743 11063 30777
rect 11063 30743 11097 30777
rect 11097 30743 11106 30777
rect 11054 30734 11106 30743
rect 11054 30617 11106 30626
rect 11054 30583 11063 30617
rect 11063 30583 11097 30617
rect 11097 30583 11106 30617
rect 11054 30574 11106 30583
rect 11054 30457 11106 30466
rect 11054 30423 11063 30457
rect 11063 30423 11097 30457
rect 11097 30423 11106 30457
rect 11054 30414 11106 30423
rect 11054 30297 11106 30306
rect 11054 30263 11063 30297
rect 11063 30263 11097 30297
rect 11097 30263 11106 30297
rect 11054 30254 11106 30263
rect 11054 29977 11106 29986
rect 11054 29943 11063 29977
rect 11063 29943 11097 29977
rect 11097 29943 11106 29977
rect 11054 29934 11106 29943
rect 11054 29817 11106 29826
rect 11054 29783 11063 29817
rect 11063 29783 11097 29817
rect 11097 29783 11106 29817
rect 11054 29774 11106 29783
rect 11054 29657 11106 29666
rect 11054 29623 11063 29657
rect 11063 29623 11097 29657
rect 11097 29623 11106 29657
rect 11054 29614 11106 29623
rect 11054 29497 11106 29506
rect 11054 29463 11063 29497
rect 11063 29463 11097 29497
rect 11097 29463 11106 29497
rect 11054 29454 11106 29463
rect 11054 29337 11106 29346
rect 11054 29303 11063 29337
rect 11063 29303 11097 29337
rect 11097 29303 11106 29337
rect 11054 29294 11106 29303
rect 11054 29177 11106 29186
rect 11054 29143 11063 29177
rect 11063 29143 11097 29177
rect 11097 29143 11106 29177
rect 11054 29134 11106 29143
rect 11054 29017 11106 29026
rect 11054 28983 11063 29017
rect 11063 28983 11097 29017
rect 11097 28983 11106 29017
rect 11054 28974 11106 28983
rect 11054 28857 11106 28866
rect 11054 28823 11063 28857
rect 11063 28823 11097 28857
rect 11097 28823 11106 28857
rect 11054 28814 11106 28823
rect 11054 28057 11106 28066
rect 11054 28023 11063 28057
rect 11063 28023 11097 28057
rect 11097 28023 11106 28057
rect 11054 28014 11106 28023
rect 11054 27897 11106 27906
rect 11054 27863 11063 27897
rect 11063 27863 11097 27897
rect 11097 27863 11106 27897
rect 11054 27854 11106 27863
rect 11054 27737 11106 27746
rect 11054 27703 11063 27737
rect 11063 27703 11097 27737
rect 11097 27703 11106 27737
rect 11054 27694 11106 27703
rect 11054 27577 11106 27586
rect 11054 27543 11063 27577
rect 11063 27543 11097 27577
rect 11097 27543 11106 27577
rect 11054 27534 11106 27543
rect 11054 27417 11106 27426
rect 11054 27383 11063 27417
rect 11063 27383 11097 27417
rect 11097 27383 11106 27417
rect 11054 27374 11106 27383
rect 11054 27257 11106 27266
rect 11054 27223 11063 27257
rect 11063 27223 11097 27257
rect 11097 27223 11106 27257
rect 11054 27214 11106 27223
rect 11054 27097 11106 27106
rect 11054 27063 11063 27097
rect 11063 27063 11097 27097
rect 11097 27063 11106 27097
rect 11054 27054 11106 27063
rect 11054 26937 11106 26946
rect 11054 26903 11063 26937
rect 11063 26903 11097 26937
rect 11097 26903 11106 26937
rect 11054 26894 11106 26903
rect 11054 26137 11106 26146
rect 11054 26103 11063 26137
rect 11063 26103 11097 26137
rect 11097 26103 11106 26137
rect 11054 26094 11106 26103
rect 11054 25977 11106 25986
rect 11054 25943 11063 25977
rect 11063 25943 11097 25977
rect 11097 25943 11106 25977
rect 11054 25934 11106 25943
rect 11054 25817 11106 25826
rect 11054 25783 11063 25817
rect 11063 25783 11097 25817
rect 11097 25783 11106 25817
rect 11054 25774 11106 25783
rect 11054 25657 11106 25666
rect 11054 25623 11063 25657
rect 11063 25623 11097 25657
rect 11097 25623 11106 25657
rect 11054 25614 11106 25623
rect 11054 25497 11106 25506
rect 11054 25463 11063 25497
rect 11063 25463 11097 25497
rect 11097 25463 11106 25497
rect 11054 25454 11106 25463
rect 11054 25337 11106 25346
rect 11054 25303 11063 25337
rect 11063 25303 11097 25337
rect 11097 25303 11106 25337
rect 11054 25294 11106 25303
rect 11054 25177 11106 25186
rect 11054 25143 11063 25177
rect 11063 25143 11097 25177
rect 11097 25143 11106 25177
rect 11054 25134 11106 25143
rect 11054 25017 11106 25026
rect 11054 24983 11063 25017
rect 11063 24983 11097 25017
rect 11097 24983 11106 25017
rect 11054 24974 11106 24983
rect 11054 24697 11106 24706
rect 11054 24663 11063 24697
rect 11063 24663 11097 24697
rect 11097 24663 11106 24697
rect 11054 24654 11106 24663
rect 11054 24537 11106 24546
rect 11054 24503 11063 24537
rect 11063 24503 11097 24537
rect 11097 24503 11106 24537
rect 11054 24494 11106 24503
rect 11054 24377 11106 24386
rect 11054 24343 11063 24377
rect 11063 24343 11097 24377
rect 11097 24343 11106 24377
rect 11054 24334 11106 24343
rect 11054 24217 11106 24226
rect 11054 24183 11063 24217
rect 11063 24183 11097 24217
rect 11097 24183 11106 24217
rect 11054 24174 11106 24183
rect 11054 24057 11106 24066
rect 11054 24023 11063 24057
rect 11063 24023 11097 24057
rect 11097 24023 11106 24057
rect 11054 24014 11106 24023
rect 11054 23897 11106 23906
rect 11054 23863 11063 23897
rect 11063 23863 11097 23897
rect 11097 23863 11106 23897
rect 11054 23854 11106 23863
rect 11054 23737 11106 23746
rect 11054 23703 11063 23737
rect 11063 23703 11097 23737
rect 11097 23703 11106 23737
rect 11054 23694 11106 23703
rect 11054 23577 11106 23586
rect 11054 23543 11063 23577
rect 11063 23543 11097 23577
rect 11097 23543 11106 23577
rect 11054 23534 11106 23543
rect 11054 23417 11106 23426
rect 11054 23383 11063 23417
rect 11063 23383 11097 23417
rect 11097 23383 11106 23417
rect 11054 23374 11106 23383
rect 11054 23257 11106 23266
rect 11054 23223 11063 23257
rect 11063 23223 11097 23257
rect 11097 23223 11106 23257
rect 11054 23214 11106 23223
rect 11054 23097 11106 23106
rect 11054 23063 11063 23097
rect 11063 23063 11097 23097
rect 11097 23063 11106 23097
rect 11054 23054 11106 23063
rect 11054 22937 11106 22946
rect 11054 22903 11063 22937
rect 11063 22903 11097 22937
rect 11097 22903 11106 22937
rect 11054 22894 11106 22903
rect 11054 22777 11106 22786
rect 11054 22743 11063 22777
rect 11063 22743 11097 22777
rect 11097 22743 11106 22777
rect 11054 22734 11106 22743
rect 11054 22617 11106 22626
rect 11054 22583 11063 22617
rect 11063 22583 11097 22617
rect 11097 22583 11106 22617
rect 11054 22574 11106 22583
rect 11054 22457 11106 22466
rect 11054 22423 11063 22457
rect 11063 22423 11097 22457
rect 11097 22423 11106 22457
rect 11054 22414 11106 22423
rect 11054 22297 11106 22306
rect 11054 22263 11063 22297
rect 11063 22263 11097 22297
rect 11097 22263 11106 22297
rect 11054 22254 11106 22263
rect 11054 22137 11106 22146
rect 11054 22103 11063 22137
rect 11063 22103 11097 22137
rect 11097 22103 11106 22137
rect 11054 22094 11106 22103
rect 11054 21817 11106 21826
rect 11054 21783 11063 21817
rect 11063 21783 11097 21817
rect 11097 21783 11106 21817
rect 11054 21774 11106 21783
rect 11054 21657 11106 21666
rect 11054 21623 11063 21657
rect 11063 21623 11097 21657
rect 11097 21623 11106 21657
rect 11054 21614 11106 21623
rect 11054 21497 11106 21506
rect 11054 21463 11063 21497
rect 11063 21463 11097 21497
rect 11097 21463 11106 21497
rect 11054 21454 11106 21463
rect 11054 21337 11106 21346
rect 11054 21303 11063 21337
rect 11063 21303 11097 21337
rect 11097 21303 11106 21337
rect 11054 21294 11106 21303
rect 11054 21177 11106 21186
rect 11054 21143 11063 21177
rect 11063 21143 11097 21177
rect 11097 21143 11106 21177
rect 11054 21134 11106 21143
rect 11054 21017 11106 21026
rect 11054 20983 11063 21017
rect 11063 20983 11097 21017
rect 11097 20983 11106 21017
rect 11054 20974 11106 20983
rect 11054 20857 11106 20866
rect 11054 20823 11063 20857
rect 11063 20823 11097 20857
rect 11097 20823 11106 20857
rect 11054 20814 11106 20823
rect 11054 20697 11106 20706
rect 11054 20663 11063 20697
rect 11063 20663 11097 20697
rect 11097 20663 11106 20697
rect 11054 20654 11106 20663
rect 11054 19897 11106 19906
rect 11054 19863 11063 19897
rect 11063 19863 11097 19897
rect 11097 19863 11106 19897
rect 11054 19854 11106 19863
rect 11054 19737 11106 19746
rect 11054 19703 11063 19737
rect 11063 19703 11097 19737
rect 11097 19703 11106 19737
rect 11054 19694 11106 19703
rect 11054 19577 11106 19586
rect 11054 19543 11063 19577
rect 11063 19543 11097 19577
rect 11097 19543 11106 19577
rect 11054 19534 11106 19543
rect 11054 19417 11106 19426
rect 11054 19383 11063 19417
rect 11063 19383 11097 19417
rect 11097 19383 11106 19417
rect 11054 19374 11106 19383
rect 11054 19257 11106 19266
rect 11054 19223 11063 19257
rect 11063 19223 11097 19257
rect 11097 19223 11106 19257
rect 11054 19214 11106 19223
rect 11054 19097 11106 19106
rect 11054 19063 11063 19097
rect 11063 19063 11097 19097
rect 11097 19063 11106 19097
rect 11054 19054 11106 19063
rect 11054 18937 11106 18946
rect 11054 18903 11063 18937
rect 11063 18903 11097 18937
rect 11097 18903 11106 18937
rect 11054 18894 11106 18903
rect 11054 18777 11106 18786
rect 11054 18743 11063 18777
rect 11063 18743 11097 18777
rect 11097 18743 11106 18777
rect 11054 18734 11106 18743
rect 11054 17977 11106 17986
rect 11054 17943 11063 17977
rect 11063 17943 11097 17977
rect 11097 17943 11106 17977
rect 11054 17934 11106 17943
rect 11054 17817 11106 17826
rect 11054 17783 11063 17817
rect 11063 17783 11097 17817
rect 11097 17783 11106 17817
rect 11054 17774 11106 17783
rect 11054 17657 11106 17666
rect 11054 17623 11063 17657
rect 11063 17623 11097 17657
rect 11097 17623 11106 17657
rect 11054 17614 11106 17623
rect 11054 17497 11106 17506
rect 11054 17463 11063 17497
rect 11063 17463 11097 17497
rect 11097 17463 11106 17497
rect 11054 17454 11106 17463
rect 11054 17337 11106 17346
rect 11054 17303 11063 17337
rect 11063 17303 11097 17337
rect 11097 17303 11106 17337
rect 11054 17294 11106 17303
rect 11054 17177 11106 17186
rect 11054 17143 11063 17177
rect 11063 17143 11097 17177
rect 11097 17143 11106 17177
rect 11054 17134 11106 17143
rect 11054 17017 11106 17026
rect 11054 16983 11063 17017
rect 11063 16983 11097 17017
rect 11097 16983 11106 17017
rect 11054 16974 11106 16983
rect 11054 16857 11106 16866
rect 11054 16823 11063 16857
rect 11063 16823 11097 16857
rect 11097 16823 11106 16857
rect 11054 16814 11106 16823
rect 11054 16537 11106 16546
rect 11054 16503 11063 16537
rect 11063 16503 11097 16537
rect 11097 16503 11106 16537
rect 11054 16494 11106 16503
rect 11054 16377 11106 16386
rect 11054 16343 11063 16377
rect 11063 16343 11097 16377
rect 11097 16343 11106 16377
rect 11054 16334 11106 16343
rect 11054 16217 11106 16226
rect 11054 16183 11063 16217
rect 11063 16183 11097 16217
rect 11097 16183 11106 16217
rect 11054 16174 11106 16183
rect 11054 16057 11106 16066
rect 11054 16023 11063 16057
rect 11063 16023 11097 16057
rect 11097 16023 11106 16057
rect 11054 16014 11106 16023
rect 11054 15897 11106 15906
rect 11054 15863 11063 15897
rect 11063 15863 11097 15897
rect 11097 15863 11106 15897
rect 11054 15854 11106 15863
rect 11054 15737 11106 15746
rect 11054 15703 11063 15737
rect 11063 15703 11097 15737
rect 11097 15703 11106 15737
rect 11054 15694 11106 15703
rect 11054 15577 11106 15586
rect 11054 15543 11063 15577
rect 11063 15543 11097 15577
rect 11097 15543 11106 15577
rect 11054 15534 11106 15543
rect 11054 15417 11106 15426
rect 11054 15383 11063 15417
rect 11063 15383 11097 15417
rect 11097 15383 11106 15417
rect 11054 15374 11106 15383
rect 11054 15257 11106 15266
rect 11054 15223 11063 15257
rect 11063 15223 11097 15257
rect 11097 15223 11106 15257
rect 11054 15214 11106 15223
rect 11054 15097 11106 15106
rect 11054 15063 11063 15097
rect 11063 15063 11097 15097
rect 11097 15063 11106 15097
rect 11054 15054 11106 15063
rect 11054 14937 11106 14946
rect 11054 14903 11063 14937
rect 11063 14903 11097 14937
rect 11097 14903 11106 14937
rect 11054 14894 11106 14903
rect 11054 14777 11106 14786
rect 11054 14743 11063 14777
rect 11063 14743 11097 14777
rect 11097 14743 11106 14777
rect 11054 14734 11106 14743
rect 11054 14617 11106 14626
rect 11054 14583 11063 14617
rect 11063 14583 11097 14617
rect 11097 14583 11106 14617
rect 11054 14574 11106 14583
rect 11054 14457 11106 14466
rect 11054 14423 11063 14457
rect 11063 14423 11097 14457
rect 11097 14423 11106 14457
rect 11054 14414 11106 14423
rect 11054 14297 11106 14306
rect 11054 14263 11063 14297
rect 11063 14263 11097 14297
rect 11097 14263 11106 14297
rect 11054 14254 11106 14263
rect 11054 14137 11106 14146
rect 11054 14103 11063 14137
rect 11063 14103 11097 14137
rect 11097 14103 11106 14137
rect 11054 14094 11106 14103
rect 11054 13977 11106 13986
rect 11054 13943 11063 13977
rect 11063 13943 11097 13977
rect 11097 13943 11106 13977
rect 11054 13934 11106 13943
rect 11054 13657 11106 13666
rect 11054 13623 11063 13657
rect 11063 13623 11097 13657
rect 11097 13623 11106 13657
rect 11054 13614 11106 13623
rect 11054 13497 11106 13506
rect 11054 13463 11063 13497
rect 11063 13463 11097 13497
rect 11097 13463 11106 13497
rect 11054 13454 11106 13463
rect 11054 13337 11106 13346
rect 11054 13303 11063 13337
rect 11063 13303 11097 13337
rect 11097 13303 11106 13337
rect 11054 13294 11106 13303
rect 11054 13177 11106 13186
rect 11054 13143 11063 13177
rect 11063 13143 11097 13177
rect 11097 13143 11106 13177
rect 11054 13134 11106 13143
rect 11054 13017 11106 13026
rect 11054 12983 11063 13017
rect 11063 12983 11097 13017
rect 11097 12983 11106 13017
rect 11054 12974 11106 12983
rect 11054 12857 11106 12866
rect 11054 12823 11063 12857
rect 11063 12823 11097 12857
rect 11097 12823 11106 12857
rect 11054 12814 11106 12823
rect 11054 12697 11106 12706
rect 11054 12663 11063 12697
rect 11063 12663 11097 12697
rect 11097 12663 11106 12697
rect 11054 12654 11106 12663
rect 11054 12537 11106 12546
rect 11054 12503 11063 12537
rect 11063 12503 11097 12537
rect 11097 12503 11106 12537
rect 11054 12494 11106 12503
rect 11054 11737 11106 11746
rect 11054 11703 11063 11737
rect 11063 11703 11097 11737
rect 11097 11703 11106 11737
rect 11054 11694 11106 11703
rect 11054 11577 11106 11586
rect 11054 11543 11063 11577
rect 11063 11543 11097 11577
rect 11097 11543 11106 11577
rect 11054 11534 11106 11543
rect 11054 11417 11106 11426
rect 11054 11383 11063 11417
rect 11063 11383 11097 11417
rect 11097 11383 11106 11417
rect 11054 11374 11106 11383
rect 11054 11257 11106 11266
rect 11054 11223 11063 11257
rect 11063 11223 11097 11257
rect 11097 11223 11106 11257
rect 11054 11214 11106 11223
rect 11054 11097 11106 11106
rect 11054 11063 11063 11097
rect 11063 11063 11097 11097
rect 11097 11063 11106 11097
rect 11054 11054 11106 11063
rect 11054 10937 11106 10946
rect 11054 10903 11063 10937
rect 11063 10903 11097 10937
rect 11097 10903 11106 10937
rect 11054 10894 11106 10903
rect 11054 10777 11106 10786
rect 11054 10743 11063 10777
rect 11063 10743 11097 10777
rect 11097 10743 11106 10777
rect 11054 10734 11106 10743
rect 11054 10617 11106 10626
rect 11054 10583 11063 10617
rect 11063 10583 11097 10617
rect 11097 10583 11106 10617
rect 11054 10574 11106 10583
rect 11054 10457 11106 10466
rect 11054 10423 11063 10457
rect 11063 10423 11097 10457
rect 11097 10423 11106 10457
rect 11054 10414 11106 10423
rect 11054 10297 11106 10306
rect 11054 10263 11063 10297
rect 11063 10263 11097 10297
rect 11097 10263 11106 10297
rect 11054 10254 11106 10263
rect 11054 10137 11106 10146
rect 11054 10103 11063 10137
rect 11063 10103 11097 10137
rect 11097 10103 11106 10137
rect 11054 10094 11106 10103
rect 11054 9977 11106 9986
rect 11054 9943 11063 9977
rect 11063 9943 11097 9977
rect 11097 9943 11106 9977
rect 11054 9934 11106 9943
rect 11054 9817 11106 9826
rect 11054 9783 11063 9817
rect 11063 9783 11097 9817
rect 11097 9783 11106 9817
rect 11054 9774 11106 9783
rect 11054 9497 11106 9506
rect 11054 9463 11063 9497
rect 11063 9463 11097 9497
rect 11097 9463 11106 9497
rect 11054 9454 11106 9463
rect 11054 9337 11106 9346
rect 11054 9303 11063 9337
rect 11063 9303 11097 9337
rect 11097 9303 11106 9337
rect 11054 9294 11106 9303
rect 11054 9017 11106 9026
rect 11054 8983 11063 9017
rect 11063 8983 11097 9017
rect 11097 8983 11106 9017
rect 11054 8974 11106 8983
rect 11054 8857 11106 8866
rect 11054 8823 11063 8857
rect 11063 8823 11097 8857
rect 11097 8823 11106 8857
rect 11054 8814 11106 8823
rect 11054 8697 11106 8706
rect 11054 8663 11063 8697
rect 11063 8663 11097 8697
rect 11097 8663 11106 8697
rect 11054 8654 11106 8663
rect 11054 8537 11106 8546
rect 11054 8503 11063 8537
rect 11063 8503 11097 8537
rect 11097 8503 11106 8537
rect 11054 8494 11106 8503
rect 11054 8377 11106 8386
rect 11054 8343 11063 8377
rect 11063 8343 11097 8377
rect 11097 8343 11106 8377
rect 11054 8334 11106 8343
rect 11054 8217 11106 8226
rect 11054 8183 11063 8217
rect 11063 8183 11097 8217
rect 11097 8183 11106 8217
rect 11054 8174 11106 8183
rect 11054 8057 11106 8066
rect 11054 8023 11063 8057
rect 11063 8023 11097 8057
rect 11097 8023 11106 8057
rect 11054 8014 11106 8023
rect 11054 7897 11106 7906
rect 11054 7863 11063 7897
rect 11063 7863 11097 7897
rect 11097 7863 11106 7897
rect 11054 7854 11106 7863
rect 11054 7737 11106 7746
rect 11054 7703 11063 7737
rect 11063 7703 11097 7737
rect 11097 7703 11106 7737
rect 11054 7694 11106 7703
rect 11054 7417 11106 7426
rect 11054 7383 11063 7417
rect 11063 7383 11097 7417
rect 11097 7383 11106 7417
rect 11054 7374 11106 7383
rect 11054 7257 11106 7266
rect 11054 7223 11063 7257
rect 11063 7223 11097 7257
rect 11097 7223 11106 7257
rect 11054 7214 11106 7223
rect 11054 6937 11106 6946
rect 11054 6903 11063 6937
rect 11063 6903 11097 6937
rect 11097 6903 11106 6937
rect 11054 6894 11106 6903
rect 11054 6777 11106 6786
rect 11054 6743 11063 6777
rect 11063 6743 11097 6777
rect 11097 6743 11106 6777
rect 11054 6734 11106 6743
rect 11054 6457 11106 6466
rect 11054 6423 11063 6457
rect 11063 6423 11097 6457
rect 11097 6423 11106 6457
rect 11054 6414 11106 6423
rect 11054 6297 11106 6306
rect 11054 6263 11063 6297
rect 11063 6263 11097 6297
rect 11097 6263 11106 6297
rect 11054 6254 11106 6263
rect 11054 6137 11106 6146
rect 11054 6103 11063 6137
rect 11063 6103 11097 6137
rect 11097 6103 11106 6137
rect 11054 6094 11106 6103
rect 11054 5977 11106 5986
rect 11054 5943 11063 5977
rect 11063 5943 11097 5977
rect 11097 5943 11106 5977
rect 11054 5934 11106 5943
rect 11054 5817 11106 5826
rect 11054 5783 11063 5817
rect 11063 5783 11097 5817
rect 11097 5783 11106 5817
rect 11054 5774 11106 5783
rect 11054 5657 11106 5666
rect 11054 5623 11063 5657
rect 11063 5623 11097 5657
rect 11097 5623 11106 5657
rect 11054 5614 11106 5623
rect 11054 5497 11106 5506
rect 11054 5463 11063 5497
rect 11063 5463 11097 5497
rect 11097 5463 11106 5497
rect 11054 5454 11106 5463
rect 11054 5337 11106 5346
rect 11054 5303 11063 5337
rect 11063 5303 11097 5337
rect 11097 5303 11106 5337
rect 11054 5294 11106 5303
rect 11054 5177 11106 5186
rect 11054 5143 11063 5177
rect 11063 5143 11097 5177
rect 11097 5143 11106 5177
rect 11054 5134 11106 5143
rect 11054 5017 11106 5026
rect 11054 4983 11063 5017
rect 11063 4983 11097 5017
rect 11097 4983 11106 5017
rect 11054 4974 11106 4983
rect 11054 4857 11106 4866
rect 11054 4823 11063 4857
rect 11063 4823 11097 4857
rect 11097 4823 11106 4857
rect 11054 4814 11106 4823
rect 11054 4697 11106 4706
rect 11054 4663 11063 4697
rect 11063 4663 11097 4697
rect 11097 4663 11106 4697
rect 11054 4654 11106 4663
rect 11054 4537 11106 4546
rect 11054 4503 11063 4537
rect 11063 4503 11097 4537
rect 11097 4503 11106 4537
rect 11054 4494 11106 4503
rect 11054 4377 11106 4386
rect 11054 4343 11063 4377
rect 11063 4343 11097 4377
rect 11097 4343 11106 4377
rect 11054 4334 11106 4343
rect 11054 4217 11106 4226
rect 11054 4183 11063 4217
rect 11063 4183 11097 4217
rect 11097 4183 11106 4217
rect 11054 4174 11106 4183
rect 11054 4057 11106 4066
rect 11054 4023 11063 4057
rect 11063 4023 11097 4057
rect 11097 4023 11106 4057
rect 11054 4014 11106 4023
rect 11054 3897 11106 3906
rect 11054 3863 11063 3897
rect 11063 3863 11097 3897
rect 11097 3863 11106 3897
rect 11054 3854 11106 3863
rect 11054 3417 11106 3426
rect 11054 3383 11063 3417
rect 11063 3383 11097 3417
rect 11097 3383 11106 3417
rect 11054 3374 11106 3383
rect 11054 3257 11106 3266
rect 11054 3223 11063 3257
rect 11063 3223 11097 3257
rect 11097 3223 11106 3257
rect 11054 3214 11106 3223
rect 11054 3097 11106 3106
rect 11054 3063 11063 3097
rect 11063 3063 11097 3097
rect 11097 3063 11106 3097
rect 11054 3054 11106 3063
rect 11054 2937 11106 2946
rect 11054 2903 11063 2937
rect 11063 2903 11097 2937
rect 11097 2903 11106 2937
rect 11054 2894 11106 2903
rect 11054 2777 11106 2786
rect 11054 2743 11063 2777
rect 11063 2743 11097 2777
rect 11097 2743 11106 2777
rect 11054 2734 11106 2743
rect 11054 2617 11106 2626
rect 11054 2583 11063 2617
rect 11063 2583 11097 2617
rect 11097 2583 11106 2617
rect 11054 2574 11106 2583
rect 11054 2457 11106 2466
rect 11054 2423 11063 2457
rect 11063 2423 11097 2457
rect 11097 2423 11106 2457
rect 11054 2414 11106 2423
rect 11054 2297 11106 2306
rect 11054 2263 11063 2297
rect 11063 2263 11097 2297
rect 11097 2263 11106 2297
rect 11054 2254 11106 2263
rect 11054 2137 11106 2146
rect 11054 2103 11063 2137
rect 11063 2103 11097 2137
rect 11097 2103 11106 2137
rect 11054 2094 11106 2103
rect 11054 1977 11106 1986
rect 11054 1943 11063 1977
rect 11063 1943 11097 1977
rect 11097 1943 11106 1977
rect 11054 1934 11106 1943
rect 11054 1657 11106 1666
rect 11054 1623 11063 1657
rect 11063 1623 11097 1657
rect 11097 1623 11106 1657
rect 11054 1614 11106 1623
rect 11054 1497 11106 1506
rect 11054 1463 11063 1497
rect 11063 1463 11097 1497
rect 11097 1463 11106 1497
rect 11054 1454 11106 1463
rect 11054 1337 11106 1346
rect 11054 1303 11063 1337
rect 11063 1303 11097 1337
rect 11097 1303 11106 1337
rect 11054 1294 11106 1303
rect 11054 1177 11106 1186
rect 11054 1143 11063 1177
rect 11063 1143 11097 1177
rect 11097 1143 11106 1177
rect 11054 1134 11106 1143
rect 11054 1017 11106 1026
rect 11054 983 11063 1017
rect 11063 983 11097 1017
rect 11097 983 11106 1017
rect 11054 974 11106 983
rect 11054 537 11106 546
rect 11054 503 11063 537
rect 11063 503 11097 537
rect 11097 503 11106 537
rect 11054 494 11106 503
rect 11054 377 11106 386
rect 11054 343 11063 377
rect 11063 343 11097 377
rect 11097 343 11106 377
rect 11054 334 11106 343
rect 11054 217 11106 226
rect 11054 183 11063 217
rect 11063 183 11097 217
rect 11097 183 11106 217
rect 11054 174 11106 183
rect 11054 57 11106 66
rect 11054 23 11063 57
rect 11063 23 11097 57
rect 11097 23 11106 57
rect 11054 14 11106 23
rect 11374 31417 11426 31426
rect 11374 31383 11383 31417
rect 11383 31383 11417 31417
rect 11417 31383 11426 31417
rect 11374 31374 11426 31383
rect 11374 31257 11426 31266
rect 11374 31223 11383 31257
rect 11383 31223 11417 31257
rect 11417 31223 11426 31257
rect 11374 31214 11426 31223
rect 11374 31097 11426 31106
rect 11374 31063 11383 31097
rect 11383 31063 11417 31097
rect 11417 31063 11426 31097
rect 11374 31054 11426 31063
rect 11374 30937 11426 30946
rect 11374 30903 11383 30937
rect 11383 30903 11417 30937
rect 11417 30903 11426 30937
rect 11374 30894 11426 30903
rect 11374 30777 11426 30786
rect 11374 30743 11383 30777
rect 11383 30743 11417 30777
rect 11417 30743 11426 30777
rect 11374 30734 11426 30743
rect 11374 30617 11426 30626
rect 11374 30583 11383 30617
rect 11383 30583 11417 30617
rect 11417 30583 11426 30617
rect 11374 30574 11426 30583
rect 11374 30457 11426 30466
rect 11374 30423 11383 30457
rect 11383 30423 11417 30457
rect 11417 30423 11426 30457
rect 11374 30414 11426 30423
rect 11374 30297 11426 30306
rect 11374 30263 11383 30297
rect 11383 30263 11417 30297
rect 11417 30263 11426 30297
rect 11374 30254 11426 30263
rect 11374 29977 11426 29986
rect 11374 29943 11383 29977
rect 11383 29943 11417 29977
rect 11417 29943 11426 29977
rect 11374 29934 11426 29943
rect 11374 29817 11426 29826
rect 11374 29783 11383 29817
rect 11383 29783 11417 29817
rect 11417 29783 11426 29817
rect 11374 29774 11426 29783
rect 11374 29657 11426 29666
rect 11374 29623 11383 29657
rect 11383 29623 11417 29657
rect 11417 29623 11426 29657
rect 11374 29614 11426 29623
rect 11374 29497 11426 29506
rect 11374 29463 11383 29497
rect 11383 29463 11417 29497
rect 11417 29463 11426 29497
rect 11374 29454 11426 29463
rect 11374 29337 11426 29346
rect 11374 29303 11383 29337
rect 11383 29303 11417 29337
rect 11417 29303 11426 29337
rect 11374 29294 11426 29303
rect 11374 29177 11426 29186
rect 11374 29143 11383 29177
rect 11383 29143 11417 29177
rect 11417 29143 11426 29177
rect 11374 29134 11426 29143
rect 11374 29017 11426 29026
rect 11374 28983 11383 29017
rect 11383 28983 11417 29017
rect 11417 28983 11426 29017
rect 11374 28974 11426 28983
rect 11374 28857 11426 28866
rect 11374 28823 11383 28857
rect 11383 28823 11417 28857
rect 11417 28823 11426 28857
rect 11374 28814 11426 28823
rect 11374 28057 11426 28066
rect 11374 28023 11383 28057
rect 11383 28023 11417 28057
rect 11417 28023 11426 28057
rect 11374 28014 11426 28023
rect 11374 27897 11426 27906
rect 11374 27863 11383 27897
rect 11383 27863 11417 27897
rect 11417 27863 11426 27897
rect 11374 27854 11426 27863
rect 11374 27737 11426 27746
rect 11374 27703 11383 27737
rect 11383 27703 11417 27737
rect 11417 27703 11426 27737
rect 11374 27694 11426 27703
rect 11374 27577 11426 27586
rect 11374 27543 11383 27577
rect 11383 27543 11417 27577
rect 11417 27543 11426 27577
rect 11374 27534 11426 27543
rect 11374 27417 11426 27426
rect 11374 27383 11383 27417
rect 11383 27383 11417 27417
rect 11417 27383 11426 27417
rect 11374 27374 11426 27383
rect 11374 27257 11426 27266
rect 11374 27223 11383 27257
rect 11383 27223 11417 27257
rect 11417 27223 11426 27257
rect 11374 27214 11426 27223
rect 11374 27097 11426 27106
rect 11374 27063 11383 27097
rect 11383 27063 11417 27097
rect 11417 27063 11426 27097
rect 11374 27054 11426 27063
rect 11374 26937 11426 26946
rect 11374 26903 11383 26937
rect 11383 26903 11417 26937
rect 11417 26903 11426 26937
rect 11374 26894 11426 26903
rect 11374 26137 11426 26146
rect 11374 26103 11383 26137
rect 11383 26103 11417 26137
rect 11417 26103 11426 26137
rect 11374 26094 11426 26103
rect 11374 25977 11426 25986
rect 11374 25943 11383 25977
rect 11383 25943 11417 25977
rect 11417 25943 11426 25977
rect 11374 25934 11426 25943
rect 11374 25817 11426 25826
rect 11374 25783 11383 25817
rect 11383 25783 11417 25817
rect 11417 25783 11426 25817
rect 11374 25774 11426 25783
rect 11374 25657 11426 25666
rect 11374 25623 11383 25657
rect 11383 25623 11417 25657
rect 11417 25623 11426 25657
rect 11374 25614 11426 25623
rect 11374 25497 11426 25506
rect 11374 25463 11383 25497
rect 11383 25463 11417 25497
rect 11417 25463 11426 25497
rect 11374 25454 11426 25463
rect 11374 25337 11426 25346
rect 11374 25303 11383 25337
rect 11383 25303 11417 25337
rect 11417 25303 11426 25337
rect 11374 25294 11426 25303
rect 11374 25177 11426 25186
rect 11374 25143 11383 25177
rect 11383 25143 11417 25177
rect 11417 25143 11426 25177
rect 11374 25134 11426 25143
rect 11374 25017 11426 25026
rect 11374 24983 11383 25017
rect 11383 24983 11417 25017
rect 11417 24983 11426 25017
rect 11374 24974 11426 24983
rect 11374 24697 11426 24706
rect 11374 24663 11383 24697
rect 11383 24663 11417 24697
rect 11417 24663 11426 24697
rect 11374 24654 11426 24663
rect 11374 24537 11426 24546
rect 11374 24503 11383 24537
rect 11383 24503 11417 24537
rect 11417 24503 11426 24537
rect 11374 24494 11426 24503
rect 11374 24377 11426 24386
rect 11374 24343 11383 24377
rect 11383 24343 11417 24377
rect 11417 24343 11426 24377
rect 11374 24334 11426 24343
rect 11374 24217 11426 24226
rect 11374 24183 11383 24217
rect 11383 24183 11417 24217
rect 11417 24183 11426 24217
rect 11374 24174 11426 24183
rect 11374 24057 11426 24066
rect 11374 24023 11383 24057
rect 11383 24023 11417 24057
rect 11417 24023 11426 24057
rect 11374 24014 11426 24023
rect 11374 23897 11426 23906
rect 11374 23863 11383 23897
rect 11383 23863 11417 23897
rect 11417 23863 11426 23897
rect 11374 23854 11426 23863
rect 11374 23737 11426 23746
rect 11374 23703 11383 23737
rect 11383 23703 11417 23737
rect 11417 23703 11426 23737
rect 11374 23694 11426 23703
rect 11374 23577 11426 23586
rect 11374 23543 11383 23577
rect 11383 23543 11417 23577
rect 11417 23543 11426 23577
rect 11374 23534 11426 23543
rect 11374 23417 11426 23426
rect 11374 23383 11383 23417
rect 11383 23383 11417 23417
rect 11417 23383 11426 23417
rect 11374 23374 11426 23383
rect 11374 23257 11426 23266
rect 11374 23223 11383 23257
rect 11383 23223 11417 23257
rect 11417 23223 11426 23257
rect 11374 23214 11426 23223
rect 11374 23097 11426 23106
rect 11374 23063 11383 23097
rect 11383 23063 11417 23097
rect 11417 23063 11426 23097
rect 11374 23054 11426 23063
rect 11374 22937 11426 22946
rect 11374 22903 11383 22937
rect 11383 22903 11417 22937
rect 11417 22903 11426 22937
rect 11374 22894 11426 22903
rect 11374 22777 11426 22786
rect 11374 22743 11383 22777
rect 11383 22743 11417 22777
rect 11417 22743 11426 22777
rect 11374 22734 11426 22743
rect 11374 22617 11426 22626
rect 11374 22583 11383 22617
rect 11383 22583 11417 22617
rect 11417 22583 11426 22617
rect 11374 22574 11426 22583
rect 11374 22457 11426 22466
rect 11374 22423 11383 22457
rect 11383 22423 11417 22457
rect 11417 22423 11426 22457
rect 11374 22414 11426 22423
rect 11374 22297 11426 22306
rect 11374 22263 11383 22297
rect 11383 22263 11417 22297
rect 11417 22263 11426 22297
rect 11374 22254 11426 22263
rect 11374 22137 11426 22146
rect 11374 22103 11383 22137
rect 11383 22103 11417 22137
rect 11417 22103 11426 22137
rect 11374 22094 11426 22103
rect 11374 21817 11426 21826
rect 11374 21783 11383 21817
rect 11383 21783 11417 21817
rect 11417 21783 11426 21817
rect 11374 21774 11426 21783
rect 11374 21657 11426 21666
rect 11374 21623 11383 21657
rect 11383 21623 11417 21657
rect 11417 21623 11426 21657
rect 11374 21614 11426 21623
rect 11374 21497 11426 21506
rect 11374 21463 11383 21497
rect 11383 21463 11417 21497
rect 11417 21463 11426 21497
rect 11374 21454 11426 21463
rect 11374 21337 11426 21346
rect 11374 21303 11383 21337
rect 11383 21303 11417 21337
rect 11417 21303 11426 21337
rect 11374 21294 11426 21303
rect 11374 21177 11426 21186
rect 11374 21143 11383 21177
rect 11383 21143 11417 21177
rect 11417 21143 11426 21177
rect 11374 21134 11426 21143
rect 11374 21017 11426 21026
rect 11374 20983 11383 21017
rect 11383 20983 11417 21017
rect 11417 20983 11426 21017
rect 11374 20974 11426 20983
rect 11374 20857 11426 20866
rect 11374 20823 11383 20857
rect 11383 20823 11417 20857
rect 11417 20823 11426 20857
rect 11374 20814 11426 20823
rect 11374 20697 11426 20706
rect 11374 20663 11383 20697
rect 11383 20663 11417 20697
rect 11417 20663 11426 20697
rect 11374 20654 11426 20663
rect 11374 19897 11426 19906
rect 11374 19863 11383 19897
rect 11383 19863 11417 19897
rect 11417 19863 11426 19897
rect 11374 19854 11426 19863
rect 11374 19737 11426 19746
rect 11374 19703 11383 19737
rect 11383 19703 11417 19737
rect 11417 19703 11426 19737
rect 11374 19694 11426 19703
rect 11374 19577 11426 19586
rect 11374 19543 11383 19577
rect 11383 19543 11417 19577
rect 11417 19543 11426 19577
rect 11374 19534 11426 19543
rect 11374 19417 11426 19426
rect 11374 19383 11383 19417
rect 11383 19383 11417 19417
rect 11417 19383 11426 19417
rect 11374 19374 11426 19383
rect 11374 19257 11426 19266
rect 11374 19223 11383 19257
rect 11383 19223 11417 19257
rect 11417 19223 11426 19257
rect 11374 19214 11426 19223
rect 11374 19097 11426 19106
rect 11374 19063 11383 19097
rect 11383 19063 11417 19097
rect 11417 19063 11426 19097
rect 11374 19054 11426 19063
rect 11374 18937 11426 18946
rect 11374 18903 11383 18937
rect 11383 18903 11417 18937
rect 11417 18903 11426 18937
rect 11374 18894 11426 18903
rect 11374 18777 11426 18786
rect 11374 18743 11383 18777
rect 11383 18743 11417 18777
rect 11417 18743 11426 18777
rect 11374 18734 11426 18743
rect 11374 17977 11426 17986
rect 11374 17943 11383 17977
rect 11383 17943 11417 17977
rect 11417 17943 11426 17977
rect 11374 17934 11426 17943
rect 11374 17817 11426 17826
rect 11374 17783 11383 17817
rect 11383 17783 11417 17817
rect 11417 17783 11426 17817
rect 11374 17774 11426 17783
rect 11374 17657 11426 17666
rect 11374 17623 11383 17657
rect 11383 17623 11417 17657
rect 11417 17623 11426 17657
rect 11374 17614 11426 17623
rect 11374 17497 11426 17506
rect 11374 17463 11383 17497
rect 11383 17463 11417 17497
rect 11417 17463 11426 17497
rect 11374 17454 11426 17463
rect 11374 17337 11426 17346
rect 11374 17303 11383 17337
rect 11383 17303 11417 17337
rect 11417 17303 11426 17337
rect 11374 17294 11426 17303
rect 11374 17177 11426 17186
rect 11374 17143 11383 17177
rect 11383 17143 11417 17177
rect 11417 17143 11426 17177
rect 11374 17134 11426 17143
rect 11374 17017 11426 17026
rect 11374 16983 11383 17017
rect 11383 16983 11417 17017
rect 11417 16983 11426 17017
rect 11374 16974 11426 16983
rect 11374 16857 11426 16866
rect 11374 16823 11383 16857
rect 11383 16823 11417 16857
rect 11417 16823 11426 16857
rect 11374 16814 11426 16823
rect 11374 16537 11426 16546
rect 11374 16503 11383 16537
rect 11383 16503 11417 16537
rect 11417 16503 11426 16537
rect 11374 16494 11426 16503
rect 11374 16377 11426 16386
rect 11374 16343 11383 16377
rect 11383 16343 11417 16377
rect 11417 16343 11426 16377
rect 11374 16334 11426 16343
rect 11374 16217 11426 16226
rect 11374 16183 11383 16217
rect 11383 16183 11417 16217
rect 11417 16183 11426 16217
rect 11374 16174 11426 16183
rect 11374 16057 11426 16066
rect 11374 16023 11383 16057
rect 11383 16023 11417 16057
rect 11417 16023 11426 16057
rect 11374 16014 11426 16023
rect 11374 15897 11426 15906
rect 11374 15863 11383 15897
rect 11383 15863 11417 15897
rect 11417 15863 11426 15897
rect 11374 15854 11426 15863
rect 11374 15737 11426 15746
rect 11374 15703 11383 15737
rect 11383 15703 11417 15737
rect 11417 15703 11426 15737
rect 11374 15694 11426 15703
rect 11374 15577 11426 15586
rect 11374 15543 11383 15577
rect 11383 15543 11417 15577
rect 11417 15543 11426 15577
rect 11374 15534 11426 15543
rect 11374 15417 11426 15426
rect 11374 15383 11383 15417
rect 11383 15383 11417 15417
rect 11417 15383 11426 15417
rect 11374 15374 11426 15383
rect 11374 15257 11426 15266
rect 11374 15223 11383 15257
rect 11383 15223 11417 15257
rect 11417 15223 11426 15257
rect 11374 15214 11426 15223
rect 11374 15097 11426 15106
rect 11374 15063 11383 15097
rect 11383 15063 11417 15097
rect 11417 15063 11426 15097
rect 11374 15054 11426 15063
rect 11374 14937 11426 14946
rect 11374 14903 11383 14937
rect 11383 14903 11417 14937
rect 11417 14903 11426 14937
rect 11374 14894 11426 14903
rect 11374 14777 11426 14786
rect 11374 14743 11383 14777
rect 11383 14743 11417 14777
rect 11417 14743 11426 14777
rect 11374 14734 11426 14743
rect 11374 14617 11426 14626
rect 11374 14583 11383 14617
rect 11383 14583 11417 14617
rect 11417 14583 11426 14617
rect 11374 14574 11426 14583
rect 11374 14457 11426 14466
rect 11374 14423 11383 14457
rect 11383 14423 11417 14457
rect 11417 14423 11426 14457
rect 11374 14414 11426 14423
rect 11374 14297 11426 14306
rect 11374 14263 11383 14297
rect 11383 14263 11417 14297
rect 11417 14263 11426 14297
rect 11374 14254 11426 14263
rect 11374 14137 11426 14146
rect 11374 14103 11383 14137
rect 11383 14103 11417 14137
rect 11417 14103 11426 14137
rect 11374 14094 11426 14103
rect 11374 13977 11426 13986
rect 11374 13943 11383 13977
rect 11383 13943 11417 13977
rect 11417 13943 11426 13977
rect 11374 13934 11426 13943
rect 11374 13657 11426 13666
rect 11374 13623 11383 13657
rect 11383 13623 11417 13657
rect 11417 13623 11426 13657
rect 11374 13614 11426 13623
rect 11374 13497 11426 13506
rect 11374 13463 11383 13497
rect 11383 13463 11417 13497
rect 11417 13463 11426 13497
rect 11374 13454 11426 13463
rect 11374 13337 11426 13346
rect 11374 13303 11383 13337
rect 11383 13303 11417 13337
rect 11417 13303 11426 13337
rect 11374 13294 11426 13303
rect 11374 13177 11426 13186
rect 11374 13143 11383 13177
rect 11383 13143 11417 13177
rect 11417 13143 11426 13177
rect 11374 13134 11426 13143
rect 11374 13017 11426 13026
rect 11374 12983 11383 13017
rect 11383 12983 11417 13017
rect 11417 12983 11426 13017
rect 11374 12974 11426 12983
rect 11374 12857 11426 12866
rect 11374 12823 11383 12857
rect 11383 12823 11417 12857
rect 11417 12823 11426 12857
rect 11374 12814 11426 12823
rect 11374 12697 11426 12706
rect 11374 12663 11383 12697
rect 11383 12663 11417 12697
rect 11417 12663 11426 12697
rect 11374 12654 11426 12663
rect 11374 12537 11426 12546
rect 11374 12503 11383 12537
rect 11383 12503 11417 12537
rect 11417 12503 11426 12537
rect 11374 12494 11426 12503
rect 11374 11737 11426 11746
rect 11374 11703 11383 11737
rect 11383 11703 11417 11737
rect 11417 11703 11426 11737
rect 11374 11694 11426 11703
rect 11374 11577 11426 11586
rect 11374 11543 11383 11577
rect 11383 11543 11417 11577
rect 11417 11543 11426 11577
rect 11374 11534 11426 11543
rect 11374 11417 11426 11426
rect 11374 11383 11383 11417
rect 11383 11383 11417 11417
rect 11417 11383 11426 11417
rect 11374 11374 11426 11383
rect 11374 11257 11426 11266
rect 11374 11223 11383 11257
rect 11383 11223 11417 11257
rect 11417 11223 11426 11257
rect 11374 11214 11426 11223
rect 11374 11097 11426 11106
rect 11374 11063 11383 11097
rect 11383 11063 11417 11097
rect 11417 11063 11426 11097
rect 11374 11054 11426 11063
rect 11374 10937 11426 10946
rect 11374 10903 11383 10937
rect 11383 10903 11417 10937
rect 11417 10903 11426 10937
rect 11374 10894 11426 10903
rect 11374 10777 11426 10786
rect 11374 10743 11383 10777
rect 11383 10743 11417 10777
rect 11417 10743 11426 10777
rect 11374 10734 11426 10743
rect 11374 10617 11426 10626
rect 11374 10583 11383 10617
rect 11383 10583 11417 10617
rect 11417 10583 11426 10617
rect 11374 10574 11426 10583
rect 11374 10457 11426 10466
rect 11374 10423 11383 10457
rect 11383 10423 11417 10457
rect 11417 10423 11426 10457
rect 11374 10414 11426 10423
rect 11374 10297 11426 10306
rect 11374 10263 11383 10297
rect 11383 10263 11417 10297
rect 11417 10263 11426 10297
rect 11374 10254 11426 10263
rect 11374 10137 11426 10146
rect 11374 10103 11383 10137
rect 11383 10103 11417 10137
rect 11417 10103 11426 10137
rect 11374 10094 11426 10103
rect 11374 9977 11426 9986
rect 11374 9943 11383 9977
rect 11383 9943 11417 9977
rect 11417 9943 11426 9977
rect 11374 9934 11426 9943
rect 11374 9817 11426 9826
rect 11374 9783 11383 9817
rect 11383 9783 11417 9817
rect 11417 9783 11426 9817
rect 11374 9774 11426 9783
rect 11374 9497 11426 9506
rect 11374 9463 11383 9497
rect 11383 9463 11417 9497
rect 11417 9463 11426 9497
rect 11374 9454 11426 9463
rect 11374 9337 11426 9346
rect 11374 9303 11383 9337
rect 11383 9303 11417 9337
rect 11417 9303 11426 9337
rect 11374 9294 11426 9303
rect 11374 9017 11426 9026
rect 11374 8983 11383 9017
rect 11383 8983 11417 9017
rect 11417 8983 11426 9017
rect 11374 8974 11426 8983
rect 11374 8857 11426 8866
rect 11374 8823 11383 8857
rect 11383 8823 11417 8857
rect 11417 8823 11426 8857
rect 11374 8814 11426 8823
rect 11374 8697 11426 8706
rect 11374 8663 11383 8697
rect 11383 8663 11417 8697
rect 11417 8663 11426 8697
rect 11374 8654 11426 8663
rect 11374 8537 11426 8546
rect 11374 8503 11383 8537
rect 11383 8503 11417 8537
rect 11417 8503 11426 8537
rect 11374 8494 11426 8503
rect 11374 8377 11426 8386
rect 11374 8343 11383 8377
rect 11383 8343 11417 8377
rect 11417 8343 11426 8377
rect 11374 8334 11426 8343
rect 11374 8217 11426 8226
rect 11374 8183 11383 8217
rect 11383 8183 11417 8217
rect 11417 8183 11426 8217
rect 11374 8174 11426 8183
rect 11374 8057 11426 8066
rect 11374 8023 11383 8057
rect 11383 8023 11417 8057
rect 11417 8023 11426 8057
rect 11374 8014 11426 8023
rect 11374 7897 11426 7906
rect 11374 7863 11383 7897
rect 11383 7863 11417 7897
rect 11417 7863 11426 7897
rect 11374 7854 11426 7863
rect 11374 7737 11426 7746
rect 11374 7703 11383 7737
rect 11383 7703 11417 7737
rect 11417 7703 11426 7737
rect 11374 7694 11426 7703
rect 11374 7417 11426 7426
rect 11374 7383 11383 7417
rect 11383 7383 11417 7417
rect 11417 7383 11426 7417
rect 11374 7374 11426 7383
rect 11374 7257 11426 7266
rect 11374 7223 11383 7257
rect 11383 7223 11417 7257
rect 11417 7223 11426 7257
rect 11374 7214 11426 7223
rect 11374 6937 11426 6946
rect 11374 6903 11383 6937
rect 11383 6903 11417 6937
rect 11417 6903 11426 6937
rect 11374 6894 11426 6903
rect 11374 6777 11426 6786
rect 11374 6743 11383 6777
rect 11383 6743 11417 6777
rect 11417 6743 11426 6777
rect 11374 6734 11426 6743
rect 11374 6457 11426 6466
rect 11374 6423 11383 6457
rect 11383 6423 11417 6457
rect 11417 6423 11426 6457
rect 11374 6414 11426 6423
rect 11374 6297 11426 6306
rect 11374 6263 11383 6297
rect 11383 6263 11417 6297
rect 11417 6263 11426 6297
rect 11374 6254 11426 6263
rect 11374 6137 11426 6146
rect 11374 6103 11383 6137
rect 11383 6103 11417 6137
rect 11417 6103 11426 6137
rect 11374 6094 11426 6103
rect 11374 5977 11426 5986
rect 11374 5943 11383 5977
rect 11383 5943 11417 5977
rect 11417 5943 11426 5977
rect 11374 5934 11426 5943
rect 11374 5817 11426 5826
rect 11374 5783 11383 5817
rect 11383 5783 11417 5817
rect 11417 5783 11426 5817
rect 11374 5774 11426 5783
rect 11374 5657 11426 5666
rect 11374 5623 11383 5657
rect 11383 5623 11417 5657
rect 11417 5623 11426 5657
rect 11374 5614 11426 5623
rect 11374 5497 11426 5506
rect 11374 5463 11383 5497
rect 11383 5463 11417 5497
rect 11417 5463 11426 5497
rect 11374 5454 11426 5463
rect 11374 5337 11426 5346
rect 11374 5303 11383 5337
rect 11383 5303 11417 5337
rect 11417 5303 11426 5337
rect 11374 5294 11426 5303
rect 11374 5177 11426 5186
rect 11374 5143 11383 5177
rect 11383 5143 11417 5177
rect 11417 5143 11426 5177
rect 11374 5134 11426 5143
rect 11374 5017 11426 5026
rect 11374 4983 11383 5017
rect 11383 4983 11417 5017
rect 11417 4983 11426 5017
rect 11374 4974 11426 4983
rect 11374 4857 11426 4866
rect 11374 4823 11383 4857
rect 11383 4823 11417 4857
rect 11417 4823 11426 4857
rect 11374 4814 11426 4823
rect 11374 4697 11426 4706
rect 11374 4663 11383 4697
rect 11383 4663 11417 4697
rect 11417 4663 11426 4697
rect 11374 4654 11426 4663
rect 11374 4537 11426 4546
rect 11374 4503 11383 4537
rect 11383 4503 11417 4537
rect 11417 4503 11426 4537
rect 11374 4494 11426 4503
rect 11374 4377 11426 4386
rect 11374 4343 11383 4377
rect 11383 4343 11417 4377
rect 11417 4343 11426 4377
rect 11374 4334 11426 4343
rect 11374 4217 11426 4226
rect 11374 4183 11383 4217
rect 11383 4183 11417 4217
rect 11417 4183 11426 4217
rect 11374 4174 11426 4183
rect 11374 4057 11426 4066
rect 11374 4023 11383 4057
rect 11383 4023 11417 4057
rect 11417 4023 11426 4057
rect 11374 4014 11426 4023
rect 11374 3897 11426 3906
rect 11374 3863 11383 3897
rect 11383 3863 11417 3897
rect 11417 3863 11426 3897
rect 11374 3854 11426 3863
rect 11374 3417 11426 3426
rect 11374 3383 11383 3417
rect 11383 3383 11417 3417
rect 11417 3383 11426 3417
rect 11374 3374 11426 3383
rect 11374 3257 11426 3266
rect 11374 3223 11383 3257
rect 11383 3223 11417 3257
rect 11417 3223 11426 3257
rect 11374 3214 11426 3223
rect 11374 3097 11426 3106
rect 11374 3063 11383 3097
rect 11383 3063 11417 3097
rect 11417 3063 11426 3097
rect 11374 3054 11426 3063
rect 11374 2937 11426 2946
rect 11374 2903 11383 2937
rect 11383 2903 11417 2937
rect 11417 2903 11426 2937
rect 11374 2894 11426 2903
rect 11374 2777 11426 2786
rect 11374 2743 11383 2777
rect 11383 2743 11417 2777
rect 11417 2743 11426 2777
rect 11374 2734 11426 2743
rect 11374 2617 11426 2626
rect 11374 2583 11383 2617
rect 11383 2583 11417 2617
rect 11417 2583 11426 2617
rect 11374 2574 11426 2583
rect 11374 2457 11426 2466
rect 11374 2423 11383 2457
rect 11383 2423 11417 2457
rect 11417 2423 11426 2457
rect 11374 2414 11426 2423
rect 11374 2297 11426 2306
rect 11374 2263 11383 2297
rect 11383 2263 11417 2297
rect 11417 2263 11426 2297
rect 11374 2254 11426 2263
rect 11374 2137 11426 2146
rect 11374 2103 11383 2137
rect 11383 2103 11417 2137
rect 11417 2103 11426 2137
rect 11374 2094 11426 2103
rect 11374 1977 11426 1986
rect 11374 1943 11383 1977
rect 11383 1943 11417 1977
rect 11417 1943 11426 1977
rect 11374 1934 11426 1943
rect 11374 1657 11426 1666
rect 11374 1623 11383 1657
rect 11383 1623 11417 1657
rect 11417 1623 11426 1657
rect 11374 1614 11426 1623
rect 11374 1497 11426 1506
rect 11374 1463 11383 1497
rect 11383 1463 11417 1497
rect 11417 1463 11426 1497
rect 11374 1454 11426 1463
rect 11374 1337 11426 1346
rect 11374 1303 11383 1337
rect 11383 1303 11417 1337
rect 11417 1303 11426 1337
rect 11374 1294 11426 1303
rect 11374 1177 11426 1186
rect 11374 1143 11383 1177
rect 11383 1143 11417 1177
rect 11417 1143 11426 1177
rect 11374 1134 11426 1143
rect 11374 1017 11426 1026
rect 11374 983 11383 1017
rect 11383 983 11417 1017
rect 11417 983 11426 1017
rect 11374 974 11426 983
rect 11374 537 11426 546
rect 11374 503 11383 537
rect 11383 503 11417 537
rect 11417 503 11426 537
rect 11374 494 11426 503
rect 11374 377 11426 386
rect 11374 343 11383 377
rect 11383 343 11417 377
rect 11417 343 11426 377
rect 11374 334 11426 343
rect 11374 217 11426 226
rect 11374 183 11383 217
rect 11383 183 11417 217
rect 11417 183 11426 217
rect 11374 174 11426 183
rect 11374 57 11426 66
rect 11374 23 11383 57
rect 11383 23 11417 57
rect 11417 23 11426 57
rect 11374 14 11426 23
rect 11534 31417 11586 31426
rect 11534 31383 11543 31417
rect 11543 31383 11577 31417
rect 11577 31383 11586 31417
rect 11534 31374 11586 31383
rect 11534 31257 11586 31266
rect 11534 31223 11543 31257
rect 11543 31223 11577 31257
rect 11577 31223 11586 31257
rect 11534 31214 11586 31223
rect 11534 31097 11586 31106
rect 11534 31063 11543 31097
rect 11543 31063 11577 31097
rect 11577 31063 11586 31097
rect 11534 31054 11586 31063
rect 11534 30937 11586 30946
rect 11534 30903 11543 30937
rect 11543 30903 11577 30937
rect 11577 30903 11586 30937
rect 11534 30894 11586 30903
rect 11534 30777 11586 30786
rect 11534 30743 11543 30777
rect 11543 30743 11577 30777
rect 11577 30743 11586 30777
rect 11534 30734 11586 30743
rect 11534 30617 11586 30626
rect 11534 30583 11543 30617
rect 11543 30583 11577 30617
rect 11577 30583 11586 30617
rect 11534 30574 11586 30583
rect 11534 30457 11586 30466
rect 11534 30423 11543 30457
rect 11543 30423 11577 30457
rect 11577 30423 11586 30457
rect 11534 30414 11586 30423
rect 11534 30297 11586 30306
rect 11534 30263 11543 30297
rect 11543 30263 11577 30297
rect 11577 30263 11586 30297
rect 11534 30254 11586 30263
rect 11534 29977 11586 29986
rect 11534 29943 11543 29977
rect 11543 29943 11577 29977
rect 11577 29943 11586 29977
rect 11534 29934 11586 29943
rect 11534 29817 11586 29826
rect 11534 29783 11543 29817
rect 11543 29783 11577 29817
rect 11577 29783 11586 29817
rect 11534 29774 11586 29783
rect 11534 29657 11586 29666
rect 11534 29623 11543 29657
rect 11543 29623 11577 29657
rect 11577 29623 11586 29657
rect 11534 29614 11586 29623
rect 11534 29497 11586 29506
rect 11534 29463 11543 29497
rect 11543 29463 11577 29497
rect 11577 29463 11586 29497
rect 11534 29454 11586 29463
rect 11534 29337 11586 29346
rect 11534 29303 11543 29337
rect 11543 29303 11577 29337
rect 11577 29303 11586 29337
rect 11534 29294 11586 29303
rect 11534 29177 11586 29186
rect 11534 29143 11543 29177
rect 11543 29143 11577 29177
rect 11577 29143 11586 29177
rect 11534 29134 11586 29143
rect 11534 29017 11586 29026
rect 11534 28983 11543 29017
rect 11543 28983 11577 29017
rect 11577 28983 11586 29017
rect 11534 28974 11586 28983
rect 11534 28857 11586 28866
rect 11534 28823 11543 28857
rect 11543 28823 11577 28857
rect 11577 28823 11586 28857
rect 11534 28814 11586 28823
rect 11534 28057 11586 28066
rect 11534 28023 11543 28057
rect 11543 28023 11577 28057
rect 11577 28023 11586 28057
rect 11534 28014 11586 28023
rect 11534 27897 11586 27906
rect 11534 27863 11543 27897
rect 11543 27863 11577 27897
rect 11577 27863 11586 27897
rect 11534 27854 11586 27863
rect 11534 27737 11586 27746
rect 11534 27703 11543 27737
rect 11543 27703 11577 27737
rect 11577 27703 11586 27737
rect 11534 27694 11586 27703
rect 11534 27577 11586 27586
rect 11534 27543 11543 27577
rect 11543 27543 11577 27577
rect 11577 27543 11586 27577
rect 11534 27534 11586 27543
rect 11534 27417 11586 27426
rect 11534 27383 11543 27417
rect 11543 27383 11577 27417
rect 11577 27383 11586 27417
rect 11534 27374 11586 27383
rect 11534 27257 11586 27266
rect 11534 27223 11543 27257
rect 11543 27223 11577 27257
rect 11577 27223 11586 27257
rect 11534 27214 11586 27223
rect 11534 27097 11586 27106
rect 11534 27063 11543 27097
rect 11543 27063 11577 27097
rect 11577 27063 11586 27097
rect 11534 27054 11586 27063
rect 11534 26937 11586 26946
rect 11534 26903 11543 26937
rect 11543 26903 11577 26937
rect 11577 26903 11586 26937
rect 11534 26894 11586 26903
rect 11534 26137 11586 26146
rect 11534 26103 11543 26137
rect 11543 26103 11577 26137
rect 11577 26103 11586 26137
rect 11534 26094 11586 26103
rect 11534 25977 11586 25986
rect 11534 25943 11543 25977
rect 11543 25943 11577 25977
rect 11577 25943 11586 25977
rect 11534 25934 11586 25943
rect 11534 25817 11586 25826
rect 11534 25783 11543 25817
rect 11543 25783 11577 25817
rect 11577 25783 11586 25817
rect 11534 25774 11586 25783
rect 11534 25657 11586 25666
rect 11534 25623 11543 25657
rect 11543 25623 11577 25657
rect 11577 25623 11586 25657
rect 11534 25614 11586 25623
rect 11534 25497 11586 25506
rect 11534 25463 11543 25497
rect 11543 25463 11577 25497
rect 11577 25463 11586 25497
rect 11534 25454 11586 25463
rect 11534 25337 11586 25346
rect 11534 25303 11543 25337
rect 11543 25303 11577 25337
rect 11577 25303 11586 25337
rect 11534 25294 11586 25303
rect 11534 25177 11586 25186
rect 11534 25143 11543 25177
rect 11543 25143 11577 25177
rect 11577 25143 11586 25177
rect 11534 25134 11586 25143
rect 11534 25017 11586 25026
rect 11534 24983 11543 25017
rect 11543 24983 11577 25017
rect 11577 24983 11586 25017
rect 11534 24974 11586 24983
rect 11534 24697 11586 24706
rect 11534 24663 11543 24697
rect 11543 24663 11577 24697
rect 11577 24663 11586 24697
rect 11534 24654 11586 24663
rect 11534 24537 11586 24546
rect 11534 24503 11543 24537
rect 11543 24503 11577 24537
rect 11577 24503 11586 24537
rect 11534 24494 11586 24503
rect 11534 24377 11586 24386
rect 11534 24343 11543 24377
rect 11543 24343 11577 24377
rect 11577 24343 11586 24377
rect 11534 24334 11586 24343
rect 11534 24217 11586 24226
rect 11534 24183 11543 24217
rect 11543 24183 11577 24217
rect 11577 24183 11586 24217
rect 11534 24174 11586 24183
rect 11534 24057 11586 24066
rect 11534 24023 11543 24057
rect 11543 24023 11577 24057
rect 11577 24023 11586 24057
rect 11534 24014 11586 24023
rect 11534 23897 11586 23906
rect 11534 23863 11543 23897
rect 11543 23863 11577 23897
rect 11577 23863 11586 23897
rect 11534 23854 11586 23863
rect 11534 23737 11586 23746
rect 11534 23703 11543 23737
rect 11543 23703 11577 23737
rect 11577 23703 11586 23737
rect 11534 23694 11586 23703
rect 11534 23577 11586 23586
rect 11534 23543 11543 23577
rect 11543 23543 11577 23577
rect 11577 23543 11586 23577
rect 11534 23534 11586 23543
rect 11534 23417 11586 23426
rect 11534 23383 11543 23417
rect 11543 23383 11577 23417
rect 11577 23383 11586 23417
rect 11534 23374 11586 23383
rect 11534 23257 11586 23266
rect 11534 23223 11543 23257
rect 11543 23223 11577 23257
rect 11577 23223 11586 23257
rect 11534 23214 11586 23223
rect 11534 23097 11586 23106
rect 11534 23063 11543 23097
rect 11543 23063 11577 23097
rect 11577 23063 11586 23097
rect 11534 23054 11586 23063
rect 11534 22937 11586 22946
rect 11534 22903 11543 22937
rect 11543 22903 11577 22937
rect 11577 22903 11586 22937
rect 11534 22894 11586 22903
rect 11534 22777 11586 22786
rect 11534 22743 11543 22777
rect 11543 22743 11577 22777
rect 11577 22743 11586 22777
rect 11534 22734 11586 22743
rect 11534 22617 11586 22626
rect 11534 22583 11543 22617
rect 11543 22583 11577 22617
rect 11577 22583 11586 22617
rect 11534 22574 11586 22583
rect 11534 22457 11586 22466
rect 11534 22423 11543 22457
rect 11543 22423 11577 22457
rect 11577 22423 11586 22457
rect 11534 22414 11586 22423
rect 11534 22297 11586 22306
rect 11534 22263 11543 22297
rect 11543 22263 11577 22297
rect 11577 22263 11586 22297
rect 11534 22254 11586 22263
rect 11534 22137 11586 22146
rect 11534 22103 11543 22137
rect 11543 22103 11577 22137
rect 11577 22103 11586 22137
rect 11534 22094 11586 22103
rect 11534 21817 11586 21826
rect 11534 21783 11543 21817
rect 11543 21783 11577 21817
rect 11577 21783 11586 21817
rect 11534 21774 11586 21783
rect 11534 21657 11586 21666
rect 11534 21623 11543 21657
rect 11543 21623 11577 21657
rect 11577 21623 11586 21657
rect 11534 21614 11586 21623
rect 11534 21497 11586 21506
rect 11534 21463 11543 21497
rect 11543 21463 11577 21497
rect 11577 21463 11586 21497
rect 11534 21454 11586 21463
rect 11534 21337 11586 21346
rect 11534 21303 11543 21337
rect 11543 21303 11577 21337
rect 11577 21303 11586 21337
rect 11534 21294 11586 21303
rect 11534 21177 11586 21186
rect 11534 21143 11543 21177
rect 11543 21143 11577 21177
rect 11577 21143 11586 21177
rect 11534 21134 11586 21143
rect 11534 21017 11586 21026
rect 11534 20983 11543 21017
rect 11543 20983 11577 21017
rect 11577 20983 11586 21017
rect 11534 20974 11586 20983
rect 11534 20857 11586 20866
rect 11534 20823 11543 20857
rect 11543 20823 11577 20857
rect 11577 20823 11586 20857
rect 11534 20814 11586 20823
rect 11534 20697 11586 20706
rect 11534 20663 11543 20697
rect 11543 20663 11577 20697
rect 11577 20663 11586 20697
rect 11534 20654 11586 20663
rect 11534 19897 11586 19906
rect 11534 19863 11543 19897
rect 11543 19863 11577 19897
rect 11577 19863 11586 19897
rect 11534 19854 11586 19863
rect 11534 19737 11586 19746
rect 11534 19703 11543 19737
rect 11543 19703 11577 19737
rect 11577 19703 11586 19737
rect 11534 19694 11586 19703
rect 11534 19577 11586 19586
rect 11534 19543 11543 19577
rect 11543 19543 11577 19577
rect 11577 19543 11586 19577
rect 11534 19534 11586 19543
rect 11534 19417 11586 19426
rect 11534 19383 11543 19417
rect 11543 19383 11577 19417
rect 11577 19383 11586 19417
rect 11534 19374 11586 19383
rect 11534 19257 11586 19266
rect 11534 19223 11543 19257
rect 11543 19223 11577 19257
rect 11577 19223 11586 19257
rect 11534 19214 11586 19223
rect 11534 19097 11586 19106
rect 11534 19063 11543 19097
rect 11543 19063 11577 19097
rect 11577 19063 11586 19097
rect 11534 19054 11586 19063
rect 11534 18937 11586 18946
rect 11534 18903 11543 18937
rect 11543 18903 11577 18937
rect 11577 18903 11586 18937
rect 11534 18894 11586 18903
rect 11534 18777 11586 18786
rect 11534 18743 11543 18777
rect 11543 18743 11577 18777
rect 11577 18743 11586 18777
rect 11534 18734 11586 18743
rect 11534 17977 11586 17986
rect 11534 17943 11543 17977
rect 11543 17943 11577 17977
rect 11577 17943 11586 17977
rect 11534 17934 11586 17943
rect 11534 17817 11586 17826
rect 11534 17783 11543 17817
rect 11543 17783 11577 17817
rect 11577 17783 11586 17817
rect 11534 17774 11586 17783
rect 11534 17657 11586 17666
rect 11534 17623 11543 17657
rect 11543 17623 11577 17657
rect 11577 17623 11586 17657
rect 11534 17614 11586 17623
rect 11534 17497 11586 17506
rect 11534 17463 11543 17497
rect 11543 17463 11577 17497
rect 11577 17463 11586 17497
rect 11534 17454 11586 17463
rect 11534 17337 11586 17346
rect 11534 17303 11543 17337
rect 11543 17303 11577 17337
rect 11577 17303 11586 17337
rect 11534 17294 11586 17303
rect 11534 17177 11586 17186
rect 11534 17143 11543 17177
rect 11543 17143 11577 17177
rect 11577 17143 11586 17177
rect 11534 17134 11586 17143
rect 11534 17017 11586 17026
rect 11534 16983 11543 17017
rect 11543 16983 11577 17017
rect 11577 16983 11586 17017
rect 11534 16974 11586 16983
rect 11534 16857 11586 16866
rect 11534 16823 11543 16857
rect 11543 16823 11577 16857
rect 11577 16823 11586 16857
rect 11534 16814 11586 16823
rect 11534 16537 11586 16546
rect 11534 16503 11543 16537
rect 11543 16503 11577 16537
rect 11577 16503 11586 16537
rect 11534 16494 11586 16503
rect 11534 16377 11586 16386
rect 11534 16343 11543 16377
rect 11543 16343 11577 16377
rect 11577 16343 11586 16377
rect 11534 16334 11586 16343
rect 11534 16217 11586 16226
rect 11534 16183 11543 16217
rect 11543 16183 11577 16217
rect 11577 16183 11586 16217
rect 11534 16174 11586 16183
rect 11534 16057 11586 16066
rect 11534 16023 11543 16057
rect 11543 16023 11577 16057
rect 11577 16023 11586 16057
rect 11534 16014 11586 16023
rect 11534 15897 11586 15906
rect 11534 15863 11543 15897
rect 11543 15863 11577 15897
rect 11577 15863 11586 15897
rect 11534 15854 11586 15863
rect 11534 15737 11586 15746
rect 11534 15703 11543 15737
rect 11543 15703 11577 15737
rect 11577 15703 11586 15737
rect 11534 15694 11586 15703
rect 11534 15577 11586 15586
rect 11534 15543 11543 15577
rect 11543 15543 11577 15577
rect 11577 15543 11586 15577
rect 11534 15534 11586 15543
rect 11534 15417 11586 15426
rect 11534 15383 11543 15417
rect 11543 15383 11577 15417
rect 11577 15383 11586 15417
rect 11534 15374 11586 15383
rect 11534 15257 11586 15266
rect 11534 15223 11543 15257
rect 11543 15223 11577 15257
rect 11577 15223 11586 15257
rect 11534 15214 11586 15223
rect 11534 15097 11586 15106
rect 11534 15063 11543 15097
rect 11543 15063 11577 15097
rect 11577 15063 11586 15097
rect 11534 15054 11586 15063
rect 11534 14937 11586 14946
rect 11534 14903 11543 14937
rect 11543 14903 11577 14937
rect 11577 14903 11586 14937
rect 11534 14894 11586 14903
rect 11534 14777 11586 14786
rect 11534 14743 11543 14777
rect 11543 14743 11577 14777
rect 11577 14743 11586 14777
rect 11534 14734 11586 14743
rect 11534 14617 11586 14626
rect 11534 14583 11543 14617
rect 11543 14583 11577 14617
rect 11577 14583 11586 14617
rect 11534 14574 11586 14583
rect 11534 14457 11586 14466
rect 11534 14423 11543 14457
rect 11543 14423 11577 14457
rect 11577 14423 11586 14457
rect 11534 14414 11586 14423
rect 11534 14297 11586 14306
rect 11534 14263 11543 14297
rect 11543 14263 11577 14297
rect 11577 14263 11586 14297
rect 11534 14254 11586 14263
rect 11534 14137 11586 14146
rect 11534 14103 11543 14137
rect 11543 14103 11577 14137
rect 11577 14103 11586 14137
rect 11534 14094 11586 14103
rect 11534 13977 11586 13986
rect 11534 13943 11543 13977
rect 11543 13943 11577 13977
rect 11577 13943 11586 13977
rect 11534 13934 11586 13943
rect 11534 13657 11586 13666
rect 11534 13623 11543 13657
rect 11543 13623 11577 13657
rect 11577 13623 11586 13657
rect 11534 13614 11586 13623
rect 11534 13497 11586 13506
rect 11534 13463 11543 13497
rect 11543 13463 11577 13497
rect 11577 13463 11586 13497
rect 11534 13454 11586 13463
rect 11534 13337 11586 13346
rect 11534 13303 11543 13337
rect 11543 13303 11577 13337
rect 11577 13303 11586 13337
rect 11534 13294 11586 13303
rect 11534 13177 11586 13186
rect 11534 13143 11543 13177
rect 11543 13143 11577 13177
rect 11577 13143 11586 13177
rect 11534 13134 11586 13143
rect 11534 13017 11586 13026
rect 11534 12983 11543 13017
rect 11543 12983 11577 13017
rect 11577 12983 11586 13017
rect 11534 12974 11586 12983
rect 11534 12857 11586 12866
rect 11534 12823 11543 12857
rect 11543 12823 11577 12857
rect 11577 12823 11586 12857
rect 11534 12814 11586 12823
rect 11534 12697 11586 12706
rect 11534 12663 11543 12697
rect 11543 12663 11577 12697
rect 11577 12663 11586 12697
rect 11534 12654 11586 12663
rect 11534 12537 11586 12546
rect 11534 12503 11543 12537
rect 11543 12503 11577 12537
rect 11577 12503 11586 12537
rect 11534 12494 11586 12503
rect 11534 11737 11586 11746
rect 11534 11703 11543 11737
rect 11543 11703 11577 11737
rect 11577 11703 11586 11737
rect 11534 11694 11586 11703
rect 11534 11577 11586 11586
rect 11534 11543 11543 11577
rect 11543 11543 11577 11577
rect 11577 11543 11586 11577
rect 11534 11534 11586 11543
rect 11534 11417 11586 11426
rect 11534 11383 11543 11417
rect 11543 11383 11577 11417
rect 11577 11383 11586 11417
rect 11534 11374 11586 11383
rect 11534 11257 11586 11266
rect 11534 11223 11543 11257
rect 11543 11223 11577 11257
rect 11577 11223 11586 11257
rect 11534 11214 11586 11223
rect 11534 11097 11586 11106
rect 11534 11063 11543 11097
rect 11543 11063 11577 11097
rect 11577 11063 11586 11097
rect 11534 11054 11586 11063
rect 11534 10937 11586 10946
rect 11534 10903 11543 10937
rect 11543 10903 11577 10937
rect 11577 10903 11586 10937
rect 11534 10894 11586 10903
rect 11534 10777 11586 10786
rect 11534 10743 11543 10777
rect 11543 10743 11577 10777
rect 11577 10743 11586 10777
rect 11534 10734 11586 10743
rect 11534 10617 11586 10626
rect 11534 10583 11543 10617
rect 11543 10583 11577 10617
rect 11577 10583 11586 10617
rect 11534 10574 11586 10583
rect 11534 10457 11586 10466
rect 11534 10423 11543 10457
rect 11543 10423 11577 10457
rect 11577 10423 11586 10457
rect 11534 10414 11586 10423
rect 11534 10297 11586 10306
rect 11534 10263 11543 10297
rect 11543 10263 11577 10297
rect 11577 10263 11586 10297
rect 11534 10254 11586 10263
rect 11534 10137 11586 10146
rect 11534 10103 11543 10137
rect 11543 10103 11577 10137
rect 11577 10103 11586 10137
rect 11534 10094 11586 10103
rect 11534 9977 11586 9986
rect 11534 9943 11543 9977
rect 11543 9943 11577 9977
rect 11577 9943 11586 9977
rect 11534 9934 11586 9943
rect 11534 9817 11586 9826
rect 11534 9783 11543 9817
rect 11543 9783 11577 9817
rect 11577 9783 11586 9817
rect 11534 9774 11586 9783
rect 11534 9497 11586 9506
rect 11534 9463 11543 9497
rect 11543 9463 11577 9497
rect 11577 9463 11586 9497
rect 11534 9454 11586 9463
rect 11534 9337 11586 9346
rect 11534 9303 11543 9337
rect 11543 9303 11577 9337
rect 11577 9303 11586 9337
rect 11534 9294 11586 9303
rect 11534 9017 11586 9026
rect 11534 8983 11543 9017
rect 11543 8983 11577 9017
rect 11577 8983 11586 9017
rect 11534 8974 11586 8983
rect 11534 8857 11586 8866
rect 11534 8823 11543 8857
rect 11543 8823 11577 8857
rect 11577 8823 11586 8857
rect 11534 8814 11586 8823
rect 11534 8697 11586 8706
rect 11534 8663 11543 8697
rect 11543 8663 11577 8697
rect 11577 8663 11586 8697
rect 11534 8654 11586 8663
rect 11534 8537 11586 8546
rect 11534 8503 11543 8537
rect 11543 8503 11577 8537
rect 11577 8503 11586 8537
rect 11534 8494 11586 8503
rect 11534 8377 11586 8386
rect 11534 8343 11543 8377
rect 11543 8343 11577 8377
rect 11577 8343 11586 8377
rect 11534 8334 11586 8343
rect 11534 8217 11586 8226
rect 11534 8183 11543 8217
rect 11543 8183 11577 8217
rect 11577 8183 11586 8217
rect 11534 8174 11586 8183
rect 11534 8057 11586 8066
rect 11534 8023 11543 8057
rect 11543 8023 11577 8057
rect 11577 8023 11586 8057
rect 11534 8014 11586 8023
rect 11534 7897 11586 7906
rect 11534 7863 11543 7897
rect 11543 7863 11577 7897
rect 11577 7863 11586 7897
rect 11534 7854 11586 7863
rect 11534 7737 11586 7746
rect 11534 7703 11543 7737
rect 11543 7703 11577 7737
rect 11577 7703 11586 7737
rect 11534 7694 11586 7703
rect 11534 7417 11586 7426
rect 11534 7383 11543 7417
rect 11543 7383 11577 7417
rect 11577 7383 11586 7417
rect 11534 7374 11586 7383
rect 11534 7257 11586 7266
rect 11534 7223 11543 7257
rect 11543 7223 11577 7257
rect 11577 7223 11586 7257
rect 11534 7214 11586 7223
rect 11534 6937 11586 6946
rect 11534 6903 11543 6937
rect 11543 6903 11577 6937
rect 11577 6903 11586 6937
rect 11534 6894 11586 6903
rect 11534 6777 11586 6786
rect 11534 6743 11543 6777
rect 11543 6743 11577 6777
rect 11577 6743 11586 6777
rect 11534 6734 11586 6743
rect 11534 6457 11586 6466
rect 11534 6423 11543 6457
rect 11543 6423 11577 6457
rect 11577 6423 11586 6457
rect 11534 6414 11586 6423
rect 11534 6297 11586 6306
rect 11534 6263 11543 6297
rect 11543 6263 11577 6297
rect 11577 6263 11586 6297
rect 11534 6254 11586 6263
rect 11534 6137 11586 6146
rect 11534 6103 11543 6137
rect 11543 6103 11577 6137
rect 11577 6103 11586 6137
rect 11534 6094 11586 6103
rect 11534 5977 11586 5986
rect 11534 5943 11543 5977
rect 11543 5943 11577 5977
rect 11577 5943 11586 5977
rect 11534 5934 11586 5943
rect 11534 5817 11586 5826
rect 11534 5783 11543 5817
rect 11543 5783 11577 5817
rect 11577 5783 11586 5817
rect 11534 5774 11586 5783
rect 11534 5657 11586 5666
rect 11534 5623 11543 5657
rect 11543 5623 11577 5657
rect 11577 5623 11586 5657
rect 11534 5614 11586 5623
rect 11534 5497 11586 5506
rect 11534 5463 11543 5497
rect 11543 5463 11577 5497
rect 11577 5463 11586 5497
rect 11534 5454 11586 5463
rect 11534 5337 11586 5346
rect 11534 5303 11543 5337
rect 11543 5303 11577 5337
rect 11577 5303 11586 5337
rect 11534 5294 11586 5303
rect 11534 5177 11586 5186
rect 11534 5143 11543 5177
rect 11543 5143 11577 5177
rect 11577 5143 11586 5177
rect 11534 5134 11586 5143
rect 11534 5017 11586 5026
rect 11534 4983 11543 5017
rect 11543 4983 11577 5017
rect 11577 4983 11586 5017
rect 11534 4974 11586 4983
rect 11534 4857 11586 4866
rect 11534 4823 11543 4857
rect 11543 4823 11577 4857
rect 11577 4823 11586 4857
rect 11534 4814 11586 4823
rect 11534 4697 11586 4706
rect 11534 4663 11543 4697
rect 11543 4663 11577 4697
rect 11577 4663 11586 4697
rect 11534 4654 11586 4663
rect 11534 4537 11586 4546
rect 11534 4503 11543 4537
rect 11543 4503 11577 4537
rect 11577 4503 11586 4537
rect 11534 4494 11586 4503
rect 11534 4377 11586 4386
rect 11534 4343 11543 4377
rect 11543 4343 11577 4377
rect 11577 4343 11586 4377
rect 11534 4334 11586 4343
rect 11534 4217 11586 4226
rect 11534 4183 11543 4217
rect 11543 4183 11577 4217
rect 11577 4183 11586 4217
rect 11534 4174 11586 4183
rect 11534 4057 11586 4066
rect 11534 4023 11543 4057
rect 11543 4023 11577 4057
rect 11577 4023 11586 4057
rect 11534 4014 11586 4023
rect 11534 3897 11586 3906
rect 11534 3863 11543 3897
rect 11543 3863 11577 3897
rect 11577 3863 11586 3897
rect 11534 3854 11586 3863
rect 11534 3417 11586 3426
rect 11534 3383 11543 3417
rect 11543 3383 11577 3417
rect 11577 3383 11586 3417
rect 11534 3374 11586 3383
rect 11534 3257 11586 3266
rect 11534 3223 11543 3257
rect 11543 3223 11577 3257
rect 11577 3223 11586 3257
rect 11534 3214 11586 3223
rect 11534 3097 11586 3106
rect 11534 3063 11543 3097
rect 11543 3063 11577 3097
rect 11577 3063 11586 3097
rect 11534 3054 11586 3063
rect 11534 2937 11586 2946
rect 11534 2903 11543 2937
rect 11543 2903 11577 2937
rect 11577 2903 11586 2937
rect 11534 2894 11586 2903
rect 11534 2777 11586 2786
rect 11534 2743 11543 2777
rect 11543 2743 11577 2777
rect 11577 2743 11586 2777
rect 11534 2734 11586 2743
rect 11534 2617 11586 2626
rect 11534 2583 11543 2617
rect 11543 2583 11577 2617
rect 11577 2583 11586 2617
rect 11534 2574 11586 2583
rect 11534 2457 11586 2466
rect 11534 2423 11543 2457
rect 11543 2423 11577 2457
rect 11577 2423 11586 2457
rect 11534 2414 11586 2423
rect 11534 2297 11586 2306
rect 11534 2263 11543 2297
rect 11543 2263 11577 2297
rect 11577 2263 11586 2297
rect 11534 2254 11586 2263
rect 11534 2137 11586 2146
rect 11534 2103 11543 2137
rect 11543 2103 11577 2137
rect 11577 2103 11586 2137
rect 11534 2094 11586 2103
rect 11534 1977 11586 1986
rect 11534 1943 11543 1977
rect 11543 1943 11577 1977
rect 11577 1943 11586 1977
rect 11534 1934 11586 1943
rect 11534 1657 11586 1666
rect 11534 1623 11543 1657
rect 11543 1623 11577 1657
rect 11577 1623 11586 1657
rect 11534 1614 11586 1623
rect 11534 1497 11586 1506
rect 11534 1463 11543 1497
rect 11543 1463 11577 1497
rect 11577 1463 11586 1497
rect 11534 1454 11586 1463
rect 11534 1337 11586 1346
rect 11534 1303 11543 1337
rect 11543 1303 11577 1337
rect 11577 1303 11586 1337
rect 11534 1294 11586 1303
rect 11534 1177 11586 1186
rect 11534 1143 11543 1177
rect 11543 1143 11577 1177
rect 11577 1143 11586 1177
rect 11534 1134 11586 1143
rect 11534 1017 11586 1026
rect 11534 983 11543 1017
rect 11543 983 11577 1017
rect 11577 983 11586 1017
rect 11534 974 11586 983
rect 11534 537 11586 546
rect 11534 503 11543 537
rect 11543 503 11577 537
rect 11577 503 11586 537
rect 11534 494 11586 503
rect 11534 377 11586 386
rect 11534 343 11543 377
rect 11543 343 11577 377
rect 11577 343 11586 377
rect 11534 334 11586 343
rect 11534 217 11586 226
rect 11534 183 11543 217
rect 11543 183 11577 217
rect 11577 183 11586 217
rect 11534 174 11586 183
rect 11534 57 11586 66
rect 11534 23 11543 57
rect 11543 23 11577 57
rect 11577 23 11586 57
rect 11534 14 11586 23
rect 11854 31417 11906 31426
rect 11854 31383 11863 31417
rect 11863 31383 11897 31417
rect 11897 31383 11906 31417
rect 11854 31374 11906 31383
rect 11854 31257 11906 31266
rect 11854 31223 11863 31257
rect 11863 31223 11897 31257
rect 11897 31223 11906 31257
rect 11854 31214 11906 31223
rect 11854 31097 11906 31106
rect 11854 31063 11863 31097
rect 11863 31063 11897 31097
rect 11897 31063 11906 31097
rect 11854 31054 11906 31063
rect 11854 30937 11906 30946
rect 11854 30903 11863 30937
rect 11863 30903 11897 30937
rect 11897 30903 11906 30937
rect 11854 30894 11906 30903
rect 11854 30777 11906 30786
rect 11854 30743 11863 30777
rect 11863 30743 11897 30777
rect 11897 30743 11906 30777
rect 11854 30734 11906 30743
rect 11854 30617 11906 30626
rect 11854 30583 11863 30617
rect 11863 30583 11897 30617
rect 11897 30583 11906 30617
rect 11854 30574 11906 30583
rect 11854 30457 11906 30466
rect 11854 30423 11863 30457
rect 11863 30423 11897 30457
rect 11897 30423 11906 30457
rect 11854 30414 11906 30423
rect 11854 30297 11906 30306
rect 11854 30263 11863 30297
rect 11863 30263 11897 30297
rect 11897 30263 11906 30297
rect 11854 30254 11906 30263
rect 11854 29977 11906 29986
rect 11854 29943 11863 29977
rect 11863 29943 11897 29977
rect 11897 29943 11906 29977
rect 11854 29934 11906 29943
rect 11854 29817 11906 29826
rect 11854 29783 11863 29817
rect 11863 29783 11897 29817
rect 11897 29783 11906 29817
rect 11854 29774 11906 29783
rect 11854 29657 11906 29666
rect 11854 29623 11863 29657
rect 11863 29623 11897 29657
rect 11897 29623 11906 29657
rect 11854 29614 11906 29623
rect 11854 29497 11906 29506
rect 11854 29463 11863 29497
rect 11863 29463 11897 29497
rect 11897 29463 11906 29497
rect 11854 29454 11906 29463
rect 11854 29337 11906 29346
rect 11854 29303 11863 29337
rect 11863 29303 11897 29337
rect 11897 29303 11906 29337
rect 11854 29294 11906 29303
rect 11854 29177 11906 29186
rect 11854 29143 11863 29177
rect 11863 29143 11897 29177
rect 11897 29143 11906 29177
rect 11854 29134 11906 29143
rect 11854 29017 11906 29026
rect 11854 28983 11863 29017
rect 11863 28983 11897 29017
rect 11897 28983 11906 29017
rect 11854 28974 11906 28983
rect 11854 28857 11906 28866
rect 11854 28823 11863 28857
rect 11863 28823 11897 28857
rect 11897 28823 11906 28857
rect 11854 28814 11906 28823
rect 11854 28057 11906 28066
rect 11854 28023 11863 28057
rect 11863 28023 11897 28057
rect 11897 28023 11906 28057
rect 11854 28014 11906 28023
rect 11854 27897 11906 27906
rect 11854 27863 11863 27897
rect 11863 27863 11897 27897
rect 11897 27863 11906 27897
rect 11854 27854 11906 27863
rect 11854 27737 11906 27746
rect 11854 27703 11863 27737
rect 11863 27703 11897 27737
rect 11897 27703 11906 27737
rect 11854 27694 11906 27703
rect 11854 27577 11906 27586
rect 11854 27543 11863 27577
rect 11863 27543 11897 27577
rect 11897 27543 11906 27577
rect 11854 27534 11906 27543
rect 11854 27417 11906 27426
rect 11854 27383 11863 27417
rect 11863 27383 11897 27417
rect 11897 27383 11906 27417
rect 11854 27374 11906 27383
rect 11854 27257 11906 27266
rect 11854 27223 11863 27257
rect 11863 27223 11897 27257
rect 11897 27223 11906 27257
rect 11854 27214 11906 27223
rect 11854 27097 11906 27106
rect 11854 27063 11863 27097
rect 11863 27063 11897 27097
rect 11897 27063 11906 27097
rect 11854 27054 11906 27063
rect 11854 26937 11906 26946
rect 11854 26903 11863 26937
rect 11863 26903 11897 26937
rect 11897 26903 11906 26937
rect 11854 26894 11906 26903
rect 11854 26137 11906 26146
rect 11854 26103 11863 26137
rect 11863 26103 11897 26137
rect 11897 26103 11906 26137
rect 11854 26094 11906 26103
rect 11854 25977 11906 25986
rect 11854 25943 11863 25977
rect 11863 25943 11897 25977
rect 11897 25943 11906 25977
rect 11854 25934 11906 25943
rect 11854 25817 11906 25826
rect 11854 25783 11863 25817
rect 11863 25783 11897 25817
rect 11897 25783 11906 25817
rect 11854 25774 11906 25783
rect 11854 25657 11906 25666
rect 11854 25623 11863 25657
rect 11863 25623 11897 25657
rect 11897 25623 11906 25657
rect 11854 25614 11906 25623
rect 11854 25497 11906 25506
rect 11854 25463 11863 25497
rect 11863 25463 11897 25497
rect 11897 25463 11906 25497
rect 11854 25454 11906 25463
rect 11854 25337 11906 25346
rect 11854 25303 11863 25337
rect 11863 25303 11897 25337
rect 11897 25303 11906 25337
rect 11854 25294 11906 25303
rect 11854 25177 11906 25186
rect 11854 25143 11863 25177
rect 11863 25143 11897 25177
rect 11897 25143 11906 25177
rect 11854 25134 11906 25143
rect 11854 25017 11906 25026
rect 11854 24983 11863 25017
rect 11863 24983 11897 25017
rect 11897 24983 11906 25017
rect 11854 24974 11906 24983
rect 11854 24697 11906 24706
rect 11854 24663 11863 24697
rect 11863 24663 11897 24697
rect 11897 24663 11906 24697
rect 11854 24654 11906 24663
rect 11854 24537 11906 24546
rect 11854 24503 11863 24537
rect 11863 24503 11897 24537
rect 11897 24503 11906 24537
rect 11854 24494 11906 24503
rect 11854 24377 11906 24386
rect 11854 24343 11863 24377
rect 11863 24343 11897 24377
rect 11897 24343 11906 24377
rect 11854 24334 11906 24343
rect 11854 24217 11906 24226
rect 11854 24183 11863 24217
rect 11863 24183 11897 24217
rect 11897 24183 11906 24217
rect 11854 24174 11906 24183
rect 11854 24057 11906 24066
rect 11854 24023 11863 24057
rect 11863 24023 11897 24057
rect 11897 24023 11906 24057
rect 11854 24014 11906 24023
rect 11854 23897 11906 23906
rect 11854 23863 11863 23897
rect 11863 23863 11897 23897
rect 11897 23863 11906 23897
rect 11854 23854 11906 23863
rect 11854 23737 11906 23746
rect 11854 23703 11863 23737
rect 11863 23703 11897 23737
rect 11897 23703 11906 23737
rect 11854 23694 11906 23703
rect 11854 23577 11906 23586
rect 11854 23543 11863 23577
rect 11863 23543 11897 23577
rect 11897 23543 11906 23577
rect 11854 23534 11906 23543
rect 11854 23417 11906 23426
rect 11854 23383 11863 23417
rect 11863 23383 11897 23417
rect 11897 23383 11906 23417
rect 11854 23374 11906 23383
rect 11854 23257 11906 23266
rect 11854 23223 11863 23257
rect 11863 23223 11897 23257
rect 11897 23223 11906 23257
rect 11854 23214 11906 23223
rect 11854 23097 11906 23106
rect 11854 23063 11863 23097
rect 11863 23063 11897 23097
rect 11897 23063 11906 23097
rect 11854 23054 11906 23063
rect 11854 22937 11906 22946
rect 11854 22903 11863 22937
rect 11863 22903 11897 22937
rect 11897 22903 11906 22937
rect 11854 22894 11906 22903
rect 11854 22777 11906 22786
rect 11854 22743 11863 22777
rect 11863 22743 11897 22777
rect 11897 22743 11906 22777
rect 11854 22734 11906 22743
rect 11854 22617 11906 22626
rect 11854 22583 11863 22617
rect 11863 22583 11897 22617
rect 11897 22583 11906 22617
rect 11854 22574 11906 22583
rect 11854 22457 11906 22466
rect 11854 22423 11863 22457
rect 11863 22423 11897 22457
rect 11897 22423 11906 22457
rect 11854 22414 11906 22423
rect 11854 22297 11906 22306
rect 11854 22263 11863 22297
rect 11863 22263 11897 22297
rect 11897 22263 11906 22297
rect 11854 22254 11906 22263
rect 11854 22137 11906 22146
rect 11854 22103 11863 22137
rect 11863 22103 11897 22137
rect 11897 22103 11906 22137
rect 11854 22094 11906 22103
rect 11854 21817 11906 21826
rect 11854 21783 11863 21817
rect 11863 21783 11897 21817
rect 11897 21783 11906 21817
rect 11854 21774 11906 21783
rect 11854 21657 11906 21666
rect 11854 21623 11863 21657
rect 11863 21623 11897 21657
rect 11897 21623 11906 21657
rect 11854 21614 11906 21623
rect 11854 21497 11906 21506
rect 11854 21463 11863 21497
rect 11863 21463 11897 21497
rect 11897 21463 11906 21497
rect 11854 21454 11906 21463
rect 11854 21337 11906 21346
rect 11854 21303 11863 21337
rect 11863 21303 11897 21337
rect 11897 21303 11906 21337
rect 11854 21294 11906 21303
rect 11854 21177 11906 21186
rect 11854 21143 11863 21177
rect 11863 21143 11897 21177
rect 11897 21143 11906 21177
rect 11854 21134 11906 21143
rect 11854 21017 11906 21026
rect 11854 20983 11863 21017
rect 11863 20983 11897 21017
rect 11897 20983 11906 21017
rect 11854 20974 11906 20983
rect 11854 20857 11906 20866
rect 11854 20823 11863 20857
rect 11863 20823 11897 20857
rect 11897 20823 11906 20857
rect 11854 20814 11906 20823
rect 11854 20697 11906 20706
rect 11854 20663 11863 20697
rect 11863 20663 11897 20697
rect 11897 20663 11906 20697
rect 11854 20654 11906 20663
rect 11854 19897 11906 19906
rect 11854 19863 11863 19897
rect 11863 19863 11897 19897
rect 11897 19863 11906 19897
rect 11854 19854 11906 19863
rect 11854 19737 11906 19746
rect 11854 19703 11863 19737
rect 11863 19703 11897 19737
rect 11897 19703 11906 19737
rect 11854 19694 11906 19703
rect 11854 19577 11906 19586
rect 11854 19543 11863 19577
rect 11863 19543 11897 19577
rect 11897 19543 11906 19577
rect 11854 19534 11906 19543
rect 11854 19417 11906 19426
rect 11854 19383 11863 19417
rect 11863 19383 11897 19417
rect 11897 19383 11906 19417
rect 11854 19374 11906 19383
rect 11854 19257 11906 19266
rect 11854 19223 11863 19257
rect 11863 19223 11897 19257
rect 11897 19223 11906 19257
rect 11854 19214 11906 19223
rect 11854 19097 11906 19106
rect 11854 19063 11863 19097
rect 11863 19063 11897 19097
rect 11897 19063 11906 19097
rect 11854 19054 11906 19063
rect 11854 18937 11906 18946
rect 11854 18903 11863 18937
rect 11863 18903 11897 18937
rect 11897 18903 11906 18937
rect 11854 18894 11906 18903
rect 11854 18777 11906 18786
rect 11854 18743 11863 18777
rect 11863 18743 11897 18777
rect 11897 18743 11906 18777
rect 11854 18734 11906 18743
rect 11854 17977 11906 17986
rect 11854 17943 11863 17977
rect 11863 17943 11897 17977
rect 11897 17943 11906 17977
rect 11854 17934 11906 17943
rect 11854 17817 11906 17826
rect 11854 17783 11863 17817
rect 11863 17783 11897 17817
rect 11897 17783 11906 17817
rect 11854 17774 11906 17783
rect 11854 17657 11906 17666
rect 11854 17623 11863 17657
rect 11863 17623 11897 17657
rect 11897 17623 11906 17657
rect 11854 17614 11906 17623
rect 11854 17497 11906 17506
rect 11854 17463 11863 17497
rect 11863 17463 11897 17497
rect 11897 17463 11906 17497
rect 11854 17454 11906 17463
rect 11854 17337 11906 17346
rect 11854 17303 11863 17337
rect 11863 17303 11897 17337
rect 11897 17303 11906 17337
rect 11854 17294 11906 17303
rect 11854 17177 11906 17186
rect 11854 17143 11863 17177
rect 11863 17143 11897 17177
rect 11897 17143 11906 17177
rect 11854 17134 11906 17143
rect 11854 17017 11906 17026
rect 11854 16983 11863 17017
rect 11863 16983 11897 17017
rect 11897 16983 11906 17017
rect 11854 16974 11906 16983
rect 11854 16857 11906 16866
rect 11854 16823 11863 16857
rect 11863 16823 11897 16857
rect 11897 16823 11906 16857
rect 11854 16814 11906 16823
rect 11854 16537 11906 16546
rect 11854 16503 11863 16537
rect 11863 16503 11897 16537
rect 11897 16503 11906 16537
rect 11854 16494 11906 16503
rect 11854 16377 11906 16386
rect 11854 16343 11863 16377
rect 11863 16343 11897 16377
rect 11897 16343 11906 16377
rect 11854 16334 11906 16343
rect 11854 16217 11906 16226
rect 11854 16183 11863 16217
rect 11863 16183 11897 16217
rect 11897 16183 11906 16217
rect 11854 16174 11906 16183
rect 11854 16057 11906 16066
rect 11854 16023 11863 16057
rect 11863 16023 11897 16057
rect 11897 16023 11906 16057
rect 11854 16014 11906 16023
rect 11854 15897 11906 15906
rect 11854 15863 11863 15897
rect 11863 15863 11897 15897
rect 11897 15863 11906 15897
rect 11854 15854 11906 15863
rect 11854 15737 11906 15746
rect 11854 15703 11863 15737
rect 11863 15703 11897 15737
rect 11897 15703 11906 15737
rect 11854 15694 11906 15703
rect 11854 15577 11906 15586
rect 11854 15543 11863 15577
rect 11863 15543 11897 15577
rect 11897 15543 11906 15577
rect 11854 15534 11906 15543
rect 11854 15417 11906 15426
rect 11854 15383 11863 15417
rect 11863 15383 11897 15417
rect 11897 15383 11906 15417
rect 11854 15374 11906 15383
rect 11854 15257 11906 15266
rect 11854 15223 11863 15257
rect 11863 15223 11897 15257
rect 11897 15223 11906 15257
rect 11854 15214 11906 15223
rect 11854 15097 11906 15106
rect 11854 15063 11863 15097
rect 11863 15063 11897 15097
rect 11897 15063 11906 15097
rect 11854 15054 11906 15063
rect 11854 14937 11906 14946
rect 11854 14903 11863 14937
rect 11863 14903 11897 14937
rect 11897 14903 11906 14937
rect 11854 14894 11906 14903
rect 11854 14777 11906 14786
rect 11854 14743 11863 14777
rect 11863 14743 11897 14777
rect 11897 14743 11906 14777
rect 11854 14734 11906 14743
rect 11854 14617 11906 14626
rect 11854 14583 11863 14617
rect 11863 14583 11897 14617
rect 11897 14583 11906 14617
rect 11854 14574 11906 14583
rect 11854 14457 11906 14466
rect 11854 14423 11863 14457
rect 11863 14423 11897 14457
rect 11897 14423 11906 14457
rect 11854 14414 11906 14423
rect 11854 14297 11906 14306
rect 11854 14263 11863 14297
rect 11863 14263 11897 14297
rect 11897 14263 11906 14297
rect 11854 14254 11906 14263
rect 11854 14137 11906 14146
rect 11854 14103 11863 14137
rect 11863 14103 11897 14137
rect 11897 14103 11906 14137
rect 11854 14094 11906 14103
rect 11854 13977 11906 13986
rect 11854 13943 11863 13977
rect 11863 13943 11897 13977
rect 11897 13943 11906 13977
rect 11854 13934 11906 13943
rect 11854 13657 11906 13666
rect 11854 13623 11863 13657
rect 11863 13623 11897 13657
rect 11897 13623 11906 13657
rect 11854 13614 11906 13623
rect 11854 13497 11906 13506
rect 11854 13463 11863 13497
rect 11863 13463 11897 13497
rect 11897 13463 11906 13497
rect 11854 13454 11906 13463
rect 11854 13337 11906 13346
rect 11854 13303 11863 13337
rect 11863 13303 11897 13337
rect 11897 13303 11906 13337
rect 11854 13294 11906 13303
rect 11854 13177 11906 13186
rect 11854 13143 11863 13177
rect 11863 13143 11897 13177
rect 11897 13143 11906 13177
rect 11854 13134 11906 13143
rect 11854 13017 11906 13026
rect 11854 12983 11863 13017
rect 11863 12983 11897 13017
rect 11897 12983 11906 13017
rect 11854 12974 11906 12983
rect 11854 12857 11906 12866
rect 11854 12823 11863 12857
rect 11863 12823 11897 12857
rect 11897 12823 11906 12857
rect 11854 12814 11906 12823
rect 11854 12697 11906 12706
rect 11854 12663 11863 12697
rect 11863 12663 11897 12697
rect 11897 12663 11906 12697
rect 11854 12654 11906 12663
rect 11854 12537 11906 12546
rect 11854 12503 11863 12537
rect 11863 12503 11897 12537
rect 11897 12503 11906 12537
rect 11854 12494 11906 12503
rect 11854 11737 11906 11746
rect 11854 11703 11863 11737
rect 11863 11703 11897 11737
rect 11897 11703 11906 11737
rect 11854 11694 11906 11703
rect 11854 11577 11906 11586
rect 11854 11543 11863 11577
rect 11863 11543 11897 11577
rect 11897 11543 11906 11577
rect 11854 11534 11906 11543
rect 11854 11417 11906 11426
rect 11854 11383 11863 11417
rect 11863 11383 11897 11417
rect 11897 11383 11906 11417
rect 11854 11374 11906 11383
rect 11854 11257 11906 11266
rect 11854 11223 11863 11257
rect 11863 11223 11897 11257
rect 11897 11223 11906 11257
rect 11854 11214 11906 11223
rect 11854 11097 11906 11106
rect 11854 11063 11863 11097
rect 11863 11063 11897 11097
rect 11897 11063 11906 11097
rect 11854 11054 11906 11063
rect 11854 10937 11906 10946
rect 11854 10903 11863 10937
rect 11863 10903 11897 10937
rect 11897 10903 11906 10937
rect 11854 10894 11906 10903
rect 11854 10777 11906 10786
rect 11854 10743 11863 10777
rect 11863 10743 11897 10777
rect 11897 10743 11906 10777
rect 11854 10734 11906 10743
rect 11854 10617 11906 10626
rect 11854 10583 11863 10617
rect 11863 10583 11897 10617
rect 11897 10583 11906 10617
rect 11854 10574 11906 10583
rect 11854 10457 11906 10466
rect 11854 10423 11863 10457
rect 11863 10423 11897 10457
rect 11897 10423 11906 10457
rect 11854 10414 11906 10423
rect 11854 10297 11906 10306
rect 11854 10263 11863 10297
rect 11863 10263 11897 10297
rect 11897 10263 11906 10297
rect 11854 10254 11906 10263
rect 11854 10137 11906 10146
rect 11854 10103 11863 10137
rect 11863 10103 11897 10137
rect 11897 10103 11906 10137
rect 11854 10094 11906 10103
rect 11854 9977 11906 9986
rect 11854 9943 11863 9977
rect 11863 9943 11897 9977
rect 11897 9943 11906 9977
rect 11854 9934 11906 9943
rect 11854 9817 11906 9826
rect 11854 9783 11863 9817
rect 11863 9783 11897 9817
rect 11897 9783 11906 9817
rect 11854 9774 11906 9783
rect 11854 9497 11906 9506
rect 11854 9463 11863 9497
rect 11863 9463 11897 9497
rect 11897 9463 11906 9497
rect 11854 9454 11906 9463
rect 11854 9337 11906 9346
rect 11854 9303 11863 9337
rect 11863 9303 11897 9337
rect 11897 9303 11906 9337
rect 11854 9294 11906 9303
rect 11854 9017 11906 9026
rect 11854 8983 11863 9017
rect 11863 8983 11897 9017
rect 11897 8983 11906 9017
rect 11854 8974 11906 8983
rect 11854 8857 11906 8866
rect 11854 8823 11863 8857
rect 11863 8823 11897 8857
rect 11897 8823 11906 8857
rect 11854 8814 11906 8823
rect 11854 8697 11906 8706
rect 11854 8663 11863 8697
rect 11863 8663 11897 8697
rect 11897 8663 11906 8697
rect 11854 8654 11906 8663
rect 11854 8537 11906 8546
rect 11854 8503 11863 8537
rect 11863 8503 11897 8537
rect 11897 8503 11906 8537
rect 11854 8494 11906 8503
rect 11854 8377 11906 8386
rect 11854 8343 11863 8377
rect 11863 8343 11897 8377
rect 11897 8343 11906 8377
rect 11854 8334 11906 8343
rect 11854 8217 11906 8226
rect 11854 8183 11863 8217
rect 11863 8183 11897 8217
rect 11897 8183 11906 8217
rect 11854 8174 11906 8183
rect 11854 8057 11906 8066
rect 11854 8023 11863 8057
rect 11863 8023 11897 8057
rect 11897 8023 11906 8057
rect 11854 8014 11906 8023
rect 11854 7897 11906 7906
rect 11854 7863 11863 7897
rect 11863 7863 11897 7897
rect 11897 7863 11906 7897
rect 11854 7854 11906 7863
rect 11854 7737 11906 7746
rect 11854 7703 11863 7737
rect 11863 7703 11897 7737
rect 11897 7703 11906 7737
rect 11854 7694 11906 7703
rect 11854 7417 11906 7426
rect 11854 7383 11863 7417
rect 11863 7383 11897 7417
rect 11897 7383 11906 7417
rect 11854 7374 11906 7383
rect 11854 7257 11906 7266
rect 11854 7223 11863 7257
rect 11863 7223 11897 7257
rect 11897 7223 11906 7257
rect 11854 7214 11906 7223
rect 11854 6937 11906 6946
rect 11854 6903 11863 6937
rect 11863 6903 11897 6937
rect 11897 6903 11906 6937
rect 11854 6894 11906 6903
rect 11854 6777 11906 6786
rect 11854 6743 11863 6777
rect 11863 6743 11897 6777
rect 11897 6743 11906 6777
rect 11854 6734 11906 6743
rect 11854 6457 11906 6466
rect 11854 6423 11863 6457
rect 11863 6423 11897 6457
rect 11897 6423 11906 6457
rect 11854 6414 11906 6423
rect 11854 6297 11906 6306
rect 11854 6263 11863 6297
rect 11863 6263 11897 6297
rect 11897 6263 11906 6297
rect 11854 6254 11906 6263
rect 11854 6137 11906 6146
rect 11854 6103 11863 6137
rect 11863 6103 11897 6137
rect 11897 6103 11906 6137
rect 11854 6094 11906 6103
rect 11854 5977 11906 5986
rect 11854 5943 11863 5977
rect 11863 5943 11897 5977
rect 11897 5943 11906 5977
rect 11854 5934 11906 5943
rect 11854 5817 11906 5826
rect 11854 5783 11863 5817
rect 11863 5783 11897 5817
rect 11897 5783 11906 5817
rect 11854 5774 11906 5783
rect 11854 5657 11906 5666
rect 11854 5623 11863 5657
rect 11863 5623 11897 5657
rect 11897 5623 11906 5657
rect 11854 5614 11906 5623
rect 11854 5497 11906 5506
rect 11854 5463 11863 5497
rect 11863 5463 11897 5497
rect 11897 5463 11906 5497
rect 11854 5454 11906 5463
rect 11854 5337 11906 5346
rect 11854 5303 11863 5337
rect 11863 5303 11897 5337
rect 11897 5303 11906 5337
rect 11854 5294 11906 5303
rect 11854 5177 11906 5186
rect 11854 5143 11863 5177
rect 11863 5143 11897 5177
rect 11897 5143 11906 5177
rect 11854 5134 11906 5143
rect 11854 5017 11906 5026
rect 11854 4983 11863 5017
rect 11863 4983 11897 5017
rect 11897 4983 11906 5017
rect 11854 4974 11906 4983
rect 11854 4857 11906 4866
rect 11854 4823 11863 4857
rect 11863 4823 11897 4857
rect 11897 4823 11906 4857
rect 11854 4814 11906 4823
rect 11854 4697 11906 4706
rect 11854 4663 11863 4697
rect 11863 4663 11897 4697
rect 11897 4663 11906 4697
rect 11854 4654 11906 4663
rect 11854 4537 11906 4546
rect 11854 4503 11863 4537
rect 11863 4503 11897 4537
rect 11897 4503 11906 4537
rect 11854 4494 11906 4503
rect 11854 4377 11906 4386
rect 11854 4343 11863 4377
rect 11863 4343 11897 4377
rect 11897 4343 11906 4377
rect 11854 4334 11906 4343
rect 11854 4217 11906 4226
rect 11854 4183 11863 4217
rect 11863 4183 11897 4217
rect 11897 4183 11906 4217
rect 11854 4174 11906 4183
rect 11854 4057 11906 4066
rect 11854 4023 11863 4057
rect 11863 4023 11897 4057
rect 11897 4023 11906 4057
rect 11854 4014 11906 4023
rect 11854 3897 11906 3906
rect 11854 3863 11863 3897
rect 11863 3863 11897 3897
rect 11897 3863 11906 3897
rect 11854 3854 11906 3863
rect 11854 3417 11906 3426
rect 11854 3383 11863 3417
rect 11863 3383 11897 3417
rect 11897 3383 11906 3417
rect 11854 3374 11906 3383
rect 11854 3257 11906 3266
rect 11854 3223 11863 3257
rect 11863 3223 11897 3257
rect 11897 3223 11906 3257
rect 11854 3214 11906 3223
rect 11854 3097 11906 3106
rect 11854 3063 11863 3097
rect 11863 3063 11897 3097
rect 11897 3063 11906 3097
rect 11854 3054 11906 3063
rect 11854 2937 11906 2946
rect 11854 2903 11863 2937
rect 11863 2903 11897 2937
rect 11897 2903 11906 2937
rect 11854 2894 11906 2903
rect 11854 2777 11906 2786
rect 11854 2743 11863 2777
rect 11863 2743 11897 2777
rect 11897 2743 11906 2777
rect 11854 2734 11906 2743
rect 11854 2617 11906 2626
rect 11854 2583 11863 2617
rect 11863 2583 11897 2617
rect 11897 2583 11906 2617
rect 11854 2574 11906 2583
rect 11854 2457 11906 2466
rect 11854 2423 11863 2457
rect 11863 2423 11897 2457
rect 11897 2423 11906 2457
rect 11854 2414 11906 2423
rect 11854 2297 11906 2306
rect 11854 2263 11863 2297
rect 11863 2263 11897 2297
rect 11897 2263 11906 2297
rect 11854 2254 11906 2263
rect 11854 2137 11906 2146
rect 11854 2103 11863 2137
rect 11863 2103 11897 2137
rect 11897 2103 11906 2137
rect 11854 2094 11906 2103
rect 11854 1977 11906 1986
rect 11854 1943 11863 1977
rect 11863 1943 11897 1977
rect 11897 1943 11906 1977
rect 11854 1934 11906 1943
rect 11854 1657 11906 1666
rect 11854 1623 11863 1657
rect 11863 1623 11897 1657
rect 11897 1623 11906 1657
rect 11854 1614 11906 1623
rect 11854 1497 11906 1506
rect 11854 1463 11863 1497
rect 11863 1463 11897 1497
rect 11897 1463 11906 1497
rect 11854 1454 11906 1463
rect 11854 1337 11906 1346
rect 11854 1303 11863 1337
rect 11863 1303 11897 1337
rect 11897 1303 11906 1337
rect 11854 1294 11906 1303
rect 11854 1177 11906 1186
rect 11854 1143 11863 1177
rect 11863 1143 11897 1177
rect 11897 1143 11906 1177
rect 11854 1134 11906 1143
rect 11854 1017 11906 1026
rect 11854 983 11863 1017
rect 11863 983 11897 1017
rect 11897 983 11906 1017
rect 11854 974 11906 983
rect 11854 537 11906 546
rect 11854 503 11863 537
rect 11863 503 11897 537
rect 11897 503 11906 537
rect 11854 494 11906 503
rect 11854 377 11906 386
rect 11854 343 11863 377
rect 11863 343 11897 377
rect 11897 343 11906 377
rect 11854 334 11906 343
rect 11854 217 11906 226
rect 11854 183 11863 217
rect 11863 183 11897 217
rect 11897 183 11906 217
rect 11854 174 11906 183
rect 11854 57 11906 66
rect 11854 23 11863 57
rect 11863 23 11897 57
rect 11897 23 11906 57
rect 11854 14 11906 23
rect 12014 31417 12066 31426
rect 12014 31383 12023 31417
rect 12023 31383 12057 31417
rect 12057 31383 12066 31417
rect 12014 31374 12066 31383
rect 12014 31257 12066 31266
rect 12014 31223 12023 31257
rect 12023 31223 12057 31257
rect 12057 31223 12066 31257
rect 12014 31214 12066 31223
rect 12014 31097 12066 31106
rect 12014 31063 12023 31097
rect 12023 31063 12057 31097
rect 12057 31063 12066 31097
rect 12014 31054 12066 31063
rect 12014 30937 12066 30946
rect 12014 30903 12023 30937
rect 12023 30903 12057 30937
rect 12057 30903 12066 30937
rect 12014 30894 12066 30903
rect 12014 30777 12066 30786
rect 12014 30743 12023 30777
rect 12023 30743 12057 30777
rect 12057 30743 12066 30777
rect 12014 30734 12066 30743
rect 12014 30617 12066 30626
rect 12014 30583 12023 30617
rect 12023 30583 12057 30617
rect 12057 30583 12066 30617
rect 12014 30574 12066 30583
rect 12014 30457 12066 30466
rect 12014 30423 12023 30457
rect 12023 30423 12057 30457
rect 12057 30423 12066 30457
rect 12014 30414 12066 30423
rect 12014 30297 12066 30306
rect 12014 30263 12023 30297
rect 12023 30263 12057 30297
rect 12057 30263 12066 30297
rect 12014 30254 12066 30263
rect 12014 29977 12066 29986
rect 12014 29943 12023 29977
rect 12023 29943 12057 29977
rect 12057 29943 12066 29977
rect 12014 29934 12066 29943
rect 12014 29817 12066 29826
rect 12014 29783 12023 29817
rect 12023 29783 12057 29817
rect 12057 29783 12066 29817
rect 12014 29774 12066 29783
rect 12014 29657 12066 29666
rect 12014 29623 12023 29657
rect 12023 29623 12057 29657
rect 12057 29623 12066 29657
rect 12014 29614 12066 29623
rect 12014 29497 12066 29506
rect 12014 29463 12023 29497
rect 12023 29463 12057 29497
rect 12057 29463 12066 29497
rect 12014 29454 12066 29463
rect 12014 29337 12066 29346
rect 12014 29303 12023 29337
rect 12023 29303 12057 29337
rect 12057 29303 12066 29337
rect 12014 29294 12066 29303
rect 12014 29177 12066 29186
rect 12014 29143 12023 29177
rect 12023 29143 12057 29177
rect 12057 29143 12066 29177
rect 12014 29134 12066 29143
rect 12014 29017 12066 29026
rect 12014 28983 12023 29017
rect 12023 28983 12057 29017
rect 12057 28983 12066 29017
rect 12014 28974 12066 28983
rect 12014 28857 12066 28866
rect 12014 28823 12023 28857
rect 12023 28823 12057 28857
rect 12057 28823 12066 28857
rect 12014 28814 12066 28823
rect 12014 28057 12066 28066
rect 12014 28023 12023 28057
rect 12023 28023 12057 28057
rect 12057 28023 12066 28057
rect 12014 28014 12066 28023
rect 12014 27897 12066 27906
rect 12014 27863 12023 27897
rect 12023 27863 12057 27897
rect 12057 27863 12066 27897
rect 12014 27854 12066 27863
rect 12014 27737 12066 27746
rect 12014 27703 12023 27737
rect 12023 27703 12057 27737
rect 12057 27703 12066 27737
rect 12014 27694 12066 27703
rect 12014 27577 12066 27586
rect 12014 27543 12023 27577
rect 12023 27543 12057 27577
rect 12057 27543 12066 27577
rect 12014 27534 12066 27543
rect 12014 27417 12066 27426
rect 12014 27383 12023 27417
rect 12023 27383 12057 27417
rect 12057 27383 12066 27417
rect 12014 27374 12066 27383
rect 12014 27257 12066 27266
rect 12014 27223 12023 27257
rect 12023 27223 12057 27257
rect 12057 27223 12066 27257
rect 12014 27214 12066 27223
rect 12014 27097 12066 27106
rect 12014 27063 12023 27097
rect 12023 27063 12057 27097
rect 12057 27063 12066 27097
rect 12014 27054 12066 27063
rect 12014 26937 12066 26946
rect 12014 26903 12023 26937
rect 12023 26903 12057 26937
rect 12057 26903 12066 26937
rect 12014 26894 12066 26903
rect 12014 26137 12066 26146
rect 12014 26103 12023 26137
rect 12023 26103 12057 26137
rect 12057 26103 12066 26137
rect 12014 26094 12066 26103
rect 12014 25977 12066 25986
rect 12014 25943 12023 25977
rect 12023 25943 12057 25977
rect 12057 25943 12066 25977
rect 12014 25934 12066 25943
rect 12014 25817 12066 25826
rect 12014 25783 12023 25817
rect 12023 25783 12057 25817
rect 12057 25783 12066 25817
rect 12014 25774 12066 25783
rect 12014 25657 12066 25666
rect 12014 25623 12023 25657
rect 12023 25623 12057 25657
rect 12057 25623 12066 25657
rect 12014 25614 12066 25623
rect 12014 25497 12066 25506
rect 12014 25463 12023 25497
rect 12023 25463 12057 25497
rect 12057 25463 12066 25497
rect 12014 25454 12066 25463
rect 12014 25337 12066 25346
rect 12014 25303 12023 25337
rect 12023 25303 12057 25337
rect 12057 25303 12066 25337
rect 12014 25294 12066 25303
rect 12014 25177 12066 25186
rect 12014 25143 12023 25177
rect 12023 25143 12057 25177
rect 12057 25143 12066 25177
rect 12014 25134 12066 25143
rect 12014 25017 12066 25026
rect 12014 24983 12023 25017
rect 12023 24983 12057 25017
rect 12057 24983 12066 25017
rect 12014 24974 12066 24983
rect 12014 24697 12066 24706
rect 12014 24663 12023 24697
rect 12023 24663 12057 24697
rect 12057 24663 12066 24697
rect 12014 24654 12066 24663
rect 12014 24537 12066 24546
rect 12014 24503 12023 24537
rect 12023 24503 12057 24537
rect 12057 24503 12066 24537
rect 12014 24494 12066 24503
rect 12014 24377 12066 24386
rect 12014 24343 12023 24377
rect 12023 24343 12057 24377
rect 12057 24343 12066 24377
rect 12014 24334 12066 24343
rect 12014 24217 12066 24226
rect 12014 24183 12023 24217
rect 12023 24183 12057 24217
rect 12057 24183 12066 24217
rect 12014 24174 12066 24183
rect 12014 24057 12066 24066
rect 12014 24023 12023 24057
rect 12023 24023 12057 24057
rect 12057 24023 12066 24057
rect 12014 24014 12066 24023
rect 12014 23897 12066 23906
rect 12014 23863 12023 23897
rect 12023 23863 12057 23897
rect 12057 23863 12066 23897
rect 12014 23854 12066 23863
rect 12014 23737 12066 23746
rect 12014 23703 12023 23737
rect 12023 23703 12057 23737
rect 12057 23703 12066 23737
rect 12014 23694 12066 23703
rect 12014 23577 12066 23586
rect 12014 23543 12023 23577
rect 12023 23543 12057 23577
rect 12057 23543 12066 23577
rect 12014 23534 12066 23543
rect 12014 23417 12066 23426
rect 12014 23383 12023 23417
rect 12023 23383 12057 23417
rect 12057 23383 12066 23417
rect 12014 23374 12066 23383
rect 12014 23257 12066 23266
rect 12014 23223 12023 23257
rect 12023 23223 12057 23257
rect 12057 23223 12066 23257
rect 12014 23214 12066 23223
rect 12014 23097 12066 23106
rect 12014 23063 12023 23097
rect 12023 23063 12057 23097
rect 12057 23063 12066 23097
rect 12014 23054 12066 23063
rect 12014 22937 12066 22946
rect 12014 22903 12023 22937
rect 12023 22903 12057 22937
rect 12057 22903 12066 22937
rect 12014 22894 12066 22903
rect 12014 22777 12066 22786
rect 12014 22743 12023 22777
rect 12023 22743 12057 22777
rect 12057 22743 12066 22777
rect 12014 22734 12066 22743
rect 12014 22617 12066 22626
rect 12014 22583 12023 22617
rect 12023 22583 12057 22617
rect 12057 22583 12066 22617
rect 12014 22574 12066 22583
rect 12014 22457 12066 22466
rect 12014 22423 12023 22457
rect 12023 22423 12057 22457
rect 12057 22423 12066 22457
rect 12014 22414 12066 22423
rect 12014 22297 12066 22306
rect 12014 22263 12023 22297
rect 12023 22263 12057 22297
rect 12057 22263 12066 22297
rect 12014 22254 12066 22263
rect 12014 22137 12066 22146
rect 12014 22103 12023 22137
rect 12023 22103 12057 22137
rect 12057 22103 12066 22137
rect 12014 22094 12066 22103
rect 12014 21817 12066 21826
rect 12014 21783 12023 21817
rect 12023 21783 12057 21817
rect 12057 21783 12066 21817
rect 12014 21774 12066 21783
rect 12014 21657 12066 21666
rect 12014 21623 12023 21657
rect 12023 21623 12057 21657
rect 12057 21623 12066 21657
rect 12014 21614 12066 21623
rect 12014 21497 12066 21506
rect 12014 21463 12023 21497
rect 12023 21463 12057 21497
rect 12057 21463 12066 21497
rect 12014 21454 12066 21463
rect 12014 21337 12066 21346
rect 12014 21303 12023 21337
rect 12023 21303 12057 21337
rect 12057 21303 12066 21337
rect 12014 21294 12066 21303
rect 12014 21177 12066 21186
rect 12014 21143 12023 21177
rect 12023 21143 12057 21177
rect 12057 21143 12066 21177
rect 12014 21134 12066 21143
rect 12014 21017 12066 21026
rect 12014 20983 12023 21017
rect 12023 20983 12057 21017
rect 12057 20983 12066 21017
rect 12014 20974 12066 20983
rect 12014 20857 12066 20866
rect 12014 20823 12023 20857
rect 12023 20823 12057 20857
rect 12057 20823 12066 20857
rect 12014 20814 12066 20823
rect 12014 20697 12066 20706
rect 12014 20663 12023 20697
rect 12023 20663 12057 20697
rect 12057 20663 12066 20697
rect 12014 20654 12066 20663
rect 12014 19897 12066 19906
rect 12014 19863 12023 19897
rect 12023 19863 12057 19897
rect 12057 19863 12066 19897
rect 12014 19854 12066 19863
rect 12014 19737 12066 19746
rect 12014 19703 12023 19737
rect 12023 19703 12057 19737
rect 12057 19703 12066 19737
rect 12014 19694 12066 19703
rect 12014 19577 12066 19586
rect 12014 19543 12023 19577
rect 12023 19543 12057 19577
rect 12057 19543 12066 19577
rect 12014 19534 12066 19543
rect 12014 19417 12066 19426
rect 12014 19383 12023 19417
rect 12023 19383 12057 19417
rect 12057 19383 12066 19417
rect 12014 19374 12066 19383
rect 12014 19257 12066 19266
rect 12014 19223 12023 19257
rect 12023 19223 12057 19257
rect 12057 19223 12066 19257
rect 12014 19214 12066 19223
rect 12014 19097 12066 19106
rect 12014 19063 12023 19097
rect 12023 19063 12057 19097
rect 12057 19063 12066 19097
rect 12014 19054 12066 19063
rect 12014 18937 12066 18946
rect 12014 18903 12023 18937
rect 12023 18903 12057 18937
rect 12057 18903 12066 18937
rect 12014 18894 12066 18903
rect 12014 18777 12066 18786
rect 12014 18743 12023 18777
rect 12023 18743 12057 18777
rect 12057 18743 12066 18777
rect 12014 18734 12066 18743
rect 12014 17977 12066 17986
rect 12014 17943 12023 17977
rect 12023 17943 12057 17977
rect 12057 17943 12066 17977
rect 12014 17934 12066 17943
rect 12014 17817 12066 17826
rect 12014 17783 12023 17817
rect 12023 17783 12057 17817
rect 12057 17783 12066 17817
rect 12014 17774 12066 17783
rect 12014 17657 12066 17666
rect 12014 17623 12023 17657
rect 12023 17623 12057 17657
rect 12057 17623 12066 17657
rect 12014 17614 12066 17623
rect 12014 17497 12066 17506
rect 12014 17463 12023 17497
rect 12023 17463 12057 17497
rect 12057 17463 12066 17497
rect 12014 17454 12066 17463
rect 12014 17337 12066 17346
rect 12014 17303 12023 17337
rect 12023 17303 12057 17337
rect 12057 17303 12066 17337
rect 12014 17294 12066 17303
rect 12014 17177 12066 17186
rect 12014 17143 12023 17177
rect 12023 17143 12057 17177
rect 12057 17143 12066 17177
rect 12014 17134 12066 17143
rect 12014 17017 12066 17026
rect 12014 16983 12023 17017
rect 12023 16983 12057 17017
rect 12057 16983 12066 17017
rect 12014 16974 12066 16983
rect 12014 16857 12066 16866
rect 12014 16823 12023 16857
rect 12023 16823 12057 16857
rect 12057 16823 12066 16857
rect 12014 16814 12066 16823
rect 12014 16537 12066 16546
rect 12014 16503 12023 16537
rect 12023 16503 12057 16537
rect 12057 16503 12066 16537
rect 12014 16494 12066 16503
rect 12014 16377 12066 16386
rect 12014 16343 12023 16377
rect 12023 16343 12057 16377
rect 12057 16343 12066 16377
rect 12014 16334 12066 16343
rect 12014 16217 12066 16226
rect 12014 16183 12023 16217
rect 12023 16183 12057 16217
rect 12057 16183 12066 16217
rect 12014 16174 12066 16183
rect 12014 16057 12066 16066
rect 12014 16023 12023 16057
rect 12023 16023 12057 16057
rect 12057 16023 12066 16057
rect 12014 16014 12066 16023
rect 12014 15897 12066 15906
rect 12014 15863 12023 15897
rect 12023 15863 12057 15897
rect 12057 15863 12066 15897
rect 12014 15854 12066 15863
rect 12014 15737 12066 15746
rect 12014 15703 12023 15737
rect 12023 15703 12057 15737
rect 12057 15703 12066 15737
rect 12014 15694 12066 15703
rect 12014 15577 12066 15586
rect 12014 15543 12023 15577
rect 12023 15543 12057 15577
rect 12057 15543 12066 15577
rect 12014 15534 12066 15543
rect 12014 15417 12066 15426
rect 12014 15383 12023 15417
rect 12023 15383 12057 15417
rect 12057 15383 12066 15417
rect 12014 15374 12066 15383
rect 12014 15257 12066 15266
rect 12014 15223 12023 15257
rect 12023 15223 12057 15257
rect 12057 15223 12066 15257
rect 12014 15214 12066 15223
rect 12014 15097 12066 15106
rect 12014 15063 12023 15097
rect 12023 15063 12057 15097
rect 12057 15063 12066 15097
rect 12014 15054 12066 15063
rect 12014 14937 12066 14946
rect 12014 14903 12023 14937
rect 12023 14903 12057 14937
rect 12057 14903 12066 14937
rect 12014 14894 12066 14903
rect 12014 14777 12066 14786
rect 12014 14743 12023 14777
rect 12023 14743 12057 14777
rect 12057 14743 12066 14777
rect 12014 14734 12066 14743
rect 12014 14617 12066 14626
rect 12014 14583 12023 14617
rect 12023 14583 12057 14617
rect 12057 14583 12066 14617
rect 12014 14574 12066 14583
rect 12014 14457 12066 14466
rect 12014 14423 12023 14457
rect 12023 14423 12057 14457
rect 12057 14423 12066 14457
rect 12014 14414 12066 14423
rect 12014 14297 12066 14306
rect 12014 14263 12023 14297
rect 12023 14263 12057 14297
rect 12057 14263 12066 14297
rect 12014 14254 12066 14263
rect 12014 14137 12066 14146
rect 12014 14103 12023 14137
rect 12023 14103 12057 14137
rect 12057 14103 12066 14137
rect 12014 14094 12066 14103
rect 12014 13977 12066 13986
rect 12014 13943 12023 13977
rect 12023 13943 12057 13977
rect 12057 13943 12066 13977
rect 12014 13934 12066 13943
rect 12014 13657 12066 13666
rect 12014 13623 12023 13657
rect 12023 13623 12057 13657
rect 12057 13623 12066 13657
rect 12014 13614 12066 13623
rect 12014 13497 12066 13506
rect 12014 13463 12023 13497
rect 12023 13463 12057 13497
rect 12057 13463 12066 13497
rect 12014 13454 12066 13463
rect 12014 13337 12066 13346
rect 12014 13303 12023 13337
rect 12023 13303 12057 13337
rect 12057 13303 12066 13337
rect 12014 13294 12066 13303
rect 12014 13177 12066 13186
rect 12014 13143 12023 13177
rect 12023 13143 12057 13177
rect 12057 13143 12066 13177
rect 12014 13134 12066 13143
rect 12014 13017 12066 13026
rect 12014 12983 12023 13017
rect 12023 12983 12057 13017
rect 12057 12983 12066 13017
rect 12014 12974 12066 12983
rect 12014 12857 12066 12866
rect 12014 12823 12023 12857
rect 12023 12823 12057 12857
rect 12057 12823 12066 12857
rect 12014 12814 12066 12823
rect 12014 12697 12066 12706
rect 12014 12663 12023 12697
rect 12023 12663 12057 12697
rect 12057 12663 12066 12697
rect 12014 12654 12066 12663
rect 12014 12537 12066 12546
rect 12014 12503 12023 12537
rect 12023 12503 12057 12537
rect 12057 12503 12066 12537
rect 12014 12494 12066 12503
rect 12014 11737 12066 11746
rect 12014 11703 12023 11737
rect 12023 11703 12057 11737
rect 12057 11703 12066 11737
rect 12014 11694 12066 11703
rect 12014 11577 12066 11586
rect 12014 11543 12023 11577
rect 12023 11543 12057 11577
rect 12057 11543 12066 11577
rect 12014 11534 12066 11543
rect 12014 11417 12066 11426
rect 12014 11383 12023 11417
rect 12023 11383 12057 11417
rect 12057 11383 12066 11417
rect 12014 11374 12066 11383
rect 12014 11257 12066 11266
rect 12014 11223 12023 11257
rect 12023 11223 12057 11257
rect 12057 11223 12066 11257
rect 12014 11214 12066 11223
rect 12014 11097 12066 11106
rect 12014 11063 12023 11097
rect 12023 11063 12057 11097
rect 12057 11063 12066 11097
rect 12014 11054 12066 11063
rect 12014 10937 12066 10946
rect 12014 10903 12023 10937
rect 12023 10903 12057 10937
rect 12057 10903 12066 10937
rect 12014 10894 12066 10903
rect 12014 10777 12066 10786
rect 12014 10743 12023 10777
rect 12023 10743 12057 10777
rect 12057 10743 12066 10777
rect 12014 10734 12066 10743
rect 12014 10617 12066 10626
rect 12014 10583 12023 10617
rect 12023 10583 12057 10617
rect 12057 10583 12066 10617
rect 12014 10574 12066 10583
rect 12014 10457 12066 10466
rect 12014 10423 12023 10457
rect 12023 10423 12057 10457
rect 12057 10423 12066 10457
rect 12014 10414 12066 10423
rect 12014 10297 12066 10306
rect 12014 10263 12023 10297
rect 12023 10263 12057 10297
rect 12057 10263 12066 10297
rect 12014 10254 12066 10263
rect 12014 10137 12066 10146
rect 12014 10103 12023 10137
rect 12023 10103 12057 10137
rect 12057 10103 12066 10137
rect 12014 10094 12066 10103
rect 12014 9977 12066 9986
rect 12014 9943 12023 9977
rect 12023 9943 12057 9977
rect 12057 9943 12066 9977
rect 12014 9934 12066 9943
rect 12014 9817 12066 9826
rect 12014 9783 12023 9817
rect 12023 9783 12057 9817
rect 12057 9783 12066 9817
rect 12014 9774 12066 9783
rect 12014 9497 12066 9506
rect 12014 9463 12023 9497
rect 12023 9463 12057 9497
rect 12057 9463 12066 9497
rect 12014 9454 12066 9463
rect 12014 9337 12066 9346
rect 12014 9303 12023 9337
rect 12023 9303 12057 9337
rect 12057 9303 12066 9337
rect 12014 9294 12066 9303
rect 12014 9017 12066 9026
rect 12014 8983 12023 9017
rect 12023 8983 12057 9017
rect 12057 8983 12066 9017
rect 12014 8974 12066 8983
rect 12014 8857 12066 8866
rect 12014 8823 12023 8857
rect 12023 8823 12057 8857
rect 12057 8823 12066 8857
rect 12014 8814 12066 8823
rect 12014 8697 12066 8706
rect 12014 8663 12023 8697
rect 12023 8663 12057 8697
rect 12057 8663 12066 8697
rect 12014 8654 12066 8663
rect 12014 8537 12066 8546
rect 12014 8503 12023 8537
rect 12023 8503 12057 8537
rect 12057 8503 12066 8537
rect 12014 8494 12066 8503
rect 12014 8377 12066 8386
rect 12014 8343 12023 8377
rect 12023 8343 12057 8377
rect 12057 8343 12066 8377
rect 12014 8334 12066 8343
rect 12014 8217 12066 8226
rect 12014 8183 12023 8217
rect 12023 8183 12057 8217
rect 12057 8183 12066 8217
rect 12014 8174 12066 8183
rect 12014 8057 12066 8066
rect 12014 8023 12023 8057
rect 12023 8023 12057 8057
rect 12057 8023 12066 8057
rect 12014 8014 12066 8023
rect 12014 7897 12066 7906
rect 12014 7863 12023 7897
rect 12023 7863 12057 7897
rect 12057 7863 12066 7897
rect 12014 7854 12066 7863
rect 12014 7737 12066 7746
rect 12014 7703 12023 7737
rect 12023 7703 12057 7737
rect 12057 7703 12066 7737
rect 12014 7694 12066 7703
rect 12014 7417 12066 7426
rect 12014 7383 12023 7417
rect 12023 7383 12057 7417
rect 12057 7383 12066 7417
rect 12014 7374 12066 7383
rect 12014 7257 12066 7266
rect 12014 7223 12023 7257
rect 12023 7223 12057 7257
rect 12057 7223 12066 7257
rect 12014 7214 12066 7223
rect 12014 6937 12066 6946
rect 12014 6903 12023 6937
rect 12023 6903 12057 6937
rect 12057 6903 12066 6937
rect 12014 6894 12066 6903
rect 12014 6777 12066 6786
rect 12014 6743 12023 6777
rect 12023 6743 12057 6777
rect 12057 6743 12066 6777
rect 12014 6734 12066 6743
rect 12014 6457 12066 6466
rect 12014 6423 12023 6457
rect 12023 6423 12057 6457
rect 12057 6423 12066 6457
rect 12014 6414 12066 6423
rect 12014 6297 12066 6306
rect 12014 6263 12023 6297
rect 12023 6263 12057 6297
rect 12057 6263 12066 6297
rect 12014 6254 12066 6263
rect 12014 6137 12066 6146
rect 12014 6103 12023 6137
rect 12023 6103 12057 6137
rect 12057 6103 12066 6137
rect 12014 6094 12066 6103
rect 12014 5977 12066 5986
rect 12014 5943 12023 5977
rect 12023 5943 12057 5977
rect 12057 5943 12066 5977
rect 12014 5934 12066 5943
rect 12014 5817 12066 5826
rect 12014 5783 12023 5817
rect 12023 5783 12057 5817
rect 12057 5783 12066 5817
rect 12014 5774 12066 5783
rect 12014 5657 12066 5666
rect 12014 5623 12023 5657
rect 12023 5623 12057 5657
rect 12057 5623 12066 5657
rect 12014 5614 12066 5623
rect 12014 5497 12066 5506
rect 12014 5463 12023 5497
rect 12023 5463 12057 5497
rect 12057 5463 12066 5497
rect 12014 5454 12066 5463
rect 12014 5337 12066 5346
rect 12014 5303 12023 5337
rect 12023 5303 12057 5337
rect 12057 5303 12066 5337
rect 12014 5294 12066 5303
rect 12014 5177 12066 5186
rect 12014 5143 12023 5177
rect 12023 5143 12057 5177
rect 12057 5143 12066 5177
rect 12014 5134 12066 5143
rect 12014 5017 12066 5026
rect 12014 4983 12023 5017
rect 12023 4983 12057 5017
rect 12057 4983 12066 5017
rect 12014 4974 12066 4983
rect 12014 4857 12066 4866
rect 12014 4823 12023 4857
rect 12023 4823 12057 4857
rect 12057 4823 12066 4857
rect 12014 4814 12066 4823
rect 12014 4697 12066 4706
rect 12014 4663 12023 4697
rect 12023 4663 12057 4697
rect 12057 4663 12066 4697
rect 12014 4654 12066 4663
rect 12014 4537 12066 4546
rect 12014 4503 12023 4537
rect 12023 4503 12057 4537
rect 12057 4503 12066 4537
rect 12014 4494 12066 4503
rect 12014 4377 12066 4386
rect 12014 4343 12023 4377
rect 12023 4343 12057 4377
rect 12057 4343 12066 4377
rect 12014 4334 12066 4343
rect 12014 4217 12066 4226
rect 12014 4183 12023 4217
rect 12023 4183 12057 4217
rect 12057 4183 12066 4217
rect 12014 4174 12066 4183
rect 12014 4057 12066 4066
rect 12014 4023 12023 4057
rect 12023 4023 12057 4057
rect 12057 4023 12066 4057
rect 12014 4014 12066 4023
rect 12014 3897 12066 3906
rect 12014 3863 12023 3897
rect 12023 3863 12057 3897
rect 12057 3863 12066 3897
rect 12014 3854 12066 3863
rect 12014 3417 12066 3426
rect 12014 3383 12023 3417
rect 12023 3383 12057 3417
rect 12057 3383 12066 3417
rect 12014 3374 12066 3383
rect 12014 3257 12066 3266
rect 12014 3223 12023 3257
rect 12023 3223 12057 3257
rect 12057 3223 12066 3257
rect 12014 3214 12066 3223
rect 12014 3097 12066 3106
rect 12014 3063 12023 3097
rect 12023 3063 12057 3097
rect 12057 3063 12066 3097
rect 12014 3054 12066 3063
rect 12014 2937 12066 2946
rect 12014 2903 12023 2937
rect 12023 2903 12057 2937
rect 12057 2903 12066 2937
rect 12014 2894 12066 2903
rect 12014 2777 12066 2786
rect 12014 2743 12023 2777
rect 12023 2743 12057 2777
rect 12057 2743 12066 2777
rect 12014 2734 12066 2743
rect 12014 2617 12066 2626
rect 12014 2583 12023 2617
rect 12023 2583 12057 2617
rect 12057 2583 12066 2617
rect 12014 2574 12066 2583
rect 12014 2457 12066 2466
rect 12014 2423 12023 2457
rect 12023 2423 12057 2457
rect 12057 2423 12066 2457
rect 12014 2414 12066 2423
rect 12014 2297 12066 2306
rect 12014 2263 12023 2297
rect 12023 2263 12057 2297
rect 12057 2263 12066 2297
rect 12014 2254 12066 2263
rect 12014 2137 12066 2146
rect 12014 2103 12023 2137
rect 12023 2103 12057 2137
rect 12057 2103 12066 2137
rect 12014 2094 12066 2103
rect 12014 1977 12066 1986
rect 12014 1943 12023 1977
rect 12023 1943 12057 1977
rect 12057 1943 12066 1977
rect 12014 1934 12066 1943
rect 12014 1657 12066 1666
rect 12014 1623 12023 1657
rect 12023 1623 12057 1657
rect 12057 1623 12066 1657
rect 12014 1614 12066 1623
rect 12014 1497 12066 1506
rect 12014 1463 12023 1497
rect 12023 1463 12057 1497
rect 12057 1463 12066 1497
rect 12014 1454 12066 1463
rect 12014 1337 12066 1346
rect 12014 1303 12023 1337
rect 12023 1303 12057 1337
rect 12057 1303 12066 1337
rect 12014 1294 12066 1303
rect 12014 1177 12066 1186
rect 12014 1143 12023 1177
rect 12023 1143 12057 1177
rect 12057 1143 12066 1177
rect 12014 1134 12066 1143
rect 12014 1017 12066 1026
rect 12014 983 12023 1017
rect 12023 983 12057 1017
rect 12057 983 12066 1017
rect 12014 974 12066 983
rect 12014 537 12066 546
rect 12014 503 12023 537
rect 12023 503 12057 537
rect 12057 503 12066 537
rect 12014 494 12066 503
rect 12014 377 12066 386
rect 12014 343 12023 377
rect 12023 343 12057 377
rect 12057 343 12066 377
rect 12014 334 12066 343
rect 12014 217 12066 226
rect 12014 183 12023 217
rect 12023 183 12057 217
rect 12057 183 12066 217
rect 12014 174 12066 183
rect 12014 57 12066 66
rect 12014 23 12023 57
rect 12023 23 12057 57
rect 12057 23 12066 57
rect 12014 14 12066 23
rect 12334 31417 12386 31426
rect 12334 31383 12343 31417
rect 12343 31383 12377 31417
rect 12377 31383 12386 31417
rect 12334 31374 12386 31383
rect 12334 31257 12386 31266
rect 12334 31223 12343 31257
rect 12343 31223 12377 31257
rect 12377 31223 12386 31257
rect 12334 31214 12386 31223
rect 12334 31097 12386 31106
rect 12334 31063 12343 31097
rect 12343 31063 12377 31097
rect 12377 31063 12386 31097
rect 12334 31054 12386 31063
rect 12334 30937 12386 30946
rect 12334 30903 12343 30937
rect 12343 30903 12377 30937
rect 12377 30903 12386 30937
rect 12334 30894 12386 30903
rect 12334 30777 12386 30786
rect 12334 30743 12343 30777
rect 12343 30743 12377 30777
rect 12377 30743 12386 30777
rect 12334 30734 12386 30743
rect 12334 30617 12386 30626
rect 12334 30583 12343 30617
rect 12343 30583 12377 30617
rect 12377 30583 12386 30617
rect 12334 30574 12386 30583
rect 12334 30457 12386 30466
rect 12334 30423 12343 30457
rect 12343 30423 12377 30457
rect 12377 30423 12386 30457
rect 12334 30414 12386 30423
rect 12334 30297 12386 30306
rect 12334 30263 12343 30297
rect 12343 30263 12377 30297
rect 12377 30263 12386 30297
rect 12334 30254 12386 30263
rect 12334 29977 12386 29986
rect 12334 29943 12343 29977
rect 12343 29943 12377 29977
rect 12377 29943 12386 29977
rect 12334 29934 12386 29943
rect 12334 29817 12386 29826
rect 12334 29783 12343 29817
rect 12343 29783 12377 29817
rect 12377 29783 12386 29817
rect 12334 29774 12386 29783
rect 12334 29657 12386 29666
rect 12334 29623 12343 29657
rect 12343 29623 12377 29657
rect 12377 29623 12386 29657
rect 12334 29614 12386 29623
rect 12334 29497 12386 29506
rect 12334 29463 12343 29497
rect 12343 29463 12377 29497
rect 12377 29463 12386 29497
rect 12334 29454 12386 29463
rect 12334 29337 12386 29346
rect 12334 29303 12343 29337
rect 12343 29303 12377 29337
rect 12377 29303 12386 29337
rect 12334 29294 12386 29303
rect 12334 29177 12386 29186
rect 12334 29143 12343 29177
rect 12343 29143 12377 29177
rect 12377 29143 12386 29177
rect 12334 29134 12386 29143
rect 12334 29017 12386 29026
rect 12334 28983 12343 29017
rect 12343 28983 12377 29017
rect 12377 28983 12386 29017
rect 12334 28974 12386 28983
rect 12334 28857 12386 28866
rect 12334 28823 12343 28857
rect 12343 28823 12377 28857
rect 12377 28823 12386 28857
rect 12334 28814 12386 28823
rect 12334 28057 12386 28066
rect 12334 28023 12343 28057
rect 12343 28023 12377 28057
rect 12377 28023 12386 28057
rect 12334 28014 12386 28023
rect 12334 27897 12386 27906
rect 12334 27863 12343 27897
rect 12343 27863 12377 27897
rect 12377 27863 12386 27897
rect 12334 27854 12386 27863
rect 12334 27737 12386 27746
rect 12334 27703 12343 27737
rect 12343 27703 12377 27737
rect 12377 27703 12386 27737
rect 12334 27694 12386 27703
rect 12334 27577 12386 27586
rect 12334 27543 12343 27577
rect 12343 27543 12377 27577
rect 12377 27543 12386 27577
rect 12334 27534 12386 27543
rect 12334 27417 12386 27426
rect 12334 27383 12343 27417
rect 12343 27383 12377 27417
rect 12377 27383 12386 27417
rect 12334 27374 12386 27383
rect 12334 27257 12386 27266
rect 12334 27223 12343 27257
rect 12343 27223 12377 27257
rect 12377 27223 12386 27257
rect 12334 27214 12386 27223
rect 12334 27097 12386 27106
rect 12334 27063 12343 27097
rect 12343 27063 12377 27097
rect 12377 27063 12386 27097
rect 12334 27054 12386 27063
rect 12334 26937 12386 26946
rect 12334 26903 12343 26937
rect 12343 26903 12377 26937
rect 12377 26903 12386 26937
rect 12334 26894 12386 26903
rect 12334 26137 12386 26146
rect 12334 26103 12343 26137
rect 12343 26103 12377 26137
rect 12377 26103 12386 26137
rect 12334 26094 12386 26103
rect 12334 25977 12386 25986
rect 12334 25943 12343 25977
rect 12343 25943 12377 25977
rect 12377 25943 12386 25977
rect 12334 25934 12386 25943
rect 12334 25817 12386 25826
rect 12334 25783 12343 25817
rect 12343 25783 12377 25817
rect 12377 25783 12386 25817
rect 12334 25774 12386 25783
rect 12334 25657 12386 25666
rect 12334 25623 12343 25657
rect 12343 25623 12377 25657
rect 12377 25623 12386 25657
rect 12334 25614 12386 25623
rect 12334 25497 12386 25506
rect 12334 25463 12343 25497
rect 12343 25463 12377 25497
rect 12377 25463 12386 25497
rect 12334 25454 12386 25463
rect 12334 25337 12386 25346
rect 12334 25303 12343 25337
rect 12343 25303 12377 25337
rect 12377 25303 12386 25337
rect 12334 25294 12386 25303
rect 12334 25177 12386 25186
rect 12334 25143 12343 25177
rect 12343 25143 12377 25177
rect 12377 25143 12386 25177
rect 12334 25134 12386 25143
rect 12334 25017 12386 25026
rect 12334 24983 12343 25017
rect 12343 24983 12377 25017
rect 12377 24983 12386 25017
rect 12334 24974 12386 24983
rect 12334 24697 12386 24706
rect 12334 24663 12343 24697
rect 12343 24663 12377 24697
rect 12377 24663 12386 24697
rect 12334 24654 12386 24663
rect 12334 24537 12386 24546
rect 12334 24503 12343 24537
rect 12343 24503 12377 24537
rect 12377 24503 12386 24537
rect 12334 24494 12386 24503
rect 12334 24377 12386 24386
rect 12334 24343 12343 24377
rect 12343 24343 12377 24377
rect 12377 24343 12386 24377
rect 12334 24334 12386 24343
rect 12334 24217 12386 24226
rect 12334 24183 12343 24217
rect 12343 24183 12377 24217
rect 12377 24183 12386 24217
rect 12334 24174 12386 24183
rect 12334 24057 12386 24066
rect 12334 24023 12343 24057
rect 12343 24023 12377 24057
rect 12377 24023 12386 24057
rect 12334 24014 12386 24023
rect 12334 23897 12386 23906
rect 12334 23863 12343 23897
rect 12343 23863 12377 23897
rect 12377 23863 12386 23897
rect 12334 23854 12386 23863
rect 12334 23737 12386 23746
rect 12334 23703 12343 23737
rect 12343 23703 12377 23737
rect 12377 23703 12386 23737
rect 12334 23694 12386 23703
rect 12334 23577 12386 23586
rect 12334 23543 12343 23577
rect 12343 23543 12377 23577
rect 12377 23543 12386 23577
rect 12334 23534 12386 23543
rect 12334 23417 12386 23426
rect 12334 23383 12343 23417
rect 12343 23383 12377 23417
rect 12377 23383 12386 23417
rect 12334 23374 12386 23383
rect 12334 23257 12386 23266
rect 12334 23223 12343 23257
rect 12343 23223 12377 23257
rect 12377 23223 12386 23257
rect 12334 23214 12386 23223
rect 12334 23097 12386 23106
rect 12334 23063 12343 23097
rect 12343 23063 12377 23097
rect 12377 23063 12386 23097
rect 12334 23054 12386 23063
rect 12334 22937 12386 22946
rect 12334 22903 12343 22937
rect 12343 22903 12377 22937
rect 12377 22903 12386 22937
rect 12334 22894 12386 22903
rect 12334 22777 12386 22786
rect 12334 22743 12343 22777
rect 12343 22743 12377 22777
rect 12377 22743 12386 22777
rect 12334 22734 12386 22743
rect 12334 22617 12386 22626
rect 12334 22583 12343 22617
rect 12343 22583 12377 22617
rect 12377 22583 12386 22617
rect 12334 22574 12386 22583
rect 12334 22457 12386 22466
rect 12334 22423 12343 22457
rect 12343 22423 12377 22457
rect 12377 22423 12386 22457
rect 12334 22414 12386 22423
rect 12334 22297 12386 22306
rect 12334 22263 12343 22297
rect 12343 22263 12377 22297
rect 12377 22263 12386 22297
rect 12334 22254 12386 22263
rect 12334 22137 12386 22146
rect 12334 22103 12343 22137
rect 12343 22103 12377 22137
rect 12377 22103 12386 22137
rect 12334 22094 12386 22103
rect 12334 21817 12386 21826
rect 12334 21783 12343 21817
rect 12343 21783 12377 21817
rect 12377 21783 12386 21817
rect 12334 21774 12386 21783
rect 12334 21657 12386 21666
rect 12334 21623 12343 21657
rect 12343 21623 12377 21657
rect 12377 21623 12386 21657
rect 12334 21614 12386 21623
rect 12334 21497 12386 21506
rect 12334 21463 12343 21497
rect 12343 21463 12377 21497
rect 12377 21463 12386 21497
rect 12334 21454 12386 21463
rect 12334 21337 12386 21346
rect 12334 21303 12343 21337
rect 12343 21303 12377 21337
rect 12377 21303 12386 21337
rect 12334 21294 12386 21303
rect 12334 21177 12386 21186
rect 12334 21143 12343 21177
rect 12343 21143 12377 21177
rect 12377 21143 12386 21177
rect 12334 21134 12386 21143
rect 12334 21017 12386 21026
rect 12334 20983 12343 21017
rect 12343 20983 12377 21017
rect 12377 20983 12386 21017
rect 12334 20974 12386 20983
rect 12334 20857 12386 20866
rect 12334 20823 12343 20857
rect 12343 20823 12377 20857
rect 12377 20823 12386 20857
rect 12334 20814 12386 20823
rect 12334 20697 12386 20706
rect 12334 20663 12343 20697
rect 12343 20663 12377 20697
rect 12377 20663 12386 20697
rect 12334 20654 12386 20663
rect 12334 19897 12386 19906
rect 12334 19863 12343 19897
rect 12343 19863 12377 19897
rect 12377 19863 12386 19897
rect 12334 19854 12386 19863
rect 12334 19737 12386 19746
rect 12334 19703 12343 19737
rect 12343 19703 12377 19737
rect 12377 19703 12386 19737
rect 12334 19694 12386 19703
rect 12334 19577 12386 19586
rect 12334 19543 12343 19577
rect 12343 19543 12377 19577
rect 12377 19543 12386 19577
rect 12334 19534 12386 19543
rect 12334 19417 12386 19426
rect 12334 19383 12343 19417
rect 12343 19383 12377 19417
rect 12377 19383 12386 19417
rect 12334 19374 12386 19383
rect 12334 19257 12386 19266
rect 12334 19223 12343 19257
rect 12343 19223 12377 19257
rect 12377 19223 12386 19257
rect 12334 19214 12386 19223
rect 12334 19097 12386 19106
rect 12334 19063 12343 19097
rect 12343 19063 12377 19097
rect 12377 19063 12386 19097
rect 12334 19054 12386 19063
rect 12334 18937 12386 18946
rect 12334 18903 12343 18937
rect 12343 18903 12377 18937
rect 12377 18903 12386 18937
rect 12334 18894 12386 18903
rect 12334 18777 12386 18786
rect 12334 18743 12343 18777
rect 12343 18743 12377 18777
rect 12377 18743 12386 18777
rect 12334 18734 12386 18743
rect 12334 17977 12386 17986
rect 12334 17943 12343 17977
rect 12343 17943 12377 17977
rect 12377 17943 12386 17977
rect 12334 17934 12386 17943
rect 12334 17817 12386 17826
rect 12334 17783 12343 17817
rect 12343 17783 12377 17817
rect 12377 17783 12386 17817
rect 12334 17774 12386 17783
rect 12334 17657 12386 17666
rect 12334 17623 12343 17657
rect 12343 17623 12377 17657
rect 12377 17623 12386 17657
rect 12334 17614 12386 17623
rect 12334 17497 12386 17506
rect 12334 17463 12343 17497
rect 12343 17463 12377 17497
rect 12377 17463 12386 17497
rect 12334 17454 12386 17463
rect 12334 17337 12386 17346
rect 12334 17303 12343 17337
rect 12343 17303 12377 17337
rect 12377 17303 12386 17337
rect 12334 17294 12386 17303
rect 12334 17177 12386 17186
rect 12334 17143 12343 17177
rect 12343 17143 12377 17177
rect 12377 17143 12386 17177
rect 12334 17134 12386 17143
rect 12334 17017 12386 17026
rect 12334 16983 12343 17017
rect 12343 16983 12377 17017
rect 12377 16983 12386 17017
rect 12334 16974 12386 16983
rect 12334 16857 12386 16866
rect 12334 16823 12343 16857
rect 12343 16823 12377 16857
rect 12377 16823 12386 16857
rect 12334 16814 12386 16823
rect 12334 16537 12386 16546
rect 12334 16503 12343 16537
rect 12343 16503 12377 16537
rect 12377 16503 12386 16537
rect 12334 16494 12386 16503
rect 12334 16377 12386 16386
rect 12334 16343 12343 16377
rect 12343 16343 12377 16377
rect 12377 16343 12386 16377
rect 12334 16334 12386 16343
rect 12334 16217 12386 16226
rect 12334 16183 12343 16217
rect 12343 16183 12377 16217
rect 12377 16183 12386 16217
rect 12334 16174 12386 16183
rect 12334 16057 12386 16066
rect 12334 16023 12343 16057
rect 12343 16023 12377 16057
rect 12377 16023 12386 16057
rect 12334 16014 12386 16023
rect 12334 15897 12386 15906
rect 12334 15863 12343 15897
rect 12343 15863 12377 15897
rect 12377 15863 12386 15897
rect 12334 15854 12386 15863
rect 12334 15737 12386 15746
rect 12334 15703 12343 15737
rect 12343 15703 12377 15737
rect 12377 15703 12386 15737
rect 12334 15694 12386 15703
rect 12334 15577 12386 15586
rect 12334 15543 12343 15577
rect 12343 15543 12377 15577
rect 12377 15543 12386 15577
rect 12334 15534 12386 15543
rect 12334 15417 12386 15426
rect 12334 15383 12343 15417
rect 12343 15383 12377 15417
rect 12377 15383 12386 15417
rect 12334 15374 12386 15383
rect 12334 15257 12386 15266
rect 12334 15223 12343 15257
rect 12343 15223 12377 15257
rect 12377 15223 12386 15257
rect 12334 15214 12386 15223
rect 12334 15097 12386 15106
rect 12334 15063 12343 15097
rect 12343 15063 12377 15097
rect 12377 15063 12386 15097
rect 12334 15054 12386 15063
rect 12334 14937 12386 14946
rect 12334 14903 12343 14937
rect 12343 14903 12377 14937
rect 12377 14903 12386 14937
rect 12334 14894 12386 14903
rect 12334 14777 12386 14786
rect 12334 14743 12343 14777
rect 12343 14743 12377 14777
rect 12377 14743 12386 14777
rect 12334 14734 12386 14743
rect 12334 14617 12386 14626
rect 12334 14583 12343 14617
rect 12343 14583 12377 14617
rect 12377 14583 12386 14617
rect 12334 14574 12386 14583
rect 12334 14457 12386 14466
rect 12334 14423 12343 14457
rect 12343 14423 12377 14457
rect 12377 14423 12386 14457
rect 12334 14414 12386 14423
rect 12334 14297 12386 14306
rect 12334 14263 12343 14297
rect 12343 14263 12377 14297
rect 12377 14263 12386 14297
rect 12334 14254 12386 14263
rect 12334 14137 12386 14146
rect 12334 14103 12343 14137
rect 12343 14103 12377 14137
rect 12377 14103 12386 14137
rect 12334 14094 12386 14103
rect 12334 13977 12386 13986
rect 12334 13943 12343 13977
rect 12343 13943 12377 13977
rect 12377 13943 12386 13977
rect 12334 13934 12386 13943
rect 12334 13657 12386 13666
rect 12334 13623 12343 13657
rect 12343 13623 12377 13657
rect 12377 13623 12386 13657
rect 12334 13614 12386 13623
rect 12334 13497 12386 13506
rect 12334 13463 12343 13497
rect 12343 13463 12377 13497
rect 12377 13463 12386 13497
rect 12334 13454 12386 13463
rect 12334 13337 12386 13346
rect 12334 13303 12343 13337
rect 12343 13303 12377 13337
rect 12377 13303 12386 13337
rect 12334 13294 12386 13303
rect 12334 13177 12386 13186
rect 12334 13143 12343 13177
rect 12343 13143 12377 13177
rect 12377 13143 12386 13177
rect 12334 13134 12386 13143
rect 12334 13017 12386 13026
rect 12334 12983 12343 13017
rect 12343 12983 12377 13017
rect 12377 12983 12386 13017
rect 12334 12974 12386 12983
rect 12334 12857 12386 12866
rect 12334 12823 12343 12857
rect 12343 12823 12377 12857
rect 12377 12823 12386 12857
rect 12334 12814 12386 12823
rect 12334 12697 12386 12706
rect 12334 12663 12343 12697
rect 12343 12663 12377 12697
rect 12377 12663 12386 12697
rect 12334 12654 12386 12663
rect 12334 12537 12386 12546
rect 12334 12503 12343 12537
rect 12343 12503 12377 12537
rect 12377 12503 12386 12537
rect 12334 12494 12386 12503
rect 12334 11737 12386 11746
rect 12334 11703 12343 11737
rect 12343 11703 12377 11737
rect 12377 11703 12386 11737
rect 12334 11694 12386 11703
rect 12334 11577 12386 11586
rect 12334 11543 12343 11577
rect 12343 11543 12377 11577
rect 12377 11543 12386 11577
rect 12334 11534 12386 11543
rect 12334 11417 12386 11426
rect 12334 11383 12343 11417
rect 12343 11383 12377 11417
rect 12377 11383 12386 11417
rect 12334 11374 12386 11383
rect 12334 11257 12386 11266
rect 12334 11223 12343 11257
rect 12343 11223 12377 11257
rect 12377 11223 12386 11257
rect 12334 11214 12386 11223
rect 12334 11097 12386 11106
rect 12334 11063 12343 11097
rect 12343 11063 12377 11097
rect 12377 11063 12386 11097
rect 12334 11054 12386 11063
rect 12334 10937 12386 10946
rect 12334 10903 12343 10937
rect 12343 10903 12377 10937
rect 12377 10903 12386 10937
rect 12334 10894 12386 10903
rect 12334 10777 12386 10786
rect 12334 10743 12343 10777
rect 12343 10743 12377 10777
rect 12377 10743 12386 10777
rect 12334 10734 12386 10743
rect 12334 10617 12386 10626
rect 12334 10583 12343 10617
rect 12343 10583 12377 10617
rect 12377 10583 12386 10617
rect 12334 10574 12386 10583
rect 12334 10457 12386 10466
rect 12334 10423 12343 10457
rect 12343 10423 12377 10457
rect 12377 10423 12386 10457
rect 12334 10414 12386 10423
rect 12334 10297 12386 10306
rect 12334 10263 12343 10297
rect 12343 10263 12377 10297
rect 12377 10263 12386 10297
rect 12334 10254 12386 10263
rect 12334 10137 12386 10146
rect 12334 10103 12343 10137
rect 12343 10103 12377 10137
rect 12377 10103 12386 10137
rect 12334 10094 12386 10103
rect 12334 9977 12386 9986
rect 12334 9943 12343 9977
rect 12343 9943 12377 9977
rect 12377 9943 12386 9977
rect 12334 9934 12386 9943
rect 12334 9817 12386 9826
rect 12334 9783 12343 9817
rect 12343 9783 12377 9817
rect 12377 9783 12386 9817
rect 12334 9774 12386 9783
rect 12334 9497 12386 9506
rect 12334 9463 12343 9497
rect 12343 9463 12377 9497
rect 12377 9463 12386 9497
rect 12334 9454 12386 9463
rect 12334 9337 12386 9346
rect 12334 9303 12343 9337
rect 12343 9303 12377 9337
rect 12377 9303 12386 9337
rect 12334 9294 12386 9303
rect 12334 9017 12386 9026
rect 12334 8983 12343 9017
rect 12343 8983 12377 9017
rect 12377 8983 12386 9017
rect 12334 8974 12386 8983
rect 12334 8857 12386 8866
rect 12334 8823 12343 8857
rect 12343 8823 12377 8857
rect 12377 8823 12386 8857
rect 12334 8814 12386 8823
rect 12334 8697 12386 8706
rect 12334 8663 12343 8697
rect 12343 8663 12377 8697
rect 12377 8663 12386 8697
rect 12334 8654 12386 8663
rect 12334 8537 12386 8546
rect 12334 8503 12343 8537
rect 12343 8503 12377 8537
rect 12377 8503 12386 8537
rect 12334 8494 12386 8503
rect 12334 8377 12386 8386
rect 12334 8343 12343 8377
rect 12343 8343 12377 8377
rect 12377 8343 12386 8377
rect 12334 8334 12386 8343
rect 12334 8217 12386 8226
rect 12334 8183 12343 8217
rect 12343 8183 12377 8217
rect 12377 8183 12386 8217
rect 12334 8174 12386 8183
rect 12334 8057 12386 8066
rect 12334 8023 12343 8057
rect 12343 8023 12377 8057
rect 12377 8023 12386 8057
rect 12334 8014 12386 8023
rect 12334 7897 12386 7906
rect 12334 7863 12343 7897
rect 12343 7863 12377 7897
rect 12377 7863 12386 7897
rect 12334 7854 12386 7863
rect 12334 7737 12386 7746
rect 12334 7703 12343 7737
rect 12343 7703 12377 7737
rect 12377 7703 12386 7737
rect 12334 7694 12386 7703
rect 12334 7417 12386 7426
rect 12334 7383 12343 7417
rect 12343 7383 12377 7417
rect 12377 7383 12386 7417
rect 12334 7374 12386 7383
rect 12334 7257 12386 7266
rect 12334 7223 12343 7257
rect 12343 7223 12377 7257
rect 12377 7223 12386 7257
rect 12334 7214 12386 7223
rect 12334 6937 12386 6946
rect 12334 6903 12343 6937
rect 12343 6903 12377 6937
rect 12377 6903 12386 6937
rect 12334 6894 12386 6903
rect 12334 6777 12386 6786
rect 12334 6743 12343 6777
rect 12343 6743 12377 6777
rect 12377 6743 12386 6777
rect 12334 6734 12386 6743
rect 12334 6457 12386 6466
rect 12334 6423 12343 6457
rect 12343 6423 12377 6457
rect 12377 6423 12386 6457
rect 12334 6414 12386 6423
rect 12334 6297 12386 6306
rect 12334 6263 12343 6297
rect 12343 6263 12377 6297
rect 12377 6263 12386 6297
rect 12334 6254 12386 6263
rect 12334 6137 12386 6146
rect 12334 6103 12343 6137
rect 12343 6103 12377 6137
rect 12377 6103 12386 6137
rect 12334 6094 12386 6103
rect 12334 5977 12386 5986
rect 12334 5943 12343 5977
rect 12343 5943 12377 5977
rect 12377 5943 12386 5977
rect 12334 5934 12386 5943
rect 12334 5817 12386 5826
rect 12334 5783 12343 5817
rect 12343 5783 12377 5817
rect 12377 5783 12386 5817
rect 12334 5774 12386 5783
rect 12334 5657 12386 5666
rect 12334 5623 12343 5657
rect 12343 5623 12377 5657
rect 12377 5623 12386 5657
rect 12334 5614 12386 5623
rect 12334 5497 12386 5506
rect 12334 5463 12343 5497
rect 12343 5463 12377 5497
rect 12377 5463 12386 5497
rect 12334 5454 12386 5463
rect 12334 5337 12386 5346
rect 12334 5303 12343 5337
rect 12343 5303 12377 5337
rect 12377 5303 12386 5337
rect 12334 5294 12386 5303
rect 12334 5177 12386 5186
rect 12334 5143 12343 5177
rect 12343 5143 12377 5177
rect 12377 5143 12386 5177
rect 12334 5134 12386 5143
rect 12334 5017 12386 5026
rect 12334 4983 12343 5017
rect 12343 4983 12377 5017
rect 12377 4983 12386 5017
rect 12334 4974 12386 4983
rect 12334 4857 12386 4866
rect 12334 4823 12343 4857
rect 12343 4823 12377 4857
rect 12377 4823 12386 4857
rect 12334 4814 12386 4823
rect 12334 4697 12386 4706
rect 12334 4663 12343 4697
rect 12343 4663 12377 4697
rect 12377 4663 12386 4697
rect 12334 4654 12386 4663
rect 12334 4537 12386 4546
rect 12334 4503 12343 4537
rect 12343 4503 12377 4537
rect 12377 4503 12386 4537
rect 12334 4494 12386 4503
rect 12334 4377 12386 4386
rect 12334 4343 12343 4377
rect 12343 4343 12377 4377
rect 12377 4343 12386 4377
rect 12334 4334 12386 4343
rect 12334 4217 12386 4226
rect 12334 4183 12343 4217
rect 12343 4183 12377 4217
rect 12377 4183 12386 4217
rect 12334 4174 12386 4183
rect 12334 4057 12386 4066
rect 12334 4023 12343 4057
rect 12343 4023 12377 4057
rect 12377 4023 12386 4057
rect 12334 4014 12386 4023
rect 12334 3897 12386 3906
rect 12334 3863 12343 3897
rect 12343 3863 12377 3897
rect 12377 3863 12386 3897
rect 12334 3854 12386 3863
rect 12334 3417 12386 3426
rect 12334 3383 12343 3417
rect 12343 3383 12377 3417
rect 12377 3383 12386 3417
rect 12334 3374 12386 3383
rect 12334 3257 12386 3266
rect 12334 3223 12343 3257
rect 12343 3223 12377 3257
rect 12377 3223 12386 3257
rect 12334 3214 12386 3223
rect 12334 3097 12386 3106
rect 12334 3063 12343 3097
rect 12343 3063 12377 3097
rect 12377 3063 12386 3097
rect 12334 3054 12386 3063
rect 12334 2937 12386 2946
rect 12334 2903 12343 2937
rect 12343 2903 12377 2937
rect 12377 2903 12386 2937
rect 12334 2894 12386 2903
rect 12334 2777 12386 2786
rect 12334 2743 12343 2777
rect 12343 2743 12377 2777
rect 12377 2743 12386 2777
rect 12334 2734 12386 2743
rect 12334 2617 12386 2626
rect 12334 2583 12343 2617
rect 12343 2583 12377 2617
rect 12377 2583 12386 2617
rect 12334 2574 12386 2583
rect 12334 2457 12386 2466
rect 12334 2423 12343 2457
rect 12343 2423 12377 2457
rect 12377 2423 12386 2457
rect 12334 2414 12386 2423
rect 12334 2297 12386 2306
rect 12334 2263 12343 2297
rect 12343 2263 12377 2297
rect 12377 2263 12386 2297
rect 12334 2254 12386 2263
rect 12334 2137 12386 2146
rect 12334 2103 12343 2137
rect 12343 2103 12377 2137
rect 12377 2103 12386 2137
rect 12334 2094 12386 2103
rect 12334 1977 12386 1986
rect 12334 1943 12343 1977
rect 12343 1943 12377 1977
rect 12377 1943 12386 1977
rect 12334 1934 12386 1943
rect 12334 1657 12386 1666
rect 12334 1623 12343 1657
rect 12343 1623 12377 1657
rect 12377 1623 12386 1657
rect 12334 1614 12386 1623
rect 12334 1497 12386 1506
rect 12334 1463 12343 1497
rect 12343 1463 12377 1497
rect 12377 1463 12386 1497
rect 12334 1454 12386 1463
rect 12334 1337 12386 1346
rect 12334 1303 12343 1337
rect 12343 1303 12377 1337
rect 12377 1303 12386 1337
rect 12334 1294 12386 1303
rect 12334 1177 12386 1186
rect 12334 1143 12343 1177
rect 12343 1143 12377 1177
rect 12377 1143 12386 1177
rect 12334 1134 12386 1143
rect 12334 1017 12386 1026
rect 12334 983 12343 1017
rect 12343 983 12377 1017
rect 12377 983 12386 1017
rect 12334 974 12386 983
rect 12334 537 12386 546
rect 12334 503 12343 537
rect 12343 503 12377 537
rect 12377 503 12386 537
rect 12334 494 12386 503
rect 12334 377 12386 386
rect 12334 343 12343 377
rect 12343 343 12377 377
rect 12377 343 12386 377
rect 12334 334 12386 343
rect 12334 217 12386 226
rect 12334 183 12343 217
rect 12343 183 12377 217
rect 12377 183 12386 217
rect 12334 174 12386 183
rect 12334 57 12386 66
rect 12334 23 12343 57
rect 12343 23 12377 57
rect 12377 23 12386 57
rect 12334 14 12386 23
<< metal2 >>
rect 8480 31428 8880 31440
rect 8480 31372 8492 31428
rect 8548 31372 8812 31428
rect 8868 31372 8880 31428
rect 8480 31360 8880 31372
rect 8960 31428 9360 31440
rect 8960 31372 8972 31428
rect 9028 31372 9292 31428
rect 9348 31372 9360 31428
rect 8960 31360 9360 31372
rect 9440 31428 11440 31440
rect 9440 31372 9452 31428
rect 9508 31372 9772 31428
rect 9828 31372 10092 31428
rect 10148 31372 10412 31428
rect 10468 31372 10732 31428
rect 10788 31372 11052 31428
rect 11108 31372 11372 31428
rect 11428 31372 11440 31428
rect 9440 31360 11440 31372
rect 11520 31428 11920 31440
rect 11520 31372 11532 31428
rect 11588 31372 11852 31428
rect 11908 31372 11920 31428
rect 11520 31360 11920 31372
rect 12000 31428 12400 31440
rect 12000 31372 12012 31428
rect 12068 31372 12332 31428
rect 12388 31372 12400 31428
rect 12000 31360 12400 31372
rect 8480 31268 8880 31280
rect 8480 31212 8492 31268
rect 8548 31212 8812 31268
rect 8868 31212 8880 31268
rect 8480 31200 8880 31212
rect 8960 31268 9360 31280
rect 8960 31212 8972 31268
rect 9028 31212 9292 31268
rect 9348 31212 9360 31268
rect 8960 31200 9360 31212
rect 9440 31268 11440 31280
rect 9440 31212 9452 31268
rect 9508 31212 9772 31268
rect 9828 31212 10092 31268
rect 10148 31212 10412 31268
rect 10468 31212 10732 31268
rect 10788 31212 11052 31268
rect 11108 31212 11372 31268
rect 11428 31212 11440 31268
rect 9440 31200 11440 31212
rect 11520 31268 11920 31280
rect 11520 31212 11532 31268
rect 11588 31212 11852 31268
rect 11908 31212 11920 31268
rect 11520 31200 11920 31212
rect 12000 31268 12400 31280
rect 12000 31212 12012 31268
rect 12068 31212 12332 31268
rect 12388 31212 12400 31268
rect 12000 31200 12400 31212
rect 8480 31108 8880 31120
rect 8480 31052 8492 31108
rect 8548 31052 8812 31108
rect 8868 31052 8880 31108
rect 8480 31040 8880 31052
rect 8960 31108 9360 31120
rect 8960 31052 8972 31108
rect 9028 31052 9292 31108
rect 9348 31052 9360 31108
rect 8960 31040 9360 31052
rect 9440 31108 11440 31120
rect 9440 31052 9452 31108
rect 9508 31052 9772 31108
rect 9828 31052 10092 31108
rect 10148 31052 10412 31108
rect 10468 31052 10732 31108
rect 10788 31052 11052 31108
rect 11108 31052 11372 31108
rect 11428 31052 11440 31108
rect 9440 31040 11440 31052
rect 11520 31108 11920 31120
rect 11520 31052 11532 31108
rect 11588 31052 11852 31108
rect 11908 31052 11920 31108
rect 11520 31040 11920 31052
rect 12000 31108 12400 31120
rect 12000 31052 12012 31108
rect 12068 31052 12332 31108
rect 12388 31052 12400 31108
rect 12000 31040 12400 31052
rect 8480 30948 8880 30960
rect 8480 30892 8492 30948
rect 8548 30892 8812 30948
rect 8868 30892 8880 30948
rect 8480 30880 8880 30892
rect 8960 30948 9360 30960
rect 8960 30892 8972 30948
rect 9028 30892 9292 30948
rect 9348 30892 9360 30948
rect 8960 30880 9360 30892
rect 9440 30948 11440 30960
rect 9440 30892 9452 30948
rect 9508 30892 9772 30948
rect 9828 30892 10092 30948
rect 10148 30892 10412 30948
rect 10468 30892 10732 30948
rect 10788 30892 11052 30948
rect 11108 30892 11372 30948
rect 11428 30892 11440 30948
rect 9440 30880 11440 30892
rect 11520 30948 11920 30960
rect 11520 30892 11532 30948
rect 11588 30892 11852 30948
rect 11908 30892 11920 30948
rect 11520 30880 11920 30892
rect 12000 30948 12400 30960
rect 12000 30892 12012 30948
rect 12068 30892 12332 30948
rect 12388 30892 12400 30948
rect 12000 30880 12400 30892
rect 8480 30788 8880 30800
rect 8480 30732 8492 30788
rect 8548 30732 8812 30788
rect 8868 30732 8880 30788
rect 8480 30720 8880 30732
rect 8960 30788 9360 30800
rect 8960 30732 8972 30788
rect 9028 30732 9292 30788
rect 9348 30732 9360 30788
rect 8960 30720 9360 30732
rect 9440 30788 11440 30800
rect 9440 30732 9452 30788
rect 9508 30732 9772 30788
rect 9828 30732 10092 30788
rect 10148 30732 10412 30788
rect 10468 30732 10732 30788
rect 10788 30732 11052 30788
rect 11108 30732 11372 30788
rect 11428 30732 11440 30788
rect 9440 30720 11440 30732
rect 11520 30788 11920 30800
rect 11520 30732 11532 30788
rect 11588 30732 11852 30788
rect 11908 30732 11920 30788
rect 11520 30720 11920 30732
rect 12000 30788 12400 30800
rect 12000 30732 12012 30788
rect 12068 30732 12332 30788
rect 12388 30732 12400 30788
rect 12000 30720 12400 30732
rect 8480 30628 8880 30640
rect 8480 30572 8492 30628
rect 8548 30572 8812 30628
rect 8868 30572 8880 30628
rect 8480 30560 8880 30572
rect 8960 30628 9360 30640
rect 8960 30572 8972 30628
rect 9028 30572 9292 30628
rect 9348 30572 9360 30628
rect 8960 30560 9360 30572
rect 9440 30628 11440 30640
rect 9440 30572 9452 30628
rect 9508 30572 9772 30628
rect 9828 30572 10092 30628
rect 10148 30572 10412 30628
rect 10468 30572 10732 30628
rect 10788 30572 11052 30628
rect 11108 30572 11372 30628
rect 11428 30572 11440 30628
rect 9440 30560 11440 30572
rect 11520 30628 11920 30640
rect 11520 30572 11532 30628
rect 11588 30572 11852 30628
rect 11908 30572 11920 30628
rect 11520 30560 11920 30572
rect 12000 30628 12400 30640
rect 12000 30572 12012 30628
rect 12068 30572 12332 30628
rect 12388 30572 12400 30628
rect 12000 30560 12400 30572
rect 8480 30468 8880 30480
rect 8480 30412 8492 30468
rect 8548 30412 8812 30468
rect 8868 30412 8880 30468
rect 8480 30400 8880 30412
rect 8960 30468 9360 30480
rect 8960 30412 8972 30468
rect 9028 30412 9292 30468
rect 9348 30412 9360 30468
rect 8960 30400 9360 30412
rect 9440 30468 11440 30480
rect 9440 30412 9452 30468
rect 9508 30412 9772 30468
rect 9828 30412 10092 30468
rect 10148 30412 10412 30468
rect 10468 30412 10732 30468
rect 10788 30412 11052 30468
rect 11108 30412 11372 30468
rect 11428 30412 11440 30468
rect 9440 30400 11440 30412
rect 11520 30468 11920 30480
rect 11520 30412 11532 30468
rect 11588 30412 11852 30468
rect 11908 30412 11920 30468
rect 11520 30400 11920 30412
rect 12000 30468 12400 30480
rect 12000 30412 12012 30468
rect 12068 30412 12332 30468
rect 12388 30412 12400 30468
rect 12000 30400 12400 30412
rect 8480 30308 8880 30320
rect 8480 30252 8492 30308
rect 8548 30252 8812 30308
rect 8868 30252 8880 30308
rect 8480 30240 8880 30252
rect 8960 30308 9360 30320
rect 8960 30252 8972 30308
rect 9028 30252 9292 30308
rect 9348 30252 9360 30308
rect 8960 30240 9360 30252
rect 9440 30308 11440 30320
rect 9440 30252 9452 30308
rect 9508 30252 9772 30308
rect 9828 30252 10092 30308
rect 10148 30252 10412 30308
rect 10468 30252 10732 30308
rect 10788 30252 11052 30308
rect 11108 30252 11372 30308
rect 11428 30252 11440 30308
rect 9440 30240 11440 30252
rect 11520 30308 11920 30320
rect 11520 30252 11532 30308
rect 11588 30252 11852 30308
rect 11908 30252 11920 30308
rect 11520 30240 11920 30252
rect 12000 30308 12400 30320
rect 12000 30252 12012 30308
rect 12068 30252 12332 30308
rect 12388 30252 12400 30308
rect 12000 30240 12400 30252
rect 0 30148 20880 30160
rect 0 30092 9132 30148
rect 9188 30092 20880 30148
rect 0 30080 20880 30092
rect 8480 29988 8880 30000
rect 8480 29932 8492 29988
rect 8548 29932 8812 29988
rect 8868 29932 8880 29988
rect 8480 29920 8880 29932
rect 8960 29988 9360 30000
rect 8960 29932 8972 29988
rect 9028 29932 9292 29988
rect 9348 29932 9360 29988
rect 8960 29920 9360 29932
rect 9440 29988 11440 30000
rect 9440 29932 9452 29988
rect 9508 29932 9772 29988
rect 9828 29932 10092 29988
rect 10148 29932 10412 29988
rect 10468 29932 10732 29988
rect 10788 29932 11052 29988
rect 11108 29932 11372 29988
rect 11428 29932 11440 29988
rect 9440 29920 11440 29932
rect 11520 29988 11920 30000
rect 11520 29932 11532 29988
rect 11588 29932 11852 29988
rect 11908 29932 11920 29988
rect 11520 29920 11920 29932
rect 12000 29988 12400 30000
rect 12000 29932 12012 29988
rect 12068 29932 12332 29988
rect 12388 29932 12400 29988
rect 12000 29920 12400 29932
rect 8480 29828 8880 29840
rect 8480 29772 8492 29828
rect 8548 29772 8812 29828
rect 8868 29772 8880 29828
rect 8480 29760 8880 29772
rect 8960 29828 9360 29840
rect 8960 29772 8972 29828
rect 9028 29772 9292 29828
rect 9348 29772 9360 29828
rect 8960 29760 9360 29772
rect 9440 29828 11440 29840
rect 9440 29772 9452 29828
rect 9508 29772 9772 29828
rect 9828 29772 10092 29828
rect 10148 29772 10412 29828
rect 10468 29772 10732 29828
rect 10788 29772 11052 29828
rect 11108 29772 11372 29828
rect 11428 29772 11440 29828
rect 9440 29760 11440 29772
rect 11520 29828 11920 29840
rect 11520 29772 11532 29828
rect 11588 29772 11852 29828
rect 11908 29772 11920 29828
rect 11520 29760 11920 29772
rect 12000 29828 12400 29840
rect 12000 29772 12012 29828
rect 12068 29772 12332 29828
rect 12388 29772 12400 29828
rect 12000 29760 12400 29772
rect 8480 29668 8880 29680
rect 8480 29612 8492 29668
rect 8548 29612 8812 29668
rect 8868 29612 8880 29668
rect 8480 29600 8880 29612
rect 8960 29668 9360 29680
rect 8960 29612 8972 29668
rect 9028 29612 9292 29668
rect 9348 29612 9360 29668
rect 8960 29600 9360 29612
rect 9440 29668 11440 29680
rect 9440 29612 9452 29668
rect 9508 29612 9772 29668
rect 9828 29612 10092 29668
rect 10148 29612 10412 29668
rect 10468 29612 10732 29668
rect 10788 29612 11052 29668
rect 11108 29612 11372 29668
rect 11428 29612 11440 29668
rect 9440 29600 11440 29612
rect 11520 29668 11920 29680
rect 11520 29612 11532 29668
rect 11588 29612 11852 29668
rect 11908 29612 11920 29668
rect 11520 29600 11920 29612
rect 12000 29668 12400 29680
rect 12000 29612 12012 29668
rect 12068 29612 12332 29668
rect 12388 29612 12400 29668
rect 12000 29600 12400 29612
rect 8480 29508 8880 29520
rect 8480 29452 8492 29508
rect 8548 29452 8812 29508
rect 8868 29452 8880 29508
rect 8480 29440 8880 29452
rect 8960 29508 9360 29520
rect 8960 29452 8972 29508
rect 9028 29452 9292 29508
rect 9348 29452 9360 29508
rect 8960 29440 9360 29452
rect 9440 29508 11440 29520
rect 9440 29452 9452 29508
rect 9508 29452 9772 29508
rect 9828 29452 10092 29508
rect 10148 29452 10412 29508
rect 10468 29452 10732 29508
rect 10788 29452 11052 29508
rect 11108 29452 11372 29508
rect 11428 29452 11440 29508
rect 9440 29440 11440 29452
rect 11520 29508 11920 29520
rect 11520 29452 11532 29508
rect 11588 29452 11852 29508
rect 11908 29452 11920 29508
rect 11520 29440 11920 29452
rect 12000 29508 12400 29520
rect 12000 29452 12012 29508
rect 12068 29452 12332 29508
rect 12388 29452 12400 29508
rect 12000 29440 12400 29452
rect 8480 29348 8880 29360
rect 8480 29292 8492 29348
rect 8548 29292 8812 29348
rect 8868 29292 8880 29348
rect 8480 29280 8880 29292
rect 8960 29348 9360 29360
rect 8960 29292 8972 29348
rect 9028 29292 9292 29348
rect 9348 29292 9360 29348
rect 8960 29280 9360 29292
rect 9440 29348 11440 29360
rect 9440 29292 9452 29348
rect 9508 29292 9772 29348
rect 9828 29292 10092 29348
rect 10148 29292 10412 29348
rect 10468 29292 10732 29348
rect 10788 29292 11052 29348
rect 11108 29292 11372 29348
rect 11428 29292 11440 29348
rect 9440 29280 11440 29292
rect 11520 29348 11920 29360
rect 11520 29292 11532 29348
rect 11588 29292 11852 29348
rect 11908 29292 11920 29348
rect 11520 29280 11920 29292
rect 12000 29348 12400 29360
rect 12000 29292 12012 29348
rect 12068 29292 12332 29348
rect 12388 29292 12400 29348
rect 12000 29280 12400 29292
rect 8480 29188 8880 29200
rect 8480 29132 8492 29188
rect 8548 29132 8812 29188
rect 8868 29132 8880 29188
rect 8480 29120 8880 29132
rect 8960 29188 9360 29200
rect 8960 29132 8972 29188
rect 9028 29132 9292 29188
rect 9348 29132 9360 29188
rect 8960 29120 9360 29132
rect 9440 29188 11440 29200
rect 9440 29132 9452 29188
rect 9508 29132 9772 29188
rect 9828 29132 10092 29188
rect 10148 29132 10412 29188
rect 10468 29132 10732 29188
rect 10788 29132 11052 29188
rect 11108 29132 11372 29188
rect 11428 29132 11440 29188
rect 9440 29120 11440 29132
rect 11520 29188 11920 29200
rect 11520 29132 11532 29188
rect 11588 29132 11852 29188
rect 11908 29132 11920 29188
rect 11520 29120 11920 29132
rect 12000 29188 12400 29200
rect 12000 29132 12012 29188
rect 12068 29132 12332 29188
rect 12388 29132 12400 29188
rect 12000 29120 12400 29132
rect 8480 29028 8880 29040
rect 8480 28972 8492 29028
rect 8548 28972 8812 29028
rect 8868 28972 8880 29028
rect 8480 28960 8880 28972
rect 8960 29028 9360 29040
rect 8960 28972 8972 29028
rect 9028 28972 9292 29028
rect 9348 28972 9360 29028
rect 8960 28960 9360 28972
rect 9440 29028 11440 29040
rect 9440 28972 9452 29028
rect 9508 28972 9772 29028
rect 9828 28972 10092 29028
rect 10148 28972 10412 29028
rect 10468 28972 10732 29028
rect 10788 28972 11052 29028
rect 11108 28972 11372 29028
rect 11428 28972 11440 29028
rect 9440 28960 11440 28972
rect 11520 29028 11920 29040
rect 11520 28972 11532 29028
rect 11588 28972 11852 29028
rect 11908 28972 11920 29028
rect 11520 28960 11920 28972
rect 12000 29028 12400 29040
rect 12000 28972 12012 29028
rect 12068 28972 12332 29028
rect 12388 28972 12400 29028
rect 12000 28960 12400 28972
rect 8480 28868 8880 28880
rect 8480 28812 8492 28868
rect 8548 28812 8812 28868
rect 8868 28812 8880 28868
rect 8480 28800 8880 28812
rect 8960 28868 9360 28880
rect 8960 28812 8972 28868
rect 9028 28812 9292 28868
rect 9348 28812 9360 28868
rect 8960 28800 9360 28812
rect 9440 28868 11440 28880
rect 9440 28812 9452 28868
rect 9508 28812 9772 28868
rect 9828 28812 10092 28868
rect 10148 28812 10412 28868
rect 10468 28812 10732 28868
rect 10788 28812 11052 28868
rect 11108 28812 11372 28868
rect 11428 28812 11440 28868
rect 9440 28800 11440 28812
rect 11520 28868 11920 28880
rect 11520 28812 11532 28868
rect 11588 28812 11852 28868
rect 11908 28812 11920 28868
rect 11520 28800 11920 28812
rect 12000 28868 12400 28880
rect 12000 28812 12012 28868
rect 12068 28812 12332 28868
rect 12388 28812 12400 28868
rect 12000 28800 12400 28812
rect 0 28628 20880 28640
rect 0 28572 10572 28628
rect 10628 28572 20880 28628
rect 0 28560 20880 28572
rect 0 28308 10000 28320
rect 0 28252 9932 28308
rect 9988 28252 10000 28308
rect 0 28240 10000 28252
rect 10880 28308 20880 28320
rect 10880 28252 10892 28308
rect 10948 28252 20880 28308
rect 10880 28240 20880 28252
rect 8480 28068 8880 28080
rect 8480 28012 8492 28068
rect 8548 28012 8812 28068
rect 8868 28012 8880 28068
rect 8480 28000 8880 28012
rect 8960 28068 9360 28080
rect 8960 28012 8972 28068
rect 9028 28012 9292 28068
rect 9348 28012 9360 28068
rect 8960 28000 9360 28012
rect 9440 28068 11440 28080
rect 9440 28012 9452 28068
rect 9508 28012 9772 28068
rect 9828 28012 10092 28068
rect 10148 28012 10412 28068
rect 10468 28012 10732 28068
rect 10788 28012 11052 28068
rect 11108 28012 11372 28068
rect 11428 28012 11440 28068
rect 9440 28000 11440 28012
rect 11520 28068 11920 28080
rect 11520 28012 11532 28068
rect 11588 28012 11852 28068
rect 11908 28012 11920 28068
rect 11520 28000 11920 28012
rect 12000 28068 12400 28080
rect 12000 28012 12012 28068
rect 12068 28012 12332 28068
rect 12388 28012 12400 28068
rect 12000 28000 12400 28012
rect 8480 27908 8880 27920
rect 8480 27852 8492 27908
rect 8548 27852 8812 27908
rect 8868 27852 8880 27908
rect 8480 27840 8880 27852
rect 8960 27908 9360 27920
rect 8960 27852 8972 27908
rect 9028 27852 9292 27908
rect 9348 27852 9360 27908
rect 8960 27840 9360 27852
rect 9440 27908 11440 27920
rect 9440 27852 9452 27908
rect 9508 27852 9772 27908
rect 9828 27852 10092 27908
rect 10148 27852 10412 27908
rect 10468 27852 10732 27908
rect 10788 27852 11052 27908
rect 11108 27852 11372 27908
rect 11428 27852 11440 27908
rect 9440 27840 11440 27852
rect 11520 27908 11920 27920
rect 11520 27852 11532 27908
rect 11588 27852 11852 27908
rect 11908 27852 11920 27908
rect 11520 27840 11920 27852
rect 12000 27908 12400 27920
rect 12000 27852 12012 27908
rect 12068 27852 12332 27908
rect 12388 27852 12400 27908
rect 12000 27840 12400 27852
rect 8480 27748 8880 27760
rect 8480 27692 8492 27748
rect 8548 27692 8812 27748
rect 8868 27692 8880 27748
rect 8480 27680 8880 27692
rect 8960 27748 9360 27760
rect 8960 27692 8972 27748
rect 9028 27692 9292 27748
rect 9348 27692 9360 27748
rect 8960 27680 9360 27692
rect 9440 27748 11440 27760
rect 9440 27692 9452 27748
rect 9508 27692 9772 27748
rect 9828 27692 10092 27748
rect 10148 27692 10412 27748
rect 10468 27692 10732 27748
rect 10788 27692 11052 27748
rect 11108 27692 11372 27748
rect 11428 27692 11440 27748
rect 9440 27680 11440 27692
rect 11520 27748 11920 27760
rect 11520 27692 11532 27748
rect 11588 27692 11852 27748
rect 11908 27692 11920 27748
rect 11520 27680 11920 27692
rect 12000 27748 12400 27760
rect 12000 27692 12012 27748
rect 12068 27692 12332 27748
rect 12388 27692 12400 27748
rect 12000 27680 12400 27692
rect 8480 27588 8880 27600
rect 8480 27532 8492 27588
rect 8548 27532 8812 27588
rect 8868 27532 8880 27588
rect 8480 27520 8880 27532
rect 8960 27588 9360 27600
rect 8960 27532 8972 27588
rect 9028 27532 9292 27588
rect 9348 27532 9360 27588
rect 8960 27520 9360 27532
rect 9440 27588 11440 27600
rect 9440 27532 9452 27588
rect 9508 27532 9772 27588
rect 9828 27532 10092 27588
rect 10148 27532 10412 27588
rect 10468 27532 10732 27588
rect 10788 27532 11052 27588
rect 11108 27532 11372 27588
rect 11428 27532 11440 27588
rect 9440 27520 11440 27532
rect 11520 27588 11920 27600
rect 11520 27532 11532 27588
rect 11588 27532 11852 27588
rect 11908 27532 11920 27588
rect 11520 27520 11920 27532
rect 12000 27588 12400 27600
rect 12000 27532 12012 27588
rect 12068 27532 12332 27588
rect 12388 27532 12400 27588
rect 12000 27520 12400 27532
rect 8480 27428 8880 27440
rect 8480 27372 8492 27428
rect 8548 27372 8812 27428
rect 8868 27372 8880 27428
rect 8480 27360 8880 27372
rect 8960 27428 9360 27440
rect 8960 27372 8972 27428
rect 9028 27372 9292 27428
rect 9348 27372 9360 27428
rect 8960 27360 9360 27372
rect 9440 27428 11440 27440
rect 9440 27372 9452 27428
rect 9508 27372 9772 27428
rect 9828 27372 10092 27428
rect 10148 27372 10412 27428
rect 10468 27372 10732 27428
rect 10788 27372 11052 27428
rect 11108 27372 11372 27428
rect 11428 27372 11440 27428
rect 9440 27360 11440 27372
rect 11520 27428 11920 27440
rect 11520 27372 11532 27428
rect 11588 27372 11852 27428
rect 11908 27372 11920 27428
rect 11520 27360 11920 27372
rect 12000 27428 12400 27440
rect 12000 27372 12012 27428
rect 12068 27372 12332 27428
rect 12388 27372 12400 27428
rect 12000 27360 12400 27372
rect 8480 27268 8880 27280
rect 8480 27212 8492 27268
rect 8548 27212 8812 27268
rect 8868 27212 8880 27268
rect 8480 27200 8880 27212
rect 8960 27268 9360 27280
rect 8960 27212 8972 27268
rect 9028 27212 9292 27268
rect 9348 27212 9360 27268
rect 8960 27200 9360 27212
rect 9440 27268 11440 27280
rect 9440 27212 9452 27268
rect 9508 27212 9772 27268
rect 9828 27212 10092 27268
rect 10148 27212 10412 27268
rect 10468 27212 10732 27268
rect 10788 27212 11052 27268
rect 11108 27212 11372 27268
rect 11428 27212 11440 27268
rect 9440 27200 11440 27212
rect 11520 27268 11920 27280
rect 11520 27212 11532 27268
rect 11588 27212 11852 27268
rect 11908 27212 11920 27268
rect 11520 27200 11920 27212
rect 12000 27268 12400 27280
rect 12000 27212 12012 27268
rect 12068 27212 12332 27268
rect 12388 27212 12400 27268
rect 12000 27200 12400 27212
rect 8480 27108 8880 27120
rect 8480 27052 8492 27108
rect 8548 27052 8812 27108
rect 8868 27052 8880 27108
rect 8480 27040 8880 27052
rect 8960 27108 9360 27120
rect 8960 27052 8972 27108
rect 9028 27052 9292 27108
rect 9348 27052 9360 27108
rect 8960 27040 9360 27052
rect 9440 27108 11440 27120
rect 9440 27052 9452 27108
rect 9508 27052 9772 27108
rect 9828 27052 10092 27108
rect 10148 27052 10412 27108
rect 10468 27052 10732 27108
rect 10788 27052 11052 27108
rect 11108 27052 11372 27108
rect 11428 27052 11440 27108
rect 9440 27040 11440 27052
rect 11520 27108 11920 27120
rect 11520 27052 11532 27108
rect 11588 27052 11852 27108
rect 11908 27052 11920 27108
rect 11520 27040 11920 27052
rect 12000 27108 12400 27120
rect 12000 27052 12012 27108
rect 12068 27052 12332 27108
rect 12388 27052 12400 27108
rect 12000 27040 12400 27052
rect 8480 26948 8880 26960
rect 8480 26892 8492 26948
rect 8548 26892 8812 26948
rect 8868 26892 8880 26948
rect 8480 26880 8880 26892
rect 8960 26948 9360 26960
rect 8960 26892 8972 26948
rect 9028 26892 9292 26948
rect 9348 26892 9360 26948
rect 8960 26880 9360 26892
rect 9440 26948 11440 26960
rect 9440 26892 9452 26948
rect 9508 26892 9772 26948
rect 9828 26892 10092 26948
rect 10148 26892 10412 26948
rect 10468 26892 10732 26948
rect 10788 26892 11052 26948
rect 11108 26892 11372 26948
rect 11428 26892 11440 26948
rect 9440 26880 11440 26892
rect 11520 26948 11920 26960
rect 11520 26892 11532 26948
rect 11588 26892 11852 26948
rect 11908 26892 11920 26948
rect 11520 26880 11920 26892
rect 12000 26948 12400 26960
rect 12000 26892 12012 26948
rect 12068 26892 12332 26948
rect 12388 26892 12400 26948
rect 12000 26880 12400 26892
rect 0 26708 20880 26720
rect 0 26652 10572 26708
rect 10628 26652 20880 26708
rect 0 26640 20880 26652
rect 0 26388 10320 26400
rect 0 26332 10252 26388
rect 10308 26332 10320 26388
rect 0 26320 10320 26332
rect 10560 26388 20880 26400
rect 10560 26332 10572 26388
rect 10628 26332 20880 26388
rect 10560 26320 20880 26332
rect 8480 26148 8880 26160
rect 8480 26092 8492 26148
rect 8548 26092 8812 26148
rect 8868 26092 8880 26148
rect 8480 26080 8880 26092
rect 8960 26148 9360 26160
rect 8960 26092 8972 26148
rect 9028 26092 9292 26148
rect 9348 26092 9360 26148
rect 8960 26080 9360 26092
rect 9440 26148 11440 26160
rect 9440 26092 9452 26148
rect 9508 26092 9772 26148
rect 9828 26092 10092 26148
rect 10148 26092 10412 26148
rect 10468 26092 10732 26148
rect 10788 26092 11052 26148
rect 11108 26092 11372 26148
rect 11428 26092 11440 26148
rect 9440 26080 11440 26092
rect 11520 26148 11920 26160
rect 11520 26092 11532 26148
rect 11588 26092 11852 26148
rect 11908 26092 11920 26148
rect 11520 26080 11920 26092
rect 12000 26148 12400 26160
rect 12000 26092 12012 26148
rect 12068 26092 12332 26148
rect 12388 26092 12400 26148
rect 12000 26080 12400 26092
rect 8480 25988 8880 26000
rect 8480 25932 8492 25988
rect 8548 25932 8812 25988
rect 8868 25932 8880 25988
rect 8480 25920 8880 25932
rect 8960 25988 9360 26000
rect 8960 25932 8972 25988
rect 9028 25932 9292 25988
rect 9348 25932 9360 25988
rect 8960 25920 9360 25932
rect 9440 25988 11440 26000
rect 9440 25932 9452 25988
rect 9508 25932 9772 25988
rect 9828 25932 10092 25988
rect 10148 25932 10412 25988
rect 10468 25932 10732 25988
rect 10788 25932 11052 25988
rect 11108 25932 11372 25988
rect 11428 25932 11440 25988
rect 9440 25920 11440 25932
rect 11520 25988 11920 26000
rect 11520 25932 11532 25988
rect 11588 25932 11852 25988
rect 11908 25932 11920 25988
rect 11520 25920 11920 25932
rect 12000 25988 12400 26000
rect 12000 25932 12012 25988
rect 12068 25932 12332 25988
rect 12388 25932 12400 25988
rect 12000 25920 12400 25932
rect 8480 25828 8880 25840
rect 8480 25772 8492 25828
rect 8548 25772 8812 25828
rect 8868 25772 8880 25828
rect 8480 25760 8880 25772
rect 8960 25828 9360 25840
rect 8960 25772 8972 25828
rect 9028 25772 9292 25828
rect 9348 25772 9360 25828
rect 8960 25760 9360 25772
rect 9440 25828 11440 25840
rect 9440 25772 9452 25828
rect 9508 25772 9772 25828
rect 9828 25772 10092 25828
rect 10148 25772 10412 25828
rect 10468 25772 10732 25828
rect 10788 25772 11052 25828
rect 11108 25772 11372 25828
rect 11428 25772 11440 25828
rect 9440 25760 11440 25772
rect 11520 25828 11920 25840
rect 11520 25772 11532 25828
rect 11588 25772 11852 25828
rect 11908 25772 11920 25828
rect 11520 25760 11920 25772
rect 12000 25828 12400 25840
rect 12000 25772 12012 25828
rect 12068 25772 12332 25828
rect 12388 25772 12400 25828
rect 12000 25760 12400 25772
rect 8480 25668 8880 25680
rect 8480 25612 8492 25668
rect 8548 25612 8812 25668
rect 8868 25612 8880 25668
rect 8480 25600 8880 25612
rect 8960 25668 9360 25680
rect 8960 25612 8972 25668
rect 9028 25612 9292 25668
rect 9348 25612 9360 25668
rect 8960 25600 9360 25612
rect 9440 25668 11440 25680
rect 9440 25612 9452 25668
rect 9508 25612 9772 25668
rect 9828 25612 10092 25668
rect 10148 25612 10412 25668
rect 10468 25612 10732 25668
rect 10788 25612 11052 25668
rect 11108 25612 11372 25668
rect 11428 25612 11440 25668
rect 9440 25600 11440 25612
rect 11520 25668 11920 25680
rect 11520 25612 11532 25668
rect 11588 25612 11852 25668
rect 11908 25612 11920 25668
rect 11520 25600 11920 25612
rect 12000 25668 12400 25680
rect 12000 25612 12012 25668
rect 12068 25612 12332 25668
rect 12388 25612 12400 25668
rect 12000 25600 12400 25612
rect 8480 25508 8880 25520
rect 8480 25452 8492 25508
rect 8548 25452 8812 25508
rect 8868 25452 8880 25508
rect 8480 25440 8880 25452
rect 8960 25508 9360 25520
rect 8960 25452 8972 25508
rect 9028 25452 9292 25508
rect 9348 25452 9360 25508
rect 8960 25440 9360 25452
rect 9440 25508 11440 25520
rect 9440 25452 9452 25508
rect 9508 25452 9772 25508
rect 9828 25452 10092 25508
rect 10148 25452 10412 25508
rect 10468 25452 10732 25508
rect 10788 25452 11052 25508
rect 11108 25452 11372 25508
rect 11428 25452 11440 25508
rect 9440 25440 11440 25452
rect 11520 25508 11920 25520
rect 11520 25452 11532 25508
rect 11588 25452 11852 25508
rect 11908 25452 11920 25508
rect 11520 25440 11920 25452
rect 12000 25508 12400 25520
rect 12000 25452 12012 25508
rect 12068 25452 12332 25508
rect 12388 25452 12400 25508
rect 12000 25440 12400 25452
rect 8480 25348 8880 25360
rect 8480 25292 8492 25348
rect 8548 25292 8812 25348
rect 8868 25292 8880 25348
rect 8480 25280 8880 25292
rect 8960 25348 9360 25360
rect 8960 25292 8972 25348
rect 9028 25292 9292 25348
rect 9348 25292 9360 25348
rect 8960 25280 9360 25292
rect 9440 25348 11440 25360
rect 9440 25292 9452 25348
rect 9508 25292 9772 25348
rect 9828 25292 10092 25348
rect 10148 25292 10412 25348
rect 10468 25292 10732 25348
rect 10788 25292 11052 25348
rect 11108 25292 11372 25348
rect 11428 25292 11440 25348
rect 9440 25280 11440 25292
rect 11520 25348 11920 25360
rect 11520 25292 11532 25348
rect 11588 25292 11852 25348
rect 11908 25292 11920 25348
rect 11520 25280 11920 25292
rect 12000 25348 12400 25360
rect 12000 25292 12012 25348
rect 12068 25292 12332 25348
rect 12388 25292 12400 25348
rect 12000 25280 12400 25292
rect 8480 25188 8880 25200
rect 8480 25132 8492 25188
rect 8548 25132 8812 25188
rect 8868 25132 8880 25188
rect 8480 25120 8880 25132
rect 8960 25188 9360 25200
rect 8960 25132 8972 25188
rect 9028 25132 9292 25188
rect 9348 25132 9360 25188
rect 8960 25120 9360 25132
rect 9440 25188 11440 25200
rect 9440 25132 9452 25188
rect 9508 25132 9772 25188
rect 9828 25132 10092 25188
rect 10148 25132 10412 25188
rect 10468 25132 10732 25188
rect 10788 25132 11052 25188
rect 11108 25132 11372 25188
rect 11428 25132 11440 25188
rect 9440 25120 11440 25132
rect 11520 25188 11920 25200
rect 11520 25132 11532 25188
rect 11588 25132 11852 25188
rect 11908 25132 11920 25188
rect 11520 25120 11920 25132
rect 12000 25188 12400 25200
rect 12000 25132 12012 25188
rect 12068 25132 12332 25188
rect 12388 25132 12400 25188
rect 12000 25120 12400 25132
rect 8480 25028 8880 25040
rect 8480 24972 8492 25028
rect 8548 24972 8812 25028
rect 8868 24972 8880 25028
rect 8480 24960 8880 24972
rect 8960 25028 9360 25040
rect 8960 24972 8972 25028
rect 9028 24972 9292 25028
rect 9348 24972 9360 25028
rect 8960 24960 9360 24972
rect 9440 25028 11440 25040
rect 9440 24972 9452 25028
rect 9508 24972 9772 25028
rect 9828 24972 10092 25028
rect 10148 24972 10412 25028
rect 10468 24972 10732 25028
rect 10788 24972 11052 25028
rect 11108 24972 11372 25028
rect 11428 24972 11440 25028
rect 9440 24960 11440 24972
rect 11520 25028 11920 25040
rect 11520 24972 11532 25028
rect 11588 24972 11852 25028
rect 11908 24972 11920 25028
rect 11520 24960 11920 24972
rect 12000 25028 12400 25040
rect 12000 24972 12012 25028
rect 12068 24972 12332 25028
rect 12388 24972 12400 25028
rect 12000 24960 12400 24972
rect 0 24868 20880 24880
rect 0 24812 9132 24868
rect 9188 24812 20880 24868
rect 0 24800 20880 24812
rect 8480 24708 8880 24720
rect 8480 24652 8492 24708
rect 8548 24652 8812 24708
rect 8868 24652 8880 24708
rect 8480 24640 8880 24652
rect 8960 24708 9360 24720
rect 8960 24652 8972 24708
rect 9028 24652 9292 24708
rect 9348 24652 9360 24708
rect 8960 24640 9360 24652
rect 9440 24708 11440 24720
rect 9440 24652 9452 24708
rect 9508 24652 9772 24708
rect 9828 24652 10092 24708
rect 10148 24652 10412 24708
rect 10468 24652 10732 24708
rect 10788 24652 11052 24708
rect 11108 24652 11372 24708
rect 11428 24652 11440 24708
rect 9440 24640 11440 24652
rect 11520 24708 11920 24720
rect 11520 24652 11532 24708
rect 11588 24652 11852 24708
rect 11908 24652 11920 24708
rect 11520 24640 11920 24652
rect 12000 24708 12400 24720
rect 12000 24652 12012 24708
rect 12068 24652 12332 24708
rect 12388 24652 12400 24708
rect 12000 24640 12400 24652
rect 8480 24548 8880 24560
rect 8480 24492 8492 24548
rect 8548 24492 8812 24548
rect 8868 24492 8880 24548
rect 8480 24480 8880 24492
rect 8960 24548 9360 24560
rect 8960 24492 8972 24548
rect 9028 24492 9292 24548
rect 9348 24492 9360 24548
rect 8960 24480 9360 24492
rect 9440 24548 11440 24560
rect 9440 24492 9452 24548
rect 9508 24492 9772 24548
rect 9828 24492 10092 24548
rect 10148 24492 10412 24548
rect 10468 24492 10732 24548
rect 10788 24492 11052 24548
rect 11108 24492 11372 24548
rect 11428 24492 11440 24548
rect 9440 24480 11440 24492
rect 11520 24548 11920 24560
rect 11520 24492 11532 24548
rect 11588 24492 11852 24548
rect 11908 24492 11920 24548
rect 11520 24480 11920 24492
rect 12000 24548 12400 24560
rect 12000 24492 12012 24548
rect 12068 24492 12332 24548
rect 12388 24492 12400 24548
rect 12000 24480 12400 24492
rect 8480 24388 8880 24400
rect 8480 24332 8492 24388
rect 8548 24332 8812 24388
rect 8868 24332 8880 24388
rect 8480 24320 8880 24332
rect 8960 24388 9360 24400
rect 8960 24332 8972 24388
rect 9028 24332 9292 24388
rect 9348 24332 9360 24388
rect 8960 24320 9360 24332
rect 9440 24388 11440 24400
rect 9440 24332 9452 24388
rect 9508 24332 9772 24388
rect 9828 24332 10092 24388
rect 10148 24332 10412 24388
rect 10468 24332 10732 24388
rect 10788 24332 11052 24388
rect 11108 24332 11372 24388
rect 11428 24332 11440 24388
rect 9440 24320 11440 24332
rect 11520 24388 11920 24400
rect 11520 24332 11532 24388
rect 11588 24332 11852 24388
rect 11908 24332 11920 24388
rect 11520 24320 11920 24332
rect 12000 24388 12400 24400
rect 12000 24332 12012 24388
rect 12068 24332 12332 24388
rect 12388 24332 12400 24388
rect 12000 24320 12400 24332
rect 8480 24228 8880 24240
rect 8480 24172 8492 24228
rect 8548 24172 8812 24228
rect 8868 24172 8880 24228
rect 8480 24160 8880 24172
rect 8960 24228 9360 24240
rect 8960 24172 8972 24228
rect 9028 24172 9292 24228
rect 9348 24172 9360 24228
rect 8960 24160 9360 24172
rect 9440 24228 11440 24240
rect 9440 24172 9452 24228
rect 9508 24172 9772 24228
rect 9828 24172 10092 24228
rect 10148 24172 10412 24228
rect 10468 24172 10732 24228
rect 10788 24172 11052 24228
rect 11108 24172 11372 24228
rect 11428 24172 11440 24228
rect 9440 24160 11440 24172
rect 11520 24228 11920 24240
rect 11520 24172 11532 24228
rect 11588 24172 11852 24228
rect 11908 24172 11920 24228
rect 11520 24160 11920 24172
rect 12000 24228 12400 24240
rect 12000 24172 12012 24228
rect 12068 24172 12332 24228
rect 12388 24172 12400 24228
rect 12000 24160 12400 24172
rect 8480 24068 8880 24080
rect 8480 24012 8492 24068
rect 8548 24012 8812 24068
rect 8868 24012 8880 24068
rect 8480 24000 8880 24012
rect 8960 24068 9360 24080
rect 8960 24012 8972 24068
rect 9028 24012 9292 24068
rect 9348 24012 9360 24068
rect 8960 24000 9360 24012
rect 9440 24068 11440 24080
rect 9440 24012 9452 24068
rect 9508 24012 9772 24068
rect 9828 24012 10092 24068
rect 10148 24012 10412 24068
rect 10468 24012 10732 24068
rect 10788 24012 11052 24068
rect 11108 24012 11372 24068
rect 11428 24012 11440 24068
rect 9440 24000 11440 24012
rect 11520 24068 11920 24080
rect 11520 24012 11532 24068
rect 11588 24012 11852 24068
rect 11908 24012 11920 24068
rect 11520 24000 11920 24012
rect 12000 24068 12400 24080
rect 12000 24012 12012 24068
rect 12068 24012 12332 24068
rect 12388 24012 12400 24068
rect 12000 24000 12400 24012
rect 8480 23908 8880 23920
rect 8480 23852 8492 23908
rect 8548 23852 8812 23908
rect 8868 23852 8880 23908
rect 8480 23840 8880 23852
rect 8960 23908 9360 23920
rect 8960 23852 8972 23908
rect 9028 23852 9292 23908
rect 9348 23852 9360 23908
rect 8960 23840 9360 23852
rect 9440 23908 11440 23920
rect 9440 23852 9452 23908
rect 9508 23852 9772 23908
rect 9828 23852 10092 23908
rect 10148 23852 10412 23908
rect 10468 23852 10732 23908
rect 10788 23852 11052 23908
rect 11108 23852 11372 23908
rect 11428 23852 11440 23908
rect 9440 23840 11440 23852
rect 11520 23908 11920 23920
rect 11520 23852 11532 23908
rect 11588 23852 11852 23908
rect 11908 23852 11920 23908
rect 11520 23840 11920 23852
rect 12000 23908 12400 23920
rect 12000 23852 12012 23908
rect 12068 23852 12332 23908
rect 12388 23852 12400 23908
rect 12000 23840 12400 23852
rect 8480 23748 8880 23760
rect 8480 23692 8492 23748
rect 8548 23692 8812 23748
rect 8868 23692 8880 23748
rect 8480 23680 8880 23692
rect 8960 23748 9360 23760
rect 8960 23692 8972 23748
rect 9028 23692 9292 23748
rect 9348 23692 9360 23748
rect 8960 23680 9360 23692
rect 9440 23748 11440 23760
rect 9440 23692 9452 23748
rect 9508 23692 9772 23748
rect 9828 23692 10092 23748
rect 10148 23692 10412 23748
rect 10468 23692 10732 23748
rect 10788 23692 11052 23748
rect 11108 23692 11372 23748
rect 11428 23692 11440 23748
rect 9440 23680 11440 23692
rect 11520 23748 11920 23760
rect 11520 23692 11532 23748
rect 11588 23692 11852 23748
rect 11908 23692 11920 23748
rect 11520 23680 11920 23692
rect 12000 23748 12400 23760
rect 12000 23692 12012 23748
rect 12068 23692 12332 23748
rect 12388 23692 12400 23748
rect 12000 23680 12400 23692
rect 8480 23588 8880 23600
rect 8480 23532 8492 23588
rect 8548 23532 8812 23588
rect 8868 23532 8880 23588
rect 8480 23520 8880 23532
rect 8960 23588 9360 23600
rect 8960 23532 8972 23588
rect 9028 23532 9292 23588
rect 9348 23532 9360 23588
rect 8960 23520 9360 23532
rect 9440 23588 11440 23600
rect 9440 23532 9452 23588
rect 9508 23532 9772 23588
rect 9828 23532 10092 23588
rect 10148 23532 10412 23588
rect 10468 23532 10732 23588
rect 10788 23532 11052 23588
rect 11108 23532 11372 23588
rect 11428 23532 11440 23588
rect 9440 23520 11440 23532
rect 11520 23588 11920 23600
rect 11520 23532 11532 23588
rect 11588 23532 11852 23588
rect 11908 23532 11920 23588
rect 11520 23520 11920 23532
rect 12000 23588 12400 23600
rect 12000 23532 12012 23588
rect 12068 23532 12332 23588
rect 12388 23532 12400 23588
rect 12000 23520 12400 23532
rect 8480 23428 8880 23440
rect 8480 23372 8492 23428
rect 8548 23372 8812 23428
rect 8868 23372 8880 23428
rect 8480 23360 8880 23372
rect 8960 23428 9360 23440
rect 8960 23372 8972 23428
rect 9028 23372 9292 23428
rect 9348 23372 9360 23428
rect 8960 23360 9360 23372
rect 9440 23428 11440 23440
rect 9440 23372 9452 23428
rect 9508 23372 9772 23428
rect 9828 23372 10092 23428
rect 10148 23372 10412 23428
rect 10468 23372 10732 23428
rect 10788 23372 11052 23428
rect 11108 23372 11372 23428
rect 11428 23372 11440 23428
rect 9440 23360 11440 23372
rect 11520 23428 11920 23440
rect 11520 23372 11532 23428
rect 11588 23372 11852 23428
rect 11908 23372 11920 23428
rect 11520 23360 11920 23372
rect 12000 23428 12400 23440
rect 12000 23372 12012 23428
rect 12068 23372 12332 23428
rect 12388 23372 12400 23428
rect 12000 23360 12400 23372
rect 8480 23268 8880 23280
rect 8480 23212 8492 23268
rect 8548 23212 8812 23268
rect 8868 23212 8880 23268
rect 8480 23200 8880 23212
rect 8960 23268 9360 23280
rect 8960 23212 8972 23268
rect 9028 23212 9292 23268
rect 9348 23212 9360 23268
rect 8960 23200 9360 23212
rect 9440 23268 11440 23280
rect 9440 23212 9452 23268
rect 9508 23212 9772 23268
rect 9828 23212 10092 23268
rect 10148 23212 10412 23268
rect 10468 23212 10732 23268
rect 10788 23212 11052 23268
rect 11108 23212 11372 23268
rect 11428 23212 11440 23268
rect 9440 23200 11440 23212
rect 11520 23268 11920 23280
rect 11520 23212 11532 23268
rect 11588 23212 11852 23268
rect 11908 23212 11920 23268
rect 11520 23200 11920 23212
rect 12000 23268 12400 23280
rect 12000 23212 12012 23268
rect 12068 23212 12332 23268
rect 12388 23212 12400 23268
rect 12000 23200 12400 23212
rect 8480 23108 8880 23120
rect 8480 23052 8492 23108
rect 8548 23052 8812 23108
rect 8868 23052 8880 23108
rect 8480 23040 8880 23052
rect 8960 23108 9360 23120
rect 8960 23052 8972 23108
rect 9028 23052 9292 23108
rect 9348 23052 9360 23108
rect 8960 23040 9360 23052
rect 9440 23108 11440 23120
rect 9440 23052 9452 23108
rect 9508 23052 9772 23108
rect 9828 23052 10092 23108
rect 10148 23052 10412 23108
rect 10468 23052 10732 23108
rect 10788 23052 11052 23108
rect 11108 23052 11372 23108
rect 11428 23052 11440 23108
rect 9440 23040 11440 23052
rect 11520 23108 11920 23120
rect 11520 23052 11532 23108
rect 11588 23052 11852 23108
rect 11908 23052 11920 23108
rect 11520 23040 11920 23052
rect 12000 23108 12400 23120
rect 12000 23052 12012 23108
rect 12068 23052 12332 23108
rect 12388 23052 12400 23108
rect 12000 23040 12400 23052
rect 8480 22948 8880 22960
rect 8480 22892 8492 22948
rect 8548 22892 8812 22948
rect 8868 22892 8880 22948
rect 8480 22880 8880 22892
rect 8960 22948 9360 22960
rect 8960 22892 8972 22948
rect 9028 22892 9292 22948
rect 9348 22892 9360 22948
rect 8960 22880 9360 22892
rect 9440 22948 11440 22960
rect 9440 22892 9452 22948
rect 9508 22892 9772 22948
rect 9828 22892 10092 22948
rect 10148 22892 10412 22948
rect 10468 22892 10732 22948
rect 10788 22892 11052 22948
rect 11108 22892 11372 22948
rect 11428 22892 11440 22948
rect 9440 22880 11440 22892
rect 11520 22948 11920 22960
rect 11520 22892 11532 22948
rect 11588 22892 11852 22948
rect 11908 22892 11920 22948
rect 11520 22880 11920 22892
rect 12000 22948 12400 22960
rect 12000 22892 12012 22948
rect 12068 22892 12332 22948
rect 12388 22892 12400 22948
rect 12000 22880 12400 22892
rect 8480 22788 8880 22800
rect 8480 22732 8492 22788
rect 8548 22732 8812 22788
rect 8868 22732 8880 22788
rect 8480 22720 8880 22732
rect 8960 22788 9360 22800
rect 8960 22732 8972 22788
rect 9028 22732 9292 22788
rect 9348 22732 9360 22788
rect 8960 22720 9360 22732
rect 9440 22788 11440 22800
rect 9440 22732 9452 22788
rect 9508 22732 9772 22788
rect 9828 22732 10092 22788
rect 10148 22732 10412 22788
rect 10468 22732 10732 22788
rect 10788 22732 11052 22788
rect 11108 22732 11372 22788
rect 11428 22732 11440 22788
rect 9440 22720 11440 22732
rect 11520 22788 11920 22800
rect 11520 22732 11532 22788
rect 11588 22732 11852 22788
rect 11908 22732 11920 22788
rect 11520 22720 11920 22732
rect 12000 22788 12400 22800
rect 12000 22732 12012 22788
rect 12068 22732 12332 22788
rect 12388 22732 12400 22788
rect 12000 22720 12400 22732
rect 8480 22628 8880 22640
rect 8480 22572 8492 22628
rect 8548 22572 8812 22628
rect 8868 22572 8880 22628
rect 8480 22560 8880 22572
rect 8960 22628 9360 22640
rect 8960 22572 8972 22628
rect 9028 22572 9292 22628
rect 9348 22572 9360 22628
rect 8960 22560 9360 22572
rect 9440 22628 11440 22640
rect 9440 22572 9452 22628
rect 9508 22572 9772 22628
rect 9828 22572 10092 22628
rect 10148 22572 10412 22628
rect 10468 22572 10732 22628
rect 10788 22572 11052 22628
rect 11108 22572 11372 22628
rect 11428 22572 11440 22628
rect 9440 22560 11440 22572
rect 11520 22628 11920 22640
rect 11520 22572 11532 22628
rect 11588 22572 11852 22628
rect 11908 22572 11920 22628
rect 11520 22560 11920 22572
rect 12000 22628 12400 22640
rect 12000 22572 12012 22628
rect 12068 22572 12332 22628
rect 12388 22572 12400 22628
rect 12000 22560 12400 22572
rect 8480 22468 8880 22480
rect 8480 22412 8492 22468
rect 8548 22412 8812 22468
rect 8868 22412 8880 22468
rect 8480 22400 8880 22412
rect 8960 22468 9360 22480
rect 8960 22412 8972 22468
rect 9028 22412 9292 22468
rect 9348 22412 9360 22468
rect 8960 22400 9360 22412
rect 9440 22468 11440 22480
rect 9440 22412 9452 22468
rect 9508 22412 9772 22468
rect 9828 22412 10092 22468
rect 10148 22412 10412 22468
rect 10468 22412 10732 22468
rect 10788 22412 11052 22468
rect 11108 22412 11372 22468
rect 11428 22412 11440 22468
rect 9440 22400 11440 22412
rect 11520 22468 11920 22480
rect 11520 22412 11532 22468
rect 11588 22412 11852 22468
rect 11908 22412 11920 22468
rect 11520 22400 11920 22412
rect 12000 22468 12400 22480
rect 12000 22412 12012 22468
rect 12068 22412 12332 22468
rect 12388 22412 12400 22468
rect 12000 22400 12400 22412
rect 8480 22308 8880 22320
rect 8480 22252 8492 22308
rect 8548 22252 8812 22308
rect 8868 22252 8880 22308
rect 8480 22240 8880 22252
rect 8960 22308 9360 22320
rect 8960 22252 8972 22308
rect 9028 22252 9292 22308
rect 9348 22252 9360 22308
rect 8960 22240 9360 22252
rect 9440 22308 11440 22320
rect 9440 22252 9452 22308
rect 9508 22252 9772 22308
rect 9828 22252 10092 22308
rect 10148 22252 10412 22308
rect 10468 22252 10732 22308
rect 10788 22252 11052 22308
rect 11108 22252 11372 22308
rect 11428 22252 11440 22308
rect 9440 22240 11440 22252
rect 11520 22308 11920 22320
rect 11520 22252 11532 22308
rect 11588 22252 11852 22308
rect 11908 22252 11920 22308
rect 11520 22240 11920 22252
rect 12000 22308 12400 22320
rect 12000 22252 12012 22308
rect 12068 22252 12332 22308
rect 12388 22252 12400 22308
rect 12000 22240 12400 22252
rect 8480 22148 8880 22160
rect 8480 22092 8492 22148
rect 8548 22092 8812 22148
rect 8868 22092 8880 22148
rect 8480 22080 8880 22092
rect 8960 22148 9360 22160
rect 8960 22092 8972 22148
rect 9028 22092 9292 22148
rect 9348 22092 9360 22148
rect 8960 22080 9360 22092
rect 9440 22148 11440 22160
rect 9440 22092 9452 22148
rect 9508 22092 9772 22148
rect 9828 22092 10092 22148
rect 10148 22092 10412 22148
rect 10468 22092 10732 22148
rect 10788 22092 11052 22148
rect 11108 22092 11372 22148
rect 11428 22092 11440 22148
rect 9440 22080 11440 22092
rect 11520 22148 11920 22160
rect 11520 22092 11532 22148
rect 11588 22092 11852 22148
rect 11908 22092 11920 22148
rect 11520 22080 11920 22092
rect 12000 22148 12400 22160
rect 12000 22092 12012 22148
rect 12068 22092 12332 22148
rect 12388 22092 12400 22148
rect 12000 22080 12400 22092
rect 0 21988 20880 22000
rect 0 21932 9132 21988
rect 9188 21932 20880 21988
rect 0 21920 20880 21932
rect 8480 21828 8880 21840
rect 8480 21772 8492 21828
rect 8548 21772 8812 21828
rect 8868 21772 8880 21828
rect 8480 21760 8880 21772
rect 8960 21828 9360 21840
rect 8960 21772 8972 21828
rect 9028 21772 9292 21828
rect 9348 21772 9360 21828
rect 8960 21760 9360 21772
rect 9440 21828 11440 21840
rect 9440 21772 9452 21828
rect 9508 21772 9772 21828
rect 9828 21772 10092 21828
rect 10148 21772 10412 21828
rect 10468 21772 10732 21828
rect 10788 21772 11052 21828
rect 11108 21772 11372 21828
rect 11428 21772 11440 21828
rect 9440 21760 11440 21772
rect 11520 21828 11920 21840
rect 11520 21772 11532 21828
rect 11588 21772 11852 21828
rect 11908 21772 11920 21828
rect 11520 21760 11920 21772
rect 12000 21828 12400 21840
rect 12000 21772 12012 21828
rect 12068 21772 12332 21828
rect 12388 21772 12400 21828
rect 12000 21760 12400 21772
rect 8480 21668 8880 21680
rect 8480 21612 8492 21668
rect 8548 21612 8812 21668
rect 8868 21612 8880 21668
rect 8480 21600 8880 21612
rect 8960 21668 9360 21680
rect 8960 21612 8972 21668
rect 9028 21612 9292 21668
rect 9348 21612 9360 21668
rect 8960 21600 9360 21612
rect 9440 21668 11440 21680
rect 9440 21612 9452 21668
rect 9508 21612 9772 21668
rect 9828 21612 10092 21668
rect 10148 21612 10412 21668
rect 10468 21612 10732 21668
rect 10788 21612 11052 21668
rect 11108 21612 11372 21668
rect 11428 21612 11440 21668
rect 9440 21600 11440 21612
rect 11520 21668 11920 21680
rect 11520 21612 11532 21668
rect 11588 21612 11852 21668
rect 11908 21612 11920 21668
rect 11520 21600 11920 21612
rect 12000 21668 12400 21680
rect 12000 21612 12012 21668
rect 12068 21612 12332 21668
rect 12388 21612 12400 21668
rect 12000 21600 12400 21612
rect 8480 21508 8880 21520
rect 8480 21452 8492 21508
rect 8548 21452 8812 21508
rect 8868 21452 8880 21508
rect 8480 21440 8880 21452
rect 8960 21508 9360 21520
rect 8960 21452 8972 21508
rect 9028 21452 9292 21508
rect 9348 21452 9360 21508
rect 8960 21440 9360 21452
rect 9440 21508 11440 21520
rect 9440 21452 9452 21508
rect 9508 21452 9772 21508
rect 9828 21452 10092 21508
rect 10148 21452 10412 21508
rect 10468 21452 10732 21508
rect 10788 21452 11052 21508
rect 11108 21452 11372 21508
rect 11428 21452 11440 21508
rect 9440 21440 11440 21452
rect 11520 21508 11920 21520
rect 11520 21452 11532 21508
rect 11588 21452 11852 21508
rect 11908 21452 11920 21508
rect 11520 21440 11920 21452
rect 12000 21508 12400 21520
rect 12000 21452 12012 21508
rect 12068 21452 12332 21508
rect 12388 21452 12400 21508
rect 12000 21440 12400 21452
rect 8480 21348 8880 21360
rect 8480 21292 8492 21348
rect 8548 21292 8812 21348
rect 8868 21292 8880 21348
rect 8480 21280 8880 21292
rect 8960 21348 9360 21360
rect 8960 21292 8972 21348
rect 9028 21292 9292 21348
rect 9348 21292 9360 21348
rect 8960 21280 9360 21292
rect 9440 21348 11440 21360
rect 9440 21292 9452 21348
rect 9508 21292 9772 21348
rect 9828 21292 10092 21348
rect 10148 21292 10412 21348
rect 10468 21292 10732 21348
rect 10788 21292 11052 21348
rect 11108 21292 11372 21348
rect 11428 21292 11440 21348
rect 9440 21280 11440 21292
rect 11520 21348 11920 21360
rect 11520 21292 11532 21348
rect 11588 21292 11852 21348
rect 11908 21292 11920 21348
rect 11520 21280 11920 21292
rect 12000 21348 12400 21360
rect 12000 21292 12012 21348
rect 12068 21292 12332 21348
rect 12388 21292 12400 21348
rect 12000 21280 12400 21292
rect 8480 21188 8880 21200
rect 8480 21132 8492 21188
rect 8548 21132 8812 21188
rect 8868 21132 8880 21188
rect 8480 21120 8880 21132
rect 8960 21188 9360 21200
rect 8960 21132 8972 21188
rect 9028 21132 9292 21188
rect 9348 21132 9360 21188
rect 8960 21120 9360 21132
rect 9440 21188 11440 21200
rect 9440 21132 9452 21188
rect 9508 21132 9772 21188
rect 9828 21132 10092 21188
rect 10148 21132 10412 21188
rect 10468 21132 10732 21188
rect 10788 21132 11052 21188
rect 11108 21132 11372 21188
rect 11428 21132 11440 21188
rect 9440 21120 11440 21132
rect 11520 21188 11920 21200
rect 11520 21132 11532 21188
rect 11588 21132 11852 21188
rect 11908 21132 11920 21188
rect 11520 21120 11920 21132
rect 12000 21188 12400 21200
rect 12000 21132 12012 21188
rect 12068 21132 12332 21188
rect 12388 21132 12400 21188
rect 12000 21120 12400 21132
rect 8480 21028 8880 21040
rect 8480 20972 8492 21028
rect 8548 20972 8812 21028
rect 8868 20972 8880 21028
rect 8480 20960 8880 20972
rect 8960 21028 9360 21040
rect 8960 20972 8972 21028
rect 9028 20972 9292 21028
rect 9348 20972 9360 21028
rect 8960 20960 9360 20972
rect 9440 21028 11440 21040
rect 9440 20972 9452 21028
rect 9508 20972 9772 21028
rect 9828 20972 10092 21028
rect 10148 20972 10412 21028
rect 10468 20972 10732 21028
rect 10788 20972 11052 21028
rect 11108 20972 11372 21028
rect 11428 20972 11440 21028
rect 9440 20960 11440 20972
rect 11520 21028 11920 21040
rect 11520 20972 11532 21028
rect 11588 20972 11852 21028
rect 11908 20972 11920 21028
rect 11520 20960 11920 20972
rect 12000 21028 12400 21040
rect 12000 20972 12012 21028
rect 12068 20972 12332 21028
rect 12388 20972 12400 21028
rect 12000 20960 12400 20972
rect 8480 20868 8880 20880
rect 8480 20812 8492 20868
rect 8548 20812 8812 20868
rect 8868 20812 8880 20868
rect 8480 20800 8880 20812
rect 8960 20868 9360 20880
rect 8960 20812 8972 20868
rect 9028 20812 9292 20868
rect 9348 20812 9360 20868
rect 8960 20800 9360 20812
rect 9440 20868 11440 20880
rect 9440 20812 9452 20868
rect 9508 20812 9772 20868
rect 9828 20812 10092 20868
rect 10148 20812 10412 20868
rect 10468 20812 10732 20868
rect 10788 20812 11052 20868
rect 11108 20812 11372 20868
rect 11428 20812 11440 20868
rect 9440 20800 11440 20812
rect 11520 20868 11920 20880
rect 11520 20812 11532 20868
rect 11588 20812 11852 20868
rect 11908 20812 11920 20868
rect 11520 20800 11920 20812
rect 12000 20868 12400 20880
rect 12000 20812 12012 20868
rect 12068 20812 12332 20868
rect 12388 20812 12400 20868
rect 12000 20800 12400 20812
rect 8480 20708 8880 20720
rect 8480 20652 8492 20708
rect 8548 20652 8812 20708
rect 8868 20652 8880 20708
rect 8480 20640 8880 20652
rect 8960 20708 9360 20720
rect 8960 20652 8972 20708
rect 9028 20652 9292 20708
rect 9348 20652 9360 20708
rect 8960 20640 9360 20652
rect 9440 20708 11440 20720
rect 9440 20652 9452 20708
rect 9508 20652 9772 20708
rect 9828 20652 10092 20708
rect 10148 20652 10412 20708
rect 10468 20652 10732 20708
rect 10788 20652 11052 20708
rect 11108 20652 11372 20708
rect 11428 20652 11440 20708
rect 9440 20640 11440 20652
rect 11520 20708 11920 20720
rect 11520 20652 11532 20708
rect 11588 20652 11852 20708
rect 11908 20652 11920 20708
rect 11520 20640 11920 20652
rect 12000 20708 12400 20720
rect 12000 20652 12012 20708
rect 12068 20652 12332 20708
rect 12388 20652 12400 20708
rect 12000 20640 12400 20652
rect 0 20468 20880 20480
rect 0 20412 10252 20468
rect 10308 20412 20880 20468
rect 0 20400 20880 20412
rect 0 20148 20880 20160
rect 0 20092 10252 20148
rect 10308 20092 20880 20148
rect 0 20080 20880 20092
rect 8480 19908 8880 19920
rect 8480 19852 8492 19908
rect 8548 19852 8812 19908
rect 8868 19852 8880 19908
rect 8480 19840 8880 19852
rect 8960 19908 9360 19920
rect 8960 19852 8972 19908
rect 9028 19852 9292 19908
rect 9348 19852 9360 19908
rect 8960 19840 9360 19852
rect 9440 19908 11440 19920
rect 9440 19852 9452 19908
rect 9508 19852 9772 19908
rect 9828 19852 10092 19908
rect 10148 19852 10412 19908
rect 10468 19852 10732 19908
rect 10788 19852 11052 19908
rect 11108 19852 11372 19908
rect 11428 19852 11440 19908
rect 9440 19840 11440 19852
rect 11520 19908 11920 19920
rect 11520 19852 11532 19908
rect 11588 19852 11852 19908
rect 11908 19852 11920 19908
rect 11520 19840 11920 19852
rect 12000 19908 12400 19920
rect 12000 19852 12012 19908
rect 12068 19852 12332 19908
rect 12388 19852 12400 19908
rect 12000 19840 12400 19852
rect 8480 19748 8880 19760
rect 8480 19692 8492 19748
rect 8548 19692 8812 19748
rect 8868 19692 8880 19748
rect 8480 19680 8880 19692
rect 8960 19748 9360 19760
rect 8960 19692 8972 19748
rect 9028 19692 9292 19748
rect 9348 19692 9360 19748
rect 8960 19680 9360 19692
rect 9440 19748 11440 19760
rect 9440 19692 9452 19748
rect 9508 19692 9772 19748
rect 9828 19692 10092 19748
rect 10148 19692 10412 19748
rect 10468 19692 10732 19748
rect 10788 19692 11052 19748
rect 11108 19692 11372 19748
rect 11428 19692 11440 19748
rect 9440 19680 11440 19692
rect 11520 19748 11920 19760
rect 11520 19692 11532 19748
rect 11588 19692 11852 19748
rect 11908 19692 11920 19748
rect 11520 19680 11920 19692
rect 12000 19748 12400 19760
rect 12000 19692 12012 19748
rect 12068 19692 12332 19748
rect 12388 19692 12400 19748
rect 12000 19680 12400 19692
rect 8480 19588 8880 19600
rect 8480 19532 8492 19588
rect 8548 19532 8812 19588
rect 8868 19532 8880 19588
rect 8480 19520 8880 19532
rect 8960 19588 9360 19600
rect 8960 19532 8972 19588
rect 9028 19532 9292 19588
rect 9348 19532 9360 19588
rect 8960 19520 9360 19532
rect 9440 19588 11440 19600
rect 9440 19532 9452 19588
rect 9508 19532 9772 19588
rect 9828 19532 10092 19588
rect 10148 19532 10412 19588
rect 10468 19532 10732 19588
rect 10788 19532 11052 19588
rect 11108 19532 11372 19588
rect 11428 19532 11440 19588
rect 9440 19520 11440 19532
rect 11520 19588 11920 19600
rect 11520 19532 11532 19588
rect 11588 19532 11852 19588
rect 11908 19532 11920 19588
rect 11520 19520 11920 19532
rect 12000 19588 12400 19600
rect 12000 19532 12012 19588
rect 12068 19532 12332 19588
rect 12388 19532 12400 19588
rect 12000 19520 12400 19532
rect 8480 19428 8880 19440
rect 8480 19372 8492 19428
rect 8548 19372 8812 19428
rect 8868 19372 8880 19428
rect 8480 19360 8880 19372
rect 8960 19428 9360 19440
rect 8960 19372 8972 19428
rect 9028 19372 9292 19428
rect 9348 19372 9360 19428
rect 8960 19360 9360 19372
rect 9440 19428 11440 19440
rect 9440 19372 9452 19428
rect 9508 19372 9772 19428
rect 9828 19372 10092 19428
rect 10148 19372 10412 19428
rect 10468 19372 10732 19428
rect 10788 19372 11052 19428
rect 11108 19372 11372 19428
rect 11428 19372 11440 19428
rect 9440 19360 11440 19372
rect 11520 19428 11920 19440
rect 11520 19372 11532 19428
rect 11588 19372 11852 19428
rect 11908 19372 11920 19428
rect 11520 19360 11920 19372
rect 12000 19428 12400 19440
rect 12000 19372 12012 19428
rect 12068 19372 12332 19428
rect 12388 19372 12400 19428
rect 12000 19360 12400 19372
rect 8480 19268 8880 19280
rect 8480 19212 8492 19268
rect 8548 19212 8812 19268
rect 8868 19212 8880 19268
rect 8480 19200 8880 19212
rect 8960 19268 9360 19280
rect 8960 19212 8972 19268
rect 9028 19212 9292 19268
rect 9348 19212 9360 19268
rect 8960 19200 9360 19212
rect 9440 19268 11440 19280
rect 9440 19212 9452 19268
rect 9508 19212 9772 19268
rect 9828 19212 10092 19268
rect 10148 19212 10412 19268
rect 10468 19212 10732 19268
rect 10788 19212 11052 19268
rect 11108 19212 11372 19268
rect 11428 19212 11440 19268
rect 9440 19200 11440 19212
rect 11520 19268 11920 19280
rect 11520 19212 11532 19268
rect 11588 19212 11852 19268
rect 11908 19212 11920 19268
rect 11520 19200 11920 19212
rect 12000 19268 12400 19280
rect 12000 19212 12012 19268
rect 12068 19212 12332 19268
rect 12388 19212 12400 19268
rect 12000 19200 12400 19212
rect 8480 19108 8880 19120
rect 8480 19052 8492 19108
rect 8548 19052 8812 19108
rect 8868 19052 8880 19108
rect 8480 19040 8880 19052
rect 8960 19108 9360 19120
rect 8960 19052 8972 19108
rect 9028 19052 9292 19108
rect 9348 19052 9360 19108
rect 8960 19040 9360 19052
rect 9440 19108 11440 19120
rect 9440 19052 9452 19108
rect 9508 19052 9772 19108
rect 9828 19052 10092 19108
rect 10148 19052 10412 19108
rect 10468 19052 10732 19108
rect 10788 19052 11052 19108
rect 11108 19052 11372 19108
rect 11428 19052 11440 19108
rect 9440 19040 11440 19052
rect 11520 19108 11920 19120
rect 11520 19052 11532 19108
rect 11588 19052 11852 19108
rect 11908 19052 11920 19108
rect 11520 19040 11920 19052
rect 12000 19108 12400 19120
rect 12000 19052 12012 19108
rect 12068 19052 12332 19108
rect 12388 19052 12400 19108
rect 12000 19040 12400 19052
rect 8480 18948 8880 18960
rect 8480 18892 8492 18948
rect 8548 18892 8812 18948
rect 8868 18892 8880 18948
rect 8480 18880 8880 18892
rect 8960 18948 9360 18960
rect 8960 18892 8972 18948
rect 9028 18892 9292 18948
rect 9348 18892 9360 18948
rect 8960 18880 9360 18892
rect 9440 18948 11440 18960
rect 9440 18892 9452 18948
rect 9508 18892 9772 18948
rect 9828 18892 10092 18948
rect 10148 18892 10412 18948
rect 10468 18892 10732 18948
rect 10788 18892 11052 18948
rect 11108 18892 11372 18948
rect 11428 18892 11440 18948
rect 9440 18880 11440 18892
rect 11520 18948 11920 18960
rect 11520 18892 11532 18948
rect 11588 18892 11852 18948
rect 11908 18892 11920 18948
rect 11520 18880 11920 18892
rect 12000 18948 12400 18960
rect 12000 18892 12012 18948
rect 12068 18892 12332 18948
rect 12388 18892 12400 18948
rect 12000 18880 12400 18892
rect 8480 18788 8880 18800
rect 8480 18732 8492 18788
rect 8548 18732 8812 18788
rect 8868 18732 8880 18788
rect 8480 18720 8880 18732
rect 8960 18788 9360 18800
rect 8960 18732 8972 18788
rect 9028 18732 9292 18788
rect 9348 18732 9360 18788
rect 8960 18720 9360 18732
rect 9440 18788 11440 18800
rect 9440 18732 9452 18788
rect 9508 18732 9772 18788
rect 9828 18732 10092 18788
rect 10148 18732 10412 18788
rect 10468 18732 10732 18788
rect 10788 18732 11052 18788
rect 11108 18732 11372 18788
rect 11428 18732 11440 18788
rect 9440 18720 11440 18732
rect 11520 18788 11920 18800
rect 11520 18732 11532 18788
rect 11588 18732 11852 18788
rect 11908 18732 11920 18788
rect 11520 18720 11920 18732
rect 12000 18788 12400 18800
rect 12000 18732 12012 18788
rect 12068 18732 12332 18788
rect 12388 18732 12400 18788
rect 12000 18720 12400 18732
rect 0 18548 20880 18560
rect 0 18492 10252 18548
rect 10308 18492 20880 18548
rect 0 18480 20880 18492
rect 0 18228 10000 18240
rect 0 18172 9932 18228
rect 9988 18172 10000 18228
rect 0 18160 10000 18172
rect 10880 18228 20880 18240
rect 10880 18172 10892 18228
rect 10948 18172 20880 18228
rect 10880 18160 20880 18172
rect 8480 17988 8880 18000
rect 8480 17932 8492 17988
rect 8548 17932 8812 17988
rect 8868 17932 8880 17988
rect 8480 17920 8880 17932
rect 8960 17988 9360 18000
rect 8960 17932 8972 17988
rect 9028 17932 9292 17988
rect 9348 17932 9360 17988
rect 8960 17920 9360 17932
rect 9440 17988 11440 18000
rect 9440 17932 9452 17988
rect 9508 17932 9772 17988
rect 9828 17932 10092 17988
rect 10148 17932 10412 17988
rect 10468 17932 10732 17988
rect 10788 17932 11052 17988
rect 11108 17932 11372 17988
rect 11428 17932 11440 17988
rect 9440 17920 11440 17932
rect 11520 17988 11920 18000
rect 11520 17932 11532 17988
rect 11588 17932 11852 17988
rect 11908 17932 11920 17988
rect 11520 17920 11920 17932
rect 12000 17988 12400 18000
rect 12000 17932 12012 17988
rect 12068 17932 12332 17988
rect 12388 17932 12400 17988
rect 12000 17920 12400 17932
rect 8480 17828 8880 17840
rect 8480 17772 8492 17828
rect 8548 17772 8812 17828
rect 8868 17772 8880 17828
rect 8480 17760 8880 17772
rect 8960 17828 9360 17840
rect 8960 17772 8972 17828
rect 9028 17772 9292 17828
rect 9348 17772 9360 17828
rect 8960 17760 9360 17772
rect 9440 17828 11440 17840
rect 9440 17772 9452 17828
rect 9508 17772 9772 17828
rect 9828 17772 10092 17828
rect 10148 17772 10412 17828
rect 10468 17772 10732 17828
rect 10788 17772 11052 17828
rect 11108 17772 11372 17828
rect 11428 17772 11440 17828
rect 9440 17760 11440 17772
rect 11520 17828 11920 17840
rect 11520 17772 11532 17828
rect 11588 17772 11852 17828
rect 11908 17772 11920 17828
rect 11520 17760 11920 17772
rect 12000 17828 12400 17840
rect 12000 17772 12012 17828
rect 12068 17772 12332 17828
rect 12388 17772 12400 17828
rect 12000 17760 12400 17772
rect 8480 17668 8880 17680
rect 8480 17612 8492 17668
rect 8548 17612 8812 17668
rect 8868 17612 8880 17668
rect 8480 17600 8880 17612
rect 8960 17668 9360 17680
rect 8960 17612 8972 17668
rect 9028 17612 9292 17668
rect 9348 17612 9360 17668
rect 8960 17600 9360 17612
rect 9440 17668 11440 17680
rect 9440 17612 9452 17668
rect 9508 17612 9772 17668
rect 9828 17612 10092 17668
rect 10148 17612 10412 17668
rect 10468 17612 10732 17668
rect 10788 17612 11052 17668
rect 11108 17612 11372 17668
rect 11428 17612 11440 17668
rect 9440 17600 11440 17612
rect 11520 17668 11920 17680
rect 11520 17612 11532 17668
rect 11588 17612 11852 17668
rect 11908 17612 11920 17668
rect 11520 17600 11920 17612
rect 12000 17668 12400 17680
rect 12000 17612 12012 17668
rect 12068 17612 12332 17668
rect 12388 17612 12400 17668
rect 12000 17600 12400 17612
rect 8480 17508 8880 17520
rect 8480 17452 8492 17508
rect 8548 17452 8812 17508
rect 8868 17452 8880 17508
rect 8480 17440 8880 17452
rect 8960 17508 9360 17520
rect 8960 17452 8972 17508
rect 9028 17452 9292 17508
rect 9348 17452 9360 17508
rect 8960 17440 9360 17452
rect 9440 17508 11440 17520
rect 9440 17452 9452 17508
rect 9508 17452 9772 17508
rect 9828 17452 10092 17508
rect 10148 17452 10412 17508
rect 10468 17452 10732 17508
rect 10788 17452 11052 17508
rect 11108 17452 11372 17508
rect 11428 17452 11440 17508
rect 9440 17440 11440 17452
rect 11520 17508 11920 17520
rect 11520 17452 11532 17508
rect 11588 17452 11852 17508
rect 11908 17452 11920 17508
rect 11520 17440 11920 17452
rect 12000 17508 12400 17520
rect 12000 17452 12012 17508
rect 12068 17452 12332 17508
rect 12388 17452 12400 17508
rect 12000 17440 12400 17452
rect 8480 17348 8880 17360
rect 8480 17292 8492 17348
rect 8548 17292 8812 17348
rect 8868 17292 8880 17348
rect 8480 17280 8880 17292
rect 8960 17348 9360 17360
rect 8960 17292 8972 17348
rect 9028 17292 9292 17348
rect 9348 17292 9360 17348
rect 8960 17280 9360 17292
rect 9440 17348 11440 17360
rect 9440 17292 9452 17348
rect 9508 17292 9772 17348
rect 9828 17292 10092 17348
rect 10148 17292 10412 17348
rect 10468 17292 10732 17348
rect 10788 17292 11052 17348
rect 11108 17292 11372 17348
rect 11428 17292 11440 17348
rect 9440 17280 11440 17292
rect 11520 17348 11920 17360
rect 11520 17292 11532 17348
rect 11588 17292 11852 17348
rect 11908 17292 11920 17348
rect 11520 17280 11920 17292
rect 12000 17348 12400 17360
rect 12000 17292 12012 17348
rect 12068 17292 12332 17348
rect 12388 17292 12400 17348
rect 12000 17280 12400 17292
rect 8480 17188 8880 17200
rect 8480 17132 8492 17188
rect 8548 17132 8812 17188
rect 8868 17132 8880 17188
rect 8480 17120 8880 17132
rect 8960 17188 9360 17200
rect 8960 17132 8972 17188
rect 9028 17132 9292 17188
rect 9348 17132 9360 17188
rect 8960 17120 9360 17132
rect 9440 17188 11440 17200
rect 9440 17132 9452 17188
rect 9508 17132 9772 17188
rect 9828 17132 10092 17188
rect 10148 17132 10412 17188
rect 10468 17132 10732 17188
rect 10788 17132 11052 17188
rect 11108 17132 11372 17188
rect 11428 17132 11440 17188
rect 9440 17120 11440 17132
rect 11520 17188 11920 17200
rect 11520 17132 11532 17188
rect 11588 17132 11852 17188
rect 11908 17132 11920 17188
rect 11520 17120 11920 17132
rect 12000 17188 12400 17200
rect 12000 17132 12012 17188
rect 12068 17132 12332 17188
rect 12388 17132 12400 17188
rect 12000 17120 12400 17132
rect 8480 17028 8880 17040
rect 8480 16972 8492 17028
rect 8548 16972 8812 17028
rect 8868 16972 8880 17028
rect 8480 16960 8880 16972
rect 8960 17028 9360 17040
rect 8960 16972 8972 17028
rect 9028 16972 9292 17028
rect 9348 16972 9360 17028
rect 8960 16960 9360 16972
rect 9440 17028 11440 17040
rect 9440 16972 9452 17028
rect 9508 16972 9772 17028
rect 9828 16972 10092 17028
rect 10148 16972 10412 17028
rect 10468 16972 10732 17028
rect 10788 16972 11052 17028
rect 11108 16972 11372 17028
rect 11428 16972 11440 17028
rect 9440 16960 11440 16972
rect 11520 17028 11920 17040
rect 11520 16972 11532 17028
rect 11588 16972 11852 17028
rect 11908 16972 11920 17028
rect 11520 16960 11920 16972
rect 12000 17028 12400 17040
rect 12000 16972 12012 17028
rect 12068 16972 12332 17028
rect 12388 16972 12400 17028
rect 12000 16960 12400 16972
rect 8480 16868 8880 16880
rect 8480 16812 8492 16868
rect 8548 16812 8812 16868
rect 8868 16812 8880 16868
rect 8480 16800 8880 16812
rect 8960 16868 9360 16880
rect 8960 16812 8972 16868
rect 9028 16812 9292 16868
rect 9348 16812 9360 16868
rect 8960 16800 9360 16812
rect 9440 16868 11440 16880
rect 9440 16812 9452 16868
rect 9508 16812 9772 16868
rect 9828 16812 10092 16868
rect 10148 16812 10412 16868
rect 10468 16812 10732 16868
rect 10788 16812 11052 16868
rect 11108 16812 11372 16868
rect 11428 16812 11440 16868
rect 9440 16800 11440 16812
rect 11520 16868 11920 16880
rect 11520 16812 11532 16868
rect 11588 16812 11852 16868
rect 11908 16812 11920 16868
rect 11520 16800 11920 16812
rect 12000 16868 12400 16880
rect 12000 16812 12012 16868
rect 12068 16812 12332 16868
rect 12388 16812 12400 16868
rect 12000 16800 12400 16812
rect 0 16708 20880 16720
rect 0 16652 9132 16708
rect 9188 16652 20880 16708
rect 0 16640 20880 16652
rect 8480 16548 8880 16560
rect 8480 16492 8492 16548
rect 8548 16492 8812 16548
rect 8868 16492 8880 16548
rect 8480 16480 8880 16492
rect 8960 16548 9360 16560
rect 8960 16492 8972 16548
rect 9028 16492 9292 16548
rect 9348 16492 9360 16548
rect 8960 16480 9360 16492
rect 9440 16548 11440 16560
rect 9440 16492 9452 16548
rect 9508 16492 9772 16548
rect 9828 16492 10092 16548
rect 10148 16492 10412 16548
rect 10468 16492 10732 16548
rect 10788 16492 11052 16548
rect 11108 16492 11372 16548
rect 11428 16492 11440 16548
rect 9440 16480 11440 16492
rect 11520 16548 11920 16560
rect 11520 16492 11532 16548
rect 11588 16492 11852 16548
rect 11908 16492 11920 16548
rect 11520 16480 11920 16492
rect 12000 16548 12400 16560
rect 12000 16492 12012 16548
rect 12068 16492 12332 16548
rect 12388 16492 12400 16548
rect 12000 16480 12400 16492
rect 8480 16388 8880 16400
rect 8480 16332 8492 16388
rect 8548 16332 8812 16388
rect 8868 16332 8880 16388
rect 8480 16320 8880 16332
rect 8960 16388 9360 16400
rect 8960 16332 8972 16388
rect 9028 16332 9292 16388
rect 9348 16332 9360 16388
rect 8960 16320 9360 16332
rect 9440 16388 11440 16400
rect 9440 16332 9452 16388
rect 9508 16332 9772 16388
rect 9828 16332 10092 16388
rect 10148 16332 10412 16388
rect 10468 16332 10732 16388
rect 10788 16332 11052 16388
rect 11108 16332 11372 16388
rect 11428 16332 11440 16388
rect 9440 16320 11440 16332
rect 11520 16388 11920 16400
rect 11520 16332 11532 16388
rect 11588 16332 11852 16388
rect 11908 16332 11920 16388
rect 11520 16320 11920 16332
rect 12000 16388 12400 16400
rect 12000 16332 12012 16388
rect 12068 16332 12332 16388
rect 12388 16332 12400 16388
rect 12000 16320 12400 16332
rect 8480 16228 8880 16240
rect 8480 16172 8492 16228
rect 8548 16172 8812 16228
rect 8868 16172 8880 16228
rect 8480 16160 8880 16172
rect 8960 16228 9360 16240
rect 8960 16172 8972 16228
rect 9028 16172 9292 16228
rect 9348 16172 9360 16228
rect 8960 16160 9360 16172
rect 9440 16228 11440 16240
rect 9440 16172 9452 16228
rect 9508 16172 9772 16228
rect 9828 16172 10092 16228
rect 10148 16172 10412 16228
rect 10468 16172 10732 16228
rect 10788 16172 11052 16228
rect 11108 16172 11372 16228
rect 11428 16172 11440 16228
rect 9440 16160 11440 16172
rect 11520 16228 11920 16240
rect 11520 16172 11532 16228
rect 11588 16172 11852 16228
rect 11908 16172 11920 16228
rect 11520 16160 11920 16172
rect 12000 16228 12400 16240
rect 12000 16172 12012 16228
rect 12068 16172 12332 16228
rect 12388 16172 12400 16228
rect 12000 16160 12400 16172
rect 8480 16068 8880 16080
rect 8480 16012 8492 16068
rect 8548 16012 8812 16068
rect 8868 16012 8880 16068
rect 8480 16000 8880 16012
rect 8960 16068 9360 16080
rect 8960 16012 8972 16068
rect 9028 16012 9292 16068
rect 9348 16012 9360 16068
rect 8960 16000 9360 16012
rect 9440 16068 11440 16080
rect 9440 16012 9452 16068
rect 9508 16012 9772 16068
rect 9828 16012 10092 16068
rect 10148 16012 10412 16068
rect 10468 16012 10732 16068
rect 10788 16012 11052 16068
rect 11108 16012 11372 16068
rect 11428 16012 11440 16068
rect 9440 16000 11440 16012
rect 11520 16068 11920 16080
rect 11520 16012 11532 16068
rect 11588 16012 11852 16068
rect 11908 16012 11920 16068
rect 11520 16000 11920 16012
rect 12000 16068 12400 16080
rect 12000 16012 12012 16068
rect 12068 16012 12332 16068
rect 12388 16012 12400 16068
rect 12000 16000 12400 16012
rect 8480 15908 8880 15920
rect 8480 15852 8492 15908
rect 8548 15852 8812 15908
rect 8868 15852 8880 15908
rect 8480 15840 8880 15852
rect 8960 15908 9360 15920
rect 8960 15852 8972 15908
rect 9028 15852 9292 15908
rect 9348 15852 9360 15908
rect 8960 15840 9360 15852
rect 9440 15908 11440 15920
rect 9440 15852 9452 15908
rect 9508 15852 9772 15908
rect 9828 15852 10092 15908
rect 10148 15852 10412 15908
rect 10468 15852 10732 15908
rect 10788 15852 11052 15908
rect 11108 15852 11372 15908
rect 11428 15852 11440 15908
rect 9440 15840 11440 15852
rect 11520 15908 11920 15920
rect 11520 15852 11532 15908
rect 11588 15852 11852 15908
rect 11908 15852 11920 15908
rect 11520 15840 11920 15852
rect 12000 15908 12400 15920
rect 12000 15852 12012 15908
rect 12068 15852 12332 15908
rect 12388 15852 12400 15908
rect 12000 15840 12400 15852
rect 8480 15748 8880 15760
rect 8480 15692 8492 15748
rect 8548 15692 8812 15748
rect 8868 15692 8880 15748
rect 8480 15680 8880 15692
rect 8960 15748 9360 15760
rect 8960 15692 8972 15748
rect 9028 15692 9292 15748
rect 9348 15692 9360 15748
rect 8960 15680 9360 15692
rect 9440 15748 11440 15760
rect 9440 15692 9452 15748
rect 9508 15692 9772 15748
rect 9828 15692 10092 15748
rect 10148 15692 10412 15748
rect 10468 15692 10732 15748
rect 10788 15692 11052 15748
rect 11108 15692 11372 15748
rect 11428 15692 11440 15748
rect 9440 15680 11440 15692
rect 11520 15748 11920 15760
rect 11520 15692 11532 15748
rect 11588 15692 11852 15748
rect 11908 15692 11920 15748
rect 11520 15680 11920 15692
rect 12000 15748 12400 15760
rect 12000 15692 12012 15748
rect 12068 15692 12332 15748
rect 12388 15692 12400 15748
rect 12000 15680 12400 15692
rect 8480 15588 8880 15600
rect 8480 15532 8492 15588
rect 8548 15532 8812 15588
rect 8868 15532 8880 15588
rect 8480 15520 8880 15532
rect 8960 15588 9360 15600
rect 8960 15532 8972 15588
rect 9028 15532 9292 15588
rect 9348 15532 9360 15588
rect 8960 15520 9360 15532
rect 9440 15588 11440 15600
rect 9440 15532 9452 15588
rect 9508 15532 9772 15588
rect 9828 15532 10092 15588
rect 10148 15532 10412 15588
rect 10468 15532 10732 15588
rect 10788 15532 11052 15588
rect 11108 15532 11372 15588
rect 11428 15532 11440 15588
rect 9440 15520 11440 15532
rect 11520 15588 11920 15600
rect 11520 15532 11532 15588
rect 11588 15532 11852 15588
rect 11908 15532 11920 15588
rect 11520 15520 11920 15532
rect 12000 15588 12400 15600
rect 12000 15532 12012 15588
rect 12068 15532 12332 15588
rect 12388 15532 12400 15588
rect 12000 15520 12400 15532
rect 8480 15428 8880 15440
rect 8480 15372 8492 15428
rect 8548 15372 8812 15428
rect 8868 15372 8880 15428
rect 8480 15360 8880 15372
rect 8960 15428 9360 15440
rect 8960 15372 8972 15428
rect 9028 15372 9292 15428
rect 9348 15372 9360 15428
rect 8960 15360 9360 15372
rect 9440 15428 11440 15440
rect 9440 15372 9452 15428
rect 9508 15372 9772 15428
rect 9828 15372 10092 15428
rect 10148 15372 10412 15428
rect 10468 15372 10732 15428
rect 10788 15372 11052 15428
rect 11108 15372 11372 15428
rect 11428 15372 11440 15428
rect 9440 15360 11440 15372
rect 11520 15428 11920 15440
rect 11520 15372 11532 15428
rect 11588 15372 11852 15428
rect 11908 15372 11920 15428
rect 11520 15360 11920 15372
rect 12000 15428 12400 15440
rect 12000 15372 12012 15428
rect 12068 15372 12332 15428
rect 12388 15372 12400 15428
rect 12000 15360 12400 15372
rect 8480 15268 8880 15280
rect 8480 15212 8492 15268
rect 8548 15212 8812 15268
rect 8868 15212 8880 15268
rect 8480 15200 8880 15212
rect 8960 15268 9360 15280
rect 8960 15212 8972 15268
rect 9028 15212 9292 15268
rect 9348 15212 9360 15268
rect 8960 15200 9360 15212
rect 9440 15268 11440 15280
rect 9440 15212 9452 15268
rect 9508 15212 9772 15268
rect 9828 15212 10092 15268
rect 10148 15212 10412 15268
rect 10468 15212 10732 15268
rect 10788 15212 11052 15268
rect 11108 15212 11372 15268
rect 11428 15212 11440 15268
rect 9440 15200 11440 15212
rect 11520 15268 11920 15280
rect 11520 15212 11532 15268
rect 11588 15212 11852 15268
rect 11908 15212 11920 15268
rect 11520 15200 11920 15212
rect 12000 15268 12400 15280
rect 12000 15212 12012 15268
rect 12068 15212 12332 15268
rect 12388 15212 12400 15268
rect 12000 15200 12400 15212
rect 8480 15108 8880 15120
rect 8480 15052 8492 15108
rect 8548 15052 8812 15108
rect 8868 15052 8880 15108
rect 8480 15040 8880 15052
rect 8960 15108 9360 15120
rect 8960 15052 8972 15108
rect 9028 15052 9292 15108
rect 9348 15052 9360 15108
rect 8960 15040 9360 15052
rect 9440 15108 11440 15120
rect 9440 15052 9452 15108
rect 9508 15052 9772 15108
rect 9828 15052 10092 15108
rect 10148 15052 10412 15108
rect 10468 15052 10732 15108
rect 10788 15052 11052 15108
rect 11108 15052 11372 15108
rect 11428 15052 11440 15108
rect 9440 15040 11440 15052
rect 11520 15108 11920 15120
rect 11520 15052 11532 15108
rect 11588 15052 11852 15108
rect 11908 15052 11920 15108
rect 11520 15040 11920 15052
rect 12000 15108 12400 15120
rect 12000 15052 12012 15108
rect 12068 15052 12332 15108
rect 12388 15052 12400 15108
rect 12000 15040 12400 15052
rect 8480 14948 8880 14960
rect 8480 14892 8492 14948
rect 8548 14892 8812 14948
rect 8868 14892 8880 14948
rect 8480 14880 8880 14892
rect 8960 14948 9360 14960
rect 8960 14892 8972 14948
rect 9028 14892 9292 14948
rect 9348 14892 9360 14948
rect 8960 14880 9360 14892
rect 9440 14948 11440 14960
rect 9440 14892 9452 14948
rect 9508 14892 9772 14948
rect 9828 14892 10092 14948
rect 10148 14892 10412 14948
rect 10468 14892 10732 14948
rect 10788 14892 11052 14948
rect 11108 14892 11372 14948
rect 11428 14892 11440 14948
rect 9440 14880 11440 14892
rect 11520 14948 11920 14960
rect 11520 14892 11532 14948
rect 11588 14892 11852 14948
rect 11908 14892 11920 14948
rect 11520 14880 11920 14892
rect 12000 14948 12400 14960
rect 12000 14892 12012 14948
rect 12068 14892 12332 14948
rect 12388 14892 12400 14948
rect 12000 14880 12400 14892
rect 8480 14788 8880 14800
rect 8480 14732 8492 14788
rect 8548 14732 8812 14788
rect 8868 14732 8880 14788
rect 8480 14720 8880 14732
rect 8960 14788 9360 14800
rect 8960 14732 8972 14788
rect 9028 14732 9292 14788
rect 9348 14732 9360 14788
rect 8960 14720 9360 14732
rect 9440 14788 11440 14800
rect 9440 14732 9452 14788
rect 9508 14732 9772 14788
rect 9828 14732 10092 14788
rect 10148 14732 10412 14788
rect 10468 14732 10732 14788
rect 10788 14732 11052 14788
rect 11108 14732 11372 14788
rect 11428 14732 11440 14788
rect 9440 14720 11440 14732
rect 11520 14788 11920 14800
rect 11520 14732 11532 14788
rect 11588 14732 11852 14788
rect 11908 14732 11920 14788
rect 11520 14720 11920 14732
rect 12000 14788 12400 14800
rect 12000 14732 12012 14788
rect 12068 14732 12332 14788
rect 12388 14732 12400 14788
rect 12000 14720 12400 14732
rect 8480 14628 8880 14640
rect 8480 14572 8492 14628
rect 8548 14572 8812 14628
rect 8868 14572 8880 14628
rect 8480 14560 8880 14572
rect 8960 14628 9360 14640
rect 8960 14572 8972 14628
rect 9028 14572 9292 14628
rect 9348 14572 9360 14628
rect 8960 14560 9360 14572
rect 9440 14628 11440 14640
rect 9440 14572 9452 14628
rect 9508 14572 9772 14628
rect 9828 14572 10092 14628
rect 10148 14572 10412 14628
rect 10468 14572 10732 14628
rect 10788 14572 11052 14628
rect 11108 14572 11372 14628
rect 11428 14572 11440 14628
rect 9440 14560 11440 14572
rect 11520 14628 11920 14640
rect 11520 14572 11532 14628
rect 11588 14572 11852 14628
rect 11908 14572 11920 14628
rect 11520 14560 11920 14572
rect 12000 14628 12400 14640
rect 12000 14572 12012 14628
rect 12068 14572 12332 14628
rect 12388 14572 12400 14628
rect 12000 14560 12400 14572
rect 8480 14468 8880 14480
rect 8480 14412 8492 14468
rect 8548 14412 8812 14468
rect 8868 14412 8880 14468
rect 8480 14400 8880 14412
rect 8960 14468 9360 14480
rect 8960 14412 8972 14468
rect 9028 14412 9292 14468
rect 9348 14412 9360 14468
rect 8960 14400 9360 14412
rect 9440 14468 11440 14480
rect 9440 14412 9452 14468
rect 9508 14412 9772 14468
rect 9828 14412 10092 14468
rect 10148 14412 10412 14468
rect 10468 14412 10732 14468
rect 10788 14412 11052 14468
rect 11108 14412 11372 14468
rect 11428 14412 11440 14468
rect 9440 14400 11440 14412
rect 11520 14468 11920 14480
rect 11520 14412 11532 14468
rect 11588 14412 11852 14468
rect 11908 14412 11920 14468
rect 11520 14400 11920 14412
rect 12000 14468 12400 14480
rect 12000 14412 12012 14468
rect 12068 14412 12332 14468
rect 12388 14412 12400 14468
rect 12000 14400 12400 14412
rect 8480 14308 8880 14320
rect 8480 14252 8492 14308
rect 8548 14252 8812 14308
rect 8868 14252 8880 14308
rect 8480 14240 8880 14252
rect 8960 14308 9360 14320
rect 8960 14252 8972 14308
rect 9028 14252 9292 14308
rect 9348 14252 9360 14308
rect 8960 14240 9360 14252
rect 9440 14308 11440 14320
rect 9440 14252 9452 14308
rect 9508 14252 9772 14308
rect 9828 14252 10092 14308
rect 10148 14252 10412 14308
rect 10468 14252 10732 14308
rect 10788 14252 11052 14308
rect 11108 14252 11372 14308
rect 11428 14252 11440 14308
rect 9440 14240 11440 14252
rect 11520 14308 11920 14320
rect 11520 14252 11532 14308
rect 11588 14252 11852 14308
rect 11908 14252 11920 14308
rect 11520 14240 11920 14252
rect 12000 14308 12400 14320
rect 12000 14252 12012 14308
rect 12068 14252 12332 14308
rect 12388 14252 12400 14308
rect 12000 14240 12400 14252
rect 8480 14148 8880 14160
rect 8480 14092 8492 14148
rect 8548 14092 8812 14148
rect 8868 14092 8880 14148
rect 8480 14080 8880 14092
rect 8960 14148 9360 14160
rect 8960 14092 8972 14148
rect 9028 14092 9292 14148
rect 9348 14092 9360 14148
rect 8960 14080 9360 14092
rect 9440 14148 11440 14160
rect 9440 14092 9452 14148
rect 9508 14092 9772 14148
rect 9828 14092 10092 14148
rect 10148 14092 10412 14148
rect 10468 14092 10732 14148
rect 10788 14092 11052 14148
rect 11108 14092 11372 14148
rect 11428 14092 11440 14148
rect 9440 14080 11440 14092
rect 11520 14148 11920 14160
rect 11520 14092 11532 14148
rect 11588 14092 11852 14148
rect 11908 14092 11920 14148
rect 11520 14080 11920 14092
rect 12000 14148 12400 14160
rect 12000 14092 12012 14148
rect 12068 14092 12332 14148
rect 12388 14092 12400 14148
rect 12000 14080 12400 14092
rect 8480 13988 8880 14000
rect 8480 13932 8492 13988
rect 8548 13932 8812 13988
rect 8868 13932 8880 13988
rect 8480 13920 8880 13932
rect 8960 13988 9360 14000
rect 8960 13932 8972 13988
rect 9028 13932 9292 13988
rect 9348 13932 9360 13988
rect 8960 13920 9360 13932
rect 9440 13988 11440 14000
rect 9440 13932 9452 13988
rect 9508 13932 9772 13988
rect 9828 13932 10092 13988
rect 10148 13932 10412 13988
rect 10468 13932 10732 13988
rect 10788 13932 11052 13988
rect 11108 13932 11372 13988
rect 11428 13932 11440 13988
rect 9440 13920 11440 13932
rect 11520 13988 11920 14000
rect 11520 13932 11532 13988
rect 11588 13932 11852 13988
rect 11908 13932 11920 13988
rect 11520 13920 11920 13932
rect 12000 13988 12400 14000
rect 12000 13932 12012 13988
rect 12068 13932 12332 13988
rect 12388 13932 12400 13988
rect 12000 13920 12400 13932
rect 0 13828 20880 13840
rect 0 13772 9132 13828
rect 9188 13772 20880 13828
rect 0 13760 20880 13772
rect 8480 13668 8880 13680
rect 8480 13612 8492 13668
rect 8548 13612 8812 13668
rect 8868 13612 8880 13668
rect 8480 13600 8880 13612
rect 8960 13668 9360 13680
rect 8960 13612 8972 13668
rect 9028 13612 9292 13668
rect 9348 13612 9360 13668
rect 8960 13600 9360 13612
rect 9440 13668 11440 13680
rect 9440 13612 9452 13668
rect 9508 13612 9772 13668
rect 9828 13612 10092 13668
rect 10148 13612 10412 13668
rect 10468 13612 10732 13668
rect 10788 13612 11052 13668
rect 11108 13612 11372 13668
rect 11428 13612 11440 13668
rect 9440 13600 11440 13612
rect 11520 13668 11920 13680
rect 11520 13612 11532 13668
rect 11588 13612 11852 13668
rect 11908 13612 11920 13668
rect 11520 13600 11920 13612
rect 12000 13668 12400 13680
rect 12000 13612 12012 13668
rect 12068 13612 12332 13668
rect 12388 13612 12400 13668
rect 12000 13600 12400 13612
rect 8480 13508 8880 13520
rect 8480 13452 8492 13508
rect 8548 13452 8812 13508
rect 8868 13452 8880 13508
rect 8480 13440 8880 13452
rect 8960 13508 9360 13520
rect 8960 13452 8972 13508
rect 9028 13452 9292 13508
rect 9348 13452 9360 13508
rect 8960 13440 9360 13452
rect 9440 13508 11440 13520
rect 9440 13452 9452 13508
rect 9508 13452 9772 13508
rect 9828 13452 10092 13508
rect 10148 13452 10412 13508
rect 10468 13452 10732 13508
rect 10788 13452 11052 13508
rect 11108 13452 11372 13508
rect 11428 13452 11440 13508
rect 9440 13440 11440 13452
rect 11520 13508 11920 13520
rect 11520 13452 11532 13508
rect 11588 13452 11852 13508
rect 11908 13452 11920 13508
rect 11520 13440 11920 13452
rect 12000 13508 12400 13520
rect 12000 13452 12012 13508
rect 12068 13452 12332 13508
rect 12388 13452 12400 13508
rect 12000 13440 12400 13452
rect 8480 13348 8880 13360
rect 8480 13292 8492 13348
rect 8548 13292 8812 13348
rect 8868 13292 8880 13348
rect 8480 13280 8880 13292
rect 8960 13348 9360 13360
rect 8960 13292 8972 13348
rect 9028 13292 9292 13348
rect 9348 13292 9360 13348
rect 8960 13280 9360 13292
rect 9440 13348 11440 13360
rect 9440 13292 9452 13348
rect 9508 13292 9772 13348
rect 9828 13292 10092 13348
rect 10148 13292 10412 13348
rect 10468 13292 10732 13348
rect 10788 13292 11052 13348
rect 11108 13292 11372 13348
rect 11428 13292 11440 13348
rect 9440 13280 11440 13292
rect 11520 13348 11920 13360
rect 11520 13292 11532 13348
rect 11588 13292 11852 13348
rect 11908 13292 11920 13348
rect 11520 13280 11920 13292
rect 12000 13348 12400 13360
rect 12000 13292 12012 13348
rect 12068 13292 12332 13348
rect 12388 13292 12400 13348
rect 12000 13280 12400 13292
rect 8480 13188 8880 13200
rect 8480 13132 8492 13188
rect 8548 13132 8812 13188
rect 8868 13132 8880 13188
rect 8480 13120 8880 13132
rect 8960 13188 9360 13200
rect 8960 13132 8972 13188
rect 9028 13132 9292 13188
rect 9348 13132 9360 13188
rect 8960 13120 9360 13132
rect 9440 13188 11440 13200
rect 9440 13132 9452 13188
rect 9508 13132 9772 13188
rect 9828 13132 10092 13188
rect 10148 13132 10412 13188
rect 10468 13132 10732 13188
rect 10788 13132 11052 13188
rect 11108 13132 11372 13188
rect 11428 13132 11440 13188
rect 9440 13120 11440 13132
rect 11520 13188 11920 13200
rect 11520 13132 11532 13188
rect 11588 13132 11852 13188
rect 11908 13132 11920 13188
rect 11520 13120 11920 13132
rect 12000 13188 12400 13200
rect 12000 13132 12012 13188
rect 12068 13132 12332 13188
rect 12388 13132 12400 13188
rect 12000 13120 12400 13132
rect 8480 13028 8880 13040
rect 8480 12972 8492 13028
rect 8548 12972 8812 13028
rect 8868 12972 8880 13028
rect 8480 12960 8880 12972
rect 8960 13028 9360 13040
rect 8960 12972 8972 13028
rect 9028 12972 9292 13028
rect 9348 12972 9360 13028
rect 8960 12960 9360 12972
rect 9440 13028 11440 13040
rect 9440 12972 9452 13028
rect 9508 12972 9772 13028
rect 9828 12972 10092 13028
rect 10148 12972 10412 13028
rect 10468 12972 10732 13028
rect 10788 12972 11052 13028
rect 11108 12972 11372 13028
rect 11428 12972 11440 13028
rect 9440 12960 11440 12972
rect 11520 13028 11920 13040
rect 11520 12972 11532 13028
rect 11588 12972 11852 13028
rect 11908 12972 11920 13028
rect 11520 12960 11920 12972
rect 12000 13028 12400 13040
rect 12000 12972 12012 13028
rect 12068 12972 12332 13028
rect 12388 12972 12400 13028
rect 12000 12960 12400 12972
rect 8480 12868 8880 12880
rect 8480 12812 8492 12868
rect 8548 12812 8812 12868
rect 8868 12812 8880 12868
rect 8480 12800 8880 12812
rect 8960 12868 9360 12880
rect 8960 12812 8972 12868
rect 9028 12812 9292 12868
rect 9348 12812 9360 12868
rect 8960 12800 9360 12812
rect 9440 12868 11440 12880
rect 9440 12812 9452 12868
rect 9508 12812 9772 12868
rect 9828 12812 10092 12868
rect 10148 12812 10412 12868
rect 10468 12812 10732 12868
rect 10788 12812 11052 12868
rect 11108 12812 11372 12868
rect 11428 12812 11440 12868
rect 9440 12800 11440 12812
rect 11520 12868 11920 12880
rect 11520 12812 11532 12868
rect 11588 12812 11852 12868
rect 11908 12812 11920 12868
rect 11520 12800 11920 12812
rect 12000 12868 12400 12880
rect 12000 12812 12012 12868
rect 12068 12812 12332 12868
rect 12388 12812 12400 12868
rect 12000 12800 12400 12812
rect 8480 12708 8880 12720
rect 8480 12652 8492 12708
rect 8548 12652 8812 12708
rect 8868 12652 8880 12708
rect 8480 12640 8880 12652
rect 8960 12708 9360 12720
rect 8960 12652 8972 12708
rect 9028 12652 9292 12708
rect 9348 12652 9360 12708
rect 8960 12640 9360 12652
rect 9440 12708 11440 12720
rect 9440 12652 9452 12708
rect 9508 12652 9772 12708
rect 9828 12652 10092 12708
rect 10148 12652 10412 12708
rect 10468 12652 10732 12708
rect 10788 12652 11052 12708
rect 11108 12652 11372 12708
rect 11428 12652 11440 12708
rect 9440 12640 11440 12652
rect 11520 12708 11920 12720
rect 11520 12652 11532 12708
rect 11588 12652 11852 12708
rect 11908 12652 11920 12708
rect 11520 12640 11920 12652
rect 12000 12708 12400 12720
rect 12000 12652 12012 12708
rect 12068 12652 12332 12708
rect 12388 12652 12400 12708
rect 12000 12640 12400 12652
rect 8480 12548 8880 12560
rect 8480 12492 8492 12548
rect 8548 12492 8812 12548
rect 8868 12492 8880 12548
rect 8480 12480 8880 12492
rect 8960 12548 9360 12560
rect 8960 12492 8972 12548
rect 9028 12492 9292 12548
rect 9348 12492 9360 12548
rect 8960 12480 9360 12492
rect 9440 12548 11440 12560
rect 9440 12492 9452 12548
rect 9508 12492 9772 12548
rect 9828 12492 10092 12548
rect 10148 12492 10412 12548
rect 10468 12492 10732 12548
rect 10788 12492 11052 12548
rect 11108 12492 11372 12548
rect 11428 12492 11440 12548
rect 9440 12480 11440 12492
rect 11520 12548 11920 12560
rect 11520 12492 11532 12548
rect 11588 12492 11852 12548
rect 11908 12492 11920 12548
rect 11520 12480 11920 12492
rect 12000 12548 12400 12560
rect 12000 12492 12012 12548
rect 12068 12492 12332 12548
rect 12388 12492 12400 12548
rect 12000 12480 12400 12492
rect 0 12308 9680 12320
rect 0 12252 9612 12308
rect 9668 12252 9680 12308
rect 0 12240 9680 12252
rect 11200 12308 20880 12320
rect 11200 12252 11212 12308
rect 11268 12252 20880 12308
rect 11200 12240 20880 12252
rect 0 11988 10000 12000
rect 0 11932 9932 11988
rect 9988 11932 10000 11988
rect 0 11920 10000 11932
rect 10880 11988 20880 12000
rect 10880 11932 10892 11988
rect 10948 11932 20880 11988
rect 10880 11920 20880 11932
rect 8480 11748 8880 11760
rect 8480 11692 8492 11748
rect 8548 11692 8812 11748
rect 8868 11692 8880 11748
rect 8480 11680 8880 11692
rect 8960 11748 9360 11760
rect 8960 11692 8972 11748
rect 9028 11692 9292 11748
rect 9348 11692 9360 11748
rect 8960 11680 9360 11692
rect 9440 11748 11440 11760
rect 9440 11692 9452 11748
rect 9508 11692 9772 11748
rect 9828 11692 10092 11748
rect 10148 11692 10412 11748
rect 10468 11692 10732 11748
rect 10788 11692 11052 11748
rect 11108 11692 11372 11748
rect 11428 11692 11440 11748
rect 9440 11680 11440 11692
rect 11520 11748 11920 11760
rect 11520 11692 11532 11748
rect 11588 11692 11852 11748
rect 11908 11692 11920 11748
rect 11520 11680 11920 11692
rect 12000 11748 12400 11760
rect 12000 11692 12012 11748
rect 12068 11692 12332 11748
rect 12388 11692 12400 11748
rect 12000 11680 12400 11692
rect 8480 11588 8880 11600
rect 8480 11532 8492 11588
rect 8548 11532 8812 11588
rect 8868 11532 8880 11588
rect 8480 11520 8880 11532
rect 8960 11588 9360 11600
rect 8960 11532 8972 11588
rect 9028 11532 9292 11588
rect 9348 11532 9360 11588
rect 8960 11520 9360 11532
rect 9440 11588 11440 11600
rect 9440 11532 9452 11588
rect 9508 11532 9772 11588
rect 9828 11532 10092 11588
rect 10148 11532 10412 11588
rect 10468 11532 10732 11588
rect 10788 11532 11052 11588
rect 11108 11532 11372 11588
rect 11428 11532 11440 11588
rect 9440 11520 11440 11532
rect 11520 11588 11920 11600
rect 11520 11532 11532 11588
rect 11588 11532 11852 11588
rect 11908 11532 11920 11588
rect 11520 11520 11920 11532
rect 12000 11588 12400 11600
rect 12000 11532 12012 11588
rect 12068 11532 12332 11588
rect 12388 11532 12400 11588
rect 12000 11520 12400 11532
rect 8480 11428 8880 11440
rect 8480 11372 8492 11428
rect 8548 11372 8812 11428
rect 8868 11372 8880 11428
rect 8480 11360 8880 11372
rect 8960 11428 9360 11440
rect 8960 11372 8972 11428
rect 9028 11372 9292 11428
rect 9348 11372 9360 11428
rect 8960 11360 9360 11372
rect 9440 11428 11440 11440
rect 9440 11372 9452 11428
rect 9508 11372 9772 11428
rect 9828 11372 10092 11428
rect 10148 11372 10412 11428
rect 10468 11372 10732 11428
rect 10788 11372 11052 11428
rect 11108 11372 11372 11428
rect 11428 11372 11440 11428
rect 9440 11360 11440 11372
rect 11520 11428 11920 11440
rect 11520 11372 11532 11428
rect 11588 11372 11852 11428
rect 11908 11372 11920 11428
rect 11520 11360 11920 11372
rect 12000 11428 12400 11440
rect 12000 11372 12012 11428
rect 12068 11372 12332 11428
rect 12388 11372 12400 11428
rect 12000 11360 12400 11372
rect 8480 11268 8880 11280
rect 8480 11212 8492 11268
rect 8548 11212 8812 11268
rect 8868 11212 8880 11268
rect 8480 11200 8880 11212
rect 8960 11268 9360 11280
rect 8960 11212 8972 11268
rect 9028 11212 9292 11268
rect 9348 11212 9360 11268
rect 8960 11200 9360 11212
rect 9440 11268 11440 11280
rect 9440 11212 9452 11268
rect 9508 11212 9772 11268
rect 9828 11212 10092 11268
rect 10148 11212 10412 11268
rect 10468 11212 10732 11268
rect 10788 11212 11052 11268
rect 11108 11212 11372 11268
rect 11428 11212 11440 11268
rect 9440 11200 11440 11212
rect 11520 11268 11920 11280
rect 11520 11212 11532 11268
rect 11588 11212 11852 11268
rect 11908 11212 11920 11268
rect 11520 11200 11920 11212
rect 12000 11268 12400 11280
rect 12000 11212 12012 11268
rect 12068 11212 12332 11268
rect 12388 11212 12400 11268
rect 12000 11200 12400 11212
rect 8480 11108 8880 11120
rect 8480 11052 8492 11108
rect 8548 11052 8812 11108
rect 8868 11052 8880 11108
rect 8480 11040 8880 11052
rect 8960 11108 9360 11120
rect 8960 11052 8972 11108
rect 9028 11052 9292 11108
rect 9348 11052 9360 11108
rect 8960 11040 9360 11052
rect 9440 11108 11440 11120
rect 9440 11052 9452 11108
rect 9508 11052 9772 11108
rect 9828 11052 10092 11108
rect 10148 11052 10412 11108
rect 10468 11052 10732 11108
rect 10788 11052 11052 11108
rect 11108 11052 11372 11108
rect 11428 11052 11440 11108
rect 9440 11040 11440 11052
rect 11520 11108 11920 11120
rect 11520 11052 11532 11108
rect 11588 11052 11852 11108
rect 11908 11052 11920 11108
rect 11520 11040 11920 11052
rect 12000 11108 12400 11120
rect 12000 11052 12012 11108
rect 12068 11052 12332 11108
rect 12388 11052 12400 11108
rect 12000 11040 12400 11052
rect 8480 10948 8880 10960
rect 8480 10892 8492 10948
rect 8548 10892 8812 10948
rect 8868 10892 8880 10948
rect 8480 10880 8880 10892
rect 8960 10948 9360 10960
rect 8960 10892 8972 10948
rect 9028 10892 9292 10948
rect 9348 10892 9360 10948
rect 8960 10880 9360 10892
rect 9440 10948 11440 10960
rect 9440 10892 9452 10948
rect 9508 10892 9772 10948
rect 9828 10892 10092 10948
rect 10148 10892 10412 10948
rect 10468 10892 10732 10948
rect 10788 10892 11052 10948
rect 11108 10892 11372 10948
rect 11428 10892 11440 10948
rect 9440 10880 11440 10892
rect 11520 10948 11920 10960
rect 11520 10892 11532 10948
rect 11588 10892 11852 10948
rect 11908 10892 11920 10948
rect 11520 10880 11920 10892
rect 12000 10948 12400 10960
rect 12000 10892 12012 10948
rect 12068 10892 12332 10948
rect 12388 10892 12400 10948
rect 12000 10880 12400 10892
rect 8480 10788 8880 10800
rect 8480 10732 8492 10788
rect 8548 10732 8812 10788
rect 8868 10732 8880 10788
rect 8480 10720 8880 10732
rect 8960 10788 9360 10800
rect 8960 10732 8972 10788
rect 9028 10732 9292 10788
rect 9348 10732 9360 10788
rect 8960 10720 9360 10732
rect 9440 10788 11440 10800
rect 9440 10732 9452 10788
rect 9508 10732 9772 10788
rect 9828 10732 10092 10788
rect 10148 10732 10412 10788
rect 10468 10732 10732 10788
rect 10788 10732 11052 10788
rect 11108 10732 11372 10788
rect 11428 10732 11440 10788
rect 9440 10720 11440 10732
rect 11520 10788 11920 10800
rect 11520 10732 11532 10788
rect 11588 10732 11852 10788
rect 11908 10732 11920 10788
rect 11520 10720 11920 10732
rect 12000 10788 12400 10800
rect 12000 10732 12012 10788
rect 12068 10732 12332 10788
rect 12388 10732 12400 10788
rect 12000 10720 12400 10732
rect 8480 10628 8880 10640
rect 8480 10572 8492 10628
rect 8548 10572 8812 10628
rect 8868 10572 8880 10628
rect 8480 10560 8880 10572
rect 8960 10628 9360 10640
rect 8960 10572 8972 10628
rect 9028 10572 9292 10628
rect 9348 10572 9360 10628
rect 8960 10560 9360 10572
rect 9440 10628 11440 10640
rect 9440 10572 9452 10628
rect 9508 10572 9772 10628
rect 9828 10572 10092 10628
rect 10148 10572 10412 10628
rect 10468 10572 10732 10628
rect 10788 10572 11052 10628
rect 11108 10572 11372 10628
rect 11428 10572 11440 10628
rect 9440 10560 11440 10572
rect 11520 10628 11920 10640
rect 11520 10572 11532 10628
rect 11588 10572 11852 10628
rect 11908 10572 11920 10628
rect 11520 10560 11920 10572
rect 12000 10628 12400 10640
rect 12000 10572 12012 10628
rect 12068 10572 12332 10628
rect 12388 10572 12400 10628
rect 12000 10560 12400 10572
rect 8480 10468 8880 10480
rect 8480 10412 8492 10468
rect 8548 10412 8812 10468
rect 8868 10412 8880 10468
rect 8480 10400 8880 10412
rect 8960 10468 9360 10480
rect 8960 10412 8972 10468
rect 9028 10412 9292 10468
rect 9348 10412 9360 10468
rect 8960 10400 9360 10412
rect 9440 10468 11440 10480
rect 9440 10412 9452 10468
rect 9508 10412 9772 10468
rect 9828 10412 10092 10468
rect 10148 10412 10412 10468
rect 10468 10412 10732 10468
rect 10788 10412 11052 10468
rect 11108 10412 11372 10468
rect 11428 10412 11440 10468
rect 9440 10400 11440 10412
rect 11520 10468 11920 10480
rect 11520 10412 11532 10468
rect 11588 10412 11852 10468
rect 11908 10412 11920 10468
rect 11520 10400 11920 10412
rect 12000 10468 12400 10480
rect 12000 10412 12012 10468
rect 12068 10412 12332 10468
rect 12388 10412 12400 10468
rect 12000 10400 12400 10412
rect 8480 10308 8880 10320
rect 8480 10252 8492 10308
rect 8548 10252 8812 10308
rect 8868 10252 8880 10308
rect 8480 10240 8880 10252
rect 8960 10308 9360 10320
rect 8960 10252 8972 10308
rect 9028 10252 9292 10308
rect 9348 10252 9360 10308
rect 8960 10240 9360 10252
rect 9440 10308 11440 10320
rect 9440 10252 9452 10308
rect 9508 10252 9772 10308
rect 9828 10252 10092 10308
rect 10148 10252 10412 10308
rect 10468 10252 10732 10308
rect 10788 10252 11052 10308
rect 11108 10252 11372 10308
rect 11428 10252 11440 10308
rect 9440 10240 11440 10252
rect 11520 10308 11920 10320
rect 11520 10252 11532 10308
rect 11588 10252 11852 10308
rect 11908 10252 11920 10308
rect 11520 10240 11920 10252
rect 12000 10308 12400 10320
rect 12000 10252 12012 10308
rect 12068 10252 12332 10308
rect 12388 10252 12400 10308
rect 12000 10240 12400 10252
rect 8480 10148 8880 10160
rect 8480 10092 8492 10148
rect 8548 10092 8812 10148
rect 8868 10092 8880 10148
rect 8480 10080 8880 10092
rect 8960 10148 9360 10160
rect 8960 10092 8972 10148
rect 9028 10092 9292 10148
rect 9348 10092 9360 10148
rect 8960 10080 9360 10092
rect 9440 10148 11440 10160
rect 9440 10092 9452 10148
rect 9508 10092 9772 10148
rect 9828 10092 10092 10148
rect 10148 10092 10412 10148
rect 10468 10092 10732 10148
rect 10788 10092 11052 10148
rect 11108 10092 11372 10148
rect 11428 10092 11440 10148
rect 9440 10080 11440 10092
rect 11520 10148 11920 10160
rect 11520 10092 11532 10148
rect 11588 10092 11852 10148
rect 11908 10092 11920 10148
rect 11520 10080 11920 10092
rect 12000 10148 12400 10160
rect 12000 10092 12012 10148
rect 12068 10092 12332 10148
rect 12388 10092 12400 10148
rect 12000 10080 12400 10092
rect 8480 9988 8880 10000
rect 8480 9932 8492 9988
rect 8548 9932 8812 9988
rect 8868 9932 8880 9988
rect 8480 9920 8880 9932
rect 8960 9988 9360 10000
rect 8960 9932 8972 9988
rect 9028 9932 9292 9988
rect 9348 9932 9360 9988
rect 8960 9920 9360 9932
rect 9440 9988 11440 10000
rect 9440 9932 9452 9988
rect 9508 9932 9772 9988
rect 9828 9932 10092 9988
rect 10148 9932 10412 9988
rect 10468 9932 10732 9988
rect 10788 9932 11052 9988
rect 11108 9932 11372 9988
rect 11428 9932 11440 9988
rect 9440 9920 11440 9932
rect 11520 9988 11920 10000
rect 11520 9932 11532 9988
rect 11588 9932 11852 9988
rect 11908 9932 11920 9988
rect 11520 9920 11920 9932
rect 12000 9988 12400 10000
rect 12000 9932 12012 9988
rect 12068 9932 12332 9988
rect 12388 9932 12400 9988
rect 12000 9920 12400 9932
rect 8480 9828 8880 9840
rect 8480 9772 8492 9828
rect 8548 9772 8812 9828
rect 8868 9772 8880 9828
rect 8480 9760 8880 9772
rect 8960 9828 9360 9840
rect 8960 9772 8972 9828
rect 9028 9772 9292 9828
rect 9348 9772 9360 9828
rect 8960 9760 9360 9772
rect 9440 9828 11440 9840
rect 9440 9772 9452 9828
rect 9508 9772 9772 9828
rect 9828 9772 10092 9828
rect 10148 9772 10412 9828
rect 10468 9772 10732 9828
rect 10788 9772 11052 9828
rect 11108 9772 11372 9828
rect 11428 9772 11440 9828
rect 9440 9760 11440 9772
rect 11520 9828 11920 9840
rect 11520 9772 11532 9828
rect 11588 9772 11852 9828
rect 11908 9772 11920 9828
rect 11520 9760 11920 9772
rect 12000 9828 12400 9840
rect 12000 9772 12012 9828
rect 12068 9772 12332 9828
rect 12388 9772 12400 9828
rect 12000 9760 12400 9772
rect 0 9668 20880 9680
rect 0 9612 11692 9668
rect 11748 9612 20880 9668
rect 0 9600 20880 9612
rect 8480 9508 8880 9520
rect 8480 9452 8492 9508
rect 8548 9452 8812 9508
rect 8868 9452 8880 9508
rect 8480 9440 8880 9452
rect 8960 9508 9360 9520
rect 8960 9452 8972 9508
rect 9028 9452 9292 9508
rect 9348 9452 9360 9508
rect 8960 9440 9360 9452
rect 9440 9508 11440 9520
rect 9440 9452 9452 9508
rect 9508 9452 9772 9508
rect 9828 9452 10092 9508
rect 10148 9452 10412 9508
rect 10468 9452 10732 9508
rect 10788 9452 11052 9508
rect 11108 9452 11372 9508
rect 11428 9452 11440 9508
rect 9440 9440 11440 9452
rect 11520 9508 11920 9520
rect 11520 9452 11532 9508
rect 11588 9452 11852 9508
rect 11908 9452 11920 9508
rect 11520 9440 11920 9452
rect 12000 9508 12400 9520
rect 12000 9452 12012 9508
rect 12068 9452 12332 9508
rect 12388 9452 12400 9508
rect 12000 9440 12400 9452
rect 8480 9348 8880 9360
rect 8480 9292 8492 9348
rect 8548 9292 8812 9348
rect 8868 9292 8880 9348
rect 8480 9280 8880 9292
rect 8960 9348 9360 9360
rect 8960 9292 8972 9348
rect 9028 9292 9292 9348
rect 9348 9292 9360 9348
rect 8960 9280 9360 9292
rect 9440 9348 11440 9360
rect 9440 9292 9452 9348
rect 9508 9292 9772 9348
rect 9828 9292 10092 9348
rect 10148 9292 10412 9348
rect 10468 9292 10732 9348
rect 10788 9292 11052 9348
rect 11108 9292 11372 9348
rect 11428 9292 11440 9348
rect 9440 9280 11440 9292
rect 11520 9348 11920 9360
rect 11520 9292 11532 9348
rect 11588 9292 11852 9348
rect 11908 9292 11920 9348
rect 11520 9280 11920 9292
rect 12000 9348 12400 9360
rect 12000 9292 12012 9348
rect 12068 9292 12332 9348
rect 12388 9292 12400 9348
rect 12000 9280 12400 9292
rect 0 9188 20880 9200
rect 0 9132 12172 9188
rect 12228 9132 20880 9188
rect 0 9120 20880 9132
rect 8480 9028 8880 9040
rect 8480 8972 8492 9028
rect 8548 8972 8812 9028
rect 8868 8972 8880 9028
rect 8480 8960 8880 8972
rect 8960 9028 9360 9040
rect 8960 8972 8972 9028
rect 9028 8972 9292 9028
rect 9348 8972 9360 9028
rect 8960 8960 9360 8972
rect 9440 9028 11440 9040
rect 9440 8972 9452 9028
rect 9508 8972 9772 9028
rect 9828 8972 10092 9028
rect 10148 8972 10412 9028
rect 10468 8972 10732 9028
rect 10788 8972 11052 9028
rect 11108 8972 11372 9028
rect 11428 8972 11440 9028
rect 9440 8960 11440 8972
rect 11520 9028 11920 9040
rect 11520 8972 11532 9028
rect 11588 8972 11852 9028
rect 11908 8972 11920 9028
rect 11520 8960 11920 8972
rect 12000 9028 12400 9040
rect 12000 8972 12012 9028
rect 12068 8972 12332 9028
rect 12388 8972 12400 9028
rect 12000 8960 12400 8972
rect 8480 8868 8880 8880
rect 8480 8812 8492 8868
rect 8548 8812 8812 8868
rect 8868 8812 8880 8868
rect 8480 8800 8880 8812
rect 8960 8868 9360 8880
rect 8960 8812 8972 8868
rect 9028 8812 9292 8868
rect 9348 8812 9360 8868
rect 8960 8800 9360 8812
rect 9440 8868 11440 8880
rect 9440 8812 9452 8868
rect 9508 8812 9772 8868
rect 9828 8812 10092 8868
rect 10148 8812 10412 8868
rect 10468 8812 10732 8868
rect 10788 8812 11052 8868
rect 11108 8812 11372 8868
rect 11428 8812 11440 8868
rect 9440 8800 11440 8812
rect 11520 8868 11920 8880
rect 11520 8812 11532 8868
rect 11588 8812 11852 8868
rect 11908 8812 11920 8868
rect 11520 8800 11920 8812
rect 12000 8868 12400 8880
rect 12000 8812 12012 8868
rect 12068 8812 12332 8868
rect 12388 8812 12400 8868
rect 12000 8800 12400 8812
rect 8480 8708 8880 8720
rect 8480 8652 8492 8708
rect 8548 8652 8812 8708
rect 8868 8652 8880 8708
rect 8480 8640 8880 8652
rect 8960 8708 9360 8720
rect 8960 8652 8972 8708
rect 9028 8652 9292 8708
rect 9348 8652 9360 8708
rect 8960 8640 9360 8652
rect 9440 8708 11440 8720
rect 9440 8652 9452 8708
rect 9508 8652 9772 8708
rect 9828 8652 10092 8708
rect 10148 8652 10412 8708
rect 10468 8652 10732 8708
rect 10788 8652 11052 8708
rect 11108 8652 11372 8708
rect 11428 8652 11440 8708
rect 9440 8640 11440 8652
rect 11520 8708 11920 8720
rect 11520 8652 11532 8708
rect 11588 8652 11852 8708
rect 11908 8652 11920 8708
rect 11520 8640 11920 8652
rect 12000 8708 12400 8720
rect 12000 8652 12012 8708
rect 12068 8652 12332 8708
rect 12388 8652 12400 8708
rect 12000 8640 12400 8652
rect 8480 8548 8880 8560
rect 8480 8492 8492 8548
rect 8548 8492 8812 8548
rect 8868 8492 8880 8548
rect 8480 8480 8880 8492
rect 8960 8548 9360 8560
rect 8960 8492 8972 8548
rect 9028 8492 9292 8548
rect 9348 8492 9360 8548
rect 8960 8480 9360 8492
rect 9440 8548 11440 8560
rect 9440 8492 9452 8548
rect 9508 8492 9772 8548
rect 9828 8492 10092 8548
rect 10148 8492 10412 8548
rect 10468 8492 10732 8548
rect 10788 8492 11052 8548
rect 11108 8492 11372 8548
rect 11428 8492 11440 8548
rect 9440 8480 11440 8492
rect 11520 8548 11920 8560
rect 11520 8492 11532 8548
rect 11588 8492 11852 8548
rect 11908 8492 11920 8548
rect 11520 8480 11920 8492
rect 12000 8548 12400 8560
rect 12000 8492 12012 8548
rect 12068 8492 12332 8548
rect 12388 8492 12400 8548
rect 12000 8480 12400 8492
rect 8480 8388 8880 8400
rect 8480 8332 8492 8388
rect 8548 8332 8812 8388
rect 8868 8332 8880 8388
rect 8480 8320 8880 8332
rect 8960 8388 9360 8400
rect 8960 8332 8972 8388
rect 9028 8332 9292 8388
rect 9348 8332 9360 8388
rect 8960 8320 9360 8332
rect 9440 8388 11440 8400
rect 9440 8332 9452 8388
rect 9508 8332 9772 8388
rect 9828 8332 10092 8388
rect 10148 8332 10412 8388
rect 10468 8332 10732 8388
rect 10788 8332 11052 8388
rect 11108 8332 11372 8388
rect 11428 8332 11440 8388
rect 9440 8320 11440 8332
rect 11520 8388 11920 8400
rect 11520 8332 11532 8388
rect 11588 8332 11852 8388
rect 11908 8332 11920 8388
rect 11520 8320 11920 8332
rect 12000 8388 12400 8400
rect 12000 8332 12012 8388
rect 12068 8332 12332 8388
rect 12388 8332 12400 8388
rect 12000 8320 12400 8332
rect 8480 8228 8880 8240
rect 8480 8172 8492 8228
rect 8548 8172 8812 8228
rect 8868 8172 8880 8228
rect 8480 8160 8880 8172
rect 8960 8228 9360 8240
rect 8960 8172 8972 8228
rect 9028 8172 9292 8228
rect 9348 8172 9360 8228
rect 8960 8160 9360 8172
rect 9440 8228 11440 8240
rect 9440 8172 9452 8228
rect 9508 8172 9772 8228
rect 9828 8172 10092 8228
rect 10148 8172 10412 8228
rect 10468 8172 10732 8228
rect 10788 8172 11052 8228
rect 11108 8172 11372 8228
rect 11428 8172 11440 8228
rect 9440 8160 11440 8172
rect 11520 8228 11920 8240
rect 11520 8172 11532 8228
rect 11588 8172 11852 8228
rect 11908 8172 11920 8228
rect 11520 8160 11920 8172
rect 12000 8228 12400 8240
rect 12000 8172 12012 8228
rect 12068 8172 12332 8228
rect 12388 8172 12400 8228
rect 12000 8160 12400 8172
rect 8480 8068 8880 8080
rect 8480 8012 8492 8068
rect 8548 8012 8812 8068
rect 8868 8012 8880 8068
rect 8480 8000 8880 8012
rect 8960 8068 9360 8080
rect 8960 8012 8972 8068
rect 9028 8012 9292 8068
rect 9348 8012 9360 8068
rect 8960 8000 9360 8012
rect 9440 8068 11440 8080
rect 9440 8012 9452 8068
rect 9508 8012 9772 8068
rect 9828 8012 10092 8068
rect 10148 8012 10412 8068
rect 10468 8012 10732 8068
rect 10788 8012 11052 8068
rect 11108 8012 11372 8068
rect 11428 8012 11440 8068
rect 9440 8000 11440 8012
rect 11520 8068 11920 8080
rect 11520 8012 11532 8068
rect 11588 8012 11852 8068
rect 11908 8012 11920 8068
rect 11520 8000 11920 8012
rect 12000 8068 12400 8080
rect 12000 8012 12012 8068
rect 12068 8012 12332 8068
rect 12388 8012 12400 8068
rect 12000 8000 12400 8012
rect 8480 7908 8880 7920
rect 8480 7852 8492 7908
rect 8548 7852 8812 7908
rect 8868 7852 8880 7908
rect 8480 7840 8880 7852
rect 8960 7908 9360 7920
rect 8960 7852 8972 7908
rect 9028 7852 9292 7908
rect 9348 7852 9360 7908
rect 8960 7840 9360 7852
rect 9440 7908 11440 7920
rect 9440 7852 9452 7908
rect 9508 7852 9772 7908
rect 9828 7852 10092 7908
rect 10148 7852 10412 7908
rect 10468 7852 10732 7908
rect 10788 7852 11052 7908
rect 11108 7852 11372 7908
rect 11428 7852 11440 7908
rect 9440 7840 11440 7852
rect 11520 7908 11920 7920
rect 11520 7852 11532 7908
rect 11588 7852 11852 7908
rect 11908 7852 11920 7908
rect 11520 7840 11920 7852
rect 12000 7908 12400 7920
rect 12000 7852 12012 7908
rect 12068 7852 12332 7908
rect 12388 7852 12400 7908
rect 12000 7840 12400 7852
rect 8480 7748 8880 7760
rect 8480 7692 8492 7748
rect 8548 7692 8812 7748
rect 8868 7692 8880 7748
rect 8480 7680 8880 7692
rect 8960 7748 9360 7760
rect 8960 7692 8972 7748
rect 9028 7692 9292 7748
rect 9348 7692 9360 7748
rect 8960 7680 9360 7692
rect 9440 7748 11440 7760
rect 9440 7692 9452 7748
rect 9508 7692 9772 7748
rect 9828 7692 10092 7748
rect 10148 7692 10412 7748
rect 10468 7692 10732 7748
rect 10788 7692 11052 7748
rect 11108 7692 11372 7748
rect 11428 7692 11440 7748
rect 9440 7680 11440 7692
rect 11520 7748 11920 7760
rect 11520 7692 11532 7748
rect 11588 7692 11852 7748
rect 11908 7692 11920 7748
rect 11520 7680 11920 7692
rect 12000 7748 12400 7760
rect 12000 7692 12012 7748
rect 12068 7692 12332 7748
rect 12388 7692 12400 7748
rect 12000 7680 12400 7692
rect 0 7588 20880 7600
rect 0 7532 8652 7588
rect 8708 7532 20880 7588
rect 0 7520 20880 7532
rect 8480 7428 8880 7440
rect 8480 7372 8492 7428
rect 8548 7372 8812 7428
rect 8868 7372 8880 7428
rect 8480 7360 8880 7372
rect 8960 7428 9360 7440
rect 8960 7372 8972 7428
rect 9028 7372 9292 7428
rect 9348 7372 9360 7428
rect 8960 7360 9360 7372
rect 9440 7428 11440 7440
rect 9440 7372 9452 7428
rect 9508 7372 9772 7428
rect 9828 7372 10092 7428
rect 10148 7372 10412 7428
rect 10468 7372 10732 7428
rect 10788 7372 11052 7428
rect 11108 7372 11372 7428
rect 11428 7372 11440 7428
rect 9440 7360 11440 7372
rect 11520 7428 11920 7440
rect 11520 7372 11532 7428
rect 11588 7372 11852 7428
rect 11908 7372 11920 7428
rect 11520 7360 11920 7372
rect 12000 7428 12400 7440
rect 12000 7372 12012 7428
rect 12068 7372 12332 7428
rect 12388 7372 12400 7428
rect 12000 7360 12400 7372
rect 8480 7268 8880 7280
rect 8480 7212 8492 7268
rect 8548 7212 8812 7268
rect 8868 7212 8880 7268
rect 8480 7200 8880 7212
rect 8960 7268 9360 7280
rect 8960 7212 8972 7268
rect 9028 7212 9292 7268
rect 9348 7212 9360 7268
rect 8960 7200 9360 7212
rect 9440 7268 11440 7280
rect 9440 7212 9452 7268
rect 9508 7212 9772 7268
rect 9828 7212 10092 7268
rect 10148 7212 10412 7268
rect 10468 7212 10732 7268
rect 10788 7212 11052 7268
rect 11108 7212 11372 7268
rect 11428 7212 11440 7268
rect 9440 7200 11440 7212
rect 11520 7268 11920 7280
rect 11520 7212 11532 7268
rect 11588 7212 11852 7268
rect 11908 7212 11920 7268
rect 11520 7200 11920 7212
rect 12000 7268 12400 7280
rect 12000 7212 12012 7268
rect 12068 7212 12332 7268
rect 12388 7212 12400 7268
rect 12000 7200 12400 7212
rect 0 7108 20880 7120
rect 0 7052 9132 7108
rect 9188 7052 20880 7108
rect 0 7040 20880 7052
rect 8480 6948 8880 6960
rect 8480 6892 8492 6948
rect 8548 6892 8812 6948
rect 8868 6892 8880 6948
rect 8480 6880 8880 6892
rect 8960 6948 9360 6960
rect 8960 6892 8972 6948
rect 9028 6892 9292 6948
rect 9348 6892 9360 6948
rect 8960 6880 9360 6892
rect 9440 6948 11440 6960
rect 9440 6892 9452 6948
rect 9508 6892 9772 6948
rect 9828 6892 10092 6948
rect 10148 6892 10412 6948
rect 10468 6892 10732 6948
rect 10788 6892 11052 6948
rect 11108 6892 11372 6948
rect 11428 6892 11440 6948
rect 9440 6880 11440 6892
rect 11520 6948 11920 6960
rect 11520 6892 11532 6948
rect 11588 6892 11852 6948
rect 11908 6892 11920 6948
rect 11520 6880 11920 6892
rect 12000 6948 12400 6960
rect 12000 6892 12012 6948
rect 12068 6892 12332 6948
rect 12388 6892 12400 6948
rect 12000 6880 12400 6892
rect 8480 6788 8880 6800
rect 8480 6732 8492 6788
rect 8548 6732 8812 6788
rect 8868 6732 8880 6788
rect 8480 6720 8880 6732
rect 8960 6788 9360 6800
rect 8960 6732 8972 6788
rect 9028 6732 9292 6788
rect 9348 6732 9360 6788
rect 8960 6720 9360 6732
rect 9440 6788 11440 6800
rect 9440 6732 9452 6788
rect 9508 6732 9772 6788
rect 9828 6732 10092 6788
rect 10148 6732 10412 6788
rect 10468 6732 10732 6788
rect 10788 6732 11052 6788
rect 11108 6732 11372 6788
rect 11428 6732 11440 6788
rect 9440 6720 11440 6732
rect 11520 6788 11920 6800
rect 11520 6732 11532 6788
rect 11588 6732 11852 6788
rect 11908 6732 11920 6788
rect 11520 6720 11920 6732
rect 12000 6788 12400 6800
rect 12000 6732 12012 6788
rect 12068 6732 12332 6788
rect 12388 6732 12400 6788
rect 12000 6720 12400 6732
rect 0 6628 20880 6640
rect 0 6572 11692 6628
rect 11748 6572 20880 6628
rect 0 6560 20880 6572
rect 8480 6468 8880 6480
rect 8480 6412 8492 6468
rect 8548 6412 8812 6468
rect 8868 6412 8880 6468
rect 8480 6400 8880 6412
rect 8960 6468 9360 6480
rect 8960 6412 8972 6468
rect 9028 6412 9292 6468
rect 9348 6412 9360 6468
rect 8960 6400 9360 6412
rect 9440 6468 11440 6480
rect 9440 6412 9452 6468
rect 9508 6412 9772 6468
rect 9828 6412 10092 6468
rect 10148 6412 10412 6468
rect 10468 6412 10732 6468
rect 10788 6412 11052 6468
rect 11108 6412 11372 6468
rect 11428 6412 11440 6468
rect 9440 6400 11440 6412
rect 11520 6468 11920 6480
rect 11520 6412 11532 6468
rect 11588 6412 11852 6468
rect 11908 6412 11920 6468
rect 11520 6400 11920 6412
rect 12000 6468 12400 6480
rect 12000 6412 12012 6468
rect 12068 6412 12332 6468
rect 12388 6412 12400 6468
rect 12000 6400 12400 6412
rect 8480 6308 8880 6320
rect 8480 6252 8492 6308
rect 8548 6252 8812 6308
rect 8868 6252 8880 6308
rect 8480 6240 8880 6252
rect 8960 6308 9360 6320
rect 8960 6252 8972 6308
rect 9028 6252 9292 6308
rect 9348 6252 9360 6308
rect 8960 6240 9360 6252
rect 9440 6308 11440 6320
rect 9440 6252 9452 6308
rect 9508 6252 9772 6308
rect 9828 6252 10092 6308
rect 10148 6252 10412 6308
rect 10468 6252 10732 6308
rect 10788 6252 11052 6308
rect 11108 6252 11372 6308
rect 11428 6252 11440 6308
rect 9440 6240 11440 6252
rect 11520 6308 11920 6320
rect 11520 6252 11532 6308
rect 11588 6252 11852 6308
rect 11908 6252 11920 6308
rect 11520 6240 11920 6252
rect 12000 6308 12400 6320
rect 12000 6252 12012 6308
rect 12068 6252 12332 6308
rect 12388 6252 12400 6308
rect 12000 6240 12400 6252
rect 8480 6148 8880 6160
rect 8480 6092 8492 6148
rect 8548 6092 8812 6148
rect 8868 6092 8880 6148
rect 8480 6080 8880 6092
rect 8960 6148 9360 6160
rect 8960 6092 8972 6148
rect 9028 6092 9292 6148
rect 9348 6092 9360 6148
rect 8960 6080 9360 6092
rect 9440 6148 11440 6160
rect 9440 6092 9452 6148
rect 9508 6092 9772 6148
rect 9828 6092 10092 6148
rect 10148 6092 10412 6148
rect 10468 6092 10732 6148
rect 10788 6092 11052 6148
rect 11108 6092 11372 6148
rect 11428 6092 11440 6148
rect 9440 6080 11440 6092
rect 11520 6148 11920 6160
rect 11520 6092 11532 6148
rect 11588 6092 11852 6148
rect 11908 6092 11920 6148
rect 11520 6080 11920 6092
rect 12000 6148 12400 6160
rect 12000 6092 12012 6148
rect 12068 6092 12332 6148
rect 12388 6092 12400 6148
rect 12000 6080 12400 6092
rect 8480 5988 8880 6000
rect 8480 5932 8492 5988
rect 8548 5932 8812 5988
rect 8868 5932 8880 5988
rect 8480 5920 8880 5932
rect 8960 5988 9360 6000
rect 8960 5932 8972 5988
rect 9028 5932 9292 5988
rect 9348 5932 9360 5988
rect 8960 5920 9360 5932
rect 9440 5988 11440 6000
rect 9440 5932 9452 5988
rect 9508 5932 9772 5988
rect 9828 5932 10092 5988
rect 10148 5932 10412 5988
rect 10468 5932 10732 5988
rect 10788 5932 11052 5988
rect 11108 5932 11372 5988
rect 11428 5932 11440 5988
rect 9440 5920 11440 5932
rect 11520 5988 11920 6000
rect 11520 5932 11532 5988
rect 11588 5932 11852 5988
rect 11908 5932 11920 5988
rect 11520 5920 11920 5932
rect 12000 5988 12400 6000
rect 12000 5932 12012 5988
rect 12068 5932 12332 5988
rect 12388 5932 12400 5988
rect 12000 5920 12400 5932
rect 8480 5828 8880 5840
rect 8480 5772 8492 5828
rect 8548 5772 8812 5828
rect 8868 5772 8880 5828
rect 8480 5760 8880 5772
rect 8960 5828 9360 5840
rect 8960 5772 8972 5828
rect 9028 5772 9292 5828
rect 9348 5772 9360 5828
rect 8960 5760 9360 5772
rect 9440 5828 11440 5840
rect 9440 5772 9452 5828
rect 9508 5772 9772 5828
rect 9828 5772 10092 5828
rect 10148 5772 10412 5828
rect 10468 5772 10732 5828
rect 10788 5772 11052 5828
rect 11108 5772 11372 5828
rect 11428 5772 11440 5828
rect 9440 5760 11440 5772
rect 11520 5828 11920 5840
rect 11520 5772 11532 5828
rect 11588 5772 11852 5828
rect 11908 5772 11920 5828
rect 11520 5760 11920 5772
rect 12000 5828 12400 5840
rect 12000 5772 12012 5828
rect 12068 5772 12332 5828
rect 12388 5772 12400 5828
rect 12000 5760 12400 5772
rect 8480 5668 8880 5680
rect 8480 5612 8492 5668
rect 8548 5612 8812 5668
rect 8868 5612 8880 5668
rect 8480 5600 8880 5612
rect 8960 5668 9360 5680
rect 8960 5612 8972 5668
rect 9028 5612 9292 5668
rect 9348 5612 9360 5668
rect 8960 5600 9360 5612
rect 9440 5668 11440 5680
rect 9440 5612 9452 5668
rect 9508 5612 9772 5668
rect 9828 5612 10092 5668
rect 10148 5612 10412 5668
rect 10468 5612 10732 5668
rect 10788 5612 11052 5668
rect 11108 5612 11372 5668
rect 11428 5612 11440 5668
rect 9440 5600 11440 5612
rect 11520 5668 11920 5680
rect 11520 5612 11532 5668
rect 11588 5612 11852 5668
rect 11908 5612 11920 5668
rect 11520 5600 11920 5612
rect 12000 5668 12400 5680
rect 12000 5612 12012 5668
rect 12068 5612 12332 5668
rect 12388 5612 12400 5668
rect 12000 5600 12400 5612
rect 8480 5508 8880 5520
rect 8480 5452 8492 5508
rect 8548 5452 8812 5508
rect 8868 5452 8880 5508
rect 8480 5440 8880 5452
rect 8960 5508 9360 5520
rect 8960 5452 8972 5508
rect 9028 5452 9292 5508
rect 9348 5452 9360 5508
rect 8960 5440 9360 5452
rect 9440 5508 11440 5520
rect 9440 5452 9452 5508
rect 9508 5452 9772 5508
rect 9828 5452 10092 5508
rect 10148 5452 10412 5508
rect 10468 5452 10732 5508
rect 10788 5452 11052 5508
rect 11108 5452 11372 5508
rect 11428 5452 11440 5508
rect 9440 5440 11440 5452
rect 11520 5508 11920 5520
rect 11520 5452 11532 5508
rect 11588 5452 11852 5508
rect 11908 5452 11920 5508
rect 11520 5440 11920 5452
rect 12000 5508 12400 5520
rect 12000 5452 12012 5508
rect 12068 5452 12332 5508
rect 12388 5452 12400 5508
rect 12000 5440 12400 5452
rect 8480 5348 8880 5360
rect 8480 5292 8492 5348
rect 8548 5292 8812 5348
rect 8868 5292 8880 5348
rect 8480 5280 8880 5292
rect 8960 5348 9360 5360
rect 8960 5292 8972 5348
rect 9028 5292 9292 5348
rect 9348 5292 9360 5348
rect 8960 5280 9360 5292
rect 9440 5348 11440 5360
rect 9440 5292 9452 5348
rect 9508 5292 9772 5348
rect 9828 5292 10092 5348
rect 10148 5292 10412 5348
rect 10468 5292 10732 5348
rect 10788 5292 11052 5348
rect 11108 5292 11372 5348
rect 11428 5292 11440 5348
rect 9440 5280 11440 5292
rect 11520 5348 11920 5360
rect 11520 5292 11532 5348
rect 11588 5292 11852 5348
rect 11908 5292 11920 5348
rect 11520 5280 11920 5292
rect 12000 5348 12400 5360
rect 12000 5292 12012 5348
rect 12068 5292 12332 5348
rect 12388 5292 12400 5348
rect 12000 5280 12400 5292
rect 8480 5188 8880 5200
rect 8480 5132 8492 5188
rect 8548 5132 8812 5188
rect 8868 5132 8880 5188
rect 8480 5120 8880 5132
rect 8960 5188 9360 5200
rect 8960 5132 8972 5188
rect 9028 5132 9292 5188
rect 9348 5132 9360 5188
rect 8960 5120 9360 5132
rect 9440 5188 11440 5200
rect 9440 5132 9452 5188
rect 9508 5132 9772 5188
rect 9828 5132 10092 5188
rect 10148 5132 10412 5188
rect 10468 5132 10732 5188
rect 10788 5132 11052 5188
rect 11108 5132 11372 5188
rect 11428 5132 11440 5188
rect 9440 5120 11440 5132
rect 11520 5188 11920 5200
rect 11520 5132 11532 5188
rect 11588 5132 11852 5188
rect 11908 5132 11920 5188
rect 11520 5120 11920 5132
rect 12000 5188 12400 5200
rect 12000 5132 12012 5188
rect 12068 5132 12332 5188
rect 12388 5132 12400 5188
rect 12000 5120 12400 5132
rect 8480 5028 8880 5040
rect 8480 4972 8492 5028
rect 8548 4972 8812 5028
rect 8868 4972 8880 5028
rect 8480 4960 8880 4972
rect 8960 5028 9360 5040
rect 8960 4972 8972 5028
rect 9028 4972 9292 5028
rect 9348 4972 9360 5028
rect 8960 4960 9360 4972
rect 9440 5028 11440 5040
rect 9440 4972 9452 5028
rect 9508 4972 9772 5028
rect 9828 4972 10092 5028
rect 10148 4972 10412 5028
rect 10468 4972 10732 5028
rect 10788 4972 11052 5028
rect 11108 4972 11372 5028
rect 11428 4972 11440 5028
rect 9440 4960 11440 4972
rect 11520 5028 11920 5040
rect 11520 4972 11532 5028
rect 11588 4972 11852 5028
rect 11908 4972 11920 5028
rect 11520 4960 11920 4972
rect 12000 5028 12400 5040
rect 12000 4972 12012 5028
rect 12068 4972 12332 5028
rect 12388 4972 12400 5028
rect 12000 4960 12400 4972
rect 8480 4868 8880 4880
rect 8480 4812 8492 4868
rect 8548 4812 8812 4868
rect 8868 4812 8880 4868
rect 8480 4800 8880 4812
rect 8960 4868 9360 4880
rect 8960 4812 8972 4868
rect 9028 4812 9292 4868
rect 9348 4812 9360 4868
rect 8960 4800 9360 4812
rect 9440 4868 11440 4880
rect 9440 4812 9452 4868
rect 9508 4812 9772 4868
rect 9828 4812 10092 4868
rect 10148 4812 10412 4868
rect 10468 4812 10732 4868
rect 10788 4812 11052 4868
rect 11108 4812 11372 4868
rect 11428 4812 11440 4868
rect 9440 4800 11440 4812
rect 11520 4868 11920 4880
rect 11520 4812 11532 4868
rect 11588 4812 11852 4868
rect 11908 4812 11920 4868
rect 11520 4800 11920 4812
rect 12000 4868 12400 4880
rect 12000 4812 12012 4868
rect 12068 4812 12332 4868
rect 12388 4812 12400 4868
rect 12000 4800 12400 4812
rect 8480 4708 8880 4720
rect 8480 4652 8492 4708
rect 8548 4652 8812 4708
rect 8868 4652 8880 4708
rect 8480 4640 8880 4652
rect 8960 4708 9360 4720
rect 8960 4652 8972 4708
rect 9028 4652 9292 4708
rect 9348 4652 9360 4708
rect 8960 4640 9360 4652
rect 9440 4708 11440 4720
rect 9440 4652 9452 4708
rect 9508 4652 9772 4708
rect 9828 4652 10092 4708
rect 10148 4652 10412 4708
rect 10468 4652 10732 4708
rect 10788 4652 11052 4708
rect 11108 4652 11372 4708
rect 11428 4652 11440 4708
rect 9440 4640 11440 4652
rect 11520 4708 11920 4720
rect 11520 4652 11532 4708
rect 11588 4652 11852 4708
rect 11908 4652 11920 4708
rect 11520 4640 11920 4652
rect 12000 4708 12400 4720
rect 12000 4652 12012 4708
rect 12068 4652 12332 4708
rect 12388 4652 12400 4708
rect 12000 4640 12400 4652
rect 8480 4548 8880 4560
rect 8480 4492 8492 4548
rect 8548 4492 8812 4548
rect 8868 4492 8880 4548
rect 8480 4480 8880 4492
rect 8960 4548 9360 4560
rect 8960 4492 8972 4548
rect 9028 4492 9292 4548
rect 9348 4492 9360 4548
rect 8960 4480 9360 4492
rect 9440 4548 11440 4560
rect 9440 4492 9452 4548
rect 9508 4492 9772 4548
rect 9828 4492 10092 4548
rect 10148 4492 10412 4548
rect 10468 4492 10732 4548
rect 10788 4492 11052 4548
rect 11108 4492 11372 4548
rect 11428 4492 11440 4548
rect 9440 4480 11440 4492
rect 11520 4548 11920 4560
rect 11520 4492 11532 4548
rect 11588 4492 11852 4548
rect 11908 4492 11920 4548
rect 11520 4480 11920 4492
rect 12000 4548 12400 4560
rect 12000 4492 12012 4548
rect 12068 4492 12332 4548
rect 12388 4492 12400 4548
rect 12000 4480 12400 4492
rect 8480 4388 8880 4400
rect 8480 4332 8492 4388
rect 8548 4332 8812 4388
rect 8868 4332 8880 4388
rect 8480 4320 8880 4332
rect 8960 4388 9360 4400
rect 8960 4332 8972 4388
rect 9028 4332 9292 4388
rect 9348 4332 9360 4388
rect 8960 4320 9360 4332
rect 9440 4388 11440 4400
rect 9440 4332 9452 4388
rect 9508 4332 9772 4388
rect 9828 4332 10092 4388
rect 10148 4332 10412 4388
rect 10468 4332 10732 4388
rect 10788 4332 11052 4388
rect 11108 4332 11372 4388
rect 11428 4332 11440 4388
rect 9440 4320 11440 4332
rect 11520 4388 11920 4400
rect 11520 4332 11532 4388
rect 11588 4332 11852 4388
rect 11908 4332 11920 4388
rect 11520 4320 11920 4332
rect 12000 4388 12400 4400
rect 12000 4332 12012 4388
rect 12068 4332 12332 4388
rect 12388 4332 12400 4388
rect 12000 4320 12400 4332
rect 8480 4228 8880 4240
rect 8480 4172 8492 4228
rect 8548 4172 8812 4228
rect 8868 4172 8880 4228
rect 8480 4160 8880 4172
rect 8960 4228 9360 4240
rect 8960 4172 8972 4228
rect 9028 4172 9292 4228
rect 9348 4172 9360 4228
rect 8960 4160 9360 4172
rect 9440 4228 11440 4240
rect 9440 4172 9452 4228
rect 9508 4172 9772 4228
rect 9828 4172 10092 4228
rect 10148 4172 10412 4228
rect 10468 4172 10732 4228
rect 10788 4172 11052 4228
rect 11108 4172 11372 4228
rect 11428 4172 11440 4228
rect 9440 4160 11440 4172
rect 11520 4228 11920 4240
rect 11520 4172 11532 4228
rect 11588 4172 11852 4228
rect 11908 4172 11920 4228
rect 11520 4160 11920 4172
rect 12000 4228 12400 4240
rect 12000 4172 12012 4228
rect 12068 4172 12332 4228
rect 12388 4172 12400 4228
rect 12000 4160 12400 4172
rect 8480 4068 8880 4080
rect 8480 4012 8492 4068
rect 8548 4012 8812 4068
rect 8868 4012 8880 4068
rect 8480 4000 8880 4012
rect 8960 4068 9360 4080
rect 8960 4012 8972 4068
rect 9028 4012 9292 4068
rect 9348 4012 9360 4068
rect 8960 4000 9360 4012
rect 9440 4068 11440 4080
rect 9440 4012 9452 4068
rect 9508 4012 9772 4068
rect 9828 4012 10092 4068
rect 10148 4012 10412 4068
rect 10468 4012 10732 4068
rect 10788 4012 11052 4068
rect 11108 4012 11372 4068
rect 11428 4012 11440 4068
rect 9440 4000 11440 4012
rect 11520 4068 11920 4080
rect 11520 4012 11532 4068
rect 11588 4012 11852 4068
rect 11908 4012 11920 4068
rect 11520 4000 11920 4012
rect 12000 4068 12400 4080
rect 12000 4012 12012 4068
rect 12068 4012 12332 4068
rect 12388 4012 12400 4068
rect 12000 4000 12400 4012
rect 8480 3908 8880 3920
rect 8480 3852 8492 3908
rect 8548 3852 8812 3908
rect 8868 3852 8880 3908
rect 8480 3840 8880 3852
rect 8960 3908 9360 3920
rect 8960 3852 8972 3908
rect 9028 3852 9292 3908
rect 9348 3852 9360 3908
rect 8960 3840 9360 3852
rect 9440 3908 11440 3920
rect 9440 3852 9452 3908
rect 9508 3852 9772 3908
rect 9828 3852 10092 3908
rect 10148 3852 10412 3908
rect 10468 3852 10732 3908
rect 10788 3852 11052 3908
rect 11108 3852 11372 3908
rect 11428 3852 11440 3908
rect 9440 3840 11440 3852
rect 11520 3908 11920 3920
rect 11520 3852 11532 3908
rect 11588 3852 11852 3908
rect 11908 3852 11920 3908
rect 11520 3840 11920 3852
rect 12000 3908 12400 3920
rect 12000 3852 12012 3908
rect 12068 3852 12332 3908
rect 12388 3852 12400 3908
rect 12000 3840 12400 3852
rect 0 3668 20880 3680
rect 0 3612 9132 3668
rect 9188 3612 20880 3668
rect 0 3600 20880 3612
rect 8480 3428 8880 3440
rect 8480 3372 8492 3428
rect 8548 3372 8812 3428
rect 8868 3372 8880 3428
rect 8480 3360 8880 3372
rect 8960 3428 9360 3440
rect 8960 3372 8972 3428
rect 9028 3372 9292 3428
rect 9348 3372 9360 3428
rect 8960 3360 9360 3372
rect 9440 3428 11440 3440
rect 9440 3372 9452 3428
rect 9508 3372 9772 3428
rect 9828 3372 10092 3428
rect 10148 3372 10412 3428
rect 10468 3372 10732 3428
rect 10788 3372 11052 3428
rect 11108 3372 11372 3428
rect 11428 3372 11440 3428
rect 9440 3360 11440 3372
rect 11520 3428 11920 3440
rect 11520 3372 11532 3428
rect 11588 3372 11852 3428
rect 11908 3372 11920 3428
rect 11520 3360 11920 3372
rect 12000 3428 12400 3440
rect 12000 3372 12012 3428
rect 12068 3372 12332 3428
rect 12388 3372 12400 3428
rect 12000 3360 12400 3372
rect 8480 3268 8880 3280
rect 8480 3212 8492 3268
rect 8548 3212 8812 3268
rect 8868 3212 8880 3268
rect 8480 3200 8880 3212
rect 8960 3268 9360 3280
rect 8960 3212 8972 3268
rect 9028 3212 9292 3268
rect 9348 3212 9360 3268
rect 8960 3200 9360 3212
rect 9440 3268 11440 3280
rect 9440 3212 9452 3268
rect 9508 3212 9772 3268
rect 9828 3212 10092 3268
rect 10148 3212 10412 3268
rect 10468 3212 10732 3268
rect 10788 3212 11052 3268
rect 11108 3212 11372 3268
rect 11428 3212 11440 3268
rect 9440 3200 11440 3212
rect 11520 3268 11920 3280
rect 11520 3212 11532 3268
rect 11588 3212 11852 3268
rect 11908 3212 11920 3268
rect 11520 3200 11920 3212
rect 12000 3268 12400 3280
rect 12000 3212 12012 3268
rect 12068 3212 12332 3268
rect 12388 3212 12400 3268
rect 12000 3200 12400 3212
rect 8480 3108 8880 3120
rect 8480 3052 8492 3108
rect 8548 3052 8812 3108
rect 8868 3052 8880 3108
rect 8480 3040 8880 3052
rect 8960 3108 9360 3120
rect 8960 3052 8972 3108
rect 9028 3052 9292 3108
rect 9348 3052 9360 3108
rect 8960 3040 9360 3052
rect 9440 3108 11440 3120
rect 9440 3052 9452 3108
rect 9508 3052 9772 3108
rect 9828 3052 10092 3108
rect 10148 3052 10412 3108
rect 10468 3052 10732 3108
rect 10788 3052 11052 3108
rect 11108 3052 11372 3108
rect 11428 3052 11440 3108
rect 9440 3040 11440 3052
rect 11520 3108 11920 3120
rect 11520 3052 11532 3108
rect 11588 3052 11852 3108
rect 11908 3052 11920 3108
rect 11520 3040 11920 3052
rect 12000 3108 12400 3120
rect 12000 3052 12012 3108
rect 12068 3052 12332 3108
rect 12388 3052 12400 3108
rect 12000 3040 12400 3052
rect 8480 2948 8880 2960
rect 8480 2892 8492 2948
rect 8548 2892 8812 2948
rect 8868 2892 8880 2948
rect 8480 2880 8880 2892
rect 8960 2948 9360 2960
rect 8960 2892 8972 2948
rect 9028 2892 9292 2948
rect 9348 2892 9360 2948
rect 8960 2880 9360 2892
rect 9440 2948 11440 2960
rect 9440 2892 9452 2948
rect 9508 2892 9772 2948
rect 9828 2892 10092 2948
rect 10148 2892 10412 2948
rect 10468 2892 10732 2948
rect 10788 2892 11052 2948
rect 11108 2892 11372 2948
rect 11428 2892 11440 2948
rect 9440 2880 11440 2892
rect 11520 2948 11920 2960
rect 11520 2892 11532 2948
rect 11588 2892 11852 2948
rect 11908 2892 11920 2948
rect 11520 2880 11920 2892
rect 12000 2948 12400 2960
rect 12000 2892 12012 2948
rect 12068 2892 12332 2948
rect 12388 2892 12400 2948
rect 12000 2880 12400 2892
rect 8480 2788 8880 2800
rect 8480 2732 8492 2788
rect 8548 2732 8812 2788
rect 8868 2732 8880 2788
rect 8480 2720 8880 2732
rect 8960 2788 9360 2800
rect 8960 2732 8972 2788
rect 9028 2732 9292 2788
rect 9348 2732 9360 2788
rect 8960 2720 9360 2732
rect 9440 2788 11440 2800
rect 9440 2732 9452 2788
rect 9508 2732 9772 2788
rect 9828 2732 10092 2788
rect 10148 2732 10412 2788
rect 10468 2732 10732 2788
rect 10788 2732 11052 2788
rect 11108 2732 11372 2788
rect 11428 2732 11440 2788
rect 9440 2720 11440 2732
rect 11520 2788 11920 2800
rect 11520 2732 11532 2788
rect 11588 2732 11852 2788
rect 11908 2732 11920 2788
rect 11520 2720 11920 2732
rect 12000 2788 12400 2800
rect 12000 2732 12012 2788
rect 12068 2732 12332 2788
rect 12388 2732 12400 2788
rect 12000 2720 12400 2732
rect 8480 2628 8880 2640
rect 8480 2572 8492 2628
rect 8548 2572 8812 2628
rect 8868 2572 8880 2628
rect 8480 2560 8880 2572
rect 8960 2628 9360 2640
rect 8960 2572 8972 2628
rect 9028 2572 9292 2628
rect 9348 2572 9360 2628
rect 8960 2560 9360 2572
rect 9440 2628 11440 2640
rect 9440 2572 9452 2628
rect 9508 2572 9772 2628
rect 9828 2572 10092 2628
rect 10148 2572 10412 2628
rect 10468 2572 10732 2628
rect 10788 2572 11052 2628
rect 11108 2572 11372 2628
rect 11428 2572 11440 2628
rect 9440 2560 11440 2572
rect 11520 2628 11920 2640
rect 11520 2572 11532 2628
rect 11588 2572 11852 2628
rect 11908 2572 11920 2628
rect 11520 2560 11920 2572
rect 12000 2628 12400 2640
rect 12000 2572 12012 2628
rect 12068 2572 12332 2628
rect 12388 2572 12400 2628
rect 12000 2560 12400 2572
rect 8480 2468 8880 2480
rect 8480 2412 8492 2468
rect 8548 2412 8812 2468
rect 8868 2412 8880 2468
rect 8480 2400 8880 2412
rect 8960 2468 9360 2480
rect 8960 2412 8972 2468
rect 9028 2412 9292 2468
rect 9348 2412 9360 2468
rect 8960 2400 9360 2412
rect 9440 2468 11440 2480
rect 9440 2412 9452 2468
rect 9508 2412 9772 2468
rect 9828 2412 10092 2468
rect 10148 2412 10412 2468
rect 10468 2412 10732 2468
rect 10788 2412 11052 2468
rect 11108 2412 11372 2468
rect 11428 2412 11440 2468
rect 9440 2400 11440 2412
rect 11520 2468 11920 2480
rect 11520 2412 11532 2468
rect 11588 2412 11852 2468
rect 11908 2412 11920 2468
rect 11520 2400 11920 2412
rect 12000 2468 12400 2480
rect 12000 2412 12012 2468
rect 12068 2412 12332 2468
rect 12388 2412 12400 2468
rect 12000 2400 12400 2412
rect 8480 2308 8880 2320
rect 8480 2252 8492 2308
rect 8548 2252 8812 2308
rect 8868 2252 8880 2308
rect 8480 2240 8880 2252
rect 8960 2308 9360 2320
rect 8960 2252 8972 2308
rect 9028 2252 9292 2308
rect 9348 2252 9360 2308
rect 8960 2240 9360 2252
rect 9440 2308 11440 2320
rect 9440 2252 9452 2308
rect 9508 2252 9772 2308
rect 9828 2252 10092 2308
rect 10148 2252 10412 2308
rect 10468 2252 10732 2308
rect 10788 2252 11052 2308
rect 11108 2252 11372 2308
rect 11428 2252 11440 2308
rect 9440 2240 11440 2252
rect 11520 2308 11920 2320
rect 11520 2252 11532 2308
rect 11588 2252 11852 2308
rect 11908 2252 11920 2308
rect 11520 2240 11920 2252
rect 12000 2308 12400 2320
rect 12000 2252 12012 2308
rect 12068 2252 12332 2308
rect 12388 2252 12400 2308
rect 12000 2240 12400 2252
rect 8480 2148 8880 2160
rect 8480 2092 8492 2148
rect 8548 2092 8812 2148
rect 8868 2092 8880 2148
rect 8480 2080 8880 2092
rect 8960 2148 9360 2160
rect 8960 2092 8972 2148
rect 9028 2092 9292 2148
rect 9348 2092 9360 2148
rect 8960 2080 9360 2092
rect 9440 2148 11440 2160
rect 9440 2092 9452 2148
rect 9508 2092 9772 2148
rect 9828 2092 10092 2148
rect 10148 2092 10412 2148
rect 10468 2092 10732 2148
rect 10788 2092 11052 2148
rect 11108 2092 11372 2148
rect 11428 2092 11440 2148
rect 9440 2080 11440 2092
rect 11520 2148 11920 2160
rect 11520 2092 11532 2148
rect 11588 2092 11852 2148
rect 11908 2092 11920 2148
rect 11520 2080 11920 2092
rect 12000 2148 12400 2160
rect 12000 2092 12012 2148
rect 12068 2092 12332 2148
rect 12388 2092 12400 2148
rect 12000 2080 12400 2092
rect 8480 1988 8880 2000
rect 8480 1932 8492 1988
rect 8548 1932 8812 1988
rect 8868 1932 8880 1988
rect 8480 1920 8880 1932
rect 8960 1988 9360 2000
rect 8960 1932 8972 1988
rect 9028 1932 9292 1988
rect 9348 1932 9360 1988
rect 8960 1920 9360 1932
rect 9440 1988 11440 2000
rect 9440 1932 9452 1988
rect 9508 1932 9772 1988
rect 9828 1932 10092 1988
rect 10148 1932 10412 1988
rect 10468 1932 10732 1988
rect 10788 1932 11052 1988
rect 11108 1932 11372 1988
rect 11428 1932 11440 1988
rect 9440 1920 11440 1932
rect 11520 1988 11920 2000
rect 11520 1932 11532 1988
rect 11588 1932 11852 1988
rect 11908 1932 11920 1988
rect 11520 1920 11920 1932
rect 12000 1988 12400 2000
rect 12000 1932 12012 1988
rect 12068 1932 12332 1988
rect 12388 1932 12400 1988
rect 12000 1920 12400 1932
rect 0 1828 20880 1840
rect 0 1772 12172 1828
rect 12228 1772 20880 1828
rect 0 1760 20880 1772
rect 8480 1668 8880 1680
rect 8480 1612 8492 1668
rect 8548 1612 8812 1668
rect 8868 1612 8880 1668
rect 8480 1600 8880 1612
rect 8960 1668 9360 1680
rect 8960 1612 8972 1668
rect 9028 1612 9292 1668
rect 9348 1612 9360 1668
rect 8960 1600 9360 1612
rect 9440 1668 11440 1680
rect 9440 1612 9452 1668
rect 9508 1612 9772 1668
rect 9828 1612 10092 1668
rect 10148 1612 10412 1668
rect 10468 1612 10732 1668
rect 10788 1612 11052 1668
rect 11108 1612 11372 1668
rect 11428 1612 11440 1668
rect 9440 1600 11440 1612
rect 11520 1668 11920 1680
rect 11520 1612 11532 1668
rect 11588 1612 11852 1668
rect 11908 1612 11920 1668
rect 11520 1600 11920 1612
rect 12000 1668 12400 1680
rect 12000 1612 12012 1668
rect 12068 1612 12332 1668
rect 12388 1612 12400 1668
rect 12000 1600 12400 1612
rect 8480 1508 8880 1520
rect 8480 1452 8492 1508
rect 8548 1452 8812 1508
rect 8868 1452 8880 1508
rect 8480 1440 8880 1452
rect 8960 1508 9360 1520
rect 8960 1452 8972 1508
rect 9028 1452 9292 1508
rect 9348 1452 9360 1508
rect 8960 1440 9360 1452
rect 9440 1508 11440 1520
rect 9440 1452 9452 1508
rect 9508 1452 9772 1508
rect 9828 1452 10092 1508
rect 10148 1452 10412 1508
rect 10468 1452 10732 1508
rect 10788 1452 11052 1508
rect 11108 1452 11372 1508
rect 11428 1452 11440 1508
rect 9440 1440 11440 1452
rect 11520 1508 11920 1520
rect 11520 1452 11532 1508
rect 11588 1452 11852 1508
rect 11908 1452 11920 1508
rect 11520 1440 11920 1452
rect 12000 1508 12400 1520
rect 12000 1452 12012 1508
rect 12068 1452 12332 1508
rect 12388 1452 12400 1508
rect 12000 1440 12400 1452
rect 8480 1348 8880 1360
rect 8480 1292 8492 1348
rect 8548 1292 8812 1348
rect 8868 1292 8880 1348
rect 8480 1280 8880 1292
rect 8960 1348 9360 1360
rect 8960 1292 8972 1348
rect 9028 1292 9292 1348
rect 9348 1292 9360 1348
rect 8960 1280 9360 1292
rect 9440 1348 11440 1360
rect 9440 1292 9452 1348
rect 9508 1292 9772 1348
rect 9828 1292 10092 1348
rect 10148 1292 10412 1348
rect 10468 1292 10732 1348
rect 10788 1292 11052 1348
rect 11108 1292 11372 1348
rect 11428 1292 11440 1348
rect 9440 1280 11440 1292
rect 11520 1348 11920 1360
rect 11520 1292 11532 1348
rect 11588 1292 11852 1348
rect 11908 1292 11920 1348
rect 11520 1280 11920 1292
rect 12000 1348 12400 1360
rect 12000 1292 12012 1348
rect 12068 1292 12332 1348
rect 12388 1292 12400 1348
rect 12000 1280 12400 1292
rect 8480 1188 8880 1200
rect 8480 1132 8492 1188
rect 8548 1132 8812 1188
rect 8868 1132 8880 1188
rect 8480 1120 8880 1132
rect 8960 1188 9360 1200
rect 8960 1132 8972 1188
rect 9028 1132 9292 1188
rect 9348 1132 9360 1188
rect 8960 1120 9360 1132
rect 9440 1188 11440 1200
rect 9440 1132 9452 1188
rect 9508 1132 9772 1188
rect 9828 1132 10092 1188
rect 10148 1132 10412 1188
rect 10468 1132 10732 1188
rect 10788 1132 11052 1188
rect 11108 1132 11372 1188
rect 11428 1132 11440 1188
rect 9440 1120 11440 1132
rect 11520 1188 11920 1200
rect 11520 1132 11532 1188
rect 11588 1132 11852 1188
rect 11908 1132 11920 1188
rect 11520 1120 11920 1132
rect 12000 1188 12400 1200
rect 12000 1132 12012 1188
rect 12068 1132 12332 1188
rect 12388 1132 12400 1188
rect 12000 1120 12400 1132
rect 8480 1028 8880 1040
rect 8480 972 8492 1028
rect 8548 972 8812 1028
rect 8868 972 8880 1028
rect 8480 960 8880 972
rect 8960 1028 9360 1040
rect 8960 972 8972 1028
rect 9028 972 9292 1028
rect 9348 972 9360 1028
rect 8960 960 9360 972
rect 9440 1028 11440 1040
rect 9440 972 9452 1028
rect 9508 972 9772 1028
rect 9828 972 10092 1028
rect 10148 972 10412 1028
rect 10468 972 10732 1028
rect 10788 972 11052 1028
rect 11108 972 11372 1028
rect 11428 972 11440 1028
rect 9440 960 11440 972
rect 11520 1028 11920 1040
rect 11520 972 11532 1028
rect 11588 972 11852 1028
rect 11908 972 11920 1028
rect 11520 960 11920 972
rect 12000 1028 12400 1040
rect 12000 972 12012 1028
rect 12068 972 12332 1028
rect 12388 972 12400 1028
rect 12000 960 12400 972
rect 0 788 20880 800
rect 0 732 8652 788
rect 8708 732 20880 788
rect 0 720 20880 732
rect 8480 548 8880 560
rect 8480 492 8492 548
rect 8548 492 8812 548
rect 8868 492 8880 548
rect 8480 480 8880 492
rect 8960 548 9360 560
rect 8960 492 8972 548
rect 9028 492 9292 548
rect 9348 492 9360 548
rect 8960 480 9360 492
rect 9440 548 11440 560
rect 9440 492 9452 548
rect 9508 492 9772 548
rect 9828 492 10092 548
rect 10148 492 10412 548
rect 10468 492 10732 548
rect 10788 492 11052 548
rect 11108 492 11372 548
rect 11428 492 11440 548
rect 9440 480 11440 492
rect 11520 548 11920 560
rect 11520 492 11532 548
rect 11588 492 11852 548
rect 11908 492 11920 548
rect 11520 480 11920 492
rect 12000 548 12400 560
rect 12000 492 12012 548
rect 12068 492 12332 548
rect 12388 492 12400 548
rect 12000 480 12400 492
rect 8480 388 8880 400
rect 8480 332 8492 388
rect 8548 332 8812 388
rect 8868 332 8880 388
rect 8480 320 8880 332
rect 8960 388 9360 400
rect 8960 332 8972 388
rect 9028 332 9292 388
rect 9348 332 9360 388
rect 8960 320 9360 332
rect 9440 388 11440 400
rect 9440 332 9452 388
rect 9508 332 9772 388
rect 9828 332 10092 388
rect 10148 332 10412 388
rect 10468 332 10732 388
rect 10788 332 11052 388
rect 11108 332 11372 388
rect 11428 332 11440 388
rect 9440 320 11440 332
rect 11520 388 11920 400
rect 11520 332 11532 388
rect 11588 332 11852 388
rect 11908 332 11920 388
rect 11520 320 11920 332
rect 12000 388 12400 400
rect 12000 332 12012 388
rect 12068 332 12332 388
rect 12388 332 12400 388
rect 12000 320 12400 332
rect 8480 228 8880 240
rect 8480 172 8492 228
rect 8548 172 8812 228
rect 8868 172 8880 228
rect 8480 160 8880 172
rect 8960 228 9360 240
rect 8960 172 8972 228
rect 9028 172 9292 228
rect 9348 172 9360 228
rect 8960 160 9360 172
rect 9440 228 11440 240
rect 9440 172 9452 228
rect 9508 172 9772 228
rect 9828 172 10092 228
rect 10148 172 10412 228
rect 10468 172 10732 228
rect 10788 172 11052 228
rect 11108 172 11372 228
rect 11428 172 11440 228
rect 9440 160 11440 172
rect 11520 228 11920 240
rect 11520 172 11532 228
rect 11588 172 11852 228
rect 11908 172 11920 228
rect 11520 160 11920 172
rect 12000 228 12400 240
rect 12000 172 12012 228
rect 12068 172 12332 228
rect 12388 172 12400 228
rect 12000 160 12400 172
rect 8480 68 8880 80
rect 8480 12 8492 68
rect 8548 12 8812 68
rect 8868 12 8880 68
rect 8480 0 8880 12
rect 8960 68 9360 80
rect 8960 12 8972 68
rect 9028 12 9292 68
rect 9348 12 9360 68
rect 8960 0 9360 12
rect 9440 68 11440 80
rect 9440 12 9452 68
rect 9508 12 9772 68
rect 9828 12 10092 68
rect 10148 12 10412 68
rect 10468 12 10732 68
rect 10788 12 11052 68
rect 11108 12 11372 68
rect 11428 12 11440 68
rect 9440 0 11440 12
rect 11520 68 11920 80
rect 11520 12 11532 68
rect 11588 12 11852 68
rect 11908 12 11920 68
rect 11520 0 11920 12
rect 12000 68 12400 80
rect 12000 12 12012 68
rect 12068 12 12332 68
rect 12388 12 12400 68
rect 12000 0 12400 12
<< via2 >>
rect 8492 31426 8548 31428
rect 8492 31374 8494 31426
rect 8494 31374 8546 31426
rect 8546 31374 8548 31426
rect 8492 31372 8548 31374
rect 8812 31426 8868 31428
rect 8812 31374 8814 31426
rect 8814 31374 8866 31426
rect 8866 31374 8868 31426
rect 8812 31372 8868 31374
rect 8972 31426 9028 31428
rect 8972 31374 8974 31426
rect 8974 31374 9026 31426
rect 9026 31374 9028 31426
rect 8972 31372 9028 31374
rect 9292 31426 9348 31428
rect 9292 31374 9294 31426
rect 9294 31374 9346 31426
rect 9346 31374 9348 31426
rect 9292 31372 9348 31374
rect 9452 31426 9508 31428
rect 9452 31374 9454 31426
rect 9454 31374 9506 31426
rect 9506 31374 9508 31426
rect 9452 31372 9508 31374
rect 9772 31426 9828 31428
rect 9772 31374 9774 31426
rect 9774 31374 9826 31426
rect 9826 31374 9828 31426
rect 9772 31372 9828 31374
rect 10092 31426 10148 31428
rect 10092 31374 10094 31426
rect 10094 31374 10146 31426
rect 10146 31374 10148 31426
rect 10092 31372 10148 31374
rect 10412 31426 10468 31428
rect 10412 31374 10414 31426
rect 10414 31374 10466 31426
rect 10466 31374 10468 31426
rect 10412 31372 10468 31374
rect 10732 31426 10788 31428
rect 10732 31374 10734 31426
rect 10734 31374 10786 31426
rect 10786 31374 10788 31426
rect 10732 31372 10788 31374
rect 11052 31426 11108 31428
rect 11052 31374 11054 31426
rect 11054 31374 11106 31426
rect 11106 31374 11108 31426
rect 11052 31372 11108 31374
rect 11372 31426 11428 31428
rect 11372 31374 11374 31426
rect 11374 31374 11426 31426
rect 11426 31374 11428 31426
rect 11372 31372 11428 31374
rect 11532 31426 11588 31428
rect 11532 31374 11534 31426
rect 11534 31374 11586 31426
rect 11586 31374 11588 31426
rect 11532 31372 11588 31374
rect 11852 31426 11908 31428
rect 11852 31374 11854 31426
rect 11854 31374 11906 31426
rect 11906 31374 11908 31426
rect 11852 31372 11908 31374
rect 12012 31426 12068 31428
rect 12012 31374 12014 31426
rect 12014 31374 12066 31426
rect 12066 31374 12068 31426
rect 12012 31372 12068 31374
rect 12332 31426 12388 31428
rect 12332 31374 12334 31426
rect 12334 31374 12386 31426
rect 12386 31374 12388 31426
rect 12332 31372 12388 31374
rect 8492 31266 8548 31268
rect 8492 31214 8494 31266
rect 8494 31214 8546 31266
rect 8546 31214 8548 31266
rect 8492 31212 8548 31214
rect 8812 31266 8868 31268
rect 8812 31214 8814 31266
rect 8814 31214 8866 31266
rect 8866 31214 8868 31266
rect 8812 31212 8868 31214
rect 8972 31266 9028 31268
rect 8972 31214 8974 31266
rect 8974 31214 9026 31266
rect 9026 31214 9028 31266
rect 8972 31212 9028 31214
rect 9292 31266 9348 31268
rect 9292 31214 9294 31266
rect 9294 31214 9346 31266
rect 9346 31214 9348 31266
rect 9292 31212 9348 31214
rect 9452 31266 9508 31268
rect 9452 31214 9454 31266
rect 9454 31214 9506 31266
rect 9506 31214 9508 31266
rect 9452 31212 9508 31214
rect 9772 31266 9828 31268
rect 9772 31214 9774 31266
rect 9774 31214 9826 31266
rect 9826 31214 9828 31266
rect 9772 31212 9828 31214
rect 10092 31266 10148 31268
rect 10092 31214 10094 31266
rect 10094 31214 10146 31266
rect 10146 31214 10148 31266
rect 10092 31212 10148 31214
rect 10412 31266 10468 31268
rect 10412 31214 10414 31266
rect 10414 31214 10466 31266
rect 10466 31214 10468 31266
rect 10412 31212 10468 31214
rect 10732 31266 10788 31268
rect 10732 31214 10734 31266
rect 10734 31214 10786 31266
rect 10786 31214 10788 31266
rect 10732 31212 10788 31214
rect 11052 31266 11108 31268
rect 11052 31214 11054 31266
rect 11054 31214 11106 31266
rect 11106 31214 11108 31266
rect 11052 31212 11108 31214
rect 11372 31266 11428 31268
rect 11372 31214 11374 31266
rect 11374 31214 11426 31266
rect 11426 31214 11428 31266
rect 11372 31212 11428 31214
rect 11532 31266 11588 31268
rect 11532 31214 11534 31266
rect 11534 31214 11586 31266
rect 11586 31214 11588 31266
rect 11532 31212 11588 31214
rect 11852 31266 11908 31268
rect 11852 31214 11854 31266
rect 11854 31214 11906 31266
rect 11906 31214 11908 31266
rect 11852 31212 11908 31214
rect 12012 31266 12068 31268
rect 12012 31214 12014 31266
rect 12014 31214 12066 31266
rect 12066 31214 12068 31266
rect 12012 31212 12068 31214
rect 12332 31266 12388 31268
rect 12332 31214 12334 31266
rect 12334 31214 12386 31266
rect 12386 31214 12388 31266
rect 12332 31212 12388 31214
rect 8492 31106 8548 31108
rect 8492 31054 8494 31106
rect 8494 31054 8546 31106
rect 8546 31054 8548 31106
rect 8492 31052 8548 31054
rect 8812 31106 8868 31108
rect 8812 31054 8814 31106
rect 8814 31054 8866 31106
rect 8866 31054 8868 31106
rect 8812 31052 8868 31054
rect 8972 31106 9028 31108
rect 8972 31054 8974 31106
rect 8974 31054 9026 31106
rect 9026 31054 9028 31106
rect 8972 31052 9028 31054
rect 9292 31106 9348 31108
rect 9292 31054 9294 31106
rect 9294 31054 9346 31106
rect 9346 31054 9348 31106
rect 9292 31052 9348 31054
rect 9452 31106 9508 31108
rect 9452 31054 9454 31106
rect 9454 31054 9506 31106
rect 9506 31054 9508 31106
rect 9452 31052 9508 31054
rect 9772 31106 9828 31108
rect 9772 31054 9774 31106
rect 9774 31054 9826 31106
rect 9826 31054 9828 31106
rect 9772 31052 9828 31054
rect 10092 31106 10148 31108
rect 10092 31054 10094 31106
rect 10094 31054 10146 31106
rect 10146 31054 10148 31106
rect 10092 31052 10148 31054
rect 10412 31106 10468 31108
rect 10412 31054 10414 31106
rect 10414 31054 10466 31106
rect 10466 31054 10468 31106
rect 10412 31052 10468 31054
rect 10732 31106 10788 31108
rect 10732 31054 10734 31106
rect 10734 31054 10786 31106
rect 10786 31054 10788 31106
rect 10732 31052 10788 31054
rect 11052 31106 11108 31108
rect 11052 31054 11054 31106
rect 11054 31054 11106 31106
rect 11106 31054 11108 31106
rect 11052 31052 11108 31054
rect 11372 31106 11428 31108
rect 11372 31054 11374 31106
rect 11374 31054 11426 31106
rect 11426 31054 11428 31106
rect 11372 31052 11428 31054
rect 11532 31106 11588 31108
rect 11532 31054 11534 31106
rect 11534 31054 11586 31106
rect 11586 31054 11588 31106
rect 11532 31052 11588 31054
rect 11852 31106 11908 31108
rect 11852 31054 11854 31106
rect 11854 31054 11906 31106
rect 11906 31054 11908 31106
rect 11852 31052 11908 31054
rect 12012 31106 12068 31108
rect 12012 31054 12014 31106
rect 12014 31054 12066 31106
rect 12066 31054 12068 31106
rect 12012 31052 12068 31054
rect 12332 31106 12388 31108
rect 12332 31054 12334 31106
rect 12334 31054 12386 31106
rect 12386 31054 12388 31106
rect 12332 31052 12388 31054
rect 8492 30946 8548 30948
rect 8492 30894 8494 30946
rect 8494 30894 8546 30946
rect 8546 30894 8548 30946
rect 8492 30892 8548 30894
rect 8812 30946 8868 30948
rect 8812 30894 8814 30946
rect 8814 30894 8866 30946
rect 8866 30894 8868 30946
rect 8812 30892 8868 30894
rect 8972 30946 9028 30948
rect 8972 30894 8974 30946
rect 8974 30894 9026 30946
rect 9026 30894 9028 30946
rect 8972 30892 9028 30894
rect 9292 30946 9348 30948
rect 9292 30894 9294 30946
rect 9294 30894 9346 30946
rect 9346 30894 9348 30946
rect 9292 30892 9348 30894
rect 9452 30946 9508 30948
rect 9452 30894 9454 30946
rect 9454 30894 9506 30946
rect 9506 30894 9508 30946
rect 9452 30892 9508 30894
rect 9772 30946 9828 30948
rect 9772 30894 9774 30946
rect 9774 30894 9826 30946
rect 9826 30894 9828 30946
rect 9772 30892 9828 30894
rect 10092 30946 10148 30948
rect 10092 30894 10094 30946
rect 10094 30894 10146 30946
rect 10146 30894 10148 30946
rect 10092 30892 10148 30894
rect 10412 30946 10468 30948
rect 10412 30894 10414 30946
rect 10414 30894 10466 30946
rect 10466 30894 10468 30946
rect 10412 30892 10468 30894
rect 10732 30946 10788 30948
rect 10732 30894 10734 30946
rect 10734 30894 10786 30946
rect 10786 30894 10788 30946
rect 10732 30892 10788 30894
rect 11052 30946 11108 30948
rect 11052 30894 11054 30946
rect 11054 30894 11106 30946
rect 11106 30894 11108 30946
rect 11052 30892 11108 30894
rect 11372 30946 11428 30948
rect 11372 30894 11374 30946
rect 11374 30894 11426 30946
rect 11426 30894 11428 30946
rect 11372 30892 11428 30894
rect 11532 30946 11588 30948
rect 11532 30894 11534 30946
rect 11534 30894 11586 30946
rect 11586 30894 11588 30946
rect 11532 30892 11588 30894
rect 11852 30946 11908 30948
rect 11852 30894 11854 30946
rect 11854 30894 11906 30946
rect 11906 30894 11908 30946
rect 11852 30892 11908 30894
rect 12012 30946 12068 30948
rect 12012 30894 12014 30946
rect 12014 30894 12066 30946
rect 12066 30894 12068 30946
rect 12012 30892 12068 30894
rect 12332 30946 12388 30948
rect 12332 30894 12334 30946
rect 12334 30894 12386 30946
rect 12386 30894 12388 30946
rect 12332 30892 12388 30894
rect 8492 30786 8548 30788
rect 8492 30734 8494 30786
rect 8494 30734 8546 30786
rect 8546 30734 8548 30786
rect 8492 30732 8548 30734
rect 8812 30786 8868 30788
rect 8812 30734 8814 30786
rect 8814 30734 8866 30786
rect 8866 30734 8868 30786
rect 8812 30732 8868 30734
rect 8972 30786 9028 30788
rect 8972 30734 8974 30786
rect 8974 30734 9026 30786
rect 9026 30734 9028 30786
rect 8972 30732 9028 30734
rect 9292 30786 9348 30788
rect 9292 30734 9294 30786
rect 9294 30734 9346 30786
rect 9346 30734 9348 30786
rect 9292 30732 9348 30734
rect 9452 30786 9508 30788
rect 9452 30734 9454 30786
rect 9454 30734 9506 30786
rect 9506 30734 9508 30786
rect 9452 30732 9508 30734
rect 9772 30786 9828 30788
rect 9772 30734 9774 30786
rect 9774 30734 9826 30786
rect 9826 30734 9828 30786
rect 9772 30732 9828 30734
rect 10092 30786 10148 30788
rect 10092 30734 10094 30786
rect 10094 30734 10146 30786
rect 10146 30734 10148 30786
rect 10092 30732 10148 30734
rect 10412 30786 10468 30788
rect 10412 30734 10414 30786
rect 10414 30734 10466 30786
rect 10466 30734 10468 30786
rect 10412 30732 10468 30734
rect 10732 30786 10788 30788
rect 10732 30734 10734 30786
rect 10734 30734 10786 30786
rect 10786 30734 10788 30786
rect 10732 30732 10788 30734
rect 11052 30786 11108 30788
rect 11052 30734 11054 30786
rect 11054 30734 11106 30786
rect 11106 30734 11108 30786
rect 11052 30732 11108 30734
rect 11372 30786 11428 30788
rect 11372 30734 11374 30786
rect 11374 30734 11426 30786
rect 11426 30734 11428 30786
rect 11372 30732 11428 30734
rect 11532 30786 11588 30788
rect 11532 30734 11534 30786
rect 11534 30734 11586 30786
rect 11586 30734 11588 30786
rect 11532 30732 11588 30734
rect 11852 30786 11908 30788
rect 11852 30734 11854 30786
rect 11854 30734 11906 30786
rect 11906 30734 11908 30786
rect 11852 30732 11908 30734
rect 12012 30786 12068 30788
rect 12012 30734 12014 30786
rect 12014 30734 12066 30786
rect 12066 30734 12068 30786
rect 12012 30732 12068 30734
rect 12332 30786 12388 30788
rect 12332 30734 12334 30786
rect 12334 30734 12386 30786
rect 12386 30734 12388 30786
rect 12332 30732 12388 30734
rect 8492 30626 8548 30628
rect 8492 30574 8494 30626
rect 8494 30574 8546 30626
rect 8546 30574 8548 30626
rect 8492 30572 8548 30574
rect 8812 30626 8868 30628
rect 8812 30574 8814 30626
rect 8814 30574 8866 30626
rect 8866 30574 8868 30626
rect 8812 30572 8868 30574
rect 8972 30626 9028 30628
rect 8972 30574 8974 30626
rect 8974 30574 9026 30626
rect 9026 30574 9028 30626
rect 8972 30572 9028 30574
rect 9292 30626 9348 30628
rect 9292 30574 9294 30626
rect 9294 30574 9346 30626
rect 9346 30574 9348 30626
rect 9292 30572 9348 30574
rect 9452 30626 9508 30628
rect 9452 30574 9454 30626
rect 9454 30574 9506 30626
rect 9506 30574 9508 30626
rect 9452 30572 9508 30574
rect 9772 30626 9828 30628
rect 9772 30574 9774 30626
rect 9774 30574 9826 30626
rect 9826 30574 9828 30626
rect 9772 30572 9828 30574
rect 10092 30626 10148 30628
rect 10092 30574 10094 30626
rect 10094 30574 10146 30626
rect 10146 30574 10148 30626
rect 10092 30572 10148 30574
rect 10412 30626 10468 30628
rect 10412 30574 10414 30626
rect 10414 30574 10466 30626
rect 10466 30574 10468 30626
rect 10412 30572 10468 30574
rect 10732 30626 10788 30628
rect 10732 30574 10734 30626
rect 10734 30574 10786 30626
rect 10786 30574 10788 30626
rect 10732 30572 10788 30574
rect 11052 30626 11108 30628
rect 11052 30574 11054 30626
rect 11054 30574 11106 30626
rect 11106 30574 11108 30626
rect 11052 30572 11108 30574
rect 11372 30626 11428 30628
rect 11372 30574 11374 30626
rect 11374 30574 11426 30626
rect 11426 30574 11428 30626
rect 11372 30572 11428 30574
rect 11532 30626 11588 30628
rect 11532 30574 11534 30626
rect 11534 30574 11586 30626
rect 11586 30574 11588 30626
rect 11532 30572 11588 30574
rect 11852 30626 11908 30628
rect 11852 30574 11854 30626
rect 11854 30574 11906 30626
rect 11906 30574 11908 30626
rect 11852 30572 11908 30574
rect 12012 30626 12068 30628
rect 12012 30574 12014 30626
rect 12014 30574 12066 30626
rect 12066 30574 12068 30626
rect 12012 30572 12068 30574
rect 12332 30626 12388 30628
rect 12332 30574 12334 30626
rect 12334 30574 12386 30626
rect 12386 30574 12388 30626
rect 12332 30572 12388 30574
rect 8492 30466 8548 30468
rect 8492 30414 8494 30466
rect 8494 30414 8546 30466
rect 8546 30414 8548 30466
rect 8492 30412 8548 30414
rect 8812 30466 8868 30468
rect 8812 30414 8814 30466
rect 8814 30414 8866 30466
rect 8866 30414 8868 30466
rect 8812 30412 8868 30414
rect 8972 30466 9028 30468
rect 8972 30414 8974 30466
rect 8974 30414 9026 30466
rect 9026 30414 9028 30466
rect 8972 30412 9028 30414
rect 9292 30466 9348 30468
rect 9292 30414 9294 30466
rect 9294 30414 9346 30466
rect 9346 30414 9348 30466
rect 9292 30412 9348 30414
rect 9452 30466 9508 30468
rect 9452 30414 9454 30466
rect 9454 30414 9506 30466
rect 9506 30414 9508 30466
rect 9452 30412 9508 30414
rect 9772 30466 9828 30468
rect 9772 30414 9774 30466
rect 9774 30414 9826 30466
rect 9826 30414 9828 30466
rect 9772 30412 9828 30414
rect 10092 30466 10148 30468
rect 10092 30414 10094 30466
rect 10094 30414 10146 30466
rect 10146 30414 10148 30466
rect 10092 30412 10148 30414
rect 10412 30466 10468 30468
rect 10412 30414 10414 30466
rect 10414 30414 10466 30466
rect 10466 30414 10468 30466
rect 10412 30412 10468 30414
rect 10732 30466 10788 30468
rect 10732 30414 10734 30466
rect 10734 30414 10786 30466
rect 10786 30414 10788 30466
rect 10732 30412 10788 30414
rect 11052 30466 11108 30468
rect 11052 30414 11054 30466
rect 11054 30414 11106 30466
rect 11106 30414 11108 30466
rect 11052 30412 11108 30414
rect 11372 30466 11428 30468
rect 11372 30414 11374 30466
rect 11374 30414 11426 30466
rect 11426 30414 11428 30466
rect 11372 30412 11428 30414
rect 11532 30466 11588 30468
rect 11532 30414 11534 30466
rect 11534 30414 11586 30466
rect 11586 30414 11588 30466
rect 11532 30412 11588 30414
rect 11852 30466 11908 30468
rect 11852 30414 11854 30466
rect 11854 30414 11906 30466
rect 11906 30414 11908 30466
rect 11852 30412 11908 30414
rect 12012 30466 12068 30468
rect 12012 30414 12014 30466
rect 12014 30414 12066 30466
rect 12066 30414 12068 30466
rect 12012 30412 12068 30414
rect 12332 30466 12388 30468
rect 12332 30414 12334 30466
rect 12334 30414 12386 30466
rect 12386 30414 12388 30466
rect 12332 30412 12388 30414
rect 8492 30306 8548 30308
rect 8492 30254 8494 30306
rect 8494 30254 8546 30306
rect 8546 30254 8548 30306
rect 8492 30252 8548 30254
rect 8812 30306 8868 30308
rect 8812 30254 8814 30306
rect 8814 30254 8866 30306
rect 8866 30254 8868 30306
rect 8812 30252 8868 30254
rect 8972 30306 9028 30308
rect 8972 30254 8974 30306
rect 8974 30254 9026 30306
rect 9026 30254 9028 30306
rect 8972 30252 9028 30254
rect 9292 30306 9348 30308
rect 9292 30254 9294 30306
rect 9294 30254 9346 30306
rect 9346 30254 9348 30306
rect 9292 30252 9348 30254
rect 9452 30306 9508 30308
rect 9452 30254 9454 30306
rect 9454 30254 9506 30306
rect 9506 30254 9508 30306
rect 9452 30252 9508 30254
rect 9772 30306 9828 30308
rect 9772 30254 9774 30306
rect 9774 30254 9826 30306
rect 9826 30254 9828 30306
rect 9772 30252 9828 30254
rect 10092 30306 10148 30308
rect 10092 30254 10094 30306
rect 10094 30254 10146 30306
rect 10146 30254 10148 30306
rect 10092 30252 10148 30254
rect 10412 30306 10468 30308
rect 10412 30254 10414 30306
rect 10414 30254 10466 30306
rect 10466 30254 10468 30306
rect 10412 30252 10468 30254
rect 10732 30306 10788 30308
rect 10732 30254 10734 30306
rect 10734 30254 10786 30306
rect 10786 30254 10788 30306
rect 10732 30252 10788 30254
rect 11052 30306 11108 30308
rect 11052 30254 11054 30306
rect 11054 30254 11106 30306
rect 11106 30254 11108 30306
rect 11052 30252 11108 30254
rect 11372 30306 11428 30308
rect 11372 30254 11374 30306
rect 11374 30254 11426 30306
rect 11426 30254 11428 30306
rect 11372 30252 11428 30254
rect 11532 30306 11588 30308
rect 11532 30254 11534 30306
rect 11534 30254 11586 30306
rect 11586 30254 11588 30306
rect 11532 30252 11588 30254
rect 11852 30306 11908 30308
rect 11852 30254 11854 30306
rect 11854 30254 11906 30306
rect 11906 30254 11908 30306
rect 11852 30252 11908 30254
rect 12012 30306 12068 30308
rect 12012 30254 12014 30306
rect 12014 30254 12066 30306
rect 12066 30254 12068 30306
rect 12012 30252 12068 30254
rect 12332 30306 12388 30308
rect 12332 30254 12334 30306
rect 12334 30254 12386 30306
rect 12386 30254 12388 30306
rect 12332 30252 12388 30254
rect 9132 30092 9188 30148
rect 8492 29986 8548 29988
rect 8492 29934 8494 29986
rect 8494 29934 8546 29986
rect 8546 29934 8548 29986
rect 8492 29932 8548 29934
rect 8812 29986 8868 29988
rect 8812 29934 8814 29986
rect 8814 29934 8866 29986
rect 8866 29934 8868 29986
rect 8812 29932 8868 29934
rect 8972 29986 9028 29988
rect 8972 29934 8974 29986
rect 8974 29934 9026 29986
rect 9026 29934 9028 29986
rect 8972 29932 9028 29934
rect 9292 29986 9348 29988
rect 9292 29934 9294 29986
rect 9294 29934 9346 29986
rect 9346 29934 9348 29986
rect 9292 29932 9348 29934
rect 9452 29986 9508 29988
rect 9452 29934 9454 29986
rect 9454 29934 9506 29986
rect 9506 29934 9508 29986
rect 9452 29932 9508 29934
rect 9772 29986 9828 29988
rect 9772 29934 9774 29986
rect 9774 29934 9826 29986
rect 9826 29934 9828 29986
rect 9772 29932 9828 29934
rect 10092 29986 10148 29988
rect 10092 29934 10094 29986
rect 10094 29934 10146 29986
rect 10146 29934 10148 29986
rect 10092 29932 10148 29934
rect 10412 29986 10468 29988
rect 10412 29934 10414 29986
rect 10414 29934 10466 29986
rect 10466 29934 10468 29986
rect 10412 29932 10468 29934
rect 10732 29986 10788 29988
rect 10732 29934 10734 29986
rect 10734 29934 10786 29986
rect 10786 29934 10788 29986
rect 10732 29932 10788 29934
rect 11052 29986 11108 29988
rect 11052 29934 11054 29986
rect 11054 29934 11106 29986
rect 11106 29934 11108 29986
rect 11052 29932 11108 29934
rect 11372 29986 11428 29988
rect 11372 29934 11374 29986
rect 11374 29934 11426 29986
rect 11426 29934 11428 29986
rect 11372 29932 11428 29934
rect 11532 29986 11588 29988
rect 11532 29934 11534 29986
rect 11534 29934 11586 29986
rect 11586 29934 11588 29986
rect 11532 29932 11588 29934
rect 11852 29986 11908 29988
rect 11852 29934 11854 29986
rect 11854 29934 11906 29986
rect 11906 29934 11908 29986
rect 11852 29932 11908 29934
rect 12012 29986 12068 29988
rect 12012 29934 12014 29986
rect 12014 29934 12066 29986
rect 12066 29934 12068 29986
rect 12012 29932 12068 29934
rect 12332 29986 12388 29988
rect 12332 29934 12334 29986
rect 12334 29934 12386 29986
rect 12386 29934 12388 29986
rect 12332 29932 12388 29934
rect 8492 29826 8548 29828
rect 8492 29774 8494 29826
rect 8494 29774 8546 29826
rect 8546 29774 8548 29826
rect 8492 29772 8548 29774
rect 8812 29826 8868 29828
rect 8812 29774 8814 29826
rect 8814 29774 8866 29826
rect 8866 29774 8868 29826
rect 8812 29772 8868 29774
rect 8972 29826 9028 29828
rect 8972 29774 8974 29826
rect 8974 29774 9026 29826
rect 9026 29774 9028 29826
rect 8972 29772 9028 29774
rect 9292 29826 9348 29828
rect 9292 29774 9294 29826
rect 9294 29774 9346 29826
rect 9346 29774 9348 29826
rect 9292 29772 9348 29774
rect 9452 29826 9508 29828
rect 9452 29774 9454 29826
rect 9454 29774 9506 29826
rect 9506 29774 9508 29826
rect 9452 29772 9508 29774
rect 9772 29826 9828 29828
rect 9772 29774 9774 29826
rect 9774 29774 9826 29826
rect 9826 29774 9828 29826
rect 9772 29772 9828 29774
rect 10092 29826 10148 29828
rect 10092 29774 10094 29826
rect 10094 29774 10146 29826
rect 10146 29774 10148 29826
rect 10092 29772 10148 29774
rect 10412 29826 10468 29828
rect 10412 29774 10414 29826
rect 10414 29774 10466 29826
rect 10466 29774 10468 29826
rect 10412 29772 10468 29774
rect 10732 29826 10788 29828
rect 10732 29774 10734 29826
rect 10734 29774 10786 29826
rect 10786 29774 10788 29826
rect 10732 29772 10788 29774
rect 11052 29826 11108 29828
rect 11052 29774 11054 29826
rect 11054 29774 11106 29826
rect 11106 29774 11108 29826
rect 11052 29772 11108 29774
rect 11372 29826 11428 29828
rect 11372 29774 11374 29826
rect 11374 29774 11426 29826
rect 11426 29774 11428 29826
rect 11372 29772 11428 29774
rect 11532 29826 11588 29828
rect 11532 29774 11534 29826
rect 11534 29774 11586 29826
rect 11586 29774 11588 29826
rect 11532 29772 11588 29774
rect 11852 29826 11908 29828
rect 11852 29774 11854 29826
rect 11854 29774 11906 29826
rect 11906 29774 11908 29826
rect 11852 29772 11908 29774
rect 12012 29826 12068 29828
rect 12012 29774 12014 29826
rect 12014 29774 12066 29826
rect 12066 29774 12068 29826
rect 12012 29772 12068 29774
rect 12332 29826 12388 29828
rect 12332 29774 12334 29826
rect 12334 29774 12386 29826
rect 12386 29774 12388 29826
rect 12332 29772 12388 29774
rect 8492 29666 8548 29668
rect 8492 29614 8494 29666
rect 8494 29614 8546 29666
rect 8546 29614 8548 29666
rect 8492 29612 8548 29614
rect 8812 29666 8868 29668
rect 8812 29614 8814 29666
rect 8814 29614 8866 29666
rect 8866 29614 8868 29666
rect 8812 29612 8868 29614
rect 8972 29666 9028 29668
rect 8972 29614 8974 29666
rect 8974 29614 9026 29666
rect 9026 29614 9028 29666
rect 8972 29612 9028 29614
rect 9292 29666 9348 29668
rect 9292 29614 9294 29666
rect 9294 29614 9346 29666
rect 9346 29614 9348 29666
rect 9292 29612 9348 29614
rect 9452 29666 9508 29668
rect 9452 29614 9454 29666
rect 9454 29614 9506 29666
rect 9506 29614 9508 29666
rect 9452 29612 9508 29614
rect 9772 29666 9828 29668
rect 9772 29614 9774 29666
rect 9774 29614 9826 29666
rect 9826 29614 9828 29666
rect 9772 29612 9828 29614
rect 10092 29666 10148 29668
rect 10092 29614 10094 29666
rect 10094 29614 10146 29666
rect 10146 29614 10148 29666
rect 10092 29612 10148 29614
rect 10412 29666 10468 29668
rect 10412 29614 10414 29666
rect 10414 29614 10466 29666
rect 10466 29614 10468 29666
rect 10412 29612 10468 29614
rect 10732 29666 10788 29668
rect 10732 29614 10734 29666
rect 10734 29614 10786 29666
rect 10786 29614 10788 29666
rect 10732 29612 10788 29614
rect 11052 29666 11108 29668
rect 11052 29614 11054 29666
rect 11054 29614 11106 29666
rect 11106 29614 11108 29666
rect 11052 29612 11108 29614
rect 11372 29666 11428 29668
rect 11372 29614 11374 29666
rect 11374 29614 11426 29666
rect 11426 29614 11428 29666
rect 11372 29612 11428 29614
rect 11532 29666 11588 29668
rect 11532 29614 11534 29666
rect 11534 29614 11586 29666
rect 11586 29614 11588 29666
rect 11532 29612 11588 29614
rect 11852 29666 11908 29668
rect 11852 29614 11854 29666
rect 11854 29614 11906 29666
rect 11906 29614 11908 29666
rect 11852 29612 11908 29614
rect 12012 29666 12068 29668
rect 12012 29614 12014 29666
rect 12014 29614 12066 29666
rect 12066 29614 12068 29666
rect 12012 29612 12068 29614
rect 12332 29666 12388 29668
rect 12332 29614 12334 29666
rect 12334 29614 12386 29666
rect 12386 29614 12388 29666
rect 12332 29612 12388 29614
rect 8492 29506 8548 29508
rect 8492 29454 8494 29506
rect 8494 29454 8546 29506
rect 8546 29454 8548 29506
rect 8492 29452 8548 29454
rect 8812 29506 8868 29508
rect 8812 29454 8814 29506
rect 8814 29454 8866 29506
rect 8866 29454 8868 29506
rect 8812 29452 8868 29454
rect 8972 29506 9028 29508
rect 8972 29454 8974 29506
rect 8974 29454 9026 29506
rect 9026 29454 9028 29506
rect 8972 29452 9028 29454
rect 9292 29506 9348 29508
rect 9292 29454 9294 29506
rect 9294 29454 9346 29506
rect 9346 29454 9348 29506
rect 9292 29452 9348 29454
rect 9452 29506 9508 29508
rect 9452 29454 9454 29506
rect 9454 29454 9506 29506
rect 9506 29454 9508 29506
rect 9452 29452 9508 29454
rect 9772 29506 9828 29508
rect 9772 29454 9774 29506
rect 9774 29454 9826 29506
rect 9826 29454 9828 29506
rect 9772 29452 9828 29454
rect 10092 29506 10148 29508
rect 10092 29454 10094 29506
rect 10094 29454 10146 29506
rect 10146 29454 10148 29506
rect 10092 29452 10148 29454
rect 10412 29506 10468 29508
rect 10412 29454 10414 29506
rect 10414 29454 10466 29506
rect 10466 29454 10468 29506
rect 10412 29452 10468 29454
rect 10732 29506 10788 29508
rect 10732 29454 10734 29506
rect 10734 29454 10786 29506
rect 10786 29454 10788 29506
rect 10732 29452 10788 29454
rect 11052 29506 11108 29508
rect 11052 29454 11054 29506
rect 11054 29454 11106 29506
rect 11106 29454 11108 29506
rect 11052 29452 11108 29454
rect 11372 29506 11428 29508
rect 11372 29454 11374 29506
rect 11374 29454 11426 29506
rect 11426 29454 11428 29506
rect 11372 29452 11428 29454
rect 11532 29506 11588 29508
rect 11532 29454 11534 29506
rect 11534 29454 11586 29506
rect 11586 29454 11588 29506
rect 11532 29452 11588 29454
rect 11852 29506 11908 29508
rect 11852 29454 11854 29506
rect 11854 29454 11906 29506
rect 11906 29454 11908 29506
rect 11852 29452 11908 29454
rect 12012 29506 12068 29508
rect 12012 29454 12014 29506
rect 12014 29454 12066 29506
rect 12066 29454 12068 29506
rect 12012 29452 12068 29454
rect 12332 29506 12388 29508
rect 12332 29454 12334 29506
rect 12334 29454 12386 29506
rect 12386 29454 12388 29506
rect 12332 29452 12388 29454
rect 8492 29346 8548 29348
rect 8492 29294 8494 29346
rect 8494 29294 8546 29346
rect 8546 29294 8548 29346
rect 8492 29292 8548 29294
rect 8812 29346 8868 29348
rect 8812 29294 8814 29346
rect 8814 29294 8866 29346
rect 8866 29294 8868 29346
rect 8812 29292 8868 29294
rect 8972 29346 9028 29348
rect 8972 29294 8974 29346
rect 8974 29294 9026 29346
rect 9026 29294 9028 29346
rect 8972 29292 9028 29294
rect 9292 29346 9348 29348
rect 9292 29294 9294 29346
rect 9294 29294 9346 29346
rect 9346 29294 9348 29346
rect 9292 29292 9348 29294
rect 9452 29346 9508 29348
rect 9452 29294 9454 29346
rect 9454 29294 9506 29346
rect 9506 29294 9508 29346
rect 9452 29292 9508 29294
rect 9772 29346 9828 29348
rect 9772 29294 9774 29346
rect 9774 29294 9826 29346
rect 9826 29294 9828 29346
rect 9772 29292 9828 29294
rect 10092 29346 10148 29348
rect 10092 29294 10094 29346
rect 10094 29294 10146 29346
rect 10146 29294 10148 29346
rect 10092 29292 10148 29294
rect 10412 29346 10468 29348
rect 10412 29294 10414 29346
rect 10414 29294 10466 29346
rect 10466 29294 10468 29346
rect 10412 29292 10468 29294
rect 10732 29346 10788 29348
rect 10732 29294 10734 29346
rect 10734 29294 10786 29346
rect 10786 29294 10788 29346
rect 10732 29292 10788 29294
rect 11052 29346 11108 29348
rect 11052 29294 11054 29346
rect 11054 29294 11106 29346
rect 11106 29294 11108 29346
rect 11052 29292 11108 29294
rect 11372 29346 11428 29348
rect 11372 29294 11374 29346
rect 11374 29294 11426 29346
rect 11426 29294 11428 29346
rect 11372 29292 11428 29294
rect 11532 29346 11588 29348
rect 11532 29294 11534 29346
rect 11534 29294 11586 29346
rect 11586 29294 11588 29346
rect 11532 29292 11588 29294
rect 11852 29346 11908 29348
rect 11852 29294 11854 29346
rect 11854 29294 11906 29346
rect 11906 29294 11908 29346
rect 11852 29292 11908 29294
rect 12012 29346 12068 29348
rect 12012 29294 12014 29346
rect 12014 29294 12066 29346
rect 12066 29294 12068 29346
rect 12012 29292 12068 29294
rect 12332 29346 12388 29348
rect 12332 29294 12334 29346
rect 12334 29294 12386 29346
rect 12386 29294 12388 29346
rect 12332 29292 12388 29294
rect 8492 29186 8548 29188
rect 8492 29134 8494 29186
rect 8494 29134 8546 29186
rect 8546 29134 8548 29186
rect 8492 29132 8548 29134
rect 8812 29186 8868 29188
rect 8812 29134 8814 29186
rect 8814 29134 8866 29186
rect 8866 29134 8868 29186
rect 8812 29132 8868 29134
rect 8972 29186 9028 29188
rect 8972 29134 8974 29186
rect 8974 29134 9026 29186
rect 9026 29134 9028 29186
rect 8972 29132 9028 29134
rect 9292 29186 9348 29188
rect 9292 29134 9294 29186
rect 9294 29134 9346 29186
rect 9346 29134 9348 29186
rect 9292 29132 9348 29134
rect 9452 29186 9508 29188
rect 9452 29134 9454 29186
rect 9454 29134 9506 29186
rect 9506 29134 9508 29186
rect 9452 29132 9508 29134
rect 9772 29186 9828 29188
rect 9772 29134 9774 29186
rect 9774 29134 9826 29186
rect 9826 29134 9828 29186
rect 9772 29132 9828 29134
rect 10092 29186 10148 29188
rect 10092 29134 10094 29186
rect 10094 29134 10146 29186
rect 10146 29134 10148 29186
rect 10092 29132 10148 29134
rect 10412 29186 10468 29188
rect 10412 29134 10414 29186
rect 10414 29134 10466 29186
rect 10466 29134 10468 29186
rect 10412 29132 10468 29134
rect 10732 29186 10788 29188
rect 10732 29134 10734 29186
rect 10734 29134 10786 29186
rect 10786 29134 10788 29186
rect 10732 29132 10788 29134
rect 11052 29186 11108 29188
rect 11052 29134 11054 29186
rect 11054 29134 11106 29186
rect 11106 29134 11108 29186
rect 11052 29132 11108 29134
rect 11372 29186 11428 29188
rect 11372 29134 11374 29186
rect 11374 29134 11426 29186
rect 11426 29134 11428 29186
rect 11372 29132 11428 29134
rect 11532 29186 11588 29188
rect 11532 29134 11534 29186
rect 11534 29134 11586 29186
rect 11586 29134 11588 29186
rect 11532 29132 11588 29134
rect 11852 29186 11908 29188
rect 11852 29134 11854 29186
rect 11854 29134 11906 29186
rect 11906 29134 11908 29186
rect 11852 29132 11908 29134
rect 12012 29186 12068 29188
rect 12012 29134 12014 29186
rect 12014 29134 12066 29186
rect 12066 29134 12068 29186
rect 12012 29132 12068 29134
rect 12332 29186 12388 29188
rect 12332 29134 12334 29186
rect 12334 29134 12386 29186
rect 12386 29134 12388 29186
rect 12332 29132 12388 29134
rect 8492 29026 8548 29028
rect 8492 28974 8494 29026
rect 8494 28974 8546 29026
rect 8546 28974 8548 29026
rect 8492 28972 8548 28974
rect 8812 29026 8868 29028
rect 8812 28974 8814 29026
rect 8814 28974 8866 29026
rect 8866 28974 8868 29026
rect 8812 28972 8868 28974
rect 8972 29026 9028 29028
rect 8972 28974 8974 29026
rect 8974 28974 9026 29026
rect 9026 28974 9028 29026
rect 8972 28972 9028 28974
rect 9292 29026 9348 29028
rect 9292 28974 9294 29026
rect 9294 28974 9346 29026
rect 9346 28974 9348 29026
rect 9292 28972 9348 28974
rect 9452 29026 9508 29028
rect 9452 28974 9454 29026
rect 9454 28974 9506 29026
rect 9506 28974 9508 29026
rect 9452 28972 9508 28974
rect 9772 29026 9828 29028
rect 9772 28974 9774 29026
rect 9774 28974 9826 29026
rect 9826 28974 9828 29026
rect 9772 28972 9828 28974
rect 10092 29026 10148 29028
rect 10092 28974 10094 29026
rect 10094 28974 10146 29026
rect 10146 28974 10148 29026
rect 10092 28972 10148 28974
rect 10412 29026 10468 29028
rect 10412 28974 10414 29026
rect 10414 28974 10466 29026
rect 10466 28974 10468 29026
rect 10412 28972 10468 28974
rect 10732 29026 10788 29028
rect 10732 28974 10734 29026
rect 10734 28974 10786 29026
rect 10786 28974 10788 29026
rect 10732 28972 10788 28974
rect 11052 29026 11108 29028
rect 11052 28974 11054 29026
rect 11054 28974 11106 29026
rect 11106 28974 11108 29026
rect 11052 28972 11108 28974
rect 11372 29026 11428 29028
rect 11372 28974 11374 29026
rect 11374 28974 11426 29026
rect 11426 28974 11428 29026
rect 11372 28972 11428 28974
rect 11532 29026 11588 29028
rect 11532 28974 11534 29026
rect 11534 28974 11586 29026
rect 11586 28974 11588 29026
rect 11532 28972 11588 28974
rect 11852 29026 11908 29028
rect 11852 28974 11854 29026
rect 11854 28974 11906 29026
rect 11906 28974 11908 29026
rect 11852 28972 11908 28974
rect 12012 29026 12068 29028
rect 12012 28974 12014 29026
rect 12014 28974 12066 29026
rect 12066 28974 12068 29026
rect 12012 28972 12068 28974
rect 12332 29026 12388 29028
rect 12332 28974 12334 29026
rect 12334 28974 12386 29026
rect 12386 28974 12388 29026
rect 12332 28972 12388 28974
rect 8492 28866 8548 28868
rect 8492 28814 8494 28866
rect 8494 28814 8546 28866
rect 8546 28814 8548 28866
rect 8492 28812 8548 28814
rect 8812 28866 8868 28868
rect 8812 28814 8814 28866
rect 8814 28814 8866 28866
rect 8866 28814 8868 28866
rect 8812 28812 8868 28814
rect 8972 28866 9028 28868
rect 8972 28814 8974 28866
rect 8974 28814 9026 28866
rect 9026 28814 9028 28866
rect 8972 28812 9028 28814
rect 9292 28866 9348 28868
rect 9292 28814 9294 28866
rect 9294 28814 9346 28866
rect 9346 28814 9348 28866
rect 9292 28812 9348 28814
rect 9452 28866 9508 28868
rect 9452 28814 9454 28866
rect 9454 28814 9506 28866
rect 9506 28814 9508 28866
rect 9452 28812 9508 28814
rect 9772 28866 9828 28868
rect 9772 28814 9774 28866
rect 9774 28814 9826 28866
rect 9826 28814 9828 28866
rect 9772 28812 9828 28814
rect 10092 28866 10148 28868
rect 10092 28814 10094 28866
rect 10094 28814 10146 28866
rect 10146 28814 10148 28866
rect 10092 28812 10148 28814
rect 10412 28866 10468 28868
rect 10412 28814 10414 28866
rect 10414 28814 10466 28866
rect 10466 28814 10468 28866
rect 10412 28812 10468 28814
rect 10732 28866 10788 28868
rect 10732 28814 10734 28866
rect 10734 28814 10786 28866
rect 10786 28814 10788 28866
rect 10732 28812 10788 28814
rect 11052 28866 11108 28868
rect 11052 28814 11054 28866
rect 11054 28814 11106 28866
rect 11106 28814 11108 28866
rect 11052 28812 11108 28814
rect 11372 28866 11428 28868
rect 11372 28814 11374 28866
rect 11374 28814 11426 28866
rect 11426 28814 11428 28866
rect 11372 28812 11428 28814
rect 11532 28866 11588 28868
rect 11532 28814 11534 28866
rect 11534 28814 11586 28866
rect 11586 28814 11588 28866
rect 11532 28812 11588 28814
rect 11852 28866 11908 28868
rect 11852 28814 11854 28866
rect 11854 28814 11906 28866
rect 11906 28814 11908 28866
rect 11852 28812 11908 28814
rect 12012 28866 12068 28868
rect 12012 28814 12014 28866
rect 12014 28814 12066 28866
rect 12066 28814 12068 28866
rect 12012 28812 12068 28814
rect 12332 28866 12388 28868
rect 12332 28814 12334 28866
rect 12334 28814 12386 28866
rect 12386 28814 12388 28866
rect 12332 28812 12388 28814
rect 10572 28572 10628 28628
rect 9932 28252 9988 28308
rect 10892 28252 10948 28308
rect 8492 28066 8548 28068
rect 8492 28014 8494 28066
rect 8494 28014 8546 28066
rect 8546 28014 8548 28066
rect 8492 28012 8548 28014
rect 8812 28066 8868 28068
rect 8812 28014 8814 28066
rect 8814 28014 8866 28066
rect 8866 28014 8868 28066
rect 8812 28012 8868 28014
rect 8972 28066 9028 28068
rect 8972 28014 8974 28066
rect 8974 28014 9026 28066
rect 9026 28014 9028 28066
rect 8972 28012 9028 28014
rect 9292 28066 9348 28068
rect 9292 28014 9294 28066
rect 9294 28014 9346 28066
rect 9346 28014 9348 28066
rect 9292 28012 9348 28014
rect 9452 28066 9508 28068
rect 9452 28014 9454 28066
rect 9454 28014 9506 28066
rect 9506 28014 9508 28066
rect 9452 28012 9508 28014
rect 9772 28066 9828 28068
rect 9772 28014 9774 28066
rect 9774 28014 9826 28066
rect 9826 28014 9828 28066
rect 9772 28012 9828 28014
rect 10092 28066 10148 28068
rect 10092 28014 10094 28066
rect 10094 28014 10146 28066
rect 10146 28014 10148 28066
rect 10092 28012 10148 28014
rect 10412 28066 10468 28068
rect 10412 28014 10414 28066
rect 10414 28014 10466 28066
rect 10466 28014 10468 28066
rect 10412 28012 10468 28014
rect 10732 28066 10788 28068
rect 10732 28014 10734 28066
rect 10734 28014 10786 28066
rect 10786 28014 10788 28066
rect 10732 28012 10788 28014
rect 11052 28066 11108 28068
rect 11052 28014 11054 28066
rect 11054 28014 11106 28066
rect 11106 28014 11108 28066
rect 11052 28012 11108 28014
rect 11372 28066 11428 28068
rect 11372 28014 11374 28066
rect 11374 28014 11426 28066
rect 11426 28014 11428 28066
rect 11372 28012 11428 28014
rect 11532 28066 11588 28068
rect 11532 28014 11534 28066
rect 11534 28014 11586 28066
rect 11586 28014 11588 28066
rect 11532 28012 11588 28014
rect 11852 28066 11908 28068
rect 11852 28014 11854 28066
rect 11854 28014 11906 28066
rect 11906 28014 11908 28066
rect 11852 28012 11908 28014
rect 12012 28066 12068 28068
rect 12012 28014 12014 28066
rect 12014 28014 12066 28066
rect 12066 28014 12068 28066
rect 12012 28012 12068 28014
rect 12332 28066 12388 28068
rect 12332 28014 12334 28066
rect 12334 28014 12386 28066
rect 12386 28014 12388 28066
rect 12332 28012 12388 28014
rect 8492 27906 8548 27908
rect 8492 27854 8494 27906
rect 8494 27854 8546 27906
rect 8546 27854 8548 27906
rect 8492 27852 8548 27854
rect 8812 27906 8868 27908
rect 8812 27854 8814 27906
rect 8814 27854 8866 27906
rect 8866 27854 8868 27906
rect 8812 27852 8868 27854
rect 8972 27906 9028 27908
rect 8972 27854 8974 27906
rect 8974 27854 9026 27906
rect 9026 27854 9028 27906
rect 8972 27852 9028 27854
rect 9292 27906 9348 27908
rect 9292 27854 9294 27906
rect 9294 27854 9346 27906
rect 9346 27854 9348 27906
rect 9292 27852 9348 27854
rect 9452 27906 9508 27908
rect 9452 27854 9454 27906
rect 9454 27854 9506 27906
rect 9506 27854 9508 27906
rect 9452 27852 9508 27854
rect 9772 27906 9828 27908
rect 9772 27854 9774 27906
rect 9774 27854 9826 27906
rect 9826 27854 9828 27906
rect 9772 27852 9828 27854
rect 10092 27906 10148 27908
rect 10092 27854 10094 27906
rect 10094 27854 10146 27906
rect 10146 27854 10148 27906
rect 10092 27852 10148 27854
rect 10412 27906 10468 27908
rect 10412 27854 10414 27906
rect 10414 27854 10466 27906
rect 10466 27854 10468 27906
rect 10412 27852 10468 27854
rect 10732 27906 10788 27908
rect 10732 27854 10734 27906
rect 10734 27854 10786 27906
rect 10786 27854 10788 27906
rect 10732 27852 10788 27854
rect 11052 27906 11108 27908
rect 11052 27854 11054 27906
rect 11054 27854 11106 27906
rect 11106 27854 11108 27906
rect 11052 27852 11108 27854
rect 11372 27906 11428 27908
rect 11372 27854 11374 27906
rect 11374 27854 11426 27906
rect 11426 27854 11428 27906
rect 11372 27852 11428 27854
rect 11532 27906 11588 27908
rect 11532 27854 11534 27906
rect 11534 27854 11586 27906
rect 11586 27854 11588 27906
rect 11532 27852 11588 27854
rect 11852 27906 11908 27908
rect 11852 27854 11854 27906
rect 11854 27854 11906 27906
rect 11906 27854 11908 27906
rect 11852 27852 11908 27854
rect 12012 27906 12068 27908
rect 12012 27854 12014 27906
rect 12014 27854 12066 27906
rect 12066 27854 12068 27906
rect 12012 27852 12068 27854
rect 12332 27906 12388 27908
rect 12332 27854 12334 27906
rect 12334 27854 12386 27906
rect 12386 27854 12388 27906
rect 12332 27852 12388 27854
rect 8492 27746 8548 27748
rect 8492 27694 8494 27746
rect 8494 27694 8546 27746
rect 8546 27694 8548 27746
rect 8492 27692 8548 27694
rect 8812 27746 8868 27748
rect 8812 27694 8814 27746
rect 8814 27694 8866 27746
rect 8866 27694 8868 27746
rect 8812 27692 8868 27694
rect 8972 27746 9028 27748
rect 8972 27694 8974 27746
rect 8974 27694 9026 27746
rect 9026 27694 9028 27746
rect 8972 27692 9028 27694
rect 9292 27746 9348 27748
rect 9292 27694 9294 27746
rect 9294 27694 9346 27746
rect 9346 27694 9348 27746
rect 9292 27692 9348 27694
rect 9452 27746 9508 27748
rect 9452 27694 9454 27746
rect 9454 27694 9506 27746
rect 9506 27694 9508 27746
rect 9452 27692 9508 27694
rect 9772 27746 9828 27748
rect 9772 27694 9774 27746
rect 9774 27694 9826 27746
rect 9826 27694 9828 27746
rect 9772 27692 9828 27694
rect 10092 27746 10148 27748
rect 10092 27694 10094 27746
rect 10094 27694 10146 27746
rect 10146 27694 10148 27746
rect 10092 27692 10148 27694
rect 10412 27746 10468 27748
rect 10412 27694 10414 27746
rect 10414 27694 10466 27746
rect 10466 27694 10468 27746
rect 10412 27692 10468 27694
rect 10732 27746 10788 27748
rect 10732 27694 10734 27746
rect 10734 27694 10786 27746
rect 10786 27694 10788 27746
rect 10732 27692 10788 27694
rect 11052 27746 11108 27748
rect 11052 27694 11054 27746
rect 11054 27694 11106 27746
rect 11106 27694 11108 27746
rect 11052 27692 11108 27694
rect 11372 27746 11428 27748
rect 11372 27694 11374 27746
rect 11374 27694 11426 27746
rect 11426 27694 11428 27746
rect 11372 27692 11428 27694
rect 11532 27746 11588 27748
rect 11532 27694 11534 27746
rect 11534 27694 11586 27746
rect 11586 27694 11588 27746
rect 11532 27692 11588 27694
rect 11852 27746 11908 27748
rect 11852 27694 11854 27746
rect 11854 27694 11906 27746
rect 11906 27694 11908 27746
rect 11852 27692 11908 27694
rect 12012 27746 12068 27748
rect 12012 27694 12014 27746
rect 12014 27694 12066 27746
rect 12066 27694 12068 27746
rect 12012 27692 12068 27694
rect 12332 27746 12388 27748
rect 12332 27694 12334 27746
rect 12334 27694 12386 27746
rect 12386 27694 12388 27746
rect 12332 27692 12388 27694
rect 8492 27586 8548 27588
rect 8492 27534 8494 27586
rect 8494 27534 8546 27586
rect 8546 27534 8548 27586
rect 8492 27532 8548 27534
rect 8812 27586 8868 27588
rect 8812 27534 8814 27586
rect 8814 27534 8866 27586
rect 8866 27534 8868 27586
rect 8812 27532 8868 27534
rect 8972 27586 9028 27588
rect 8972 27534 8974 27586
rect 8974 27534 9026 27586
rect 9026 27534 9028 27586
rect 8972 27532 9028 27534
rect 9292 27586 9348 27588
rect 9292 27534 9294 27586
rect 9294 27534 9346 27586
rect 9346 27534 9348 27586
rect 9292 27532 9348 27534
rect 9452 27586 9508 27588
rect 9452 27534 9454 27586
rect 9454 27534 9506 27586
rect 9506 27534 9508 27586
rect 9452 27532 9508 27534
rect 9772 27586 9828 27588
rect 9772 27534 9774 27586
rect 9774 27534 9826 27586
rect 9826 27534 9828 27586
rect 9772 27532 9828 27534
rect 10092 27586 10148 27588
rect 10092 27534 10094 27586
rect 10094 27534 10146 27586
rect 10146 27534 10148 27586
rect 10092 27532 10148 27534
rect 10412 27586 10468 27588
rect 10412 27534 10414 27586
rect 10414 27534 10466 27586
rect 10466 27534 10468 27586
rect 10412 27532 10468 27534
rect 10732 27586 10788 27588
rect 10732 27534 10734 27586
rect 10734 27534 10786 27586
rect 10786 27534 10788 27586
rect 10732 27532 10788 27534
rect 11052 27586 11108 27588
rect 11052 27534 11054 27586
rect 11054 27534 11106 27586
rect 11106 27534 11108 27586
rect 11052 27532 11108 27534
rect 11372 27586 11428 27588
rect 11372 27534 11374 27586
rect 11374 27534 11426 27586
rect 11426 27534 11428 27586
rect 11372 27532 11428 27534
rect 11532 27586 11588 27588
rect 11532 27534 11534 27586
rect 11534 27534 11586 27586
rect 11586 27534 11588 27586
rect 11532 27532 11588 27534
rect 11852 27586 11908 27588
rect 11852 27534 11854 27586
rect 11854 27534 11906 27586
rect 11906 27534 11908 27586
rect 11852 27532 11908 27534
rect 12012 27586 12068 27588
rect 12012 27534 12014 27586
rect 12014 27534 12066 27586
rect 12066 27534 12068 27586
rect 12012 27532 12068 27534
rect 12332 27586 12388 27588
rect 12332 27534 12334 27586
rect 12334 27534 12386 27586
rect 12386 27534 12388 27586
rect 12332 27532 12388 27534
rect 8492 27426 8548 27428
rect 8492 27374 8494 27426
rect 8494 27374 8546 27426
rect 8546 27374 8548 27426
rect 8492 27372 8548 27374
rect 8812 27426 8868 27428
rect 8812 27374 8814 27426
rect 8814 27374 8866 27426
rect 8866 27374 8868 27426
rect 8812 27372 8868 27374
rect 8972 27426 9028 27428
rect 8972 27374 8974 27426
rect 8974 27374 9026 27426
rect 9026 27374 9028 27426
rect 8972 27372 9028 27374
rect 9292 27426 9348 27428
rect 9292 27374 9294 27426
rect 9294 27374 9346 27426
rect 9346 27374 9348 27426
rect 9292 27372 9348 27374
rect 9452 27426 9508 27428
rect 9452 27374 9454 27426
rect 9454 27374 9506 27426
rect 9506 27374 9508 27426
rect 9452 27372 9508 27374
rect 9772 27426 9828 27428
rect 9772 27374 9774 27426
rect 9774 27374 9826 27426
rect 9826 27374 9828 27426
rect 9772 27372 9828 27374
rect 10092 27426 10148 27428
rect 10092 27374 10094 27426
rect 10094 27374 10146 27426
rect 10146 27374 10148 27426
rect 10092 27372 10148 27374
rect 10412 27426 10468 27428
rect 10412 27374 10414 27426
rect 10414 27374 10466 27426
rect 10466 27374 10468 27426
rect 10412 27372 10468 27374
rect 10732 27426 10788 27428
rect 10732 27374 10734 27426
rect 10734 27374 10786 27426
rect 10786 27374 10788 27426
rect 10732 27372 10788 27374
rect 11052 27426 11108 27428
rect 11052 27374 11054 27426
rect 11054 27374 11106 27426
rect 11106 27374 11108 27426
rect 11052 27372 11108 27374
rect 11372 27426 11428 27428
rect 11372 27374 11374 27426
rect 11374 27374 11426 27426
rect 11426 27374 11428 27426
rect 11372 27372 11428 27374
rect 11532 27426 11588 27428
rect 11532 27374 11534 27426
rect 11534 27374 11586 27426
rect 11586 27374 11588 27426
rect 11532 27372 11588 27374
rect 11852 27426 11908 27428
rect 11852 27374 11854 27426
rect 11854 27374 11906 27426
rect 11906 27374 11908 27426
rect 11852 27372 11908 27374
rect 12012 27426 12068 27428
rect 12012 27374 12014 27426
rect 12014 27374 12066 27426
rect 12066 27374 12068 27426
rect 12012 27372 12068 27374
rect 12332 27426 12388 27428
rect 12332 27374 12334 27426
rect 12334 27374 12386 27426
rect 12386 27374 12388 27426
rect 12332 27372 12388 27374
rect 8492 27266 8548 27268
rect 8492 27214 8494 27266
rect 8494 27214 8546 27266
rect 8546 27214 8548 27266
rect 8492 27212 8548 27214
rect 8812 27266 8868 27268
rect 8812 27214 8814 27266
rect 8814 27214 8866 27266
rect 8866 27214 8868 27266
rect 8812 27212 8868 27214
rect 8972 27266 9028 27268
rect 8972 27214 8974 27266
rect 8974 27214 9026 27266
rect 9026 27214 9028 27266
rect 8972 27212 9028 27214
rect 9292 27266 9348 27268
rect 9292 27214 9294 27266
rect 9294 27214 9346 27266
rect 9346 27214 9348 27266
rect 9292 27212 9348 27214
rect 9452 27266 9508 27268
rect 9452 27214 9454 27266
rect 9454 27214 9506 27266
rect 9506 27214 9508 27266
rect 9452 27212 9508 27214
rect 9772 27266 9828 27268
rect 9772 27214 9774 27266
rect 9774 27214 9826 27266
rect 9826 27214 9828 27266
rect 9772 27212 9828 27214
rect 10092 27266 10148 27268
rect 10092 27214 10094 27266
rect 10094 27214 10146 27266
rect 10146 27214 10148 27266
rect 10092 27212 10148 27214
rect 10412 27266 10468 27268
rect 10412 27214 10414 27266
rect 10414 27214 10466 27266
rect 10466 27214 10468 27266
rect 10412 27212 10468 27214
rect 10732 27266 10788 27268
rect 10732 27214 10734 27266
rect 10734 27214 10786 27266
rect 10786 27214 10788 27266
rect 10732 27212 10788 27214
rect 11052 27266 11108 27268
rect 11052 27214 11054 27266
rect 11054 27214 11106 27266
rect 11106 27214 11108 27266
rect 11052 27212 11108 27214
rect 11372 27266 11428 27268
rect 11372 27214 11374 27266
rect 11374 27214 11426 27266
rect 11426 27214 11428 27266
rect 11372 27212 11428 27214
rect 11532 27266 11588 27268
rect 11532 27214 11534 27266
rect 11534 27214 11586 27266
rect 11586 27214 11588 27266
rect 11532 27212 11588 27214
rect 11852 27266 11908 27268
rect 11852 27214 11854 27266
rect 11854 27214 11906 27266
rect 11906 27214 11908 27266
rect 11852 27212 11908 27214
rect 12012 27266 12068 27268
rect 12012 27214 12014 27266
rect 12014 27214 12066 27266
rect 12066 27214 12068 27266
rect 12012 27212 12068 27214
rect 12332 27266 12388 27268
rect 12332 27214 12334 27266
rect 12334 27214 12386 27266
rect 12386 27214 12388 27266
rect 12332 27212 12388 27214
rect 8492 27106 8548 27108
rect 8492 27054 8494 27106
rect 8494 27054 8546 27106
rect 8546 27054 8548 27106
rect 8492 27052 8548 27054
rect 8812 27106 8868 27108
rect 8812 27054 8814 27106
rect 8814 27054 8866 27106
rect 8866 27054 8868 27106
rect 8812 27052 8868 27054
rect 8972 27106 9028 27108
rect 8972 27054 8974 27106
rect 8974 27054 9026 27106
rect 9026 27054 9028 27106
rect 8972 27052 9028 27054
rect 9292 27106 9348 27108
rect 9292 27054 9294 27106
rect 9294 27054 9346 27106
rect 9346 27054 9348 27106
rect 9292 27052 9348 27054
rect 9452 27106 9508 27108
rect 9452 27054 9454 27106
rect 9454 27054 9506 27106
rect 9506 27054 9508 27106
rect 9452 27052 9508 27054
rect 9772 27106 9828 27108
rect 9772 27054 9774 27106
rect 9774 27054 9826 27106
rect 9826 27054 9828 27106
rect 9772 27052 9828 27054
rect 10092 27106 10148 27108
rect 10092 27054 10094 27106
rect 10094 27054 10146 27106
rect 10146 27054 10148 27106
rect 10092 27052 10148 27054
rect 10412 27106 10468 27108
rect 10412 27054 10414 27106
rect 10414 27054 10466 27106
rect 10466 27054 10468 27106
rect 10412 27052 10468 27054
rect 10732 27106 10788 27108
rect 10732 27054 10734 27106
rect 10734 27054 10786 27106
rect 10786 27054 10788 27106
rect 10732 27052 10788 27054
rect 11052 27106 11108 27108
rect 11052 27054 11054 27106
rect 11054 27054 11106 27106
rect 11106 27054 11108 27106
rect 11052 27052 11108 27054
rect 11372 27106 11428 27108
rect 11372 27054 11374 27106
rect 11374 27054 11426 27106
rect 11426 27054 11428 27106
rect 11372 27052 11428 27054
rect 11532 27106 11588 27108
rect 11532 27054 11534 27106
rect 11534 27054 11586 27106
rect 11586 27054 11588 27106
rect 11532 27052 11588 27054
rect 11852 27106 11908 27108
rect 11852 27054 11854 27106
rect 11854 27054 11906 27106
rect 11906 27054 11908 27106
rect 11852 27052 11908 27054
rect 12012 27106 12068 27108
rect 12012 27054 12014 27106
rect 12014 27054 12066 27106
rect 12066 27054 12068 27106
rect 12012 27052 12068 27054
rect 12332 27106 12388 27108
rect 12332 27054 12334 27106
rect 12334 27054 12386 27106
rect 12386 27054 12388 27106
rect 12332 27052 12388 27054
rect 8492 26946 8548 26948
rect 8492 26894 8494 26946
rect 8494 26894 8546 26946
rect 8546 26894 8548 26946
rect 8492 26892 8548 26894
rect 8812 26946 8868 26948
rect 8812 26894 8814 26946
rect 8814 26894 8866 26946
rect 8866 26894 8868 26946
rect 8812 26892 8868 26894
rect 8972 26946 9028 26948
rect 8972 26894 8974 26946
rect 8974 26894 9026 26946
rect 9026 26894 9028 26946
rect 8972 26892 9028 26894
rect 9292 26946 9348 26948
rect 9292 26894 9294 26946
rect 9294 26894 9346 26946
rect 9346 26894 9348 26946
rect 9292 26892 9348 26894
rect 9452 26946 9508 26948
rect 9452 26894 9454 26946
rect 9454 26894 9506 26946
rect 9506 26894 9508 26946
rect 9452 26892 9508 26894
rect 9772 26946 9828 26948
rect 9772 26894 9774 26946
rect 9774 26894 9826 26946
rect 9826 26894 9828 26946
rect 9772 26892 9828 26894
rect 10092 26946 10148 26948
rect 10092 26894 10094 26946
rect 10094 26894 10146 26946
rect 10146 26894 10148 26946
rect 10092 26892 10148 26894
rect 10412 26946 10468 26948
rect 10412 26894 10414 26946
rect 10414 26894 10466 26946
rect 10466 26894 10468 26946
rect 10412 26892 10468 26894
rect 10732 26946 10788 26948
rect 10732 26894 10734 26946
rect 10734 26894 10786 26946
rect 10786 26894 10788 26946
rect 10732 26892 10788 26894
rect 11052 26946 11108 26948
rect 11052 26894 11054 26946
rect 11054 26894 11106 26946
rect 11106 26894 11108 26946
rect 11052 26892 11108 26894
rect 11372 26946 11428 26948
rect 11372 26894 11374 26946
rect 11374 26894 11426 26946
rect 11426 26894 11428 26946
rect 11372 26892 11428 26894
rect 11532 26946 11588 26948
rect 11532 26894 11534 26946
rect 11534 26894 11586 26946
rect 11586 26894 11588 26946
rect 11532 26892 11588 26894
rect 11852 26946 11908 26948
rect 11852 26894 11854 26946
rect 11854 26894 11906 26946
rect 11906 26894 11908 26946
rect 11852 26892 11908 26894
rect 12012 26946 12068 26948
rect 12012 26894 12014 26946
rect 12014 26894 12066 26946
rect 12066 26894 12068 26946
rect 12012 26892 12068 26894
rect 12332 26946 12388 26948
rect 12332 26894 12334 26946
rect 12334 26894 12386 26946
rect 12386 26894 12388 26946
rect 12332 26892 12388 26894
rect 10572 26652 10628 26708
rect 10252 26332 10308 26388
rect 10572 26332 10628 26388
rect 8492 26146 8548 26148
rect 8492 26094 8494 26146
rect 8494 26094 8546 26146
rect 8546 26094 8548 26146
rect 8492 26092 8548 26094
rect 8812 26146 8868 26148
rect 8812 26094 8814 26146
rect 8814 26094 8866 26146
rect 8866 26094 8868 26146
rect 8812 26092 8868 26094
rect 8972 26146 9028 26148
rect 8972 26094 8974 26146
rect 8974 26094 9026 26146
rect 9026 26094 9028 26146
rect 8972 26092 9028 26094
rect 9292 26146 9348 26148
rect 9292 26094 9294 26146
rect 9294 26094 9346 26146
rect 9346 26094 9348 26146
rect 9292 26092 9348 26094
rect 9452 26146 9508 26148
rect 9452 26094 9454 26146
rect 9454 26094 9506 26146
rect 9506 26094 9508 26146
rect 9452 26092 9508 26094
rect 9772 26146 9828 26148
rect 9772 26094 9774 26146
rect 9774 26094 9826 26146
rect 9826 26094 9828 26146
rect 9772 26092 9828 26094
rect 10092 26146 10148 26148
rect 10092 26094 10094 26146
rect 10094 26094 10146 26146
rect 10146 26094 10148 26146
rect 10092 26092 10148 26094
rect 10412 26146 10468 26148
rect 10412 26094 10414 26146
rect 10414 26094 10466 26146
rect 10466 26094 10468 26146
rect 10412 26092 10468 26094
rect 10732 26146 10788 26148
rect 10732 26094 10734 26146
rect 10734 26094 10786 26146
rect 10786 26094 10788 26146
rect 10732 26092 10788 26094
rect 11052 26146 11108 26148
rect 11052 26094 11054 26146
rect 11054 26094 11106 26146
rect 11106 26094 11108 26146
rect 11052 26092 11108 26094
rect 11372 26146 11428 26148
rect 11372 26094 11374 26146
rect 11374 26094 11426 26146
rect 11426 26094 11428 26146
rect 11372 26092 11428 26094
rect 11532 26146 11588 26148
rect 11532 26094 11534 26146
rect 11534 26094 11586 26146
rect 11586 26094 11588 26146
rect 11532 26092 11588 26094
rect 11852 26146 11908 26148
rect 11852 26094 11854 26146
rect 11854 26094 11906 26146
rect 11906 26094 11908 26146
rect 11852 26092 11908 26094
rect 12012 26146 12068 26148
rect 12012 26094 12014 26146
rect 12014 26094 12066 26146
rect 12066 26094 12068 26146
rect 12012 26092 12068 26094
rect 12332 26146 12388 26148
rect 12332 26094 12334 26146
rect 12334 26094 12386 26146
rect 12386 26094 12388 26146
rect 12332 26092 12388 26094
rect 8492 25986 8548 25988
rect 8492 25934 8494 25986
rect 8494 25934 8546 25986
rect 8546 25934 8548 25986
rect 8492 25932 8548 25934
rect 8812 25986 8868 25988
rect 8812 25934 8814 25986
rect 8814 25934 8866 25986
rect 8866 25934 8868 25986
rect 8812 25932 8868 25934
rect 8972 25986 9028 25988
rect 8972 25934 8974 25986
rect 8974 25934 9026 25986
rect 9026 25934 9028 25986
rect 8972 25932 9028 25934
rect 9292 25986 9348 25988
rect 9292 25934 9294 25986
rect 9294 25934 9346 25986
rect 9346 25934 9348 25986
rect 9292 25932 9348 25934
rect 9452 25986 9508 25988
rect 9452 25934 9454 25986
rect 9454 25934 9506 25986
rect 9506 25934 9508 25986
rect 9452 25932 9508 25934
rect 9772 25986 9828 25988
rect 9772 25934 9774 25986
rect 9774 25934 9826 25986
rect 9826 25934 9828 25986
rect 9772 25932 9828 25934
rect 10092 25986 10148 25988
rect 10092 25934 10094 25986
rect 10094 25934 10146 25986
rect 10146 25934 10148 25986
rect 10092 25932 10148 25934
rect 10412 25986 10468 25988
rect 10412 25934 10414 25986
rect 10414 25934 10466 25986
rect 10466 25934 10468 25986
rect 10412 25932 10468 25934
rect 10732 25986 10788 25988
rect 10732 25934 10734 25986
rect 10734 25934 10786 25986
rect 10786 25934 10788 25986
rect 10732 25932 10788 25934
rect 11052 25986 11108 25988
rect 11052 25934 11054 25986
rect 11054 25934 11106 25986
rect 11106 25934 11108 25986
rect 11052 25932 11108 25934
rect 11372 25986 11428 25988
rect 11372 25934 11374 25986
rect 11374 25934 11426 25986
rect 11426 25934 11428 25986
rect 11372 25932 11428 25934
rect 11532 25986 11588 25988
rect 11532 25934 11534 25986
rect 11534 25934 11586 25986
rect 11586 25934 11588 25986
rect 11532 25932 11588 25934
rect 11852 25986 11908 25988
rect 11852 25934 11854 25986
rect 11854 25934 11906 25986
rect 11906 25934 11908 25986
rect 11852 25932 11908 25934
rect 12012 25986 12068 25988
rect 12012 25934 12014 25986
rect 12014 25934 12066 25986
rect 12066 25934 12068 25986
rect 12012 25932 12068 25934
rect 12332 25986 12388 25988
rect 12332 25934 12334 25986
rect 12334 25934 12386 25986
rect 12386 25934 12388 25986
rect 12332 25932 12388 25934
rect 8492 25826 8548 25828
rect 8492 25774 8494 25826
rect 8494 25774 8546 25826
rect 8546 25774 8548 25826
rect 8492 25772 8548 25774
rect 8812 25826 8868 25828
rect 8812 25774 8814 25826
rect 8814 25774 8866 25826
rect 8866 25774 8868 25826
rect 8812 25772 8868 25774
rect 8972 25826 9028 25828
rect 8972 25774 8974 25826
rect 8974 25774 9026 25826
rect 9026 25774 9028 25826
rect 8972 25772 9028 25774
rect 9292 25826 9348 25828
rect 9292 25774 9294 25826
rect 9294 25774 9346 25826
rect 9346 25774 9348 25826
rect 9292 25772 9348 25774
rect 9452 25826 9508 25828
rect 9452 25774 9454 25826
rect 9454 25774 9506 25826
rect 9506 25774 9508 25826
rect 9452 25772 9508 25774
rect 9772 25826 9828 25828
rect 9772 25774 9774 25826
rect 9774 25774 9826 25826
rect 9826 25774 9828 25826
rect 9772 25772 9828 25774
rect 10092 25826 10148 25828
rect 10092 25774 10094 25826
rect 10094 25774 10146 25826
rect 10146 25774 10148 25826
rect 10092 25772 10148 25774
rect 10412 25826 10468 25828
rect 10412 25774 10414 25826
rect 10414 25774 10466 25826
rect 10466 25774 10468 25826
rect 10412 25772 10468 25774
rect 10732 25826 10788 25828
rect 10732 25774 10734 25826
rect 10734 25774 10786 25826
rect 10786 25774 10788 25826
rect 10732 25772 10788 25774
rect 11052 25826 11108 25828
rect 11052 25774 11054 25826
rect 11054 25774 11106 25826
rect 11106 25774 11108 25826
rect 11052 25772 11108 25774
rect 11372 25826 11428 25828
rect 11372 25774 11374 25826
rect 11374 25774 11426 25826
rect 11426 25774 11428 25826
rect 11372 25772 11428 25774
rect 11532 25826 11588 25828
rect 11532 25774 11534 25826
rect 11534 25774 11586 25826
rect 11586 25774 11588 25826
rect 11532 25772 11588 25774
rect 11852 25826 11908 25828
rect 11852 25774 11854 25826
rect 11854 25774 11906 25826
rect 11906 25774 11908 25826
rect 11852 25772 11908 25774
rect 12012 25826 12068 25828
rect 12012 25774 12014 25826
rect 12014 25774 12066 25826
rect 12066 25774 12068 25826
rect 12012 25772 12068 25774
rect 12332 25826 12388 25828
rect 12332 25774 12334 25826
rect 12334 25774 12386 25826
rect 12386 25774 12388 25826
rect 12332 25772 12388 25774
rect 8492 25666 8548 25668
rect 8492 25614 8494 25666
rect 8494 25614 8546 25666
rect 8546 25614 8548 25666
rect 8492 25612 8548 25614
rect 8812 25666 8868 25668
rect 8812 25614 8814 25666
rect 8814 25614 8866 25666
rect 8866 25614 8868 25666
rect 8812 25612 8868 25614
rect 8972 25666 9028 25668
rect 8972 25614 8974 25666
rect 8974 25614 9026 25666
rect 9026 25614 9028 25666
rect 8972 25612 9028 25614
rect 9292 25666 9348 25668
rect 9292 25614 9294 25666
rect 9294 25614 9346 25666
rect 9346 25614 9348 25666
rect 9292 25612 9348 25614
rect 9452 25666 9508 25668
rect 9452 25614 9454 25666
rect 9454 25614 9506 25666
rect 9506 25614 9508 25666
rect 9452 25612 9508 25614
rect 9772 25666 9828 25668
rect 9772 25614 9774 25666
rect 9774 25614 9826 25666
rect 9826 25614 9828 25666
rect 9772 25612 9828 25614
rect 10092 25666 10148 25668
rect 10092 25614 10094 25666
rect 10094 25614 10146 25666
rect 10146 25614 10148 25666
rect 10092 25612 10148 25614
rect 10412 25666 10468 25668
rect 10412 25614 10414 25666
rect 10414 25614 10466 25666
rect 10466 25614 10468 25666
rect 10412 25612 10468 25614
rect 10732 25666 10788 25668
rect 10732 25614 10734 25666
rect 10734 25614 10786 25666
rect 10786 25614 10788 25666
rect 10732 25612 10788 25614
rect 11052 25666 11108 25668
rect 11052 25614 11054 25666
rect 11054 25614 11106 25666
rect 11106 25614 11108 25666
rect 11052 25612 11108 25614
rect 11372 25666 11428 25668
rect 11372 25614 11374 25666
rect 11374 25614 11426 25666
rect 11426 25614 11428 25666
rect 11372 25612 11428 25614
rect 11532 25666 11588 25668
rect 11532 25614 11534 25666
rect 11534 25614 11586 25666
rect 11586 25614 11588 25666
rect 11532 25612 11588 25614
rect 11852 25666 11908 25668
rect 11852 25614 11854 25666
rect 11854 25614 11906 25666
rect 11906 25614 11908 25666
rect 11852 25612 11908 25614
rect 12012 25666 12068 25668
rect 12012 25614 12014 25666
rect 12014 25614 12066 25666
rect 12066 25614 12068 25666
rect 12012 25612 12068 25614
rect 12332 25666 12388 25668
rect 12332 25614 12334 25666
rect 12334 25614 12386 25666
rect 12386 25614 12388 25666
rect 12332 25612 12388 25614
rect 8492 25506 8548 25508
rect 8492 25454 8494 25506
rect 8494 25454 8546 25506
rect 8546 25454 8548 25506
rect 8492 25452 8548 25454
rect 8812 25506 8868 25508
rect 8812 25454 8814 25506
rect 8814 25454 8866 25506
rect 8866 25454 8868 25506
rect 8812 25452 8868 25454
rect 8972 25506 9028 25508
rect 8972 25454 8974 25506
rect 8974 25454 9026 25506
rect 9026 25454 9028 25506
rect 8972 25452 9028 25454
rect 9292 25506 9348 25508
rect 9292 25454 9294 25506
rect 9294 25454 9346 25506
rect 9346 25454 9348 25506
rect 9292 25452 9348 25454
rect 9452 25506 9508 25508
rect 9452 25454 9454 25506
rect 9454 25454 9506 25506
rect 9506 25454 9508 25506
rect 9452 25452 9508 25454
rect 9772 25506 9828 25508
rect 9772 25454 9774 25506
rect 9774 25454 9826 25506
rect 9826 25454 9828 25506
rect 9772 25452 9828 25454
rect 10092 25506 10148 25508
rect 10092 25454 10094 25506
rect 10094 25454 10146 25506
rect 10146 25454 10148 25506
rect 10092 25452 10148 25454
rect 10412 25506 10468 25508
rect 10412 25454 10414 25506
rect 10414 25454 10466 25506
rect 10466 25454 10468 25506
rect 10412 25452 10468 25454
rect 10732 25506 10788 25508
rect 10732 25454 10734 25506
rect 10734 25454 10786 25506
rect 10786 25454 10788 25506
rect 10732 25452 10788 25454
rect 11052 25506 11108 25508
rect 11052 25454 11054 25506
rect 11054 25454 11106 25506
rect 11106 25454 11108 25506
rect 11052 25452 11108 25454
rect 11372 25506 11428 25508
rect 11372 25454 11374 25506
rect 11374 25454 11426 25506
rect 11426 25454 11428 25506
rect 11372 25452 11428 25454
rect 11532 25506 11588 25508
rect 11532 25454 11534 25506
rect 11534 25454 11586 25506
rect 11586 25454 11588 25506
rect 11532 25452 11588 25454
rect 11852 25506 11908 25508
rect 11852 25454 11854 25506
rect 11854 25454 11906 25506
rect 11906 25454 11908 25506
rect 11852 25452 11908 25454
rect 12012 25506 12068 25508
rect 12012 25454 12014 25506
rect 12014 25454 12066 25506
rect 12066 25454 12068 25506
rect 12012 25452 12068 25454
rect 12332 25506 12388 25508
rect 12332 25454 12334 25506
rect 12334 25454 12386 25506
rect 12386 25454 12388 25506
rect 12332 25452 12388 25454
rect 8492 25346 8548 25348
rect 8492 25294 8494 25346
rect 8494 25294 8546 25346
rect 8546 25294 8548 25346
rect 8492 25292 8548 25294
rect 8812 25346 8868 25348
rect 8812 25294 8814 25346
rect 8814 25294 8866 25346
rect 8866 25294 8868 25346
rect 8812 25292 8868 25294
rect 8972 25346 9028 25348
rect 8972 25294 8974 25346
rect 8974 25294 9026 25346
rect 9026 25294 9028 25346
rect 8972 25292 9028 25294
rect 9292 25346 9348 25348
rect 9292 25294 9294 25346
rect 9294 25294 9346 25346
rect 9346 25294 9348 25346
rect 9292 25292 9348 25294
rect 9452 25346 9508 25348
rect 9452 25294 9454 25346
rect 9454 25294 9506 25346
rect 9506 25294 9508 25346
rect 9452 25292 9508 25294
rect 9772 25346 9828 25348
rect 9772 25294 9774 25346
rect 9774 25294 9826 25346
rect 9826 25294 9828 25346
rect 9772 25292 9828 25294
rect 10092 25346 10148 25348
rect 10092 25294 10094 25346
rect 10094 25294 10146 25346
rect 10146 25294 10148 25346
rect 10092 25292 10148 25294
rect 10412 25346 10468 25348
rect 10412 25294 10414 25346
rect 10414 25294 10466 25346
rect 10466 25294 10468 25346
rect 10412 25292 10468 25294
rect 10732 25346 10788 25348
rect 10732 25294 10734 25346
rect 10734 25294 10786 25346
rect 10786 25294 10788 25346
rect 10732 25292 10788 25294
rect 11052 25346 11108 25348
rect 11052 25294 11054 25346
rect 11054 25294 11106 25346
rect 11106 25294 11108 25346
rect 11052 25292 11108 25294
rect 11372 25346 11428 25348
rect 11372 25294 11374 25346
rect 11374 25294 11426 25346
rect 11426 25294 11428 25346
rect 11372 25292 11428 25294
rect 11532 25346 11588 25348
rect 11532 25294 11534 25346
rect 11534 25294 11586 25346
rect 11586 25294 11588 25346
rect 11532 25292 11588 25294
rect 11852 25346 11908 25348
rect 11852 25294 11854 25346
rect 11854 25294 11906 25346
rect 11906 25294 11908 25346
rect 11852 25292 11908 25294
rect 12012 25346 12068 25348
rect 12012 25294 12014 25346
rect 12014 25294 12066 25346
rect 12066 25294 12068 25346
rect 12012 25292 12068 25294
rect 12332 25346 12388 25348
rect 12332 25294 12334 25346
rect 12334 25294 12386 25346
rect 12386 25294 12388 25346
rect 12332 25292 12388 25294
rect 8492 25186 8548 25188
rect 8492 25134 8494 25186
rect 8494 25134 8546 25186
rect 8546 25134 8548 25186
rect 8492 25132 8548 25134
rect 8812 25186 8868 25188
rect 8812 25134 8814 25186
rect 8814 25134 8866 25186
rect 8866 25134 8868 25186
rect 8812 25132 8868 25134
rect 8972 25186 9028 25188
rect 8972 25134 8974 25186
rect 8974 25134 9026 25186
rect 9026 25134 9028 25186
rect 8972 25132 9028 25134
rect 9292 25186 9348 25188
rect 9292 25134 9294 25186
rect 9294 25134 9346 25186
rect 9346 25134 9348 25186
rect 9292 25132 9348 25134
rect 9452 25186 9508 25188
rect 9452 25134 9454 25186
rect 9454 25134 9506 25186
rect 9506 25134 9508 25186
rect 9452 25132 9508 25134
rect 9772 25186 9828 25188
rect 9772 25134 9774 25186
rect 9774 25134 9826 25186
rect 9826 25134 9828 25186
rect 9772 25132 9828 25134
rect 10092 25186 10148 25188
rect 10092 25134 10094 25186
rect 10094 25134 10146 25186
rect 10146 25134 10148 25186
rect 10092 25132 10148 25134
rect 10412 25186 10468 25188
rect 10412 25134 10414 25186
rect 10414 25134 10466 25186
rect 10466 25134 10468 25186
rect 10412 25132 10468 25134
rect 10732 25186 10788 25188
rect 10732 25134 10734 25186
rect 10734 25134 10786 25186
rect 10786 25134 10788 25186
rect 10732 25132 10788 25134
rect 11052 25186 11108 25188
rect 11052 25134 11054 25186
rect 11054 25134 11106 25186
rect 11106 25134 11108 25186
rect 11052 25132 11108 25134
rect 11372 25186 11428 25188
rect 11372 25134 11374 25186
rect 11374 25134 11426 25186
rect 11426 25134 11428 25186
rect 11372 25132 11428 25134
rect 11532 25186 11588 25188
rect 11532 25134 11534 25186
rect 11534 25134 11586 25186
rect 11586 25134 11588 25186
rect 11532 25132 11588 25134
rect 11852 25186 11908 25188
rect 11852 25134 11854 25186
rect 11854 25134 11906 25186
rect 11906 25134 11908 25186
rect 11852 25132 11908 25134
rect 12012 25186 12068 25188
rect 12012 25134 12014 25186
rect 12014 25134 12066 25186
rect 12066 25134 12068 25186
rect 12012 25132 12068 25134
rect 12332 25186 12388 25188
rect 12332 25134 12334 25186
rect 12334 25134 12386 25186
rect 12386 25134 12388 25186
rect 12332 25132 12388 25134
rect 8492 25026 8548 25028
rect 8492 24974 8494 25026
rect 8494 24974 8546 25026
rect 8546 24974 8548 25026
rect 8492 24972 8548 24974
rect 8812 25026 8868 25028
rect 8812 24974 8814 25026
rect 8814 24974 8866 25026
rect 8866 24974 8868 25026
rect 8812 24972 8868 24974
rect 8972 25026 9028 25028
rect 8972 24974 8974 25026
rect 8974 24974 9026 25026
rect 9026 24974 9028 25026
rect 8972 24972 9028 24974
rect 9292 25026 9348 25028
rect 9292 24974 9294 25026
rect 9294 24974 9346 25026
rect 9346 24974 9348 25026
rect 9292 24972 9348 24974
rect 9452 25026 9508 25028
rect 9452 24974 9454 25026
rect 9454 24974 9506 25026
rect 9506 24974 9508 25026
rect 9452 24972 9508 24974
rect 9772 25026 9828 25028
rect 9772 24974 9774 25026
rect 9774 24974 9826 25026
rect 9826 24974 9828 25026
rect 9772 24972 9828 24974
rect 10092 25026 10148 25028
rect 10092 24974 10094 25026
rect 10094 24974 10146 25026
rect 10146 24974 10148 25026
rect 10092 24972 10148 24974
rect 10412 25026 10468 25028
rect 10412 24974 10414 25026
rect 10414 24974 10466 25026
rect 10466 24974 10468 25026
rect 10412 24972 10468 24974
rect 10732 25026 10788 25028
rect 10732 24974 10734 25026
rect 10734 24974 10786 25026
rect 10786 24974 10788 25026
rect 10732 24972 10788 24974
rect 11052 25026 11108 25028
rect 11052 24974 11054 25026
rect 11054 24974 11106 25026
rect 11106 24974 11108 25026
rect 11052 24972 11108 24974
rect 11372 25026 11428 25028
rect 11372 24974 11374 25026
rect 11374 24974 11426 25026
rect 11426 24974 11428 25026
rect 11372 24972 11428 24974
rect 11532 25026 11588 25028
rect 11532 24974 11534 25026
rect 11534 24974 11586 25026
rect 11586 24974 11588 25026
rect 11532 24972 11588 24974
rect 11852 25026 11908 25028
rect 11852 24974 11854 25026
rect 11854 24974 11906 25026
rect 11906 24974 11908 25026
rect 11852 24972 11908 24974
rect 12012 25026 12068 25028
rect 12012 24974 12014 25026
rect 12014 24974 12066 25026
rect 12066 24974 12068 25026
rect 12012 24972 12068 24974
rect 12332 25026 12388 25028
rect 12332 24974 12334 25026
rect 12334 24974 12386 25026
rect 12386 24974 12388 25026
rect 12332 24972 12388 24974
rect 9132 24812 9188 24868
rect 8492 24706 8548 24708
rect 8492 24654 8494 24706
rect 8494 24654 8546 24706
rect 8546 24654 8548 24706
rect 8492 24652 8548 24654
rect 8812 24706 8868 24708
rect 8812 24654 8814 24706
rect 8814 24654 8866 24706
rect 8866 24654 8868 24706
rect 8812 24652 8868 24654
rect 8972 24706 9028 24708
rect 8972 24654 8974 24706
rect 8974 24654 9026 24706
rect 9026 24654 9028 24706
rect 8972 24652 9028 24654
rect 9292 24706 9348 24708
rect 9292 24654 9294 24706
rect 9294 24654 9346 24706
rect 9346 24654 9348 24706
rect 9292 24652 9348 24654
rect 9452 24706 9508 24708
rect 9452 24654 9454 24706
rect 9454 24654 9506 24706
rect 9506 24654 9508 24706
rect 9452 24652 9508 24654
rect 9772 24706 9828 24708
rect 9772 24654 9774 24706
rect 9774 24654 9826 24706
rect 9826 24654 9828 24706
rect 9772 24652 9828 24654
rect 10092 24706 10148 24708
rect 10092 24654 10094 24706
rect 10094 24654 10146 24706
rect 10146 24654 10148 24706
rect 10092 24652 10148 24654
rect 10412 24706 10468 24708
rect 10412 24654 10414 24706
rect 10414 24654 10466 24706
rect 10466 24654 10468 24706
rect 10412 24652 10468 24654
rect 10732 24706 10788 24708
rect 10732 24654 10734 24706
rect 10734 24654 10786 24706
rect 10786 24654 10788 24706
rect 10732 24652 10788 24654
rect 11052 24706 11108 24708
rect 11052 24654 11054 24706
rect 11054 24654 11106 24706
rect 11106 24654 11108 24706
rect 11052 24652 11108 24654
rect 11372 24706 11428 24708
rect 11372 24654 11374 24706
rect 11374 24654 11426 24706
rect 11426 24654 11428 24706
rect 11372 24652 11428 24654
rect 11532 24706 11588 24708
rect 11532 24654 11534 24706
rect 11534 24654 11586 24706
rect 11586 24654 11588 24706
rect 11532 24652 11588 24654
rect 11852 24706 11908 24708
rect 11852 24654 11854 24706
rect 11854 24654 11906 24706
rect 11906 24654 11908 24706
rect 11852 24652 11908 24654
rect 12012 24706 12068 24708
rect 12012 24654 12014 24706
rect 12014 24654 12066 24706
rect 12066 24654 12068 24706
rect 12012 24652 12068 24654
rect 12332 24706 12388 24708
rect 12332 24654 12334 24706
rect 12334 24654 12386 24706
rect 12386 24654 12388 24706
rect 12332 24652 12388 24654
rect 8492 24546 8548 24548
rect 8492 24494 8494 24546
rect 8494 24494 8546 24546
rect 8546 24494 8548 24546
rect 8492 24492 8548 24494
rect 8812 24546 8868 24548
rect 8812 24494 8814 24546
rect 8814 24494 8866 24546
rect 8866 24494 8868 24546
rect 8812 24492 8868 24494
rect 8972 24546 9028 24548
rect 8972 24494 8974 24546
rect 8974 24494 9026 24546
rect 9026 24494 9028 24546
rect 8972 24492 9028 24494
rect 9292 24546 9348 24548
rect 9292 24494 9294 24546
rect 9294 24494 9346 24546
rect 9346 24494 9348 24546
rect 9292 24492 9348 24494
rect 9452 24546 9508 24548
rect 9452 24494 9454 24546
rect 9454 24494 9506 24546
rect 9506 24494 9508 24546
rect 9452 24492 9508 24494
rect 9772 24546 9828 24548
rect 9772 24494 9774 24546
rect 9774 24494 9826 24546
rect 9826 24494 9828 24546
rect 9772 24492 9828 24494
rect 10092 24546 10148 24548
rect 10092 24494 10094 24546
rect 10094 24494 10146 24546
rect 10146 24494 10148 24546
rect 10092 24492 10148 24494
rect 10412 24546 10468 24548
rect 10412 24494 10414 24546
rect 10414 24494 10466 24546
rect 10466 24494 10468 24546
rect 10412 24492 10468 24494
rect 10732 24546 10788 24548
rect 10732 24494 10734 24546
rect 10734 24494 10786 24546
rect 10786 24494 10788 24546
rect 10732 24492 10788 24494
rect 11052 24546 11108 24548
rect 11052 24494 11054 24546
rect 11054 24494 11106 24546
rect 11106 24494 11108 24546
rect 11052 24492 11108 24494
rect 11372 24546 11428 24548
rect 11372 24494 11374 24546
rect 11374 24494 11426 24546
rect 11426 24494 11428 24546
rect 11372 24492 11428 24494
rect 11532 24546 11588 24548
rect 11532 24494 11534 24546
rect 11534 24494 11586 24546
rect 11586 24494 11588 24546
rect 11532 24492 11588 24494
rect 11852 24546 11908 24548
rect 11852 24494 11854 24546
rect 11854 24494 11906 24546
rect 11906 24494 11908 24546
rect 11852 24492 11908 24494
rect 12012 24546 12068 24548
rect 12012 24494 12014 24546
rect 12014 24494 12066 24546
rect 12066 24494 12068 24546
rect 12012 24492 12068 24494
rect 12332 24546 12388 24548
rect 12332 24494 12334 24546
rect 12334 24494 12386 24546
rect 12386 24494 12388 24546
rect 12332 24492 12388 24494
rect 8492 24386 8548 24388
rect 8492 24334 8494 24386
rect 8494 24334 8546 24386
rect 8546 24334 8548 24386
rect 8492 24332 8548 24334
rect 8812 24386 8868 24388
rect 8812 24334 8814 24386
rect 8814 24334 8866 24386
rect 8866 24334 8868 24386
rect 8812 24332 8868 24334
rect 8972 24386 9028 24388
rect 8972 24334 8974 24386
rect 8974 24334 9026 24386
rect 9026 24334 9028 24386
rect 8972 24332 9028 24334
rect 9292 24386 9348 24388
rect 9292 24334 9294 24386
rect 9294 24334 9346 24386
rect 9346 24334 9348 24386
rect 9292 24332 9348 24334
rect 9452 24386 9508 24388
rect 9452 24334 9454 24386
rect 9454 24334 9506 24386
rect 9506 24334 9508 24386
rect 9452 24332 9508 24334
rect 9772 24386 9828 24388
rect 9772 24334 9774 24386
rect 9774 24334 9826 24386
rect 9826 24334 9828 24386
rect 9772 24332 9828 24334
rect 10092 24386 10148 24388
rect 10092 24334 10094 24386
rect 10094 24334 10146 24386
rect 10146 24334 10148 24386
rect 10092 24332 10148 24334
rect 10412 24386 10468 24388
rect 10412 24334 10414 24386
rect 10414 24334 10466 24386
rect 10466 24334 10468 24386
rect 10412 24332 10468 24334
rect 10732 24386 10788 24388
rect 10732 24334 10734 24386
rect 10734 24334 10786 24386
rect 10786 24334 10788 24386
rect 10732 24332 10788 24334
rect 11052 24386 11108 24388
rect 11052 24334 11054 24386
rect 11054 24334 11106 24386
rect 11106 24334 11108 24386
rect 11052 24332 11108 24334
rect 11372 24386 11428 24388
rect 11372 24334 11374 24386
rect 11374 24334 11426 24386
rect 11426 24334 11428 24386
rect 11372 24332 11428 24334
rect 11532 24386 11588 24388
rect 11532 24334 11534 24386
rect 11534 24334 11586 24386
rect 11586 24334 11588 24386
rect 11532 24332 11588 24334
rect 11852 24386 11908 24388
rect 11852 24334 11854 24386
rect 11854 24334 11906 24386
rect 11906 24334 11908 24386
rect 11852 24332 11908 24334
rect 12012 24386 12068 24388
rect 12012 24334 12014 24386
rect 12014 24334 12066 24386
rect 12066 24334 12068 24386
rect 12012 24332 12068 24334
rect 12332 24386 12388 24388
rect 12332 24334 12334 24386
rect 12334 24334 12386 24386
rect 12386 24334 12388 24386
rect 12332 24332 12388 24334
rect 8492 24226 8548 24228
rect 8492 24174 8494 24226
rect 8494 24174 8546 24226
rect 8546 24174 8548 24226
rect 8492 24172 8548 24174
rect 8812 24226 8868 24228
rect 8812 24174 8814 24226
rect 8814 24174 8866 24226
rect 8866 24174 8868 24226
rect 8812 24172 8868 24174
rect 8972 24226 9028 24228
rect 8972 24174 8974 24226
rect 8974 24174 9026 24226
rect 9026 24174 9028 24226
rect 8972 24172 9028 24174
rect 9292 24226 9348 24228
rect 9292 24174 9294 24226
rect 9294 24174 9346 24226
rect 9346 24174 9348 24226
rect 9292 24172 9348 24174
rect 9452 24226 9508 24228
rect 9452 24174 9454 24226
rect 9454 24174 9506 24226
rect 9506 24174 9508 24226
rect 9452 24172 9508 24174
rect 9772 24226 9828 24228
rect 9772 24174 9774 24226
rect 9774 24174 9826 24226
rect 9826 24174 9828 24226
rect 9772 24172 9828 24174
rect 10092 24226 10148 24228
rect 10092 24174 10094 24226
rect 10094 24174 10146 24226
rect 10146 24174 10148 24226
rect 10092 24172 10148 24174
rect 10412 24226 10468 24228
rect 10412 24174 10414 24226
rect 10414 24174 10466 24226
rect 10466 24174 10468 24226
rect 10412 24172 10468 24174
rect 10732 24226 10788 24228
rect 10732 24174 10734 24226
rect 10734 24174 10786 24226
rect 10786 24174 10788 24226
rect 10732 24172 10788 24174
rect 11052 24226 11108 24228
rect 11052 24174 11054 24226
rect 11054 24174 11106 24226
rect 11106 24174 11108 24226
rect 11052 24172 11108 24174
rect 11372 24226 11428 24228
rect 11372 24174 11374 24226
rect 11374 24174 11426 24226
rect 11426 24174 11428 24226
rect 11372 24172 11428 24174
rect 11532 24226 11588 24228
rect 11532 24174 11534 24226
rect 11534 24174 11586 24226
rect 11586 24174 11588 24226
rect 11532 24172 11588 24174
rect 11852 24226 11908 24228
rect 11852 24174 11854 24226
rect 11854 24174 11906 24226
rect 11906 24174 11908 24226
rect 11852 24172 11908 24174
rect 12012 24226 12068 24228
rect 12012 24174 12014 24226
rect 12014 24174 12066 24226
rect 12066 24174 12068 24226
rect 12012 24172 12068 24174
rect 12332 24226 12388 24228
rect 12332 24174 12334 24226
rect 12334 24174 12386 24226
rect 12386 24174 12388 24226
rect 12332 24172 12388 24174
rect 8492 24066 8548 24068
rect 8492 24014 8494 24066
rect 8494 24014 8546 24066
rect 8546 24014 8548 24066
rect 8492 24012 8548 24014
rect 8812 24066 8868 24068
rect 8812 24014 8814 24066
rect 8814 24014 8866 24066
rect 8866 24014 8868 24066
rect 8812 24012 8868 24014
rect 8972 24066 9028 24068
rect 8972 24014 8974 24066
rect 8974 24014 9026 24066
rect 9026 24014 9028 24066
rect 8972 24012 9028 24014
rect 9292 24066 9348 24068
rect 9292 24014 9294 24066
rect 9294 24014 9346 24066
rect 9346 24014 9348 24066
rect 9292 24012 9348 24014
rect 9452 24066 9508 24068
rect 9452 24014 9454 24066
rect 9454 24014 9506 24066
rect 9506 24014 9508 24066
rect 9452 24012 9508 24014
rect 9772 24066 9828 24068
rect 9772 24014 9774 24066
rect 9774 24014 9826 24066
rect 9826 24014 9828 24066
rect 9772 24012 9828 24014
rect 10092 24066 10148 24068
rect 10092 24014 10094 24066
rect 10094 24014 10146 24066
rect 10146 24014 10148 24066
rect 10092 24012 10148 24014
rect 10412 24066 10468 24068
rect 10412 24014 10414 24066
rect 10414 24014 10466 24066
rect 10466 24014 10468 24066
rect 10412 24012 10468 24014
rect 10732 24066 10788 24068
rect 10732 24014 10734 24066
rect 10734 24014 10786 24066
rect 10786 24014 10788 24066
rect 10732 24012 10788 24014
rect 11052 24066 11108 24068
rect 11052 24014 11054 24066
rect 11054 24014 11106 24066
rect 11106 24014 11108 24066
rect 11052 24012 11108 24014
rect 11372 24066 11428 24068
rect 11372 24014 11374 24066
rect 11374 24014 11426 24066
rect 11426 24014 11428 24066
rect 11372 24012 11428 24014
rect 11532 24066 11588 24068
rect 11532 24014 11534 24066
rect 11534 24014 11586 24066
rect 11586 24014 11588 24066
rect 11532 24012 11588 24014
rect 11852 24066 11908 24068
rect 11852 24014 11854 24066
rect 11854 24014 11906 24066
rect 11906 24014 11908 24066
rect 11852 24012 11908 24014
rect 12012 24066 12068 24068
rect 12012 24014 12014 24066
rect 12014 24014 12066 24066
rect 12066 24014 12068 24066
rect 12012 24012 12068 24014
rect 12332 24066 12388 24068
rect 12332 24014 12334 24066
rect 12334 24014 12386 24066
rect 12386 24014 12388 24066
rect 12332 24012 12388 24014
rect 8492 23906 8548 23908
rect 8492 23854 8494 23906
rect 8494 23854 8546 23906
rect 8546 23854 8548 23906
rect 8492 23852 8548 23854
rect 8812 23906 8868 23908
rect 8812 23854 8814 23906
rect 8814 23854 8866 23906
rect 8866 23854 8868 23906
rect 8812 23852 8868 23854
rect 8972 23906 9028 23908
rect 8972 23854 8974 23906
rect 8974 23854 9026 23906
rect 9026 23854 9028 23906
rect 8972 23852 9028 23854
rect 9292 23906 9348 23908
rect 9292 23854 9294 23906
rect 9294 23854 9346 23906
rect 9346 23854 9348 23906
rect 9292 23852 9348 23854
rect 9452 23906 9508 23908
rect 9452 23854 9454 23906
rect 9454 23854 9506 23906
rect 9506 23854 9508 23906
rect 9452 23852 9508 23854
rect 9772 23906 9828 23908
rect 9772 23854 9774 23906
rect 9774 23854 9826 23906
rect 9826 23854 9828 23906
rect 9772 23852 9828 23854
rect 10092 23906 10148 23908
rect 10092 23854 10094 23906
rect 10094 23854 10146 23906
rect 10146 23854 10148 23906
rect 10092 23852 10148 23854
rect 10412 23906 10468 23908
rect 10412 23854 10414 23906
rect 10414 23854 10466 23906
rect 10466 23854 10468 23906
rect 10412 23852 10468 23854
rect 10732 23906 10788 23908
rect 10732 23854 10734 23906
rect 10734 23854 10786 23906
rect 10786 23854 10788 23906
rect 10732 23852 10788 23854
rect 11052 23906 11108 23908
rect 11052 23854 11054 23906
rect 11054 23854 11106 23906
rect 11106 23854 11108 23906
rect 11052 23852 11108 23854
rect 11372 23906 11428 23908
rect 11372 23854 11374 23906
rect 11374 23854 11426 23906
rect 11426 23854 11428 23906
rect 11372 23852 11428 23854
rect 11532 23906 11588 23908
rect 11532 23854 11534 23906
rect 11534 23854 11586 23906
rect 11586 23854 11588 23906
rect 11532 23852 11588 23854
rect 11852 23906 11908 23908
rect 11852 23854 11854 23906
rect 11854 23854 11906 23906
rect 11906 23854 11908 23906
rect 11852 23852 11908 23854
rect 12012 23906 12068 23908
rect 12012 23854 12014 23906
rect 12014 23854 12066 23906
rect 12066 23854 12068 23906
rect 12012 23852 12068 23854
rect 12332 23906 12388 23908
rect 12332 23854 12334 23906
rect 12334 23854 12386 23906
rect 12386 23854 12388 23906
rect 12332 23852 12388 23854
rect 8492 23746 8548 23748
rect 8492 23694 8494 23746
rect 8494 23694 8546 23746
rect 8546 23694 8548 23746
rect 8492 23692 8548 23694
rect 8812 23746 8868 23748
rect 8812 23694 8814 23746
rect 8814 23694 8866 23746
rect 8866 23694 8868 23746
rect 8812 23692 8868 23694
rect 8972 23746 9028 23748
rect 8972 23694 8974 23746
rect 8974 23694 9026 23746
rect 9026 23694 9028 23746
rect 8972 23692 9028 23694
rect 9292 23746 9348 23748
rect 9292 23694 9294 23746
rect 9294 23694 9346 23746
rect 9346 23694 9348 23746
rect 9292 23692 9348 23694
rect 9452 23746 9508 23748
rect 9452 23694 9454 23746
rect 9454 23694 9506 23746
rect 9506 23694 9508 23746
rect 9452 23692 9508 23694
rect 9772 23746 9828 23748
rect 9772 23694 9774 23746
rect 9774 23694 9826 23746
rect 9826 23694 9828 23746
rect 9772 23692 9828 23694
rect 10092 23746 10148 23748
rect 10092 23694 10094 23746
rect 10094 23694 10146 23746
rect 10146 23694 10148 23746
rect 10092 23692 10148 23694
rect 10412 23746 10468 23748
rect 10412 23694 10414 23746
rect 10414 23694 10466 23746
rect 10466 23694 10468 23746
rect 10412 23692 10468 23694
rect 10732 23746 10788 23748
rect 10732 23694 10734 23746
rect 10734 23694 10786 23746
rect 10786 23694 10788 23746
rect 10732 23692 10788 23694
rect 11052 23746 11108 23748
rect 11052 23694 11054 23746
rect 11054 23694 11106 23746
rect 11106 23694 11108 23746
rect 11052 23692 11108 23694
rect 11372 23746 11428 23748
rect 11372 23694 11374 23746
rect 11374 23694 11426 23746
rect 11426 23694 11428 23746
rect 11372 23692 11428 23694
rect 11532 23746 11588 23748
rect 11532 23694 11534 23746
rect 11534 23694 11586 23746
rect 11586 23694 11588 23746
rect 11532 23692 11588 23694
rect 11852 23746 11908 23748
rect 11852 23694 11854 23746
rect 11854 23694 11906 23746
rect 11906 23694 11908 23746
rect 11852 23692 11908 23694
rect 12012 23746 12068 23748
rect 12012 23694 12014 23746
rect 12014 23694 12066 23746
rect 12066 23694 12068 23746
rect 12012 23692 12068 23694
rect 12332 23746 12388 23748
rect 12332 23694 12334 23746
rect 12334 23694 12386 23746
rect 12386 23694 12388 23746
rect 12332 23692 12388 23694
rect 8492 23586 8548 23588
rect 8492 23534 8494 23586
rect 8494 23534 8546 23586
rect 8546 23534 8548 23586
rect 8492 23532 8548 23534
rect 8812 23586 8868 23588
rect 8812 23534 8814 23586
rect 8814 23534 8866 23586
rect 8866 23534 8868 23586
rect 8812 23532 8868 23534
rect 8972 23586 9028 23588
rect 8972 23534 8974 23586
rect 8974 23534 9026 23586
rect 9026 23534 9028 23586
rect 8972 23532 9028 23534
rect 9292 23586 9348 23588
rect 9292 23534 9294 23586
rect 9294 23534 9346 23586
rect 9346 23534 9348 23586
rect 9292 23532 9348 23534
rect 9452 23586 9508 23588
rect 9452 23534 9454 23586
rect 9454 23534 9506 23586
rect 9506 23534 9508 23586
rect 9452 23532 9508 23534
rect 9772 23586 9828 23588
rect 9772 23534 9774 23586
rect 9774 23534 9826 23586
rect 9826 23534 9828 23586
rect 9772 23532 9828 23534
rect 10092 23586 10148 23588
rect 10092 23534 10094 23586
rect 10094 23534 10146 23586
rect 10146 23534 10148 23586
rect 10092 23532 10148 23534
rect 10412 23586 10468 23588
rect 10412 23534 10414 23586
rect 10414 23534 10466 23586
rect 10466 23534 10468 23586
rect 10412 23532 10468 23534
rect 10732 23586 10788 23588
rect 10732 23534 10734 23586
rect 10734 23534 10786 23586
rect 10786 23534 10788 23586
rect 10732 23532 10788 23534
rect 11052 23586 11108 23588
rect 11052 23534 11054 23586
rect 11054 23534 11106 23586
rect 11106 23534 11108 23586
rect 11052 23532 11108 23534
rect 11372 23586 11428 23588
rect 11372 23534 11374 23586
rect 11374 23534 11426 23586
rect 11426 23534 11428 23586
rect 11372 23532 11428 23534
rect 11532 23586 11588 23588
rect 11532 23534 11534 23586
rect 11534 23534 11586 23586
rect 11586 23534 11588 23586
rect 11532 23532 11588 23534
rect 11852 23586 11908 23588
rect 11852 23534 11854 23586
rect 11854 23534 11906 23586
rect 11906 23534 11908 23586
rect 11852 23532 11908 23534
rect 12012 23586 12068 23588
rect 12012 23534 12014 23586
rect 12014 23534 12066 23586
rect 12066 23534 12068 23586
rect 12012 23532 12068 23534
rect 12332 23586 12388 23588
rect 12332 23534 12334 23586
rect 12334 23534 12386 23586
rect 12386 23534 12388 23586
rect 12332 23532 12388 23534
rect 8492 23426 8548 23428
rect 8492 23374 8494 23426
rect 8494 23374 8546 23426
rect 8546 23374 8548 23426
rect 8492 23372 8548 23374
rect 8812 23426 8868 23428
rect 8812 23374 8814 23426
rect 8814 23374 8866 23426
rect 8866 23374 8868 23426
rect 8812 23372 8868 23374
rect 8972 23426 9028 23428
rect 8972 23374 8974 23426
rect 8974 23374 9026 23426
rect 9026 23374 9028 23426
rect 8972 23372 9028 23374
rect 9292 23426 9348 23428
rect 9292 23374 9294 23426
rect 9294 23374 9346 23426
rect 9346 23374 9348 23426
rect 9292 23372 9348 23374
rect 9452 23426 9508 23428
rect 9452 23374 9454 23426
rect 9454 23374 9506 23426
rect 9506 23374 9508 23426
rect 9452 23372 9508 23374
rect 9772 23426 9828 23428
rect 9772 23374 9774 23426
rect 9774 23374 9826 23426
rect 9826 23374 9828 23426
rect 9772 23372 9828 23374
rect 10092 23426 10148 23428
rect 10092 23374 10094 23426
rect 10094 23374 10146 23426
rect 10146 23374 10148 23426
rect 10092 23372 10148 23374
rect 10412 23426 10468 23428
rect 10412 23374 10414 23426
rect 10414 23374 10466 23426
rect 10466 23374 10468 23426
rect 10412 23372 10468 23374
rect 10732 23426 10788 23428
rect 10732 23374 10734 23426
rect 10734 23374 10786 23426
rect 10786 23374 10788 23426
rect 10732 23372 10788 23374
rect 11052 23426 11108 23428
rect 11052 23374 11054 23426
rect 11054 23374 11106 23426
rect 11106 23374 11108 23426
rect 11052 23372 11108 23374
rect 11372 23426 11428 23428
rect 11372 23374 11374 23426
rect 11374 23374 11426 23426
rect 11426 23374 11428 23426
rect 11372 23372 11428 23374
rect 11532 23426 11588 23428
rect 11532 23374 11534 23426
rect 11534 23374 11586 23426
rect 11586 23374 11588 23426
rect 11532 23372 11588 23374
rect 11852 23426 11908 23428
rect 11852 23374 11854 23426
rect 11854 23374 11906 23426
rect 11906 23374 11908 23426
rect 11852 23372 11908 23374
rect 12012 23426 12068 23428
rect 12012 23374 12014 23426
rect 12014 23374 12066 23426
rect 12066 23374 12068 23426
rect 12012 23372 12068 23374
rect 12332 23426 12388 23428
rect 12332 23374 12334 23426
rect 12334 23374 12386 23426
rect 12386 23374 12388 23426
rect 12332 23372 12388 23374
rect 8492 23266 8548 23268
rect 8492 23214 8494 23266
rect 8494 23214 8546 23266
rect 8546 23214 8548 23266
rect 8492 23212 8548 23214
rect 8812 23266 8868 23268
rect 8812 23214 8814 23266
rect 8814 23214 8866 23266
rect 8866 23214 8868 23266
rect 8812 23212 8868 23214
rect 8972 23266 9028 23268
rect 8972 23214 8974 23266
rect 8974 23214 9026 23266
rect 9026 23214 9028 23266
rect 8972 23212 9028 23214
rect 9292 23266 9348 23268
rect 9292 23214 9294 23266
rect 9294 23214 9346 23266
rect 9346 23214 9348 23266
rect 9292 23212 9348 23214
rect 9452 23266 9508 23268
rect 9452 23214 9454 23266
rect 9454 23214 9506 23266
rect 9506 23214 9508 23266
rect 9452 23212 9508 23214
rect 9772 23266 9828 23268
rect 9772 23214 9774 23266
rect 9774 23214 9826 23266
rect 9826 23214 9828 23266
rect 9772 23212 9828 23214
rect 10092 23266 10148 23268
rect 10092 23214 10094 23266
rect 10094 23214 10146 23266
rect 10146 23214 10148 23266
rect 10092 23212 10148 23214
rect 10412 23266 10468 23268
rect 10412 23214 10414 23266
rect 10414 23214 10466 23266
rect 10466 23214 10468 23266
rect 10412 23212 10468 23214
rect 10732 23266 10788 23268
rect 10732 23214 10734 23266
rect 10734 23214 10786 23266
rect 10786 23214 10788 23266
rect 10732 23212 10788 23214
rect 11052 23266 11108 23268
rect 11052 23214 11054 23266
rect 11054 23214 11106 23266
rect 11106 23214 11108 23266
rect 11052 23212 11108 23214
rect 11372 23266 11428 23268
rect 11372 23214 11374 23266
rect 11374 23214 11426 23266
rect 11426 23214 11428 23266
rect 11372 23212 11428 23214
rect 11532 23266 11588 23268
rect 11532 23214 11534 23266
rect 11534 23214 11586 23266
rect 11586 23214 11588 23266
rect 11532 23212 11588 23214
rect 11852 23266 11908 23268
rect 11852 23214 11854 23266
rect 11854 23214 11906 23266
rect 11906 23214 11908 23266
rect 11852 23212 11908 23214
rect 12012 23266 12068 23268
rect 12012 23214 12014 23266
rect 12014 23214 12066 23266
rect 12066 23214 12068 23266
rect 12012 23212 12068 23214
rect 12332 23266 12388 23268
rect 12332 23214 12334 23266
rect 12334 23214 12386 23266
rect 12386 23214 12388 23266
rect 12332 23212 12388 23214
rect 8492 23106 8548 23108
rect 8492 23054 8494 23106
rect 8494 23054 8546 23106
rect 8546 23054 8548 23106
rect 8492 23052 8548 23054
rect 8812 23106 8868 23108
rect 8812 23054 8814 23106
rect 8814 23054 8866 23106
rect 8866 23054 8868 23106
rect 8812 23052 8868 23054
rect 8972 23106 9028 23108
rect 8972 23054 8974 23106
rect 8974 23054 9026 23106
rect 9026 23054 9028 23106
rect 8972 23052 9028 23054
rect 9292 23106 9348 23108
rect 9292 23054 9294 23106
rect 9294 23054 9346 23106
rect 9346 23054 9348 23106
rect 9292 23052 9348 23054
rect 9452 23106 9508 23108
rect 9452 23054 9454 23106
rect 9454 23054 9506 23106
rect 9506 23054 9508 23106
rect 9452 23052 9508 23054
rect 9772 23106 9828 23108
rect 9772 23054 9774 23106
rect 9774 23054 9826 23106
rect 9826 23054 9828 23106
rect 9772 23052 9828 23054
rect 10092 23106 10148 23108
rect 10092 23054 10094 23106
rect 10094 23054 10146 23106
rect 10146 23054 10148 23106
rect 10092 23052 10148 23054
rect 10412 23106 10468 23108
rect 10412 23054 10414 23106
rect 10414 23054 10466 23106
rect 10466 23054 10468 23106
rect 10412 23052 10468 23054
rect 10732 23106 10788 23108
rect 10732 23054 10734 23106
rect 10734 23054 10786 23106
rect 10786 23054 10788 23106
rect 10732 23052 10788 23054
rect 11052 23106 11108 23108
rect 11052 23054 11054 23106
rect 11054 23054 11106 23106
rect 11106 23054 11108 23106
rect 11052 23052 11108 23054
rect 11372 23106 11428 23108
rect 11372 23054 11374 23106
rect 11374 23054 11426 23106
rect 11426 23054 11428 23106
rect 11372 23052 11428 23054
rect 11532 23106 11588 23108
rect 11532 23054 11534 23106
rect 11534 23054 11586 23106
rect 11586 23054 11588 23106
rect 11532 23052 11588 23054
rect 11852 23106 11908 23108
rect 11852 23054 11854 23106
rect 11854 23054 11906 23106
rect 11906 23054 11908 23106
rect 11852 23052 11908 23054
rect 12012 23106 12068 23108
rect 12012 23054 12014 23106
rect 12014 23054 12066 23106
rect 12066 23054 12068 23106
rect 12012 23052 12068 23054
rect 12332 23106 12388 23108
rect 12332 23054 12334 23106
rect 12334 23054 12386 23106
rect 12386 23054 12388 23106
rect 12332 23052 12388 23054
rect 8492 22946 8548 22948
rect 8492 22894 8494 22946
rect 8494 22894 8546 22946
rect 8546 22894 8548 22946
rect 8492 22892 8548 22894
rect 8812 22946 8868 22948
rect 8812 22894 8814 22946
rect 8814 22894 8866 22946
rect 8866 22894 8868 22946
rect 8812 22892 8868 22894
rect 8972 22946 9028 22948
rect 8972 22894 8974 22946
rect 8974 22894 9026 22946
rect 9026 22894 9028 22946
rect 8972 22892 9028 22894
rect 9292 22946 9348 22948
rect 9292 22894 9294 22946
rect 9294 22894 9346 22946
rect 9346 22894 9348 22946
rect 9292 22892 9348 22894
rect 9452 22946 9508 22948
rect 9452 22894 9454 22946
rect 9454 22894 9506 22946
rect 9506 22894 9508 22946
rect 9452 22892 9508 22894
rect 9772 22946 9828 22948
rect 9772 22894 9774 22946
rect 9774 22894 9826 22946
rect 9826 22894 9828 22946
rect 9772 22892 9828 22894
rect 10092 22946 10148 22948
rect 10092 22894 10094 22946
rect 10094 22894 10146 22946
rect 10146 22894 10148 22946
rect 10092 22892 10148 22894
rect 10412 22946 10468 22948
rect 10412 22894 10414 22946
rect 10414 22894 10466 22946
rect 10466 22894 10468 22946
rect 10412 22892 10468 22894
rect 10732 22946 10788 22948
rect 10732 22894 10734 22946
rect 10734 22894 10786 22946
rect 10786 22894 10788 22946
rect 10732 22892 10788 22894
rect 11052 22946 11108 22948
rect 11052 22894 11054 22946
rect 11054 22894 11106 22946
rect 11106 22894 11108 22946
rect 11052 22892 11108 22894
rect 11372 22946 11428 22948
rect 11372 22894 11374 22946
rect 11374 22894 11426 22946
rect 11426 22894 11428 22946
rect 11372 22892 11428 22894
rect 11532 22946 11588 22948
rect 11532 22894 11534 22946
rect 11534 22894 11586 22946
rect 11586 22894 11588 22946
rect 11532 22892 11588 22894
rect 11852 22946 11908 22948
rect 11852 22894 11854 22946
rect 11854 22894 11906 22946
rect 11906 22894 11908 22946
rect 11852 22892 11908 22894
rect 12012 22946 12068 22948
rect 12012 22894 12014 22946
rect 12014 22894 12066 22946
rect 12066 22894 12068 22946
rect 12012 22892 12068 22894
rect 12332 22946 12388 22948
rect 12332 22894 12334 22946
rect 12334 22894 12386 22946
rect 12386 22894 12388 22946
rect 12332 22892 12388 22894
rect 8492 22786 8548 22788
rect 8492 22734 8494 22786
rect 8494 22734 8546 22786
rect 8546 22734 8548 22786
rect 8492 22732 8548 22734
rect 8812 22786 8868 22788
rect 8812 22734 8814 22786
rect 8814 22734 8866 22786
rect 8866 22734 8868 22786
rect 8812 22732 8868 22734
rect 8972 22786 9028 22788
rect 8972 22734 8974 22786
rect 8974 22734 9026 22786
rect 9026 22734 9028 22786
rect 8972 22732 9028 22734
rect 9292 22786 9348 22788
rect 9292 22734 9294 22786
rect 9294 22734 9346 22786
rect 9346 22734 9348 22786
rect 9292 22732 9348 22734
rect 9452 22786 9508 22788
rect 9452 22734 9454 22786
rect 9454 22734 9506 22786
rect 9506 22734 9508 22786
rect 9452 22732 9508 22734
rect 9772 22786 9828 22788
rect 9772 22734 9774 22786
rect 9774 22734 9826 22786
rect 9826 22734 9828 22786
rect 9772 22732 9828 22734
rect 10092 22786 10148 22788
rect 10092 22734 10094 22786
rect 10094 22734 10146 22786
rect 10146 22734 10148 22786
rect 10092 22732 10148 22734
rect 10412 22786 10468 22788
rect 10412 22734 10414 22786
rect 10414 22734 10466 22786
rect 10466 22734 10468 22786
rect 10412 22732 10468 22734
rect 10732 22786 10788 22788
rect 10732 22734 10734 22786
rect 10734 22734 10786 22786
rect 10786 22734 10788 22786
rect 10732 22732 10788 22734
rect 11052 22786 11108 22788
rect 11052 22734 11054 22786
rect 11054 22734 11106 22786
rect 11106 22734 11108 22786
rect 11052 22732 11108 22734
rect 11372 22786 11428 22788
rect 11372 22734 11374 22786
rect 11374 22734 11426 22786
rect 11426 22734 11428 22786
rect 11372 22732 11428 22734
rect 11532 22786 11588 22788
rect 11532 22734 11534 22786
rect 11534 22734 11586 22786
rect 11586 22734 11588 22786
rect 11532 22732 11588 22734
rect 11852 22786 11908 22788
rect 11852 22734 11854 22786
rect 11854 22734 11906 22786
rect 11906 22734 11908 22786
rect 11852 22732 11908 22734
rect 12012 22786 12068 22788
rect 12012 22734 12014 22786
rect 12014 22734 12066 22786
rect 12066 22734 12068 22786
rect 12012 22732 12068 22734
rect 12332 22786 12388 22788
rect 12332 22734 12334 22786
rect 12334 22734 12386 22786
rect 12386 22734 12388 22786
rect 12332 22732 12388 22734
rect 8492 22626 8548 22628
rect 8492 22574 8494 22626
rect 8494 22574 8546 22626
rect 8546 22574 8548 22626
rect 8492 22572 8548 22574
rect 8812 22626 8868 22628
rect 8812 22574 8814 22626
rect 8814 22574 8866 22626
rect 8866 22574 8868 22626
rect 8812 22572 8868 22574
rect 8972 22626 9028 22628
rect 8972 22574 8974 22626
rect 8974 22574 9026 22626
rect 9026 22574 9028 22626
rect 8972 22572 9028 22574
rect 9292 22626 9348 22628
rect 9292 22574 9294 22626
rect 9294 22574 9346 22626
rect 9346 22574 9348 22626
rect 9292 22572 9348 22574
rect 9452 22626 9508 22628
rect 9452 22574 9454 22626
rect 9454 22574 9506 22626
rect 9506 22574 9508 22626
rect 9452 22572 9508 22574
rect 9772 22626 9828 22628
rect 9772 22574 9774 22626
rect 9774 22574 9826 22626
rect 9826 22574 9828 22626
rect 9772 22572 9828 22574
rect 10092 22626 10148 22628
rect 10092 22574 10094 22626
rect 10094 22574 10146 22626
rect 10146 22574 10148 22626
rect 10092 22572 10148 22574
rect 10412 22626 10468 22628
rect 10412 22574 10414 22626
rect 10414 22574 10466 22626
rect 10466 22574 10468 22626
rect 10412 22572 10468 22574
rect 10732 22626 10788 22628
rect 10732 22574 10734 22626
rect 10734 22574 10786 22626
rect 10786 22574 10788 22626
rect 10732 22572 10788 22574
rect 11052 22626 11108 22628
rect 11052 22574 11054 22626
rect 11054 22574 11106 22626
rect 11106 22574 11108 22626
rect 11052 22572 11108 22574
rect 11372 22626 11428 22628
rect 11372 22574 11374 22626
rect 11374 22574 11426 22626
rect 11426 22574 11428 22626
rect 11372 22572 11428 22574
rect 11532 22626 11588 22628
rect 11532 22574 11534 22626
rect 11534 22574 11586 22626
rect 11586 22574 11588 22626
rect 11532 22572 11588 22574
rect 11852 22626 11908 22628
rect 11852 22574 11854 22626
rect 11854 22574 11906 22626
rect 11906 22574 11908 22626
rect 11852 22572 11908 22574
rect 12012 22626 12068 22628
rect 12012 22574 12014 22626
rect 12014 22574 12066 22626
rect 12066 22574 12068 22626
rect 12012 22572 12068 22574
rect 12332 22626 12388 22628
rect 12332 22574 12334 22626
rect 12334 22574 12386 22626
rect 12386 22574 12388 22626
rect 12332 22572 12388 22574
rect 8492 22466 8548 22468
rect 8492 22414 8494 22466
rect 8494 22414 8546 22466
rect 8546 22414 8548 22466
rect 8492 22412 8548 22414
rect 8812 22466 8868 22468
rect 8812 22414 8814 22466
rect 8814 22414 8866 22466
rect 8866 22414 8868 22466
rect 8812 22412 8868 22414
rect 8972 22466 9028 22468
rect 8972 22414 8974 22466
rect 8974 22414 9026 22466
rect 9026 22414 9028 22466
rect 8972 22412 9028 22414
rect 9292 22466 9348 22468
rect 9292 22414 9294 22466
rect 9294 22414 9346 22466
rect 9346 22414 9348 22466
rect 9292 22412 9348 22414
rect 9452 22466 9508 22468
rect 9452 22414 9454 22466
rect 9454 22414 9506 22466
rect 9506 22414 9508 22466
rect 9452 22412 9508 22414
rect 9772 22466 9828 22468
rect 9772 22414 9774 22466
rect 9774 22414 9826 22466
rect 9826 22414 9828 22466
rect 9772 22412 9828 22414
rect 10092 22466 10148 22468
rect 10092 22414 10094 22466
rect 10094 22414 10146 22466
rect 10146 22414 10148 22466
rect 10092 22412 10148 22414
rect 10412 22466 10468 22468
rect 10412 22414 10414 22466
rect 10414 22414 10466 22466
rect 10466 22414 10468 22466
rect 10412 22412 10468 22414
rect 10732 22466 10788 22468
rect 10732 22414 10734 22466
rect 10734 22414 10786 22466
rect 10786 22414 10788 22466
rect 10732 22412 10788 22414
rect 11052 22466 11108 22468
rect 11052 22414 11054 22466
rect 11054 22414 11106 22466
rect 11106 22414 11108 22466
rect 11052 22412 11108 22414
rect 11372 22466 11428 22468
rect 11372 22414 11374 22466
rect 11374 22414 11426 22466
rect 11426 22414 11428 22466
rect 11372 22412 11428 22414
rect 11532 22466 11588 22468
rect 11532 22414 11534 22466
rect 11534 22414 11586 22466
rect 11586 22414 11588 22466
rect 11532 22412 11588 22414
rect 11852 22466 11908 22468
rect 11852 22414 11854 22466
rect 11854 22414 11906 22466
rect 11906 22414 11908 22466
rect 11852 22412 11908 22414
rect 12012 22466 12068 22468
rect 12012 22414 12014 22466
rect 12014 22414 12066 22466
rect 12066 22414 12068 22466
rect 12012 22412 12068 22414
rect 12332 22466 12388 22468
rect 12332 22414 12334 22466
rect 12334 22414 12386 22466
rect 12386 22414 12388 22466
rect 12332 22412 12388 22414
rect 8492 22306 8548 22308
rect 8492 22254 8494 22306
rect 8494 22254 8546 22306
rect 8546 22254 8548 22306
rect 8492 22252 8548 22254
rect 8812 22306 8868 22308
rect 8812 22254 8814 22306
rect 8814 22254 8866 22306
rect 8866 22254 8868 22306
rect 8812 22252 8868 22254
rect 8972 22306 9028 22308
rect 8972 22254 8974 22306
rect 8974 22254 9026 22306
rect 9026 22254 9028 22306
rect 8972 22252 9028 22254
rect 9292 22306 9348 22308
rect 9292 22254 9294 22306
rect 9294 22254 9346 22306
rect 9346 22254 9348 22306
rect 9292 22252 9348 22254
rect 9452 22306 9508 22308
rect 9452 22254 9454 22306
rect 9454 22254 9506 22306
rect 9506 22254 9508 22306
rect 9452 22252 9508 22254
rect 9772 22306 9828 22308
rect 9772 22254 9774 22306
rect 9774 22254 9826 22306
rect 9826 22254 9828 22306
rect 9772 22252 9828 22254
rect 10092 22306 10148 22308
rect 10092 22254 10094 22306
rect 10094 22254 10146 22306
rect 10146 22254 10148 22306
rect 10092 22252 10148 22254
rect 10412 22306 10468 22308
rect 10412 22254 10414 22306
rect 10414 22254 10466 22306
rect 10466 22254 10468 22306
rect 10412 22252 10468 22254
rect 10732 22306 10788 22308
rect 10732 22254 10734 22306
rect 10734 22254 10786 22306
rect 10786 22254 10788 22306
rect 10732 22252 10788 22254
rect 11052 22306 11108 22308
rect 11052 22254 11054 22306
rect 11054 22254 11106 22306
rect 11106 22254 11108 22306
rect 11052 22252 11108 22254
rect 11372 22306 11428 22308
rect 11372 22254 11374 22306
rect 11374 22254 11426 22306
rect 11426 22254 11428 22306
rect 11372 22252 11428 22254
rect 11532 22306 11588 22308
rect 11532 22254 11534 22306
rect 11534 22254 11586 22306
rect 11586 22254 11588 22306
rect 11532 22252 11588 22254
rect 11852 22306 11908 22308
rect 11852 22254 11854 22306
rect 11854 22254 11906 22306
rect 11906 22254 11908 22306
rect 11852 22252 11908 22254
rect 12012 22306 12068 22308
rect 12012 22254 12014 22306
rect 12014 22254 12066 22306
rect 12066 22254 12068 22306
rect 12012 22252 12068 22254
rect 12332 22306 12388 22308
rect 12332 22254 12334 22306
rect 12334 22254 12386 22306
rect 12386 22254 12388 22306
rect 12332 22252 12388 22254
rect 8492 22146 8548 22148
rect 8492 22094 8494 22146
rect 8494 22094 8546 22146
rect 8546 22094 8548 22146
rect 8492 22092 8548 22094
rect 8812 22146 8868 22148
rect 8812 22094 8814 22146
rect 8814 22094 8866 22146
rect 8866 22094 8868 22146
rect 8812 22092 8868 22094
rect 8972 22146 9028 22148
rect 8972 22094 8974 22146
rect 8974 22094 9026 22146
rect 9026 22094 9028 22146
rect 8972 22092 9028 22094
rect 9292 22146 9348 22148
rect 9292 22094 9294 22146
rect 9294 22094 9346 22146
rect 9346 22094 9348 22146
rect 9292 22092 9348 22094
rect 9452 22146 9508 22148
rect 9452 22094 9454 22146
rect 9454 22094 9506 22146
rect 9506 22094 9508 22146
rect 9452 22092 9508 22094
rect 9772 22146 9828 22148
rect 9772 22094 9774 22146
rect 9774 22094 9826 22146
rect 9826 22094 9828 22146
rect 9772 22092 9828 22094
rect 10092 22146 10148 22148
rect 10092 22094 10094 22146
rect 10094 22094 10146 22146
rect 10146 22094 10148 22146
rect 10092 22092 10148 22094
rect 10412 22146 10468 22148
rect 10412 22094 10414 22146
rect 10414 22094 10466 22146
rect 10466 22094 10468 22146
rect 10412 22092 10468 22094
rect 10732 22146 10788 22148
rect 10732 22094 10734 22146
rect 10734 22094 10786 22146
rect 10786 22094 10788 22146
rect 10732 22092 10788 22094
rect 11052 22146 11108 22148
rect 11052 22094 11054 22146
rect 11054 22094 11106 22146
rect 11106 22094 11108 22146
rect 11052 22092 11108 22094
rect 11372 22146 11428 22148
rect 11372 22094 11374 22146
rect 11374 22094 11426 22146
rect 11426 22094 11428 22146
rect 11372 22092 11428 22094
rect 11532 22146 11588 22148
rect 11532 22094 11534 22146
rect 11534 22094 11586 22146
rect 11586 22094 11588 22146
rect 11532 22092 11588 22094
rect 11852 22146 11908 22148
rect 11852 22094 11854 22146
rect 11854 22094 11906 22146
rect 11906 22094 11908 22146
rect 11852 22092 11908 22094
rect 12012 22146 12068 22148
rect 12012 22094 12014 22146
rect 12014 22094 12066 22146
rect 12066 22094 12068 22146
rect 12012 22092 12068 22094
rect 12332 22146 12388 22148
rect 12332 22094 12334 22146
rect 12334 22094 12386 22146
rect 12386 22094 12388 22146
rect 12332 22092 12388 22094
rect 9132 21932 9188 21988
rect 8492 21826 8548 21828
rect 8492 21774 8494 21826
rect 8494 21774 8546 21826
rect 8546 21774 8548 21826
rect 8492 21772 8548 21774
rect 8812 21826 8868 21828
rect 8812 21774 8814 21826
rect 8814 21774 8866 21826
rect 8866 21774 8868 21826
rect 8812 21772 8868 21774
rect 8972 21826 9028 21828
rect 8972 21774 8974 21826
rect 8974 21774 9026 21826
rect 9026 21774 9028 21826
rect 8972 21772 9028 21774
rect 9292 21826 9348 21828
rect 9292 21774 9294 21826
rect 9294 21774 9346 21826
rect 9346 21774 9348 21826
rect 9292 21772 9348 21774
rect 9452 21826 9508 21828
rect 9452 21774 9454 21826
rect 9454 21774 9506 21826
rect 9506 21774 9508 21826
rect 9452 21772 9508 21774
rect 9772 21826 9828 21828
rect 9772 21774 9774 21826
rect 9774 21774 9826 21826
rect 9826 21774 9828 21826
rect 9772 21772 9828 21774
rect 10092 21826 10148 21828
rect 10092 21774 10094 21826
rect 10094 21774 10146 21826
rect 10146 21774 10148 21826
rect 10092 21772 10148 21774
rect 10412 21826 10468 21828
rect 10412 21774 10414 21826
rect 10414 21774 10466 21826
rect 10466 21774 10468 21826
rect 10412 21772 10468 21774
rect 10732 21826 10788 21828
rect 10732 21774 10734 21826
rect 10734 21774 10786 21826
rect 10786 21774 10788 21826
rect 10732 21772 10788 21774
rect 11052 21826 11108 21828
rect 11052 21774 11054 21826
rect 11054 21774 11106 21826
rect 11106 21774 11108 21826
rect 11052 21772 11108 21774
rect 11372 21826 11428 21828
rect 11372 21774 11374 21826
rect 11374 21774 11426 21826
rect 11426 21774 11428 21826
rect 11372 21772 11428 21774
rect 11532 21826 11588 21828
rect 11532 21774 11534 21826
rect 11534 21774 11586 21826
rect 11586 21774 11588 21826
rect 11532 21772 11588 21774
rect 11852 21826 11908 21828
rect 11852 21774 11854 21826
rect 11854 21774 11906 21826
rect 11906 21774 11908 21826
rect 11852 21772 11908 21774
rect 12012 21826 12068 21828
rect 12012 21774 12014 21826
rect 12014 21774 12066 21826
rect 12066 21774 12068 21826
rect 12012 21772 12068 21774
rect 12332 21826 12388 21828
rect 12332 21774 12334 21826
rect 12334 21774 12386 21826
rect 12386 21774 12388 21826
rect 12332 21772 12388 21774
rect 8492 21666 8548 21668
rect 8492 21614 8494 21666
rect 8494 21614 8546 21666
rect 8546 21614 8548 21666
rect 8492 21612 8548 21614
rect 8812 21666 8868 21668
rect 8812 21614 8814 21666
rect 8814 21614 8866 21666
rect 8866 21614 8868 21666
rect 8812 21612 8868 21614
rect 8972 21666 9028 21668
rect 8972 21614 8974 21666
rect 8974 21614 9026 21666
rect 9026 21614 9028 21666
rect 8972 21612 9028 21614
rect 9292 21666 9348 21668
rect 9292 21614 9294 21666
rect 9294 21614 9346 21666
rect 9346 21614 9348 21666
rect 9292 21612 9348 21614
rect 9452 21666 9508 21668
rect 9452 21614 9454 21666
rect 9454 21614 9506 21666
rect 9506 21614 9508 21666
rect 9452 21612 9508 21614
rect 9772 21666 9828 21668
rect 9772 21614 9774 21666
rect 9774 21614 9826 21666
rect 9826 21614 9828 21666
rect 9772 21612 9828 21614
rect 10092 21666 10148 21668
rect 10092 21614 10094 21666
rect 10094 21614 10146 21666
rect 10146 21614 10148 21666
rect 10092 21612 10148 21614
rect 10412 21666 10468 21668
rect 10412 21614 10414 21666
rect 10414 21614 10466 21666
rect 10466 21614 10468 21666
rect 10412 21612 10468 21614
rect 10732 21666 10788 21668
rect 10732 21614 10734 21666
rect 10734 21614 10786 21666
rect 10786 21614 10788 21666
rect 10732 21612 10788 21614
rect 11052 21666 11108 21668
rect 11052 21614 11054 21666
rect 11054 21614 11106 21666
rect 11106 21614 11108 21666
rect 11052 21612 11108 21614
rect 11372 21666 11428 21668
rect 11372 21614 11374 21666
rect 11374 21614 11426 21666
rect 11426 21614 11428 21666
rect 11372 21612 11428 21614
rect 11532 21666 11588 21668
rect 11532 21614 11534 21666
rect 11534 21614 11586 21666
rect 11586 21614 11588 21666
rect 11532 21612 11588 21614
rect 11852 21666 11908 21668
rect 11852 21614 11854 21666
rect 11854 21614 11906 21666
rect 11906 21614 11908 21666
rect 11852 21612 11908 21614
rect 12012 21666 12068 21668
rect 12012 21614 12014 21666
rect 12014 21614 12066 21666
rect 12066 21614 12068 21666
rect 12012 21612 12068 21614
rect 12332 21666 12388 21668
rect 12332 21614 12334 21666
rect 12334 21614 12386 21666
rect 12386 21614 12388 21666
rect 12332 21612 12388 21614
rect 8492 21506 8548 21508
rect 8492 21454 8494 21506
rect 8494 21454 8546 21506
rect 8546 21454 8548 21506
rect 8492 21452 8548 21454
rect 8812 21506 8868 21508
rect 8812 21454 8814 21506
rect 8814 21454 8866 21506
rect 8866 21454 8868 21506
rect 8812 21452 8868 21454
rect 8972 21506 9028 21508
rect 8972 21454 8974 21506
rect 8974 21454 9026 21506
rect 9026 21454 9028 21506
rect 8972 21452 9028 21454
rect 9292 21506 9348 21508
rect 9292 21454 9294 21506
rect 9294 21454 9346 21506
rect 9346 21454 9348 21506
rect 9292 21452 9348 21454
rect 9452 21506 9508 21508
rect 9452 21454 9454 21506
rect 9454 21454 9506 21506
rect 9506 21454 9508 21506
rect 9452 21452 9508 21454
rect 9772 21506 9828 21508
rect 9772 21454 9774 21506
rect 9774 21454 9826 21506
rect 9826 21454 9828 21506
rect 9772 21452 9828 21454
rect 10092 21506 10148 21508
rect 10092 21454 10094 21506
rect 10094 21454 10146 21506
rect 10146 21454 10148 21506
rect 10092 21452 10148 21454
rect 10412 21506 10468 21508
rect 10412 21454 10414 21506
rect 10414 21454 10466 21506
rect 10466 21454 10468 21506
rect 10412 21452 10468 21454
rect 10732 21506 10788 21508
rect 10732 21454 10734 21506
rect 10734 21454 10786 21506
rect 10786 21454 10788 21506
rect 10732 21452 10788 21454
rect 11052 21506 11108 21508
rect 11052 21454 11054 21506
rect 11054 21454 11106 21506
rect 11106 21454 11108 21506
rect 11052 21452 11108 21454
rect 11372 21506 11428 21508
rect 11372 21454 11374 21506
rect 11374 21454 11426 21506
rect 11426 21454 11428 21506
rect 11372 21452 11428 21454
rect 11532 21506 11588 21508
rect 11532 21454 11534 21506
rect 11534 21454 11586 21506
rect 11586 21454 11588 21506
rect 11532 21452 11588 21454
rect 11852 21506 11908 21508
rect 11852 21454 11854 21506
rect 11854 21454 11906 21506
rect 11906 21454 11908 21506
rect 11852 21452 11908 21454
rect 12012 21506 12068 21508
rect 12012 21454 12014 21506
rect 12014 21454 12066 21506
rect 12066 21454 12068 21506
rect 12012 21452 12068 21454
rect 12332 21506 12388 21508
rect 12332 21454 12334 21506
rect 12334 21454 12386 21506
rect 12386 21454 12388 21506
rect 12332 21452 12388 21454
rect 8492 21346 8548 21348
rect 8492 21294 8494 21346
rect 8494 21294 8546 21346
rect 8546 21294 8548 21346
rect 8492 21292 8548 21294
rect 8812 21346 8868 21348
rect 8812 21294 8814 21346
rect 8814 21294 8866 21346
rect 8866 21294 8868 21346
rect 8812 21292 8868 21294
rect 8972 21346 9028 21348
rect 8972 21294 8974 21346
rect 8974 21294 9026 21346
rect 9026 21294 9028 21346
rect 8972 21292 9028 21294
rect 9292 21346 9348 21348
rect 9292 21294 9294 21346
rect 9294 21294 9346 21346
rect 9346 21294 9348 21346
rect 9292 21292 9348 21294
rect 9452 21346 9508 21348
rect 9452 21294 9454 21346
rect 9454 21294 9506 21346
rect 9506 21294 9508 21346
rect 9452 21292 9508 21294
rect 9772 21346 9828 21348
rect 9772 21294 9774 21346
rect 9774 21294 9826 21346
rect 9826 21294 9828 21346
rect 9772 21292 9828 21294
rect 10092 21346 10148 21348
rect 10092 21294 10094 21346
rect 10094 21294 10146 21346
rect 10146 21294 10148 21346
rect 10092 21292 10148 21294
rect 10412 21346 10468 21348
rect 10412 21294 10414 21346
rect 10414 21294 10466 21346
rect 10466 21294 10468 21346
rect 10412 21292 10468 21294
rect 10732 21346 10788 21348
rect 10732 21294 10734 21346
rect 10734 21294 10786 21346
rect 10786 21294 10788 21346
rect 10732 21292 10788 21294
rect 11052 21346 11108 21348
rect 11052 21294 11054 21346
rect 11054 21294 11106 21346
rect 11106 21294 11108 21346
rect 11052 21292 11108 21294
rect 11372 21346 11428 21348
rect 11372 21294 11374 21346
rect 11374 21294 11426 21346
rect 11426 21294 11428 21346
rect 11372 21292 11428 21294
rect 11532 21346 11588 21348
rect 11532 21294 11534 21346
rect 11534 21294 11586 21346
rect 11586 21294 11588 21346
rect 11532 21292 11588 21294
rect 11852 21346 11908 21348
rect 11852 21294 11854 21346
rect 11854 21294 11906 21346
rect 11906 21294 11908 21346
rect 11852 21292 11908 21294
rect 12012 21346 12068 21348
rect 12012 21294 12014 21346
rect 12014 21294 12066 21346
rect 12066 21294 12068 21346
rect 12012 21292 12068 21294
rect 12332 21346 12388 21348
rect 12332 21294 12334 21346
rect 12334 21294 12386 21346
rect 12386 21294 12388 21346
rect 12332 21292 12388 21294
rect 8492 21186 8548 21188
rect 8492 21134 8494 21186
rect 8494 21134 8546 21186
rect 8546 21134 8548 21186
rect 8492 21132 8548 21134
rect 8812 21186 8868 21188
rect 8812 21134 8814 21186
rect 8814 21134 8866 21186
rect 8866 21134 8868 21186
rect 8812 21132 8868 21134
rect 8972 21186 9028 21188
rect 8972 21134 8974 21186
rect 8974 21134 9026 21186
rect 9026 21134 9028 21186
rect 8972 21132 9028 21134
rect 9292 21186 9348 21188
rect 9292 21134 9294 21186
rect 9294 21134 9346 21186
rect 9346 21134 9348 21186
rect 9292 21132 9348 21134
rect 9452 21186 9508 21188
rect 9452 21134 9454 21186
rect 9454 21134 9506 21186
rect 9506 21134 9508 21186
rect 9452 21132 9508 21134
rect 9772 21186 9828 21188
rect 9772 21134 9774 21186
rect 9774 21134 9826 21186
rect 9826 21134 9828 21186
rect 9772 21132 9828 21134
rect 10092 21186 10148 21188
rect 10092 21134 10094 21186
rect 10094 21134 10146 21186
rect 10146 21134 10148 21186
rect 10092 21132 10148 21134
rect 10412 21186 10468 21188
rect 10412 21134 10414 21186
rect 10414 21134 10466 21186
rect 10466 21134 10468 21186
rect 10412 21132 10468 21134
rect 10732 21186 10788 21188
rect 10732 21134 10734 21186
rect 10734 21134 10786 21186
rect 10786 21134 10788 21186
rect 10732 21132 10788 21134
rect 11052 21186 11108 21188
rect 11052 21134 11054 21186
rect 11054 21134 11106 21186
rect 11106 21134 11108 21186
rect 11052 21132 11108 21134
rect 11372 21186 11428 21188
rect 11372 21134 11374 21186
rect 11374 21134 11426 21186
rect 11426 21134 11428 21186
rect 11372 21132 11428 21134
rect 11532 21186 11588 21188
rect 11532 21134 11534 21186
rect 11534 21134 11586 21186
rect 11586 21134 11588 21186
rect 11532 21132 11588 21134
rect 11852 21186 11908 21188
rect 11852 21134 11854 21186
rect 11854 21134 11906 21186
rect 11906 21134 11908 21186
rect 11852 21132 11908 21134
rect 12012 21186 12068 21188
rect 12012 21134 12014 21186
rect 12014 21134 12066 21186
rect 12066 21134 12068 21186
rect 12012 21132 12068 21134
rect 12332 21186 12388 21188
rect 12332 21134 12334 21186
rect 12334 21134 12386 21186
rect 12386 21134 12388 21186
rect 12332 21132 12388 21134
rect 8492 21026 8548 21028
rect 8492 20974 8494 21026
rect 8494 20974 8546 21026
rect 8546 20974 8548 21026
rect 8492 20972 8548 20974
rect 8812 21026 8868 21028
rect 8812 20974 8814 21026
rect 8814 20974 8866 21026
rect 8866 20974 8868 21026
rect 8812 20972 8868 20974
rect 8972 21026 9028 21028
rect 8972 20974 8974 21026
rect 8974 20974 9026 21026
rect 9026 20974 9028 21026
rect 8972 20972 9028 20974
rect 9292 21026 9348 21028
rect 9292 20974 9294 21026
rect 9294 20974 9346 21026
rect 9346 20974 9348 21026
rect 9292 20972 9348 20974
rect 9452 21026 9508 21028
rect 9452 20974 9454 21026
rect 9454 20974 9506 21026
rect 9506 20974 9508 21026
rect 9452 20972 9508 20974
rect 9772 21026 9828 21028
rect 9772 20974 9774 21026
rect 9774 20974 9826 21026
rect 9826 20974 9828 21026
rect 9772 20972 9828 20974
rect 10092 21026 10148 21028
rect 10092 20974 10094 21026
rect 10094 20974 10146 21026
rect 10146 20974 10148 21026
rect 10092 20972 10148 20974
rect 10412 21026 10468 21028
rect 10412 20974 10414 21026
rect 10414 20974 10466 21026
rect 10466 20974 10468 21026
rect 10412 20972 10468 20974
rect 10732 21026 10788 21028
rect 10732 20974 10734 21026
rect 10734 20974 10786 21026
rect 10786 20974 10788 21026
rect 10732 20972 10788 20974
rect 11052 21026 11108 21028
rect 11052 20974 11054 21026
rect 11054 20974 11106 21026
rect 11106 20974 11108 21026
rect 11052 20972 11108 20974
rect 11372 21026 11428 21028
rect 11372 20974 11374 21026
rect 11374 20974 11426 21026
rect 11426 20974 11428 21026
rect 11372 20972 11428 20974
rect 11532 21026 11588 21028
rect 11532 20974 11534 21026
rect 11534 20974 11586 21026
rect 11586 20974 11588 21026
rect 11532 20972 11588 20974
rect 11852 21026 11908 21028
rect 11852 20974 11854 21026
rect 11854 20974 11906 21026
rect 11906 20974 11908 21026
rect 11852 20972 11908 20974
rect 12012 21026 12068 21028
rect 12012 20974 12014 21026
rect 12014 20974 12066 21026
rect 12066 20974 12068 21026
rect 12012 20972 12068 20974
rect 12332 21026 12388 21028
rect 12332 20974 12334 21026
rect 12334 20974 12386 21026
rect 12386 20974 12388 21026
rect 12332 20972 12388 20974
rect 8492 20866 8548 20868
rect 8492 20814 8494 20866
rect 8494 20814 8546 20866
rect 8546 20814 8548 20866
rect 8492 20812 8548 20814
rect 8812 20866 8868 20868
rect 8812 20814 8814 20866
rect 8814 20814 8866 20866
rect 8866 20814 8868 20866
rect 8812 20812 8868 20814
rect 8972 20866 9028 20868
rect 8972 20814 8974 20866
rect 8974 20814 9026 20866
rect 9026 20814 9028 20866
rect 8972 20812 9028 20814
rect 9292 20866 9348 20868
rect 9292 20814 9294 20866
rect 9294 20814 9346 20866
rect 9346 20814 9348 20866
rect 9292 20812 9348 20814
rect 9452 20866 9508 20868
rect 9452 20814 9454 20866
rect 9454 20814 9506 20866
rect 9506 20814 9508 20866
rect 9452 20812 9508 20814
rect 9772 20866 9828 20868
rect 9772 20814 9774 20866
rect 9774 20814 9826 20866
rect 9826 20814 9828 20866
rect 9772 20812 9828 20814
rect 10092 20866 10148 20868
rect 10092 20814 10094 20866
rect 10094 20814 10146 20866
rect 10146 20814 10148 20866
rect 10092 20812 10148 20814
rect 10412 20866 10468 20868
rect 10412 20814 10414 20866
rect 10414 20814 10466 20866
rect 10466 20814 10468 20866
rect 10412 20812 10468 20814
rect 10732 20866 10788 20868
rect 10732 20814 10734 20866
rect 10734 20814 10786 20866
rect 10786 20814 10788 20866
rect 10732 20812 10788 20814
rect 11052 20866 11108 20868
rect 11052 20814 11054 20866
rect 11054 20814 11106 20866
rect 11106 20814 11108 20866
rect 11052 20812 11108 20814
rect 11372 20866 11428 20868
rect 11372 20814 11374 20866
rect 11374 20814 11426 20866
rect 11426 20814 11428 20866
rect 11372 20812 11428 20814
rect 11532 20866 11588 20868
rect 11532 20814 11534 20866
rect 11534 20814 11586 20866
rect 11586 20814 11588 20866
rect 11532 20812 11588 20814
rect 11852 20866 11908 20868
rect 11852 20814 11854 20866
rect 11854 20814 11906 20866
rect 11906 20814 11908 20866
rect 11852 20812 11908 20814
rect 12012 20866 12068 20868
rect 12012 20814 12014 20866
rect 12014 20814 12066 20866
rect 12066 20814 12068 20866
rect 12012 20812 12068 20814
rect 12332 20866 12388 20868
rect 12332 20814 12334 20866
rect 12334 20814 12386 20866
rect 12386 20814 12388 20866
rect 12332 20812 12388 20814
rect 8492 20706 8548 20708
rect 8492 20654 8494 20706
rect 8494 20654 8546 20706
rect 8546 20654 8548 20706
rect 8492 20652 8548 20654
rect 8812 20706 8868 20708
rect 8812 20654 8814 20706
rect 8814 20654 8866 20706
rect 8866 20654 8868 20706
rect 8812 20652 8868 20654
rect 8972 20706 9028 20708
rect 8972 20654 8974 20706
rect 8974 20654 9026 20706
rect 9026 20654 9028 20706
rect 8972 20652 9028 20654
rect 9292 20706 9348 20708
rect 9292 20654 9294 20706
rect 9294 20654 9346 20706
rect 9346 20654 9348 20706
rect 9292 20652 9348 20654
rect 9452 20706 9508 20708
rect 9452 20654 9454 20706
rect 9454 20654 9506 20706
rect 9506 20654 9508 20706
rect 9452 20652 9508 20654
rect 9772 20706 9828 20708
rect 9772 20654 9774 20706
rect 9774 20654 9826 20706
rect 9826 20654 9828 20706
rect 9772 20652 9828 20654
rect 10092 20706 10148 20708
rect 10092 20654 10094 20706
rect 10094 20654 10146 20706
rect 10146 20654 10148 20706
rect 10092 20652 10148 20654
rect 10412 20706 10468 20708
rect 10412 20654 10414 20706
rect 10414 20654 10466 20706
rect 10466 20654 10468 20706
rect 10412 20652 10468 20654
rect 10732 20706 10788 20708
rect 10732 20654 10734 20706
rect 10734 20654 10786 20706
rect 10786 20654 10788 20706
rect 10732 20652 10788 20654
rect 11052 20706 11108 20708
rect 11052 20654 11054 20706
rect 11054 20654 11106 20706
rect 11106 20654 11108 20706
rect 11052 20652 11108 20654
rect 11372 20706 11428 20708
rect 11372 20654 11374 20706
rect 11374 20654 11426 20706
rect 11426 20654 11428 20706
rect 11372 20652 11428 20654
rect 11532 20706 11588 20708
rect 11532 20654 11534 20706
rect 11534 20654 11586 20706
rect 11586 20654 11588 20706
rect 11532 20652 11588 20654
rect 11852 20706 11908 20708
rect 11852 20654 11854 20706
rect 11854 20654 11906 20706
rect 11906 20654 11908 20706
rect 11852 20652 11908 20654
rect 12012 20706 12068 20708
rect 12012 20654 12014 20706
rect 12014 20654 12066 20706
rect 12066 20654 12068 20706
rect 12012 20652 12068 20654
rect 12332 20706 12388 20708
rect 12332 20654 12334 20706
rect 12334 20654 12386 20706
rect 12386 20654 12388 20706
rect 12332 20652 12388 20654
rect 10252 20412 10308 20468
rect 10252 20092 10308 20148
rect 8492 19906 8548 19908
rect 8492 19854 8494 19906
rect 8494 19854 8546 19906
rect 8546 19854 8548 19906
rect 8492 19852 8548 19854
rect 8812 19906 8868 19908
rect 8812 19854 8814 19906
rect 8814 19854 8866 19906
rect 8866 19854 8868 19906
rect 8812 19852 8868 19854
rect 8972 19906 9028 19908
rect 8972 19854 8974 19906
rect 8974 19854 9026 19906
rect 9026 19854 9028 19906
rect 8972 19852 9028 19854
rect 9292 19906 9348 19908
rect 9292 19854 9294 19906
rect 9294 19854 9346 19906
rect 9346 19854 9348 19906
rect 9292 19852 9348 19854
rect 9452 19906 9508 19908
rect 9452 19854 9454 19906
rect 9454 19854 9506 19906
rect 9506 19854 9508 19906
rect 9452 19852 9508 19854
rect 9772 19906 9828 19908
rect 9772 19854 9774 19906
rect 9774 19854 9826 19906
rect 9826 19854 9828 19906
rect 9772 19852 9828 19854
rect 10092 19906 10148 19908
rect 10092 19854 10094 19906
rect 10094 19854 10146 19906
rect 10146 19854 10148 19906
rect 10092 19852 10148 19854
rect 10412 19906 10468 19908
rect 10412 19854 10414 19906
rect 10414 19854 10466 19906
rect 10466 19854 10468 19906
rect 10412 19852 10468 19854
rect 10732 19906 10788 19908
rect 10732 19854 10734 19906
rect 10734 19854 10786 19906
rect 10786 19854 10788 19906
rect 10732 19852 10788 19854
rect 11052 19906 11108 19908
rect 11052 19854 11054 19906
rect 11054 19854 11106 19906
rect 11106 19854 11108 19906
rect 11052 19852 11108 19854
rect 11372 19906 11428 19908
rect 11372 19854 11374 19906
rect 11374 19854 11426 19906
rect 11426 19854 11428 19906
rect 11372 19852 11428 19854
rect 11532 19906 11588 19908
rect 11532 19854 11534 19906
rect 11534 19854 11586 19906
rect 11586 19854 11588 19906
rect 11532 19852 11588 19854
rect 11852 19906 11908 19908
rect 11852 19854 11854 19906
rect 11854 19854 11906 19906
rect 11906 19854 11908 19906
rect 11852 19852 11908 19854
rect 12012 19906 12068 19908
rect 12012 19854 12014 19906
rect 12014 19854 12066 19906
rect 12066 19854 12068 19906
rect 12012 19852 12068 19854
rect 12332 19906 12388 19908
rect 12332 19854 12334 19906
rect 12334 19854 12386 19906
rect 12386 19854 12388 19906
rect 12332 19852 12388 19854
rect 8492 19746 8548 19748
rect 8492 19694 8494 19746
rect 8494 19694 8546 19746
rect 8546 19694 8548 19746
rect 8492 19692 8548 19694
rect 8812 19746 8868 19748
rect 8812 19694 8814 19746
rect 8814 19694 8866 19746
rect 8866 19694 8868 19746
rect 8812 19692 8868 19694
rect 8972 19746 9028 19748
rect 8972 19694 8974 19746
rect 8974 19694 9026 19746
rect 9026 19694 9028 19746
rect 8972 19692 9028 19694
rect 9292 19746 9348 19748
rect 9292 19694 9294 19746
rect 9294 19694 9346 19746
rect 9346 19694 9348 19746
rect 9292 19692 9348 19694
rect 9452 19746 9508 19748
rect 9452 19694 9454 19746
rect 9454 19694 9506 19746
rect 9506 19694 9508 19746
rect 9452 19692 9508 19694
rect 9772 19746 9828 19748
rect 9772 19694 9774 19746
rect 9774 19694 9826 19746
rect 9826 19694 9828 19746
rect 9772 19692 9828 19694
rect 10092 19746 10148 19748
rect 10092 19694 10094 19746
rect 10094 19694 10146 19746
rect 10146 19694 10148 19746
rect 10092 19692 10148 19694
rect 10412 19746 10468 19748
rect 10412 19694 10414 19746
rect 10414 19694 10466 19746
rect 10466 19694 10468 19746
rect 10412 19692 10468 19694
rect 10732 19746 10788 19748
rect 10732 19694 10734 19746
rect 10734 19694 10786 19746
rect 10786 19694 10788 19746
rect 10732 19692 10788 19694
rect 11052 19746 11108 19748
rect 11052 19694 11054 19746
rect 11054 19694 11106 19746
rect 11106 19694 11108 19746
rect 11052 19692 11108 19694
rect 11372 19746 11428 19748
rect 11372 19694 11374 19746
rect 11374 19694 11426 19746
rect 11426 19694 11428 19746
rect 11372 19692 11428 19694
rect 11532 19746 11588 19748
rect 11532 19694 11534 19746
rect 11534 19694 11586 19746
rect 11586 19694 11588 19746
rect 11532 19692 11588 19694
rect 11852 19746 11908 19748
rect 11852 19694 11854 19746
rect 11854 19694 11906 19746
rect 11906 19694 11908 19746
rect 11852 19692 11908 19694
rect 12012 19746 12068 19748
rect 12012 19694 12014 19746
rect 12014 19694 12066 19746
rect 12066 19694 12068 19746
rect 12012 19692 12068 19694
rect 12332 19746 12388 19748
rect 12332 19694 12334 19746
rect 12334 19694 12386 19746
rect 12386 19694 12388 19746
rect 12332 19692 12388 19694
rect 8492 19586 8548 19588
rect 8492 19534 8494 19586
rect 8494 19534 8546 19586
rect 8546 19534 8548 19586
rect 8492 19532 8548 19534
rect 8812 19586 8868 19588
rect 8812 19534 8814 19586
rect 8814 19534 8866 19586
rect 8866 19534 8868 19586
rect 8812 19532 8868 19534
rect 8972 19586 9028 19588
rect 8972 19534 8974 19586
rect 8974 19534 9026 19586
rect 9026 19534 9028 19586
rect 8972 19532 9028 19534
rect 9292 19586 9348 19588
rect 9292 19534 9294 19586
rect 9294 19534 9346 19586
rect 9346 19534 9348 19586
rect 9292 19532 9348 19534
rect 9452 19586 9508 19588
rect 9452 19534 9454 19586
rect 9454 19534 9506 19586
rect 9506 19534 9508 19586
rect 9452 19532 9508 19534
rect 9772 19586 9828 19588
rect 9772 19534 9774 19586
rect 9774 19534 9826 19586
rect 9826 19534 9828 19586
rect 9772 19532 9828 19534
rect 10092 19586 10148 19588
rect 10092 19534 10094 19586
rect 10094 19534 10146 19586
rect 10146 19534 10148 19586
rect 10092 19532 10148 19534
rect 10412 19586 10468 19588
rect 10412 19534 10414 19586
rect 10414 19534 10466 19586
rect 10466 19534 10468 19586
rect 10412 19532 10468 19534
rect 10732 19586 10788 19588
rect 10732 19534 10734 19586
rect 10734 19534 10786 19586
rect 10786 19534 10788 19586
rect 10732 19532 10788 19534
rect 11052 19586 11108 19588
rect 11052 19534 11054 19586
rect 11054 19534 11106 19586
rect 11106 19534 11108 19586
rect 11052 19532 11108 19534
rect 11372 19586 11428 19588
rect 11372 19534 11374 19586
rect 11374 19534 11426 19586
rect 11426 19534 11428 19586
rect 11372 19532 11428 19534
rect 11532 19586 11588 19588
rect 11532 19534 11534 19586
rect 11534 19534 11586 19586
rect 11586 19534 11588 19586
rect 11532 19532 11588 19534
rect 11852 19586 11908 19588
rect 11852 19534 11854 19586
rect 11854 19534 11906 19586
rect 11906 19534 11908 19586
rect 11852 19532 11908 19534
rect 12012 19586 12068 19588
rect 12012 19534 12014 19586
rect 12014 19534 12066 19586
rect 12066 19534 12068 19586
rect 12012 19532 12068 19534
rect 12332 19586 12388 19588
rect 12332 19534 12334 19586
rect 12334 19534 12386 19586
rect 12386 19534 12388 19586
rect 12332 19532 12388 19534
rect 8492 19426 8548 19428
rect 8492 19374 8494 19426
rect 8494 19374 8546 19426
rect 8546 19374 8548 19426
rect 8492 19372 8548 19374
rect 8812 19426 8868 19428
rect 8812 19374 8814 19426
rect 8814 19374 8866 19426
rect 8866 19374 8868 19426
rect 8812 19372 8868 19374
rect 8972 19426 9028 19428
rect 8972 19374 8974 19426
rect 8974 19374 9026 19426
rect 9026 19374 9028 19426
rect 8972 19372 9028 19374
rect 9292 19426 9348 19428
rect 9292 19374 9294 19426
rect 9294 19374 9346 19426
rect 9346 19374 9348 19426
rect 9292 19372 9348 19374
rect 9452 19426 9508 19428
rect 9452 19374 9454 19426
rect 9454 19374 9506 19426
rect 9506 19374 9508 19426
rect 9452 19372 9508 19374
rect 9772 19426 9828 19428
rect 9772 19374 9774 19426
rect 9774 19374 9826 19426
rect 9826 19374 9828 19426
rect 9772 19372 9828 19374
rect 10092 19426 10148 19428
rect 10092 19374 10094 19426
rect 10094 19374 10146 19426
rect 10146 19374 10148 19426
rect 10092 19372 10148 19374
rect 10412 19426 10468 19428
rect 10412 19374 10414 19426
rect 10414 19374 10466 19426
rect 10466 19374 10468 19426
rect 10412 19372 10468 19374
rect 10732 19426 10788 19428
rect 10732 19374 10734 19426
rect 10734 19374 10786 19426
rect 10786 19374 10788 19426
rect 10732 19372 10788 19374
rect 11052 19426 11108 19428
rect 11052 19374 11054 19426
rect 11054 19374 11106 19426
rect 11106 19374 11108 19426
rect 11052 19372 11108 19374
rect 11372 19426 11428 19428
rect 11372 19374 11374 19426
rect 11374 19374 11426 19426
rect 11426 19374 11428 19426
rect 11372 19372 11428 19374
rect 11532 19426 11588 19428
rect 11532 19374 11534 19426
rect 11534 19374 11586 19426
rect 11586 19374 11588 19426
rect 11532 19372 11588 19374
rect 11852 19426 11908 19428
rect 11852 19374 11854 19426
rect 11854 19374 11906 19426
rect 11906 19374 11908 19426
rect 11852 19372 11908 19374
rect 12012 19426 12068 19428
rect 12012 19374 12014 19426
rect 12014 19374 12066 19426
rect 12066 19374 12068 19426
rect 12012 19372 12068 19374
rect 12332 19426 12388 19428
rect 12332 19374 12334 19426
rect 12334 19374 12386 19426
rect 12386 19374 12388 19426
rect 12332 19372 12388 19374
rect 8492 19266 8548 19268
rect 8492 19214 8494 19266
rect 8494 19214 8546 19266
rect 8546 19214 8548 19266
rect 8492 19212 8548 19214
rect 8812 19266 8868 19268
rect 8812 19214 8814 19266
rect 8814 19214 8866 19266
rect 8866 19214 8868 19266
rect 8812 19212 8868 19214
rect 8972 19266 9028 19268
rect 8972 19214 8974 19266
rect 8974 19214 9026 19266
rect 9026 19214 9028 19266
rect 8972 19212 9028 19214
rect 9292 19266 9348 19268
rect 9292 19214 9294 19266
rect 9294 19214 9346 19266
rect 9346 19214 9348 19266
rect 9292 19212 9348 19214
rect 9452 19266 9508 19268
rect 9452 19214 9454 19266
rect 9454 19214 9506 19266
rect 9506 19214 9508 19266
rect 9452 19212 9508 19214
rect 9772 19266 9828 19268
rect 9772 19214 9774 19266
rect 9774 19214 9826 19266
rect 9826 19214 9828 19266
rect 9772 19212 9828 19214
rect 10092 19266 10148 19268
rect 10092 19214 10094 19266
rect 10094 19214 10146 19266
rect 10146 19214 10148 19266
rect 10092 19212 10148 19214
rect 10412 19266 10468 19268
rect 10412 19214 10414 19266
rect 10414 19214 10466 19266
rect 10466 19214 10468 19266
rect 10412 19212 10468 19214
rect 10732 19266 10788 19268
rect 10732 19214 10734 19266
rect 10734 19214 10786 19266
rect 10786 19214 10788 19266
rect 10732 19212 10788 19214
rect 11052 19266 11108 19268
rect 11052 19214 11054 19266
rect 11054 19214 11106 19266
rect 11106 19214 11108 19266
rect 11052 19212 11108 19214
rect 11372 19266 11428 19268
rect 11372 19214 11374 19266
rect 11374 19214 11426 19266
rect 11426 19214 11428 19266
rect 11372 19212 11428 19214
rect 11532 19266 11588 19268
rect 11532 19214 11534 19266
rect 11534 19214 11586 19266
rect 11586 19214 11588 19266
rect 11532 19212 11588 19214
rect 11852 19266 11908 19268
rect 11852 19214 11854 19266
rect 11854 19214 11906 19266
rect 11906 19214 11908 19266
rect 11852 19212 11908 19214
rect 12012 19266 12068 19268
rect 12012 19214 12014 19266
rect 12014 19214 12066 19266
rect 12066 19214 12068 19266
rect 12012 19212 12068 19214
rect 12332 19266 12388 19268
rect 12332 19214 12334 19266
rect 12334 19214 12386 19266
rect 12386 19214 12388 19266
rect 12332 19212 12388 19214
rect 8492 19106 8548 19108
rect 8492 19054 8494 19106
rect 8494 19054 8546 19106
rect 8546 19054 8548 19106
rect 8492 19052 8548 19054
rect 8812 19106 8868 19108
rect 8812 19054 8814 19106
rect 8814 19054 8866 19106
rect 8866 19054 8868 19106
rect 8812 19052 8868 19054
rect 8972 19106 9028 19108
rect 8972 19054 8974 19106
rect 8974 19054 9026 19106
rect 9026 19054 9028 19106
rect 8972 19052 9028 19054
rect 9292 19106 9348 19108
rect 9292 19054 9294 19106
rect 9294 19054 9346 19106
rect 9346 19054 9348 19106
rect 9292 19052 9348 19054
rect 9452 19106 9508 19108
rect 9452 19054 9454 19106
rect 9454 19054 9506 19106
rect 9506 19054 9508 19106
rect 9452 19052 9508 19054
rect 9772 19106 9828 19108
rect 9772 19054 9774 19106
rect 9774 19054 9826 19106
rect 9826 19054 9828 19106
rect 9772 19052 9828 19054
rect 10092 19106 10148 19108
rect 10092 19054 10094 19106
rect 10094 19054 10146 19106
rect 10146 19054 10148 19106
rect 10092 19052 10148 19054
rect 10412 19106 10468 19108
rect 10412 19054 10414 19106
rect 10414 19054 10466 19106
rect 10466 19054 10468 19106
rect 10412 19052 10468 19054
rect 10732 19106 10788 19108
rect 10732 19054 10734 19106
rect 10734 19054 10786 19106
rect 10786 19054 10788 19106
rect 10732 19052 10788 19054
rect 11052 19106 11108 19108
rect 11052 19054 11054 19106
rect 11054 19054 11106 19106
rect 11106 19054 11108 19106
rect 11052 19052 11108 19054
rect 11372 19106 11428 19108
rect 11372 19054 11374 19106
rect 11374 19054 11426 19106
rect 11426 19054 11428 19106
rect 11372 19052 11428 19054
rect 11532 19106 11588 19108
rect 11532 19054 11534 19106
rect 11534 19054 11586 19106
rect 11586 19054 11588 19106
rect 11532 19052 11588 19054
rect 11852 19106 11908 19108
rect 11852 19054 11854 19106
rect 11854 19054 11906 19106
rect 11906 19054 11908 19106
rect 11852 19052 11908 19054
rect 12012 19106 12068 19108
rect 12012 19054 12014 19106
rect 12014 19054 12066 19106
rect 12066 19054 12068 19106
rect 12012 19052 12068 19054
rect 12332 19106 12388 19108
rect 12332 19054 12334 19106
rect 12334 19054 12386 19106
rect 12386 19054 12388 19106
rect 12332 19052 12388 19054
rect 8492 18946 8548 18948
rect 8492 18894 8494 18946
rect 8494 18894 8546 18946
rect 8546 18894 8548 18946
rect 8492 18892 8548 18894
rect 8812 18946 8868 18948
rect 8812 18894 8814 18946
rect 8814 18894 8866 18946
rect 8866 18894 8868 18946
rect 8812 18892 8868 18894
rect 8972 18946 9028 18948
rect 8972 18894 8974 18946
rect 8974 18894 9026 18946
rect 9026 18894 9028 18946
rect 8972 18892 9028 18894
rect 9292 18946 9348 18948
rect 9292 18894 9294 18946
rect 9294 18894 9346 18946
rect 9346 18894 9348 18946
rect 9292 18892 9348 18894
rect 9452 18946 9508 18948
rect 9452 18894 9454 18946
rect 9454 18894 9506 18946
rect 9506 18894 9508 18946
rect 9452 18892 9508 18894
rect 9772 18946 9828 18948
rect 9772 18894 9774 18946
rect 9774 18894 9826 18946
rect 9826 18894 9828 18946
rect 9772 18892 9828 18894
rect 10092 18946 10148 18948
rect 10092 18894 10094 18946
rect 10094 18894 10146 18946
rect 10146 18894 10148 18946
rect 10092 18892 10148 18894
rect 10412 18946 10468 18948
rect 10412 18894 10414 18946
rect 10414 18894 10466 18946
rect 10466 18894 10468 18946
rect 10412 18892 10468 18894
rect 10732 18946 10788 18948
rect 10732 18894 10734 18946
rect 10734 18894 10786 18946
rect 10786 18894 10788 18946
rect 10732 18892 10788 18894
rect 11052 18946 11108 18948
rect 11052 18894 11054 18946
rect 11054 18894 11106 18946
rect 11106 18894 11108 18946
rect 11052 18892 11108 18894
rect 11372 18946 11428 18948
rect 11372 18894 11374 18946
rect 11374 18894 11426 18946
rect 11426 18894 11428 18946
rect 11372 18892 11428 18894
rect 11532 18946 11588 18948
rect 11532 18894 11534 18946
rect 11534 18894 11586 18946
rect 11586 18894 11588 18946
rect 11532 18892 11588 18894
rect 11852 18946 11908 18948
rect 11852 18894 11854 18946
rect 11854 18894 11906 18946
rect 11906 18894 11908 18946
rect 11852 18892 11908 18894
rect 12012 18946 12068 18948
rect 12012 18894 12014 18946
rect 12014 18894 12066 18946
rect 12066 18894 12068 18946
rect 12012 18892 12068 18894
rect 12332 18946 12388 18948
rect 12332 18894 12334 18946
rect 12334 18894 12386 18946
rect 12386 18894 12388 18946
rect 12332 18892 12388 18894
rect 8492 18786 8548 18788
rect 8492 18734 8494 18786
rect 8494 18734 8546 18786
rect 8546 18734 8548 18786
rect 8492 18732 8548 18734
rect 8812 18786 8868 18788
rect 8812 18734 8814 18786
rect 8814 18734 8866 18786
rect 8866 18734 8868 18786
rect 8812 18732 8868 18734
rect 8972 18786 9028 18788
rect 8972 18734 8974 18786
rect 8974 18734 9026 18786
rect 9026 18734 9028 18786
rect 8972 18732 9028 18734
rect 9292 18786 9348 18788
rect 9292 18734 9294 18786
rect 9294 18734 9346 18786
rect 9346 18734 9348 18786
rect 9292 18732 9348 18734
rect 9452 18786 9508 18788
rect 9452 18734 9454 18786
rect 9454 18734 9506 18786
rect 9506 18734 9508 18786
rect 9452 18732 9508 18734
rect 9772 18786 9828 18788
rect 9772 18734 9774 18786
rect 9774 18734 9826 18786
rect 9826 18734 9828 18786
rect 9772 18732 9828 18734
rect 10092 18786 10148 18788
rect 10092 18734 10094 18786
rect 10094 18734 10146 18786
rect 10146 18734 10148 18786
rect 10092 18732 10148 18734
rect 10412 18786 10468 18788
rect 10412 18734 10414 18786
rect 10414 18734 10466 18786
rect 10466 18734 10468 18786
rect 10412 18732 10468 18734
rect 10732 18786 10788 18788
rect 10732 18734 10734 18786
rect 10734 18734 10786 18786
rect 10786 18734 10788 18786
rect 10732 18732 10788 18734
rect 11052 18786 11108 18788
rect 11052 18734 11054 18786
rect 11054 18734 11106 18786
rect 11106 18734 11108 18786
rect 11052 18732 11108 18734
rect 11372 18786 11428 18788
rect 11372 18734 11374 18786
rect 11374 18734 11426 18786
rect 11426 18734 11428 18786
rect 11372 18732 11428 18734
rect 11532 18786 11588 18788
rect 11532 18734 11534 18786
rect 11534 18734 11586 18786
rect 11586 18734 11588 18786
rect 11532 18732 11588 18734
rect 11852 18786 11908 18788
rect 11852 18734 11854 18786
rect 11854 18734 11906 18786
rect 11906 18734 11908 18786
rect 11852 18732 11908 18734
rect 12012 18786 12068 18788
rect 12012 18734 12014 18786
rect 12014 18734 12066 18786
rect 12066 18734 12068 18786
rect 12012 18732 12068 18734
rect 12332 18786 12388 18788
rect 12332 18734 12334 18786
rect 12334 18734 12386 18786
rect 12386 18734 12388 18786
rect 12332 18732 12388 18734
rect 10252 18492 10308 18548
rect 9932 18172 9988 18228
rect 10892 18172 10948 18228
rect 8492 17986 8548 17988
rect 8492 17934 8494 17986
rect 8494 17934 8546 17986
rect 8546 17934 8548 17986
rect 8492 17932 8548 17934
rect 8812 17986 8868 17988
rect 8812 17934 8814 17986
rect 8814 17934 8866 17986
rect 8866 17934 8868 17986
rect 8812 17932 8868 17934
rect 8972 17986 9028 17988
rect 8972 17934 8974 17986
rect 8974 17934 9026 17986
rect 9026 17934 9028 17986
rect 8972 17932 9028 17934
rect 9292 17986 9348 17988
rect 9292 17934 9294 17986
rect 9294 17934 9346 17986
rect 9346 17934 9348 17986
rect 9292 17932 9348 17934
rect 9452 17986 9508 17988
rect 9452 17934 9454 17986
rect 9454 17934 9506 17986
rect 9506 17934 9508 17986
rect 9452 17932 9508 17934
rect 9772 17986 9828 17988
rect 9772 17934 9774 17986
rect 9774 17934 9826 17986
rect 9826 17934 9828 17986
rect 9772 17932 9828 17934
rect 10092 17986 10148 17988
rect 10092 17934 10094 17986
rect 10094 17934 10146 17986
rect 10146 17934 10148 17986
rect 10092 17932 10148 17934
rect 10412 17986 10468 17988
rect 10412 17934 10414 17986
rect 10414 17934 10466 17986
rect 10466 17934 10468 17986
rect 10412 17932 10468 17934
rect 10732 17986 10788 17988
rect 10732 17934 10734 17986
rect 10734 17934 10786 17986
rect 10786 17934 10788 17986
rect 10732 17932 10788 17934
rect 11052 17986 11108 17988
rect 11052 17934 11054 17986
rect 11054 17934 11106 17986
rect 11106 17934 11108 17986
rect 11052 17932 11108 17934
rect 11372 17986 11428 17988
rect 11372 17934 11374 17986
rect 11374 17934 11426 17986
rect 11426 17934 11428 17986
rect 11372 17932 11428 17934
rect 11532 17986 11588 17988
rect 11532 17934 11534 17986
rect 11534 17934 11586 17986
rect 11586 17934 11588 17986
rect 11532 17932 11588 17934
rect 11852 17986 11908 17988
rect 11852 17934 11854 17986
rect 11854 17934 11906 17986
rect 11906 17934 11908 17986
rect 11852 17932 11908 17934
rect 12012 17986 12068 17988
rect 12012 17934 12014 17986
rect 12014 17934 12066 17986
rect 12066 17934 12068 17986
rect 12012 17932 12068 17934
rect 12332 17986 12388 17988
rect 12332 17934 12334 17986
rect 12334 17934 12386 17986
rect 12386 17934 12388 17986
rect 12332 17932 12388 17934
rect 8492 17826 8548 17828
rect 8492 17774 8494 17826
rect 8494 17774 8546 17826
rect 8546 17774 8548 17826
rect 8492 17772 8548 17774
rect 8812 17826 8868 17828
rect 8812 17774 8814 17826
rect 8814 17774 8866 17826
rect 8866 17774 8868 17826
rect 8812 17772 8868 17774
rect 8972 17826 9028 17828
rect 8972 17774 8974 17826
rect 8974 17774 9026 17826
rect 9026 17774 9028 17826
rect 8972 17772 9028 17774
rect 9292 17826 9348 17828
rect 9292 17774 9294 17826
rect 9294 17774 9346 17826
rect 9346 17774 9348 17826
rect 9292 17772 9348 17774
rect 9452 17826 9508 17828
rect 9452 17774 9454 17826
rect 9454 17774 9506 17826
rect 9506 17774 9508 17826
rect 9452 17772 9508 17774
rect 9772 17826 9828 17828
rect 9772 17774 9774 17826
rect 9774 17774 9826 17826
rect 9826 17774 9828 17826
rect 9772 17772 9828 17774
rect 10092 17826 10148 17828
rect 10092 17774 10094 17826
rect 10094 17774 10146 17826
rect 10146 17774 10148 17826
rect 10092 17772 10148 17774
rect 10412 17826 10468 17828
rect 10412 17774 10414 17826
rect 10414 17774 10466 17826
rect 10466 17774 10468 17826
rect 10412 17772 10468 17774
rect 10732 17826 10788 17828
rect 10732 17774 10734 17826
rect 10734 17774 10786 17826
rect 10786 17774 10788 17826
rect 10732 17772 10788 17774
rect 11052 17826 11108 17828
rect 11052 17774 11054 17826
rect 11054 17774 11106 17826
rect 11106 17774 11108 17826
rect 11052 17772 11108 17774
rect 11372 17826 11428 17828
rect 11372 17774 11374 17826
rect 11374 17774 11426 17826
rect 11426 17774 11428 17826
rect 11372 17772 11428 17774
rect 11532 17826 11588 17828
rect 11532 17774 11534 17826
rect 11534 17774 11586 17826
rect 11586 17774 11588 17826
rect 11532 17772 11588 17774
rect 11852 17826 11908 17828
rect 11852 17774 11854 17826
rect 11854 17774 11906 17826
rect 11906 17774 11908 17826
rect 11852 17772 11908 17774
rect 12012 17826 12068 17828
rect 12012 17774 12014 17826
rect 12014 17774 12066 17826
rect 12066 17774 12068 17826
rect 12012 17772 12068 17774
rect 12332 17826 12388 17828
rect 12332 17774 12334 17826
rect 12334 17774 12386 17826
rect 12386 17774 12388 17826
rect 12332 17772 12388 17774
rect 8492 17666 8548 17668
rect 8492 17614 8494 17666
rect 8494 17614 8546 17666
rect 8546 17614 8548 17666
rect 8492 17612 8548 17614
rect 8812 17666 8868 17668
rect 8812 17614 8814 17666
rect 8814 17614 8866 17666
rect 8866 17614 8868 17666
rect 8812 17612 8868 17614
rect 8972 17666 9028 17668
rect 8972 17614 8974 17666
rect 8974 17614 9026 17666
rect 9026 17614 9028 17666
rect 8972 17612 9028 17614
rect 9292 17666 9348 17668
rect 9292 17614 9294 17666
rect 9294 17614 9346 17666
rect 9346 17614 9348 17666
rect 9292 17612 9348 17614
rect 9452 17666 9508 17668
rect 9452 17614 9454 17666
rect 9454 17614 9506 17666
rect 9506 17614 9508 17666
rect 9452 17612 9508 17614
rect 9772 17666 9828 17668
rect 9772 17614 9774 17666
rect 9774 17614 9826 17666
rect 9826 17614 9828 17666
rect 9772 17612 9828 17614
rect 10092 17666 10148 17668
rect 10092 17614 10094 17666
rect 10094 17614 10146 17666
rect 10146 17614 10148 17666
rect 10092 17612 10148 17614
rect 10412 17666 10468 17668
rect 10412 17614 10414 17666
rect 10414 17614 10466 17666
rect 10466 17614 10468 17666
rect 10412 17612 10468 17614
rect 10732 17666 10788 17668
rect 10732 17614 10734 17666
rect 10734 17614 10786 17666
rect 10786 17614 10788 17666
rect 10732 17612 10788 17614
rect 11052 17666 11108 17668
rect 11052 17614 11054 17666
rect 11054 17614 11106 17666
rect 11106 17614 11108 17666
rect 11052 17612 11108 17614
rect 11372 17666 11428 17668
rect 11372 17614 11374 17666
rect 11374 17614 11426 17666
rect 11426 17614 11428 17666
rect 11372 17612 11428 17614
rect 11532 17666 11588 17668
rect 11532 17614 11534 17666
rect 11534 17614 11586 17666
rect 11586 17614 11588 17666
rect 11532 17612 11588 17614
rect 11852 17666 11908 17668
rect 11852 17614 11854 17666
rect 11854 17614 11906 17666
rect 11906 17614 11908 17666
rect 11852 17612 11908 17614
rect 12012 17666 12068 17668
rect 12012 17614 12014 17666
rect 12014 17614 12066 17666
rect 12066 17614 12068 17666
rect 12012 17612 12068 17614
rect 12332 17666 12388 17668
rect 12332 17614 12334 17666
rect 12334 17614 12386 17666
rect 12386 17614 12388 17666
rect 12332 17612 12388 17614
rect 8492 17506 8548 17508
rect 8492 17454 8494 17506
rect 8494 17454 8546 17506
rect 8546 17454 8548 17506
rect 8492 17452 8548 17454
rect 8812 17506 8868 17508
rect 8812 17454 8814 17506
rect 8814 17454 8866 17506
rect 8866 17454 8868 17506
rect 8812 17452 8868 17454
rect 8972 17506 9028 17508
rect 8972 17454 8974 17506
rect 8974 17454 9026 17506
rect 9026 17454 9028 17506
rect 8972 17452 9028 17454
rect 9292 17506 9348 17508
rect 9292 17454 9294 17506
rect 9294 17454 9346 17506
rect 9346 17454 9348 17506
rect 9292 17452 9348 17454
rect 9452 17506 9508 17508
rect 9452 17454 9454 17506
rect 9454 17454 9506 17506
rect 9506 17454 9508 17506
rect 9452 17452 9508 17454
rect 9772 17506 9828 17508
rect 9772 17454 9774 17506
rect 9774 17454 9826 17506
rect 9826 17454 9828 17506
rect 9772 17452 9828 17454
rect 10092 17506 10148 17508
rect 10092 17454 10094 17506
rect 10094 17454 10146 17506
rect 10146 17454 10148 17506
rect 10092 17452 10148 17454
rect 10412 17506 10468 17508
rect 10412 17454 10414 17506
rect 10414 17454 10466 17506
rect 10466 17454 10468 17506
rect 10412 17452 10468 17454
rect 10732 17506 10788 17508
rect 10732 17454 10734 17506
rect 10734 17454 10786 17506
rect 10786 17454 10788 17506
rect 10732 17452 10788 17454
rect 11052 17506 11108 17508
rect 11052 17454 11054 17506
rect 11054 17454 11106 17506
rect 11106 17454 11108 17506
rect 11052 17452 11108 17454
rect 11372 17506 11428 17508
rect 11372 17454 11374 17506
rect 11374 17454 11426 17506
rect 11426 17454 11428 17506
rect 11372 17452 11428 17454
rect 11532 17506 11588 17508
rect 11532 17454 11534 17506
rect 11534 17454 11586 17506
rect 11586 17454 11588 17506
rect 11532 17452 11588 17454
rect 11852 17506 11908 17508
rect 11852 17454 11854 17506
rect 11854 17454 11906 17506
rect 11906 17454 11908 17506
rect 11852 17452 11908 17454
rect 12012 17506 12068 17508
rect 12012 17454 12014 17506
rect 12014 17454 12066 17506
rect 12066 17454 12068 17506
rect 12012 17452 12068 17454
rect 12332 17506 12388 17508
rect 12332 17454 12334 17506
rect 12334 17454 12386 17506
rect 12386 17454 12388 17506
rect 12332 17452 12388 17454
rect 8492 17346 8548 17348
rect 8492 17294 8494 17346
rect 8494 17294 8546 17346
rect 8546 17294 8548 17346
rect 8492 17292 8548 17294
rect 8812 17346 8868 17348
rect 8812 17294 8814 17346
rect 8814 17294 8866 17346
rect 8866 17294 8868 17346
rect 8812 17292 8868 17294
rect 8972 17346 9028 17348
rect 8972 17294 8974 17346
rect 8974 17294 9026 17346
rect 9026 17294 9028 17346
rect 8972 17292 9028 17294
rect 9292 17346 9348 17348
rect 9292 17294 9294 17346
rect 9294 17294 9346 17346
rect 9346 17294 9348 17346
rect 9292 17292 9348 17294
rect 9452 17346 9508 17348
rect 9452 17294 9454 17346
rect 9454 17294 9506 17346
rect 9506 17294 9508 17346
rect 9452 17292 9508 17294
rect 9772 17346 9828 17348
rect 9772 17294 9774 17346
rect 9774 17294 9826 17346
rect 9826 17294 9828 17346
rect 9772 17292 9828 17294
rect 10092 17346 10148 17348
rect 10092 17294 10094 17346
rect 10094 17294 10146 17346
rect 10146 17294 10148 17346
rect 10092 17292 10148 17294
rect 10412 17346 10468 17348
rect 10412 17294 10414 17346
rect 10414 17294 10466 17346
rect 10466 17294 10468 17346
rect 10412 17292 10468 17294
rect 10732 17346 10788 17348
rect 10732 17294 10734 17346
rect 10734 17294 10786 17346
rect 10786 17294 10788 17346
rect 10732 17292 10788 17294
rect 11052 17346 11108 17348
rect 11052 17294 11054 17346
rect 11054 17294 11106 17346
rect 11106 17294 11108 17346
rect 11052 17292 11108 17294
rect 11372 17346 11428 17348
rect 11372 17294 11374 17346
rect 11374 17294 11426 17346
rect 11426 17294 11428 17346
rect 11372 17292 11428 17294
rect 11532 17346 11588 17348
rect 11532 17294 11534 17346
rect 11534 17294 11586 17346
rect 11586 17294 11588 17346
rect 11532 17292 11588 17294
rect 11852 17346 11908 17348
rect 11852 17294 11854 17346
rect 11854 17294 11906 17346
rect 11906 17294 11908 17346
rect 11852 17292 11908 17294
rect 12012 17346 12068 17348
rect 12012 17294 12014 17346
rect 12014 17294 12066 17346
rect 12066 17294 12068 17346
rect 12012 17292 12068 17294
rect 12332 17346 12388 17348
rect 12332 17294 12334 17346
rect 12334 17294 12386 17346
rect 12386 17294 12388 17346
rect 12332 17292 12388 17294
rect 8492 17186 8548 17188
rect 8492 17134 8494 17186
rect 8494 17134 8546 17186
rect 8546 17134 8548 17186
rect 8492 17132 8548 17134
rect 8812 17186 8868 17188
rect 8812 17134 8814 17186
rect 8814 17134 8866 17186
rect 8866 17134 8868 17186
rect 8812 17132 8868 17134
rect 8972 17186 9028 17188
rect 8972 17134 8974 17186
rect 8974 17134 9026 17186
rect 9026 17134 9028 17186
rect 8972 17132 9028 17134
rect 9292 17186 9348 17188
rect 9292 17134 9294 17186
rect 9294 17134 9346 17186
rect 9346 17134 9348 17186
rect 9292 17132 9348 17134
rect 9452 17186 9508 17188
rect 9452 17134 9454 17186
rect 9454 17134 9506 17186
rect 9506 17134 9508 17186
rect 9452 17132 9508 17134
rect 9772 17186 9828 17188
rect 9772 17134 9774 17186
rect 9774 17134 9826 17186
rect 9826 17134 9828 17186
rect 9772 17132 9828 17134
rect 10092 17186 10148 17188
rect 10092 17134 10094 17186
rect 10094 17134 10146 17186
rect 10146 17134 10148 17186
rect 10092 17132 10148 17134
rect 10412 17186 10468 17188
rect 10412 17134 10414 17186
rect 10414 17134 10466 17186
rect 10466 17134 10468 17186
rect 10412 17132 10468 17134
rect 10732 17186 10788 17188
rect 10732 17134 10734 17186
rect 10734 17134 10786 17186
rect 10786 17134 10788 17186
rect 10732 17132 10788 17134
rect 11052 17186 11108 17188
rect 11052 17134 11054 17186
rect 11054 17134 11106 17186
rect 11106 17134 11108 17186
rect 11052 17132 11108 17134
rect 11372 17186 11428 17188
rect 11372 17134 11374 17186
rect 11374 17134 11426 17186
rect 11426 17134 11428 17186
rect 11372 17132 11428 17134
rect 11532 17186 11588 17188
rect 11532 17134 11534 17186
rect 11534 17134 11586 17186
rect 11586 17134 11588 17186
rect 11532 17132 11588 17134
rect 11852 17186 11908 17188
rect 11852 17134 11854 17186
rect 11854 17134 11906 17186
rect 11906 17134 11908 17186
rect 11852 17132 11908 17134
rect 12012 17186 12068 17188
rect 12012 17134 12014 17186
rect 12014 17134 12066 17186
rect 12066 17134 12068 17186
rect 12012 17132 12068 17134
rect 12332 17186 12388 17188
rect 12332 17134 12334 17186
rect 12334 17134 12386 17186
rect 12386 17134 12388 17186
rect 12332 17132 12388 17134
rect 8492 17026 8548 17028
rect 8492 16974 8494 17026
rect 8494 16974 8546 17026
rect 8546 16974 8548 17026
rect 8492 16972 8548 16974
rect 8812 17026 8868 17028
rect 8812 16974 8814 17026
rect 8814 16974 8866 17026
rect 8866 16974 8868 17026
rect 8812 16972 8868 16974
rect 8972 17026 9028 17028
rect 8972 16974 8974 17026
rect 8974 16974 9026 17026
rect 9026 16974 9028 17026
rect 8972 16972 9028 16974
rect 9292 17026 9348 17028
rect 9292 16974 9294 17026
rect 9294 16974 9346 17026
rect 9346 16974 9348 17026
rect 9292 16972 9348 16974
rect 9452 17026 9508 17028
rect 9452 16974 9454 17026
rect 9454 16974 9506 17026
rect 9506 16974 9508 17026
rect 9452 16972 9508 16974
rect 9772 17026 9828 17028
rect 9772 16974 9774 17026
rect 9774 16974 9826 17026
rect 9826 16974 9828 17026
rect 9772 16972 9828 16974
rect 10092 17026 10148 17028
rect 10092 16974 10094 17026
rect 10094 16974 10146 17026
rect 10146 16974 10148 17026
rect 10092 16972 10148 16974
rect 10412 17026 10468 17028
rect 10412 16974 10414 17026
rect 10414 16974 10466 17026
rect 10466 16974 10468 17026
rect 10412 16972 10468 16974
rect 10732 17026 10788 17028
rect 10732 16974 10734 17026
rect 10734 16974 10786 17026
rect 10786 16974 10788 17026
rect 10732 16972 10788 16974
rect 11052 17026 11108 17028
rect 11052 16974 11054 17026
rect 11054 16974 11106 17026
rect 11106 16974 11108 17026
rect 11052 16972 11108 16974
rect 11372 17026 11428 17028
rect 11372 16974 11374 17026
rect 11374 16974 11426 17026
rect 11426 16974 11428 17026
rect 11372 16972 11428 16974
rect 11532 17026 11588 17028
rect 11532 16974 11534 17026
rect 11534 16974 11586 17026
rect 11586 16974 11588 17026
rect 11532 16972 11588 16974
rect 11852 17026 11908 17028
rect 11852 16974 11854 17026
rect 11854 16974 11906 17026
rect 11906 16974 11908 17026
rect 11852 16972 11908 16974
rect 12012 17026 12068 17028
rect 12012 16974 12014 17026
rect 12014 16974 12066 17026
rect 12066 16974 12068 17026
rect 12012 16972 12068 16974
rect 12332 17026 12388 17028
rect 12332 16974 12334 17026
rect 12334 16974 12386 17026
rect 12386 16974 12388 17026
rect 12332 16972 12388 16974
rect 8492 16866 8548 16868
rect 8492 16814 8494 16866
rect 8494 16814 8546 16866
rect 8546 16814 8548 16866
rect 8492 16812 8548 16814
rect 8812 16866 8868 16868
rect 8812 16814 8814 16866
rect 8814 16814 8866 16866
rect 8866 16814 8868 16866
rect 8812 16812 8868 16814
rect 8972 16866 9028 16868
rect 8972 16814 8974 16866
rect 8974 16814 9026 16866
rect 9026 16814 9028 16866
rect 8972 16812 9028 16814
rect 9292 16866 9348 16868
rect 9292 16814 9294 16866
rect 9294 16814 9346 16866
rect 9346 16814 9348 16866
rect 9292 16812 9348 16814
rect 9452 16866 9508 16868
rect 9452 16814 9454 16866
rect 9454 16814 9506 16866
rect 9506 16814 9508 16866
rect 9452 16812 9508 16814
rect 9772 16866 9828 16868
rect 9772 16814 9774 16866
rect 9774 16814 9826 16866
rect 9826 16814 9828 16866
rect 9772 16812 9828 16814
rect 10092 16866 10148 16868
rect 10092 16814 10094 16866
rect 10094 16814 10146 16866
rect 10146 16814 10148 16866
rect 10092 16812 10148 16814
rect 10412 16866 10468 16868
rect 10412 16814 10414 16866
rect 10414 16814 10466 16866
rect 10466 16814 10468 16866
rect 10412 16812 10468 16814
rect 10732 16866 10788 16868
rect 10732 16814 10734 16866
rect 10734 16814 10786 16866
rect 10786 16814 10788 16866
rect 10732 16812 10788 16814
rect 11052 16866 11108 16868
rect 11052 16814 11054 16866
rect 11054 16814 11106 16866
rect 11106 16814 11108 16866
rect 11052 16812 11108 16814
rect 11372 16866 11428 16868
rect 11372 16814 11374 16866
rect 11374 16814 11426 16866
rect 11426 16814 11428 16866
rect 11372 16812 11428 16814
rect 11532 16866 11588 16868
rect 11532 16814 11534 16866
rect 11534 16814 11586 16866
rect 11586 16814 11588 16866
rect 11532 16812 11588 16814
rect 11852 16866 11908 16868
rect 11852 16814 11854 16866
rect 11854 16814 11906 16866
rect 11906 16814 11908 16866
rect 11852 16812 11908 16814
rect 12012 16866 12068 16868
rect 12012 16814 12014 16866
rect 12014 16814 12066 16866
rect 12066 16814 12068 16866
rect 12012 16812 12068 16814
rect 12332 16866 12388 16868
rect 12332 16814 12334 16866
rect 12334 16814 12386 16866
rect 12386 16814 12388 16866
rect 12332 16812 12388 16814
rect 9132 16652 9188 16708
rect 8492 16546 8548 16548
rect 8492 16494 8494 16546
rect 8494 16494 8546 16546
rect 8546 16494 8548 16546
rect 8492 16492 8548 16494
rect 8812 16546 8868 16548
rect 8812 16494 8814 16546
rect 8814 16494 8866 16546
rect 8866 16494 8868 16546
rect 8812 16492 8868 16494
rect 8972 16546 9028 16548
rect 8972 16494 8974 16546
rect 8974 16494 9026 16546
rect 9026 16494 9028 16546
rect 8972 16492 9028 16494
rect 9292 16546 9348 16548
rect 9292 16494 9294 16546
rect 9294 16494 9346 16546
rect 9346 16494 9348 16546
rect 9292 16492 9348 16494
rect 9452 16546 9508 16548
rect 9452 16494 9454 16546
rect 9454 16494 9506 16546
rect 9506 16494 9508 16546
rect 9452 16492 9508 16494
rect 9772 16546 9828 16548
rect 9772 16494 9774 16546
rect 9774 16494 9826 16546
rect 9826 16494 9828 16546
rect 9772 16492 9828 16494
rect 10092 16546 10148 16548
rect 10092 16494 10094 16546
rect 10094 16494 10146 16546
rect 10146 16494 10148 16546
rect 10092 16492 10148 16494
rect 10412 16546 10468 16548
rect 10412 16494 10414 16546
rect 10414 16494 10466 16546
rect 10466 16494 10468 16546
rect 10412 16492 10468 16494
rect 10732 16546 10788 16548
rect 10732 16494 10734 16546
rect 10734 16494 10786 16546
rect 10786 16494 10788 16546
rect 10732 16492 10788 16494
rect 11052 16546 11108 16548
rect 11052 16494 11054 16546
rect 11054 16494 11106 16546
rect 11106 16494 11108 16546
rect 11052 16492 11108 16494
rect 11372 16546 11428 16548
rect 11372 16494 11374 16546
rect 11374 16494 11426 16546
rect 11426 16494 11428 16546
rect 11372 16492 11428 16494
rect 11532 16546 11588 16548
rect 11532 16494 11534 16546
rect 11534 16494 11586 16546
rect 11586 16494 11588 16546
rect 11532 16492 11588 16494
rect 11852 16546 11908 16548
rect 11852 16494 11854 16546
rect 11854 16494 11906 16546
rect 11906 16494 11908 16546
rect 11852 16492 11908 16494
rect 12012 16546 12068 16548
rect 12012 16494 12014 16546
rect 12014 16494 12066 16546
rect 12066 16494 12068 16546
rect 12012 16492 12068 16494
rect 12332 16546 12388 16548
rect 12332 16494 12334 16546
rect 12334 16494 12386 16546
rect 12386 16494 12388 16546
rect 12332 16492 12388 16494
rect 8492 16386 8548 16388
rect 8492 16334 8494 16386
rect 8494 16334 8546 16386
rect 8546 16334 8548 16386
rect 8492 16332 8548 16334
rect 8812 16386 8868 16388
rect 8812 16334 8814 16386
rect 8814 16334 8866 16386
rect 8866 16334 8868 16386
rect 8812 16332 8868 16334
rect 8972 16386 9028 16388
rect 8972 16334 8974 16386
rect 8974 16334 9026 16386
rect 9026 16334 9028 16386
rect 8972 16332 9028 16334
rect 9292 16386 9348 16388
rect 9292 16334 9294 16386
rect 9294 16334 9346 16386
rect 9346 16334 9348 16386
rect 9292 16332 9348 16334
rect 9452 16386 9508 16388
rect 9452 16334 9454 16386
rect 9454 16334 9506 16386
rect 9506 16334 9508 16386
rect 9452 16332 9508 16334
rect 9772 16386 9828 16388
rect 9772 16334 9774 16386
rect 9774 16334 9826 16386
rect 9826 16334 9828 16386
rect 9772 16332 9828 16334
rect 10092 16386 10148 16388
rect 10092 16334 10094 16386
rect 10094 16334 10146 16386
rect 10146 16334 10148 16386
rect 10092 16332 10148 16334
rect 10412 16386 10468 16388
rect 10412 16334 10414 16386
rect 10414 16334 10466 16386
rect 10466 16334 10468 16386
rect 10412 16332 10468 16334
rect 10732 16386 10788 16388
rect 10732 16334 10734 16386
rect 10734 16334 10786 16386
rect 10786 16334 10788 16386
rect 10732 16332 10788 16334
rect 11052 16386 11108 16388
rect 11052 16334 11054 16386
rect 11054 16334 11106 16386
rect 11106 16334 11108 16386
rect 11052 16332 11108 16334
rect 11372 16386 11428 16388
rect 11372 16334 11374 16386
rect 11374 16334 11426 16386
rect 11426 16334 11428 16386
rect 11372 16332 11428 16334
rect 11532 16386 11588 16388
rect 11532 16334 11534 16386
rect 11534 16334 11586 16386
rect 11586 16334 11588 16386
rect 11532 16332 11588 16334
rect 11852 16386 11908 16388
rect 11852 16334 11854 16386
rect 11854 16334 11906 16386
rect 11906 16334 11908 16386
rect 11852 16332 11908 16334
rect 12012 16386 12068 16388
rect 12012 16334 12014 16386
rect 12014 16334 12066 16386
rect 12066 16334 12068 16386
rect 12012 16332 12068 16334
rect 12332 16386 12388 16388
rect 12332 16334 12334 16386
rect 12334 16334 12386 16386
rect 12386 16334 12388 16386
rect 12332 16332 12388 16334
rect 8492 16226 8548 16228
rect 8492 16174 8494 16226
rect 8494 16174 8546 16226
rect 8546 16174 8548 16226
rect 8492 16172 8548 16174
rect 8812 16226 8868 16228
rect 8812 16174 8814 16226
rect 8814 16174 8866 16226
rect 8866 16174 8868 16226
rect 8812 16172 8868 16174
rect 8972 16226 9028 16228
rect 8972 16174 8974 16226
rect 8974 16174 9026 16226
rect 9026 16174 9028 16226
rect 8972 16172 9028 16174
rect 9292 16226 9348 16228
rect 9292 16174 9294 16226
rect 9294 16174 9346 16226
rect 9346 16174 9348 16226
rect 9292 16172 9348 16174
rect 9452 16226 9508 16228
rect 9452 16174 9454 16226
rect 9454 16174 9506 16226
rect 9506 16174 9508 16226
rect 9452 16172 9508 16174
rect 9772 16226 9828 16228
rect 9772 16174 9774 16226
rect 9774 16174 9826 16226
rect 9826 16174 9828 16226
rect 9772 16172 9828 16174
rect 10092 16226 10148 16228
rect 10092 16174 10094 16226
rect 10094 16174 10146 16226
rect 10146 16174 10148 16226
rect 10092 16172 10148 16174
rect 10412 16226 10468 16228
rect 10412 16174 10414 16226
rect 10414 16174 10466 16226
rect 10466 16174 10468 16226
rect 10412 16172 10468 16174
rect 10732 16226 10788 16228
rect 10732 16174 10734 16226
rect 10734 16174 10786 16226
rect 10786 16174 10788 16226
rect 10732 16172 10788 16174
rect 11052 16226 11108 16228
rect 11052 16174 11054 16226
rect 11054 16174 11106 16226
rect 11106 16174 11108 16226
rect 11052 16172 11108 16174
rect 11372 16226 11428 16228
rect 11372 16174 11374 16226
rect 11374 16174 11426 16226
rect 11426 16174 11428 16226
rect 11372 16172 11428 16174
rect 11532 16226 11588 16228
rect 11532 16174 11534 16226
rect 11534 16174 11586 16226
rect 11586 16174 11588 16226
rect 11532 16172 11588 16174
rect 11852 16226 11908 16228
rect 11852 16174 11854 16226
rect 11854 16174 11906 16226
rect 11906 16174 11908 16226
rect 11852 16172 11908 16174
rect 12012 16226 12068 16228
rect 12012 16174 12014 16226
rect 12014 16174 12066 16226
rect 12066 16174 12068 16226
rect 12012 16172 12068 16174
rect 12332 16226 12388 16228
rect 12332 16174 12334 16226
rect 12334 16174 12386 16226
rect 12386 16174 12388 16226
rect 12332 16172 12388 16174
rect 8492 16066 8548 16068
rect 8492 16014 8494 16066
rect 8494 16014 8546 16066
rect 8546 16014 8548 16066
rect 8492 16012 8548 16014
rect 8812 16066 8868 16068
rect 8812 16014 8814 16066
rect 8814 16014 8866 16066
rect 8866 16014 8868 16066
rect 8812 16012 8868 16014
rect 8972 16066 9028 16068
rect 8972 16014 8974 16066
rect 8974 16014 9026 16066
rect 9026 16014 9028 16066
rect 8972 16012 9028 16014
rect 9292 16066 9348 16068
rect 9292 16014 9294 16066
rect 9294 16014 9346 16066
rect 9346 16014 9348 16066
rect 9292 16012 9348 16014
rect 9452 16066 9508 16068
rect 9452 16014 9454 16066
rect 9454 16014 9506 16066
rect 9506 16014 9508 16066
rect 9452 16012 9508 16014
rect 9772 16066 9828 16068
rect 9772 16014 9774 16066
rect 9774 16014 9826 16066
rect 9826 16014 9828 16066
rect 9772 16012 9828 16014
rect 10092 16066 10148 16068
rect 10092 16014 10094 16066
rect 10094 16014 10146 16066
rect 10146 16014 10148 16066
rect 10092 16012 10148 16014
rect 10412 16066 10468 16068
rect 10412 16014 10414 16066
rect 10414 16014 10466 16066
rect 10466 16014 10468 16066
rect 10412 16012 10468 16014
rect 10732 16066 10788 16068
rect 10732 16014 10734 16066
rect 10734 16014 10786 16066
rect 10786 16014 10788 16066
rect 10732 16012 10788 16014
rect 11052 16066 11108 16068
rect 11052 16014 11054 16066
rect 11054 16014 11106 16066
rect 11106 16014 11108 16066
rect 11052 16012 11108 16014
rect 11372 16066 11428 16068
rect 11372 16014 11374 16066
rect 11374 16014 11426 16066
rect 11426 16014 11428 16066
rect 11372 16012 11428 16014
rect 11532 16066 11588 16068
rect 11532 16014 11534 16066
rect 11534 16014 11586 16066
rect 11586 16014 11588 16066
rect 11532 16012 11588 16014
rect 11852 16066 11908 16068
rect 11852 16014 11854 16066
rect 11854 16014 11906 16066
rect 11906 16014 11908 16066
rect 11852 16012 11908 16014
rect 12012 16066 12068 16068
rect 12012 16014 12014 16066
rect 12014 16014 12066 16066
rect 12066 16014 12068 16066
rect 12012 16012 12068 16014
rect 12332 16066 12388 16068
rect 12332 16014 12334 16066
rect 12334 16014 12386 16066
rect 12386 16014 12388 16066
rect 12332 16012 12388 16014
rect 8492 15906 8548 15908
rect 8492 15854 8494 15906
rect 8494 15854 8546 15906
rect 8546 15854 8548 15906
rect 8492 15852 8548 15854
rect 8812 15906 8868 15908
rect 8812 15854 8814 15906
rect 8814 15854 8866 15906
rect 8866 15854 8868 15906
rect 8812 15852 8868 15854
rect 8972 15906 9028 15908
rect 8972 15854 8974 15906
rect 8974 15854 9026 15906
rect 9026 15854 9028 15906
rect 8972 15852 9028 15854
rect 9292 15906 9348 15908
rect 9292 15854 9294 15906
rect 9294 15854 9346 15906
rect 9346 15854 9348 15906
rect 9292 15852 9348 15854
rect 9452 15906 9508 15908
rect 9452 15854 9454 15906
rect 9454 15854 9506 15906
rect 9506 15854 9508 15906
rect 9452 15852 9508 15854
rect 9772 15906 9828 15908
rect 9772 15854 9774 15906
rect 9774 15854 9826 15906
rect 9826 15854 9828 15906
rect 9772 15852 9828 15854
rect 10092 15906 10148 15908
rect 10092 15854 10094 15906
rect 10094 15854 10146 15906
rect 10146 15854 10148 15906
rect 10092 15852 10148 15854
rect 10412 15906 10468 15908
rect 10412 15854 10414 15906
rect 10414 15854 10466 15906
rect 10466 15854 10468 15906
rect 10412 15852 10468 15854
rect 10732 15906 10788 15908
rect 10732 15854 10734 15906
rect 10734 15854 10786 15906
rect 10786 15854 10788 15906
rect 10732 15852 10788 15854
rect 11052 15906 11108 15908
rect 11052 15854 11054 15906
rect 11054 15854 11106 15906
rect 11106 15854 11108 15906
rect 11052 15852 11108 15854
rect 11372 15906 11428 15908
rect 11372 15854 11374 15906
rect 11374 15854 11426 15906
rect 11426 15854 11428 15906
rect 11372 15852 11428 15854
rect 11532 15906 11588 15908
rect 11532 15854 11534 15906
rect 11534 15854 11586 15906
rect 11586 15854 11588 15906
rect 11532 15852 11588 15854
rect 11852 15906 11908 15908
rect 11852 15854 11854 15906
rect 11854 15854 11906 15906
rect 11906 15854 11908 15906
rect 11852 15852 11908 15854
rect 12012 15906 12068 15908
rect 12012 15854 12014 15906
rect 12014 15854 12066 15906
rect 12066 15854 12068 15906
rect 12012 15852 12068 15854
rect 12332 15906 12388 15908
rect 12332 15854 12334 15906
rect 12334 15854 12386 15906
rect 12386 15854 12388 15906
rect 12332 15852 12388 15854
rect 8492 15746 8548 15748
rect 8492 15694 8494 15746
rect 8494 15694 8546 15746
rect 8546 15694 8548 15746
rect 8492 15692 8548 15694
rect 8812 15746 8868 15748
rect 8812 15694 8814 15746
rect 8814 15694 8866 15746
rect 8866 15694 8868 15746
rect 8812 15692 8868 15694
rect 8972 15746 9028 15748
rect 8972 15694 8974 15746
rect 8974 15694 9026 15746
rect 9026 15694 9028 15746
rect 8972 15692 9028 15694
rect 9292 15746 9348 15748
rect 9292 15694 9294 15746
rect 9294 15694 9346 15746
rect 9346 15694 9348 15746
rect 9292 15692 9348 15694
rect 9452 15746 9508 15748
rect 9452 15694 9454 15746
rect 9454 15694 9506 15746
rect 9506 15694 9508 15746
rect 9452 15692 9508 15694
rect 9772 15746 9828 15748
rect 9772 15694 9774 15746
rect 9774 15694 9826 15746
rect 9826 15694 9828 15746
rect 9772 15692 9828 15694
rect 10092 15746 10148 15748
rect 10092 15694 10094 15746
rect 10094 15694 10146 15746
rect 10146 15694 10148 15746
rect 10092 15692 10148 15694
rect 10412 15746 10468 15748
rect 10412 15694 10414 15746
rect 10414 15694 10466 15746
rect 10466 15694 10468 15746
rect 10412 15692 10468 15694
rect 10732 15746 10788 15748
rect 10732 15694 10734 15746
rect 10734 15694 10786 15746
rect 10786 15694 10788 15746
rect 10732 15692 10788 15694
rect 11052 15746 11108 15748
rect 11052 15694 11054 15746
rect 11054 15694 11106 15746
rect 11106 15694 11108 15746
rect 11052 15692 11108 15694
rect 11372 15746 11428 15748
rect 11372 15694 11374 15746
rect 11374 15694 11426 15746
rect 11426 15694 11428 15746
rect 11372 15692 11428 15694
rect 11532 15746 11588 15748
rect 11532 15694 11534 15746
rect 11534 15694 11586 15746
rect 11586 15694 11588 15746
rect 11532 15692 11588 15694
rect 11852 15746 11908 15748
rect 11852 15694 11854 15746
rect 11854 15694 11906 15746
rect 11906 15694 11908 15746
rect 11852 15692 11908 15694
rect 12012 15746 12068 15748
rect 12012 15694 12014 15746
rect 12014 15694 12066 15746
rect 12066 15694 12068 15746
rect 12012 15692 12068 15694
rect 12332 15746 12388 15748
rect 12332 15694 12334 15746
rect 12334 15694 12386 15746
rect 12386 15694 12388 15746
rect 12332 15692 12388 15694
rect 8492 15586 8548 15588
rect 8492 15534 8494 15586
rect 8494 15534 8546 15586
rect 8546 15534 8548 15586
rect 8492 15532 8548 15534
rect 8812 15586 8868 15588
rect 8812 15534 8814 15586
rect 8814 15534 8866 15586
rect 8866 15534 8868 15586
rect 8812 15532 8868 15534
rect 8972 15586 9028 15588
rect 8972 15534 8974 15586
rect 8974 15534 9026 15586
rect 9026 15534 9028 15586
rect 8972 15532 9028 15534
rect 9292 15586 9348 15588
rect 9292 15534 9294 15586
rect 9294 15534 9346 15586
rect 9346 15534 9348 15586
rect 9292 15532 9348 15534
rect 9452 15586 9508 15588
rect 9452 15534 9454 15586
rect 9454 15534 9506 15586
rect 9506 15534 9508 15586
rect 9452 15532 9508 15534
rect 9772 15586 9828 15588
rect 9772 15534 9774 15586
rect 9774 15534 9826 15586
rect 9826 15534 9828 15586
rect 9772 15532 9828 15534
rect 10092 15586 10148 15588
rect 10092 15534 10094 15586
rect 10094 15534 10146 15586
rect 10146 15534 10148 15586
rect 10092 15532 10148 15534
rect 10412 15586 10468 15588
rect 10412 15534 10414 15586
rect 10414 15534 10466 15586
rect 10466 15534 10468 15586
rect 10412 15532 10468 15534
rect 10732 15586 10788 15588
rect 10732 15534 10734 15586
rect 10734 15534 10786 15586
rect 10786 15534 10788 15586
rect 10732 15532 10788 15534
rect 11052 15586 11108 15588
rect 11052 15534 11054 15586
rect 11054 15534 11106 15586
rect 11106 15534 11108 15586
rect 11052 15532 11108 15534
rect 11372 15586 11428 15588
rect 11372 15534 11374 15586
rect 11374 15534 11426 15586
rect 11426 15534 11428 15586
rect 11372 15532 11428 15534
rect 11532 15586 11588 15588
rect 11532 15534 11534 15586
rect 11534 15534 11586 15586
rect 11586 15534 11588 15586
rect 11532 15532 11588 15534
rect 11852 15586 11908 15588
rect 11852 15534 11854 15586
rect 11854 15534 11906 15586
rect 11906 15534 11908 15586
rect 11852 15532 11908 15534
rect 12012 15586 12068 15588
rect 12012 15534 12014 15586
rect 12014 15534 12066 15586
rect 12066 15534 12068 15586
rect 12012 15532 12068 15534
rect 12332 15586 12388 15588
rect 12332 15534 12334 15586
rect 12334 15534 12386 15586
rect 12386 15534 12388 15586
rect 12332 15532 12388 15534
rect 8492 15426 8548 15428
rect 8492 15374 8494 15426
rect 8494 15374 8546 15426
rect 8546 15374 8548 15426
rect 8492 15372 8548 15374
rect 8812 15426 8868 15428
rect 8812 15374 8814 15426
rect 8814 15374 8866 15426
rect 8866 15374 8868 15426
rect 8812 15372 8868 15374
rect 8972 15426 9028 15428
rect 8972 15374 8974 15426
rect 8974 15374 9026 15426
rect 9026 15374 9028 15426
rect 8972 15372 9028 15374
rect 9292 15426 9348 15428
rect 9292 15374 9294 15426
rect 9294 15374 9346 15426
rect 9346 15374 9348 15426
rect 9292 15372 9348 15374
rect 9452 15426 9508 15428
rect 9452 15374 9454 15426
rect 9454 15374 9506 15426
rect 9506 15374 9508 15426
rect 9452 15372 9508 15374
rect 9772 15426 9828 15428
rect 9772 15374 9774 15426
rect 9774 15374 9826 15426
rect 9826 15374 9828 15426
rect 9772 15372 9828 15374
rect 10092 15426 10148 15428
rect 10092 15374 10094 15426
rect 10094 15374 10146 15426
rect 10146 15374 10148 15426
rect 10092 15372 10148 15374
rect 10412 15426 10468 15428
rect 10412 15374 10414 15426
rect 10414 15374 10466 15426
rect 10466 15374 10468 15426
rect 10412 15372 10468 15374
rect 10732 15426 10788 15428
rect 10732 15374 10734 15426
rect 10734 15374 10786 15426
rect 10786 15374 10788 15426
rect 10732 15372 10788 15374
rect 11052 15426 11108 15428
rect 11052 15374 11054 15426
rect 11054 15374 11106 15426
rect 11106 15374 11108 15426
rect 11052 15372 11108 15374
rect 11372 15426 11428 15428
rect 11372 15374 11374 15426
rect 11374 15374 11426 15426
rect 11426 15374 11428 15426
rect 11372 15372 11428 15374
rect 11532 15426 11588 15428
rect 11532 15374 11534 15426
rect 11534 15374 11586 15426
rect 11586 15374 11588 15426
rect 11532 15372 11588 15374
rect 11852 15426 11908 15428
rect 11852 15374 11854 15426
rect 11854 15374 11906 15426
rect 11906 15374 11908 15426
rect 11852 15372 11908 15374
rect 12012 15426 12068 15428
rect 12012 15374 12014 15426
rect 12014 15374 12066 15426
rect 12066 15374 12068 15426
rect 12012 15372 12068 15374
rect 12332 15426 12388 15428
rect 12332 15374 12334 15426
rect 12334 15374 12386 15426
rect 12386 15374 12388 15426
rect 12332 15372 12388 15374
rect 8492 15266 8548 15268
rect 8492 15214 8494 15266
rect 8494 15214 8546 15266
rect 8546 15214 8548 15266
rect 8492 15212 8548 15214
rect 8812 15266 8868 15268
rect 8812 15214 8814 15266
rect 8814 15214 8866 15266
rect 8866 15214 8868 15266
rect 8812 15212 8868 15214
rect 8972 15266 9028 15268
rect 8972 15214 8974 15266
rect 8974 15214 9026 15266
rect 9026 15214 9028 15266
rect 8972 15212 9028 15214
rect 9292 15266 9348 15268
rect 9292 15214 9294 15266
rect 9294 15214 9346 15266
rect 9346 15214 9348 15266
rect 9292 15212 9348 15214
rect 9452 15266 9508 15268
rect 9452 15214 9454 15266
rect 9454 15214 9506 15266
rect 9506 15214 9508 15266
rect 9452 15212 9508 15214
rect 9772 15266 9828 15268
rect 9772 15214 9774 15266
rect 9774 15214 9826 15266
rect 9826 15214 9828 15266
rect 9772 15212 9828 15214
rect 10092 15266 10148 15268
rect 10092 15214 10094 15266
rect 10094 15214 10146 15266
rect 10146 15214 10148 15266
rect 10092 15212 10148 15214
rect 10412 15266 10468 15268
rect 10412 15214 10414 15266
rect 10414 15214 10466 15266
rect 10466 15214 10468 15266
rect 10412 15212 10468 15214
rect 10732 15266 10788 15268
rect 10732 15214 10734 15266
rect 10734 15214 10786 15266
rect 10786 15214 10788 15266
rect 10732 15212 10788 15214
rect 11052 15266 11108 15268
rect 11052 15214 11054 15266
rect 11054 15214 11106 15266
rect 11106 15214 11108 15266
rect 11052 15212 11108 15214
rect 11372 15266 11428 15268
rect 11372 15214 11374 15266
rect 11374 15214 11426 15266
rect 11426 15214 11428 15266
rect 11372 15212 11428 15214
rect 11532 15266 11588 15268
rect 11532 15214 11534 15266
rect 11534 15214 11586 15266
rect 11586 15214 11588 15266
rect 11532 15212 11588 15214
rect 11852 15266 11908 15268
rect 11852 15214 11854 15266
rect 11854 15214 11906 15266
rect 11906 15214 11908 15266
rect 11852 15212 11908 15214
rect 12012 15266 12068 15268
rect 12012 15214 12014 15266
rect 12014 15214 12066 15266
rect 12066 15214 12068 15266
rect 12012 15212 12068 15214
rect 12332 15266 12388 15268
rect 12332 15214 12334 15266
rect 12334 15214 12386 15266
rect 12386 15214 12388 15266
rect 12332 15212 12388 15214
rect 8492 15106 8548 15108
rect 8492 15054 8494 15106
rect 8494 15054 8546 15106
rect 8546 15054 8548 15106
rect 8492 15052 8548 15054
rect 8812 15106 8868 15108
rect 8812 15054 8814 15106
rect 8814 15054 8866 15106
rect 8866 15054 8868 15106
rect 8812 15052 8868 15054
rect 8972 15106 9028 15108
rect 8972 15054 8974 15106
rect 8974 15054 9026 15106
rect 9026 15054 9028 15106
rect 8972 15052 9028 15054
rect 9292 15106 9348 15108
rect 9292 15054 9294 15106
rect 9294 15054 9346 15106
rect 9346 15054 9348 15106
rect 9292 15052 9348 15054
rect 9452 15106 9508 15108
rect 9452 15054 9454 15106
rect 9454 15054 9506 15106
rect 9506 15054 9508 15106
rect 9452 15052 9508 15054
rect 9772 15106 9828 15108
rect 9772 15054 9774 15106
rect 9774 15054 9826 15106
rect 9826 15054 9828 15106
rect 9772 15052 9828 15054
rect 10092 15106 10148 15108
rect 10092 15054 10094 15106
rect 10094 15054 10146 15106
rect 10146 15054 10148 15106
rect 10092 15052 10148 15054
rect 10412 15106 10468 15108
rect 10412 15054 10414 15106
rect 10414 15054 10466 15106
rect 10466 15054 10468 15106
rect 10412 15052 10468 15054
rect 10732 15106 10788 15108
rect 10732 15054 10734 15106
rect 10734 15054 10786 15106
rect 10786 15054 10788 15106
rect 10732 15052 10788 15054
rect 11052 15106 11108 15108
rect 11052 15054 11054 15106
rect 11054 15054 11106 15106
rect 11106 15054 11108 15106
rect 11052 15052 11108 15054
rect 11372 15106 11428 15108
rect 11372 15054 11374 15106
rect 11374 15054 11426 15106
rect 11426 15054 11428 15106
rect 11372 15052 11428 15054
rect 11532 15106 11588 15108
rect 11532 15054 11534 15106
rect 11534 15054 11586 15106
rect 11586 15054 11588 15106
rect 11532 15052 11588 15054
rect 11852 15106 11908 15108
rect 11852 15054 11854 15106
rect 11854 15054 11906 15106
rect 11906 15054 11908 15106
rect 11852 15052 11908 15054
rect 12012 15106 12068 15108
rect 12012 15054 12014 15106
rect 12014 15054 12066 15106
rect 12066 15054 12068 15106
rect 12012 15052 12068 15054
rect 12332 15106 12388 15108
rect 12332 15054 12334 15106
rect 12334 15054 12386 15106
rect 12386 15054 12388 15106
rect 12332 15052 12388 15054
rect 8492 14946 8548 14948
rect 8492 14894 8494 14946
rect 8494 14894 8546 14946
rect 8546 14894 8548 14946
rect 8492 14892 8548 14894
rect 8812 14946 8868 14948
rect 8812 14894 8814 14946
rect 8814 14894 8866 14946
rect 8866 14894 8868 14946
rect 8812 14892 8868 14894
rect 8972 14946 9028 14948
rect 8972 14894 8974 14946
rect 8974 14894 9026 14946
rect 9026 14894 9028 14946
rect 8972 14892 9028 14894
rect 9292 14946 9348 14948
rect 9292 14894 9294 14946
rect 9294 14894 9346 14946
rect 9346 14894 9348 14946
rect 9292 14892 9348 14894
rect 9452 14946 9508 14948
rect 9452 14894 9454 14946
rect 9454 14894 9506 14946
rect 9506 14894 9508 14946
rect 9452 14892 9508 14894
rect 9772 14946 9828 14948
rect 9772 14894 9774 14946
rect 9774 14894 9826 14946
rect 9826 14894 9828 14946
rect 9772 14892 9828 14894
rect 10092 14946 10148 14948
rect 10092 14894 10094 14946
rect 10094 14894 10146 14946
rect 10146 14894 10148 14946
rect 10092 14892 10148 14894
rect 10412 14946 10468 14948
rect 10412 14894 10414 14946
rect 10414 14894 10466 14946
rect 10466 14894 10468 14946
rect 10412 14892 10468 14894
rect 10732 14946 10788 14948
rect 10732 14894 10734 14946
rect 10734 14894 10786 14946
rect 10786 14894 10788 14946
rect 10732 14892 10788 14894
rect 11052 14946 11108 14948
rect 11052 14894 11054 14946
rect 11054 14894 11106 14946
rect 11106 14894 11108 14946
rect 11052 14892 11108 14894
rect 11372 14946 11428 14948
rect 11372 14894 11374 14946
rect 11374 14894 11426 14946
rect 11426 14894 11428 14946
rect 11372 14892 11428 14894
rect 11532 14946 11588 14948
rect 11532 14894 11534 14946
rect 11534 14894 11586 14946
rect 11586 14894 11588 14946
rect 11532 14892 11588 14894
rect 11852 14946 11908 14948
rect 11852 14894 11854 14946
rect 11854 14894 11906 14946
rect 11906 14894 11908 14946
rect 11852 14892 11908 14894
rect 12012 14946 12068 14948
rect 12012 14894 12014 14946
rect 12014 14894 12066 14946
rect 12066 14894 12068 14946
rect 12012 14892 12068 14894
rect 12332 14946 12388 14948
rect 12332 14894 12334 14946
rect 12334 14894 12386 14946
rect 12386 14894 12388 14946
rect 12332 14892 12388 14894
rect 8492 14786 8548 14788
rect 8492 14734 8494 14786
rect 8494 14734 8546 14786
rect 8546 14734 8548 14786
rect 8492 14732 8548 14734
rect 8812 14786 8868 14788
rect 8812 14734 8814 14786
rect 8814 14734 8866 14786
rect 8866 14734 8868 14786
rect 8812 14732 8868 14734
rect 8972 14786 9028 14788
rect 8972 14734 8974 14786
rect 8974 14734 9026 14786
rect 9026 14734 9028 14786
rect 8972 14732 9028 14734
rect 9292 14786 9348 14788
rect 9292 14734 9294 14786
rect 9294 14734 9346 14786
rect 9346 14734 9348 14786
rect 9292 14732 9348 14734
rect 9452 14786 9508 14788
rect 9452 14734 9454 14786
rect 9454 14734 9506 14786
rect 9506 14734 9508 14786
rect 9452 14732 9508 14734
rect 9772 14786 9828 14788
rect 9772 14734 9774 14786
rect 9774 14734 9826 14786
rect 9826 14734 9828 14786
rect 9772 14732 9828 14734
rect 10092 14786 10148 14788
rect 10092 14734 10094 14786
rect 10094 14734 10146 14786
rect 10146 14734 10148 14786
rect 10092 14732 10148 14734
rect 10412 14786 10468 14788
rect 10412 14734 10414 14786
rect 10414 14734 10466 14786
rect 10466 14734 10468 14786
rect 10412 14732 10468 14734
rect 10732 14786 10788 14788
rect 10732 14734 10734 14786
rect 10734 14734 10786 14786
rect 10786 14734 10788 14786
rect 10732 14732 10788 14734
rect 11052 14786 11108 14788
rect 11052 14734 11054 14786
rect 11054 14734 11106 14786
rect 11106 14734 11108 14786
rect 11052 14732 11108 14734
rect 11372 14786 11428 14788
rect 11372 14734 11374 14786
rect 11374 14734 11426 14786
rect 11426 14734 11428 14786
rect 11372 14732 11428 14734
rect 11532 14786 11588 14788
rect 11532 14734 11534 14786
rect 11534 14734 11586 14786
rect 11586 14734 11588 14786
rect 11532 14732 11588 14734
rect 11852 14786 11908 14788
rect 11852 14734 11854 14786
rect 11854 14734 11906 14786
rect 11906 14734 11908 14786
rect 11852 14732 11908 14734
rect 12012 14786 12068 14788
rect 12012 14734 12014 14786
rect 12014 14734 12066 14786
rect 12066 14734 12068 14786
rect 12012 14732 12068 14734
rect 12332 14786 12388 14788
rect 12332 14734 12334 14786
rect 12334 14734 12386 14786
rect 12386 14734 12388 14786
rect 12332 14732 12388 14734
rect 8492 14626 8548 14628
rect 8492 14574 8494 14626
rect 8494 14574 8546 14626
rect 8546 14574 8548 14626
rect 8492 14572 8548 14574
rect 8812 14626 8868 14628
rect 8812 14574 8814 14626
rect 8814 14574 8866 14626
rect 8866 14574 8868 14626
rect 8812 14572 8868 14574
rect 8972 14626 9028 14628
rect 8972 14574 8974 14626
rect 8974 14574 9026 14626
rect 9026 14574 9028 14626
rect 8972 14572 9028 14574
rect 9292 14626 9348 14628
rect 9292 14574 9294 14626
rect 9294 14574 9346 14626
rect 9346 14574 9348 14626
rect 9292 14572 9348 14574
rect 9452 14626 9508 14628
rect 9452 14574 9454 14626
rect 9454 14574 9506 14626
rect 9506 14574 9508 14626
rect 9452 14572 9508 14574
rect 9772 14626 9828 14628
rect 9772 14574 9774 14626
rect 9774 14574 9826 14626
rect 9826 14574 9828 14626
rect 9772 14572 9828 14574
rect 10092 14626 10148 14628
rect 10092 14574 10094 14626
rect 10094 14574 10146 14626
rect 10146 14574 10148 14626
rect 10092 14572 10148 14574
rect 10412 14626 10468 14628
rect 10412 14574 10414 14626
rect 10414 14574 10466 14626
rect 10466 14574 10468 14626
rect 10412 14572 10468 14574
rect 10732 14626 10788 14628
rect 10732 14574 10734 14626
rect 10734 14574 10786 14626
rect 10786 14574 10788 14626
rect 10732 14572 10788 14574
rect 11052 14626 11108 14628
rect 11052 14574 11054 14626
rect 11054 14574 11106 14626
rect 11106 14574 11108 14626
rect 11052 14572 11108 14574
rect 11372 14626 11428 14628
rect 11372 14574 11374 14626
rect 11374 14574 11426 14626
rect 11426 14574 11428 14626
rect 11372 14572 11428 14574
rect 11532 14626 11588 14628
rect 11532 14574 11534 14626
rect 11534 14574 11586 14626
rect 11586 14574 11588 14626
rect 11532 14572 11588 14574
rect 11852 14626 11908 14628
rect 11852 14574 11854 14626
rect 11854 14574 11906 14626
rect 11906 14574 11908 14626
rect 11852 14572 11908 14574
rect 12012 14626 12068 14628
rect 12012 14574 12014 14626
rect 12014 14574 12066 14626
rect 12066 14574 12068 14626
rect 12012 14572 12068 14574
rect 12332 14626 12388 14628
rect 12332 14574 12334 14626
rect 12334 14574 12386 14626
rect 12386 14574 12388 14626
rect 12332 14572 12388 14574
rect 8492 14466 8548 14468
rect 8492 14414 8494 14466
rect 8494 14414 8546 14466
rect 8546 14414 8548 14466
rect 8492 14412 8548 14414
rect 8812 14466 8868 14468
rect 8812 14414 8814 14466
rect 8814 14414 8866 14466
rect 8866 14414 8868 14466
rect 8812 14412 8868 14414
rect 8972 14466 9028 14468
rect 8972 14414 8974 14466
rect 8974 14414 9026 14466
rect 9026 14414 9028 14466
rect 8972 14412 9028 14414
rect 9292 14466 9348 14468
rect 9292 14414 9294 14466
rect 9294 14414 9346 14466
rect 9346 14414 9348 14466
rect 9292 14412 9348 14414
rect 9452 14466 9508 14468
rect 9452 14414 9454 14466
rect 9454 14414 9506 14466
rect 9506 14414 9508 14466
rect 9452 14412 9508 14414
rect 9772 14466 9828 14468
rect 9772 14414 9774 14466
rect 9774 14414 9826 14466
rect 9826 14414 9828 14466
rect 9772 14412 9828 14414
rect 10092 14466 10148 14468
rect 10092 14414 10094 14466
rect 10094 14414 10146 14466
rect 10146 14414 10148 14466
rect 10092 14412 10148 14414
rect 10412 14466 10468 14468
rect 10412 14414 10414 14466
rect 10414 14414 10466 14466
rect 10466 14414 10468 14466
rect 10412 14412 10468 14414
rect 10732 14466 10788 14468
rect 10732 14414 10734 14466
rect 10734 14414 10786 14466
rect 10786 14414 10788 14466
rect 10732 14412 10788 14414
rect 11052 14466 11108 14468
rect 11052 14414 11054 14466
rect 11054 14414 11106 14466
rect 11106 14414 11108 14466
rect 11052 14412 11108 14414
rect 11372 14466 11428 14468
rect 11372 14414 11374 14466
rect 11374 14414 11426 14466
rect 11426 14414 11428 14466
rect 11372 14412 11428 14414
rect 11532 14466 11588 14468
rect 11532 14414 11534 14466
rect 11534 14414 11586 14466
rect 11586 14414 11588 14466
rect 11532 14412 11588 14414
rect 11852 14466 11908 14468
rect 11852 14414 11854 14466
rect 11854 14414 11906 14466
rect 11906 14414 11908 14466
rect 11852 14412 11908 14414
rect 12012 14466 12068 14468
rect 12012 14414 12014 14466
rect 12014 14414 12066 14466
rect 12066 14414 12068 14466
rect 12012 14412 12068 14414
rect 12332 14466 12388 14468
rect 12332 14414 12334 14466
rect 12334 14414 12386 14466
rect 12386 14414 12388 14466
rect 12332 14412 12388 14414
rect 8492 14306 8548 14308
rect 8492 14254 8494 14306
rect 8494 14254 8546 14306
rect 8546 14254 8548 14306
rect 8492 14252 8548 14254
rect 8812 14306 8868 14308
rect 8812 14254 8814 14306
rect 8814 14254 8866 14306
rect 8866 14254 8868 14306
rect 8812 14252 8868 14254
rect 8972 14306 9028 14308
rect 8972 14254 8974 14306
rect 8974 14254 9026 14306
rect 9026 14254 9028 14306
rect 8972 14252 9028 14254
rect 9292 14306 9348 14308
rect 9292 14254 9294 14306
rect 9294 14254 9346 14306
rect 9346 14254 9348 14306
rect 9292 14252 9348 14254
rect 9452 14306 9508 14308
rect 9452 14254 9454 14306
rect 9454 14254 9506 14306
rect 9506 14254 9508 14306
rect 9452 14252 9508 14254
rect 9772 14306 9828 14308
rect 9772 14254 9774 14306
rect 9774 14254 9826 14306
rect 9826 14254 9828 14306
rect 9772 14252 9828 14254
rect 10092 14306 10148 14308
rect 10092 14254 10094 14306
rect 10094 14254 10146 14306
rect 10146 14254 10148 14306
rect 10092 14252 10148 14254
rect 10412 14306 10468 14308
rect 10412 14254 10414 14306
rect 10414 14254 10466 14306
rect 10466 14254 10468 14306
rect 10412 14252 10468 14254
rect 10732 14306 10788 14308
rect 10732 14254 10734 14306
rect 10734 14254 10786 14306
rect 10786 14254 10788 14306
rect 10732 14252 10788 14254
rect 11052 14306 11108 14308
rect 11052 14254 11054 14306
rect 11054 14254 11106 14306
rect 11106 14254 11108 14306
rect 11052 14252 11108 14254
rect 11372 14306 11428 14308
rect 11372 14254 11374 14306
rect 11374 14254 11426 14306
rect 11426 14254 11428 14306
rect 11372 14252 11428 14254
rect 11532 14306 11588 14308
rect 11532 14254 11534 14306
rect 11534 14254 11586 14306
rect 11586 14254 11588 14306
rect 11532 14252 11588 14254
rect 11852 14306 11908 14308
rect 11852 14254 11854 14306
rect 11854 14254 11906 14306
rect 11906 14254 11908 14306
rect 11852 14252 11908 14254
rect 12012 14306 12068 14308
rect 12012 14254 12014 14306
rect 12014 14254 12066 14306
rect 12066 14254 12068 14306
rect 12012 14252 12068 14254
rect 12332 14306 12388 14308
rect 12332 14254 12334 14306
rect 12334 14254 12386 14306
rect 12386 14254 12388 14306
rect 12332 14252 12388 14254
rect 8492 14146 8548 14148
rect 8492 14094 8494 14146
rect 8494 14094 8546 14146
rect 8546 14094 8548 14146
rect 8492 14092 8548 14094
rect 8812 14146 8868 14148
rect 8812 14094 8814 14146
rect 8814 14094 8866 14146
rect 8866 14094 8868 14146
rect 8812 14092 8868 14094
rect 8972 14146 9028 14148
rect 8972 14094 8974 14146
rect 8974 14094 9026 14146
rect 9026 14094 9028 14146
rect 8972 14092 9028 14094
rect 9292 14146 9348 14148
rect 9292 14094 9294 14146
rect 9294 14094 9346 14146
rect 9346 14094 9348 14146
rect 9292 14092 9348 14094
rect 9452 14146 9508 14148
rect 9452 14094 9454 14146
rect 9454 14094 9506 14146
rect 9506 14094 9508 14146
rect 9452 14092 9508 14094
rect 9772 14146 9828 14148
rect 9772 14094 9774 14146
rect 9774 14094 9826 14146
rect 9826 14094 9828 14146
rect 9772 14092 9828 14094
rect 10092 14146 10148 14148
rect 10092 14094 10094 14146
rect 10094 14094 10146 14146
rect 10146 14094 10148 14146
rect 10092 14092 10148 14094
rect 10412 14146 10468 14148
rect 10412 14094 10414 14146
rect 10414 14094 10466 14146
rect 10466 14094 10468 14146
rect 10412 14092 10468 14094
rect 10732 14146 10788 14148
rect 10732 14094 10734 14146
rect 10734 14094 10786 14146
rect 10786 14094 10788 14146
rect 10732 14092 10788 14094
rect 11052 14146 11108 14148
rect 11052 14094 11054 14146
rect 11054 14094 11106 14146
rect 11106 14094 11108 14146
rect 11052 14092 11108 14094
rect 11372 14146 11428 14148
rect 11372 14094 11374 14146
rect 11374 14094 11426 14146
rect 11426 14094 11428 14146
rect 11372 14092 11428 14094
rect 11532 14146 11588 14148
rect 11532 14094 11534 14146
rect 11534 14094 11586 14146
rect 11586 14094 11588 14146
rect 11532 14092 11588 14094
rect 11852 14146 11908 14148
rect 11852 14094 11854 14146
rect 11854 14094 11906 14146
rect 11906 14094 11908 14146
rect 11852 14092 11908 14094
rect 12012 14146 12068 14148
rect 12012 14094 12014 14146
rect 12014 14094 12066 14146
rect 12066 14094 12068 14146
rect 12012 14092 12068 14094
rect 12332 14146 12388 14148
rect 12332 14094 12334 14146
rect 12334 14094 12386 14146
rect 12386 14094 12388 14146
rect 12332 14092 12388 14094
rect 8492 13986 8548 13988
rect 8492 13934 8494 13986
rect 8494 13934 8546 13986
rect 8546 13934 8548 13986
rect 8492 13932 8548 13934
rect 8812 13986 8868 13988
rect 8812 13934 8814 13986
rect 8814 13934 8866 13986
rect 8866 13934 8868 13986
rect 8812 13932 8868 13934
rect 8972 13986 9028 13988
rect 8972 13934 8974 13986
rect 8974 13934 9026 13986
rect 9026 13934 9028 13986
rect 8972 13932 9028 13934
rect 9292 13986 9348 13988
rect 9292 13934 9294 13986
rect 9294 13934 9346 13986
rect 9346 13934 9348 13986
rect 9292 13932 9348 13934
rect 9452 13986 9508 13988
rect 9452 13934 9454 13986
rect 9454 13934 9506 13986
rect 9506 13934 9508 13986
rect 9452 13932 9508 13934
rect 9772 13986 9828 13988
rect 9772 13934 9774 13986
rect 9774 13934 9826 13986
rect 9826 13934 9828 13986
rect 9772 13932 9828 13934
rect 10092 13986 10148 13988
rect 10092 13934 10094 13986
rect 10094 13934 10146 13986
rect 10146 13934 10148 13986
rect 10092 13932 10148 13934
rect 10412 13986 10468 13988
rect 10412 13934 10414 13986
rect 10414 13934 10466 13986
rect 10466 13934 10468 13986
rect 10412 13932 10468 13934
rect 10732 13986 10788 13988
rect 10732 13934 10734 13986
rect 10734 13934 10786 13986
rect 10786 13934 10788 13986
rect 10732 13932 10788 13934
rect 11052 13986 11108 13988
rect 11052 13934 11054 13986
rect 11054 13934 11106 13986
rect 11106 13934 11108 13986
rect 11052 13932 11108 13934
rect 11372 13986 11428 13988
rect 11372 13934 11374 13986
rect 11374 13934 11426 13986
rect 11426 13934 11428 13986
rect 11372 13932 11428 13934
rect 11532 13986 11588 13988
rect 11532 13934 11534 13986
rect 11534 13934 11586 13986
rect 11586 13934 11588 13986
rect 11532 13932 11588 13934
rect 11852 13986 11908 13988
rect 11852 13934 11854 13986
rect 11854 13934 11906 13986
rect 11906 13934 11908 13986
rect 11852 13932 11908 13934
rect 12012 13986 12068 13988
rect 12012 13934 12014 13986
rect 12014 13934 12066 13986
rect 12066 13934 12068 13986
rect 12012 13932 12068 13934
rect 12332 13986 12388 13988
rect 12332 13934 12334 13986
rect 12334 13934 12386 13986
rect 12386 13934 12388 13986
rect 12332 13932 12388 13934
rect 9132 13772 9188 13828
rect 8492 13666 8548 13668
rect 8492 13614 8494 13666
rect 8494 13614 8546 13666
rect 8546 13614 8548 13666
rect 8492 13612 8548 13614
rect 8812 13666 8868 13668
rect 8812 13614 8814 13666
rect 8814 13614 8866 13666
rect 8866 13614 8868 13666
rect 8812 13612 8868 13614
rect 8972 13666 9028 13668
rect 8972 13614 8974 13666
rect 8974 13614 9026 13666
rect 9026 13614 9028 13666
rect 8972 13612 9028 13614
rect 9292 13666 9348 13668
rect 9292 13614 9294 13666
rect 9294 13614 9346 13666
rect 9346 13614 9348 13666
rect 9292 13612 9348 13614
rect 9452 13666 9508 13668
rect 9452 13614 9454 13666
rect 9454 13614 9506 13666
rect 9506 13614 9508 13666
rect 9452 13612 9508 13614
rect 9772 13666 9828 13668
rect 9772 13614 9774 13666
rect 9774 13614 9826 13666
rect 9826 13614 9828 13666
rect 9772 13612 9828 13614
rect 10092 13666 10148 13668
rect 10092 13614 10094 13666
rect 10094 13614 10146 13666
rect 10146 13614 10148 13666
rect 10092 13612 10148 13614
rect 10412 13666 10468 13668
rect 10412 13614 10414 13666
rect 10414 13614 10466 13666
rect 10466 13614 10468 13666
rect 10412 13612 10468 13614
rect 10732 13666 10788 13668
rect 10732 13614 10734 13666
rect 10734 13614 10786 13666
rect 10786 13614 10788 13666
rect 10732 13612 10788 13614
rect 11052 13666 11108 13668
rect 11052 13614 11054 13666
rect 11054 13614 11106 13666
rect 11106 13614 11108 13666
rect 11052 13612 11108 13614
rect 11372 13666 11428 13668
rect 11372 13614 11374 13666
rect 11374 13614 11426 13666
rect 11426 13614 11428 13666
rect 11372 13612 11428 13614
rect 11532 13666 11588 13668
rect 11532 13614 11534 13666
rect 11534 13614 11586 13666
rect 11586 13614 11588 13666
rect 11532 13612 11588 13614
rect 11852 13666 11908 13668
rect 11852 13614 11854 13666
rect 11854 13614 11906 13666
rect 11906 13614 11908 13666
rect 11852 13612 11908 13614
rect 12012 13666 12068 13668
rect 12012 13614 12014 13666
rect 12014 13614 12066 13666
rect 12066 13614 12068 13666
rect 12012 13612 12068 13614
rect 12332 13666 12388 13668
rect 12332 13614 12334 13666
rect 12334 13614 12386 13666
rect 12386 13614 12388 13666
rect 12332 13612 12388 13614
rect 8492 13506 8548 13508
rect 8492 13454 8494 13506
rect 8494 13454 8546 13506
rect 8546 13454 8548 13506
rect 8492 13452 8548 13454
rect 8812 13506 8868 13508
rect 8812 13454 8814 13506
rect 8814 13454 8866 13506
rect 8866 13454 8868 13506
rect 8812 13452 8868 13454
rect 8972 13506 9028 13508
rect 8972 13454 8974 13506
rect 8974 13454 9026 13506
rect 9026 13454 9028 13506
rect 8972 13452 9028 13454
rect 9292 13506 9348 13508
rect 9292 13454 9294 13506
rect 9294 13454 9346 13506
rect 9346 13454 9348 13506
rect 9292 13452 9348 13454
rect 9452 13506 9508 13508
rect 9452 13454 9454 13506
rect 9454 13454 9506 13506
rect 9506 13454 9508 13506
rect 9452 13452 9508 13454
rect 9772 13506 9828 13508
rect 9772 13454 9774 13506
rect 9774 13454 9826 13506
rect 9826 13454 9828 13506
rect 9772 13452 9828 13454
rect 10092 13506 10148 13508
rect 10092 13454 10094 13506
rect 10094 13454 10146 13506
rect 10146 13454 10148 13506
rect 10092 13452 10148 13454
rect 10412 13506 10468 13508
rect 10412 13454 10414 13506
rect 10414 13454 10466 13506
rect 10466 13454 10468 13506
rect 10412 13452 10468 13454
rect 10732 13506 10788 13508
rect 10732 13454 10734 13506
rect 10734 13454 10786 13506
rect 10786 13454 10788 13506
rect 10732 13452 10788 13454
rect 11052 13506 11108 13508
rect 11052 13454 11054 13506
rect 11054 13454 11106 13506
rect 11106 13454 11108 13506
rect 11052 13452 11108 13454
rect 11372 13506 11428 13508
rect 11372 13454 11374 13506
rect 11374 13454 11426 13506
rect 11426 13454 11428 13506
rect 11372 13452 11428 13454
rect 11532 13506 11588 13508
rect 11532 13454 11534 13506
rect 11534 13454 11586 13506
rect 11586 13454 11588 13506
rect 11532 13452 11588 13454
rect 11852 13506 11908 13508
rect 11852 13454 11854 13506
rect 11854 13454 11906 13506
rect 11906 13454 11908 13506
rect 11852 13452 11908 13454
rect 12012 13506 12068 13508
rect 12012 13454 12014 13506
rect 12014 13454 12066 13506
rect 12066 13454 12068 13506
rect 12012 13452 12068 13454
rect 12332 13506 12388 13508
rect 12332 13454 12334 13506
rect 12334 13454 12386 13506
rect 12386 13454 12388 13506
rect 12332 13452 12388 13454
rect 8492 13346 8548 13348
rect 8492 13294 8494 13346
rect 8494 13294 8546 13346
rect 8546 13294 8548 13346
rect 8492 13292 8548 13294
rect 8812 13346 8868 13348
rect 8812 13294 8814 13346
rect 8814 13294 8866 13346
rect 8866 13294 8868 13346
rect 8812 13292 8868 13294
rect 8972 13346 9028 13348
rect 8972 13294 8974 13346
rect 8974 13294 9026 13346
rect 9026 13294 9028 13346
rect 8972 13292 9028 13294
rect 9292 13346 9348 13348
rect 9292 13294 9294 13346
rect 9294 13294 9346 13346
rect 9346 13294 9348 13346
rect 9292 13292 9348 13294
rect 9452 13346 9508 13348
rect 9452 13294 9454 13346
rect 9454 13294 9506 13346
rect 9506 13294 9508 13346
rect 9452 13292 9508 13294
rect 9772 13346 9828 13348
rect 9772 13294 9774 13346
rect 9774 13294 9826 13346
rect 9826 13294 9828 13346
rect 9772 13292 9828 13294
rect 10092 13346 10148 13348
rect 10092 13294 10094 13346
rect 10094 13294 10146 13346
rect 10146 13294 10148 13346
rect 10092 13292 10148 13294
rect 10412 13346 10468 13348
rect 10412 13294 10414 13346
rect 10414 13294 10466 13346
rect 10466 13294 10468 13346
rect 10412 13292 10468 13294
rect 10732 13346 10788 13348
rect 10732 13294 10734 13346
rect 10734 13294 10786 13346
rect 10786 13294 10788 13346
rect 10732 13292 10788 13294
rect 11052 13346 11108 13348
rect 11052 13294 11054 13346
rect 11054 13294 11106 13346
rect 11106 13294 11108 13346
rect 11052 13292 11108 13294
rect 11372 13346 11428 13348
rect 11372 13294 11374 13346
rect 11374 13294 11426 13346
rect 11426 13294 11428 13346
rect 11372 13292 11428 13294
rect 11532 13346 11588 13348
rect 11532 13294 11534 13346
rect 11534 13294 11586 13346
rect 11586 13294 11588 13346
rect 11532 13292 11588 13294
rect 11852 13346 11908 13348
rect 11852 13294 11854 13346
rect 11854 13294 11906 13346
rect 11906 13294 11908 13346
rect 11852 13292 11908 13294
rect 12012 13346 12068 13348
rect 12012 13294 12014 13346
rect 12014 13294 12066 13346
rect 12066 13294 12068 13346
rect 12012 13292 12068 13294
rect 12332 13346 12388 13348
rect 12332 13294 12334 13346
rect 12334 13294 12386 13346
rect 12386 13294 12388 13346
rect 12332 13292 12388 13294
rect 8492 13186 8548 13188
rect 8492 13134 8494 13186
rect 8494 13134 8546 13186
rect 8546 13134 8548 13186
rect 8492 13132 8548 13134
rect 8812 13186 8868 13188
rect 8812 13134 8814 13186
rect 8814 13134 8866 13186
rect 8866 13134 8868 13186
rect 8812 13132 8868 13134
rect 8972 13186 9028 13188
rect 8972 13134 8974 13186
rect 8974 13134 9026 13186
rect 9026 13134 9028 13186
rect 8972 13132 9028 13134
rect 9292 13186 9348 13188
rect 9292 13134 9294 13186
rect 9294 13134 9346 13186
rect 9346 13134 9348 13186
rect 9292 13132 9348 13134
rect 9452 13186 9508 13188
rect 9452 13134 9454 13186
rect 9454 13134 9506 13186
rect 9506 13134 9508 13186
rect 9452 13132 9508 13134
rect 9772 13186 9828 13188
rect 9772 13134 9774 13186
rect 9774 13134 9826 13186
rect 9826 13134 9828 13186
rect 9772 13132 9828 13134
rect 10092 13186 10148 13188
rect 10092 13134 10094 13186
rect 10094 13134 10146 13186
rect 10146 13134 10148 13186
rect 10092 13132 10148 13134
rect 10412 13186 10468 13188
rect 10412 13134 10414 13186
rect 10414 13134 10466 13186
rect 10466 13134 10468 13186
rect 10412 13132 10468 13134
rect 10732 13186 10788 13188
rect 10732 13134 10734 13186
rect 10734 13134 10786 13186
rect 10786 13134 10788 13186
rect 10732 13132 10788 13134
rect 11052 13186 11108 13188
rect 11052 13134 11054 13186
rect 11054 13134 11106 13186
rect 11106 13134 11108 13186
rect 11052 13132 11108 13134
rect 11372 13186 11428 13188
rect 11372 13134 11374 13186
rect 11374 13134 11426 13186
rect 11426 13134 11428 13186
rect 11372 13132 11428 13134
rect 11532 13186 11588 13188
rect 11532 13134 11534 13186
rect 11534 13134 11586 13186
rect 11586 13134 11588 13186
rect 11532 13132 11588 13134
rect 11852 13186 11908 13188
rect 11852 13134 11854 13186
rect 11854 13134 11906 13186
rect 11906 13134 11908 13186
rect 11852 13132 11908 13134
rect 12012 13186 12068 13188
rect 12012 13134 12014 13186
rect 12014 13134 12066 13186
rect 12066 13134 12068 13186
rect 12012 13132 12068 13134
rect 12332 13186 12388 13188
rect 12332 13134 12334 13186
rect 12334 13134 12386 13186
rect 12386 13134 12388 13186
rect 12332 13132 12388 13134
rect 8492 13026 8548 13028
rect 8492 12974 8494 13026
rect 8494 12974 8546 13026
rect 8546 12974 8548 13026
rect 8492 12972 8548 12974
rect 8812 13026 8868 13028
rect 8812 12974 8814 13026
rect 8814 12974 8866 13026
rect 8866 12974 8868 13026
rect 8812 12972 8868 12974
rect 8972 13026 9028 13028
rect 8972 12974 8974 13026
rect 8974 12974 9026 13026
rect 9026 12974 9028 13026
rect 8972 12972 9028 12974
rect 9292 13026 9348 13028
rect 9292 12974 9294 13026
rect 9294 12974 9346 13026
rect 9346 12974 9348 13026
rect 9292 12972 9348 12974
rect 9452 13026 9508 13028
rect 9452 12974 9454 13026
rect 9454 12974 9506 13026
rect 9506 12974 9508 13026
rect 9452 12972 9508 12974
rect 9772 13026 9828 13028
rect 9772 12974 9774 13026
rect 9774 12974 9826 13026
rect 9826 12974 9828 13026
rect 9772 12972 9828 12974
rect 10092 13026 10148 13028
rect 10092 12974 10094 13026
rect 10094 12974 10146 13026
rect 10146 12974 10148 13026
rect 10092 12972 10148 12974
rect 10412 13026 10468 13028
rect 10412 12974 10414 13026
rect 10414 12974 10466 13026
rect 10466 12974 10468 13026
rect 10412 12972 10468 12974
rect 10732 13026 10788 13028
rect 10732 12974 10734 13026
rect 10734 12974 10786 13026
rect 10786 12974 10788 13026
rect 10732 12972 10788 12974
rect 11052 13026 11108 13028
rect 11052 12974 11054 13026
rect 11054 12974 11106 13026
rect 11106 12974 11108 13026
rect 11052 12972 11108 12974
rect 11372 13026 11428 13028
rect 11372 12974 11374 13026
rect 11374 12974 11426 13026
rect 11426 12974 11428 13026
rect 11372 12972 11428 12974
rect 11532 13026 11588 13028
rect 11532 12974 11534 13026
rect 11534 12974 11586 13026
rect 11586 12974 11588 13026
rect 11532 12972 11588 12974
rect 11852 13026 11908 13028
rect 11852 12974 11854 13026
rect 11854 12974 11906 13026
rect 11906 12974 11908 13026
rect 11852 12972 11908 12974
rect 12012 13026 12068 13028
rect 12012 12974 12014 13026
rect 12014 12974 12066 13026
rect 12066 12974 12068 13026
rect 12012 12972 12068 12974
rect 12332 13026 12388 13028
rect 12332 12974 12334 13026
rect 12334 12974 12386 13026
rect 12386 12974 12388 13026
rect 12332 12972 12388 12974
rect 8492 12866 8548 12868
rect 8492 12814 8494 12866
rect 8494 12814 8546 12866
rect 8546 12814 8548 12866
rect 8492 12812 8548 12814
rect 8812 12866 8868 12868
rect 8812 12814 8814 12866
rect 8814 12814 8866 12866
rect 8866 12814 8868 12866
rect 8812 12812 8868 12814
rect 8972 12866 9028 12868
rect 8972 12814 8974 12866
rect 8974 12814 9026 12866
rect 9026 12814 9028 12866
rect 8972 12812 9028 12814
rect 9292 12866 9348 12868
rect 9292 12814 9294 12866
rect 9294 12814 9346 12866
rect 9346 12814 9348 12866
rect 9292 12812 9348 12814
rect 9452 12866 9508 12868
rect 9452 12814 9454 12866
rect 9454 12814 9506 12866
rect 9506 12814 9508 12866
rect 9452 12812 9508 12814
rect 9772 12866 9828 12868
rect 9772 12814 9774 12866
rect 9774 12814 9826 12866
rect 9826 12814 9828 12866
rect 9772 12812 9828 12814
rect 10092 12866 10148 12868
rect 10092 12814 10094 12866
rect 10094 12814 10146 12866
rect 10146 12814 10148 12866
rect 10092 12812 10148 12814
rect 10412 12866 10468 12868
rect 10412 12814 10414 12866
rect 10414 12814 10466 12866
rect 10466 12814 10468 12866
rect 10412 12812 10468 12814
rect 10732 12866 10788 12868
rect 10732 12814 10734 12866
rect 10734 12814 10786 12866
rect 10786 12814 10788 12866
rect 10732 12812 10788 12814
rect 11052 12866 11108 12868
rect 11052 12814 11054 12866
rect 11054 12814 11106 12866
rect 11106 12814 11108 12866
rect 11052 12812 11108 12814
rect 11372 12866 11428 12868
rect 11372 12814 11374 12866
rect 11374 12814 11426 12866
rect 11426 12814 11428 12866
rect 11372 12812 11428 12814
rect 11532 12866 11588 12868
rect 11532 12814 11534 12866
rect 11534 12814 11586 12866
rect 11586 12814 11588 12866
rect 11532 12812 11588 12814
rect 11852 12866 11908 12868
rect 11852 12814 11854 12866
rect 11854 12814 11906 12866
rect 11906 12814 11908 12866
rect 11852 12812 11908 12814
rect 12012 12866 12068 12868
rect 12012 12814 12014 12866
rect 12014 12814 12066 12866
rect 12066 12814 12068 12866
rect 12012 12812 12068 12814
rect 12332 12866 12388 12868
rect 12332 12814 12334 12866
rect 12334 12814 12386 12866
rect 12386 12814 12388 12866
rect 12332 12812 12388 12814
rect 8492 12706 8548 12708
rect 8492 12654 8494 12706
rect 8494 12654 8546 12706
rect 8546 12654 8548 12706
rect 8492 12652 8548 12654
rect 8812 12706 8868 12708
rect 8812 12654 8814 12706
rect 8814 12654 8866 12706
rect 8866 12654 8868 12706
rect 8812 12652 8868 12654
rect 8972 12706 9028 12708
rect 8972 12654 8974 12706
rect 8974 12654 9026 12706
rect 9026 12654 9028 12706
rect 8972 12652 9028 12654
rect 9292 12706 9348 12708
rect 9292 12654 9294 12706
rect 9294 12654 9346 12706
rect 9346 12654 9348 12706
rect 9292 12652 9348 12654
rect 9452 12706 9508 12708
rect 9452 12654 9454 12706
rect 9454 12654 9506 12706
rect 9506 12654 9508 12706
rect 9452 12652 9508 12654
rect 9772 12706 9828 12708
rect 9772 12654 9774 12706
rect 9774 12654 9826 12706
rect 9826 12654 9828 12706
rect 9772 12652 9828 12654
rect 10092 12706 10148 12708
rect 10092 12654 10094 12706
rect 10094 12654 10146 12706
rect 10146 12654 10148 12706
rect 10092 12652 10148 12654
rect 10412 12706 10468 12708
rect 10412 12654 10414 12706
rect 10414 12654 10466 12706
rect 10466 12654 10468 12706
rect 10412 12652 10468 12654
rect 10732 12706 10788 12708
rect 10732 12654 10734 12706
rect 10734 12654 10786 12706
rect 10786 12654 10788 12706
rect 10732 12652 10788 12654
rect 11052 12706 11108 12708
rect 11052 12654 11054 12706
rect 11054 12654 11106 12706
rect 11106 12654 11108 12706
rect 11052 12652 11108 12654
rect 11372 12706 11428 12708
rect 11372 12654 11374 12706
rect 11374 12654 11426 12706
rect 11426 12654 11428 12706
rect 11372 12652 11428 12654
rect 11532 12706 11588 12708
rect 11532 12654 11534 12706
rect 11534 12654 11586 12706
rect 11586 12654 11588 12706
rect 11532 12652 11588 12654
rect 11852 12706 11908 12708
rect 11852 12654 11854 12706
rect 11854 12654 11906 12706
rect 11906 12654 11908 12706
rect 11852 12652 11908 12654
rect 12012 12706 12068 12708
rect 12012 12654 12014 12706
rect 12014 12654 12066 12706
rect 12066 12654 12068 12706
rect 12012 12652 12068 12654
rect 12332 12706 12388 12708
rect 12332 12654 12334 12706
rect 12334 12654 12386 12706
rect 12386 12654 12388 12706
rect 12332 12652 12388 12654
rect 8492 12546 8548 12548
rect 8492 12494 8494 12546
rect 8494 12494 8546 12546
rect 8546 12494 8548 12546
rect 8492 12492 8548 12494
rect 8812 12546 8868 12548
rect 8812 12494 8814 12546
rect 8814 12494 8866 12546
rect 8866 12494 8868 12546
rect 8812 12492 8868 12494
rect 8972 12546 9028 12548
rect 8972 12494 8974 12546
rect 8974 12494 9026 12546
rect 9026 12494 9028 12546
rect 8972 12492 9028 12494
rect 9292 12546 9348 12548
rect 9292 12494 9294 12546
rect 9294 12494 9346 12546
rect 9346 12494 9348 12546
rect 9292 12492 9348 12494
rect 9452 12546 9508 12548
rect 9452 12494 9454 12546
rect 9454 12494 9506 12546
rect 9506 12494 9508 12546
rect 9452 12492 9508 12494
rect 9772 12546 9828 12548
rect 9772 12494 9774 12546
rect 9774 12494 9826 12546
rect 9826 12494 9828 12546
rect 9772 12492 9828 12494
rect 10092 12546 10148 12548
rect 10092 12494 10094 12546
rect 10094 12494 10146 12546
rect 10146 12494 10148 12546
rect 10092 12492 10148 12494
rect 10412 12546 10468 12548
rect 10412 12494 10414 12546
rect 10414 12494 10466 12546
rect 10466 12494 10468 12546
rect 10412 12492 10468 12494
rect 10732 12546 10788 12548
rect 10732 12494 10734 12546
rect 10734 12494 10786 12546
rect 10786 12494 10788 12546
rect 10732 12492 10788 12494
rect 11052 12546 11108 12548
rect 11052 12494 11054 12546
rect 11054 12494 11106 12546
rect 11106 12494 11108 12546
rect 11052 12492 11108 12494
rect 11372 12546 11428 12548
rect 11372 12494 11374 12546
rect 11374 12494 11426 12546
rect 11426 12494 11428 12546
rect 11372 12492 11428 12494
rect 11532 12546 11588 12548
rect 11532 12494 11534 12546
rect 11534 12494 11586 12546
rect 11586 12494 11588 12546
rect 11532 12492 11588 12494
rect 11852 12546 11908 12548
rect 11852 12494 11854 12546
rect 11854 12494 11906 12546
rect 11906 12494 11908 12546
rect 11852 12492 11908 12494
rect 12012 12546 12068 12548
rect 12012 12494 12014 12546
rect 12014 12494 12066 12546
rect 12066 12494 12068 12546
rect 12012 12492 12068 12494
rect 12332 12546 12388 12548
rect 12332 12494 12334 12546
rect 12334 12494 12386 12546
rect 12386 12494 12388 12546
rect 12332 12492 12388 12494
rect 9612 12252 9668 12308
rect 11212 12252 11268 12308
rect 9932 11932 9988 11988
rect 10892 11932 10948 11988
rect 8492 11746 8548 11748
rect 8492 11694 8494 11746
rect 8494 11694 8546 11746
rect 8546 11694 8548 11746
rect 8492 11692 8548 11694
rect 8812 11746 8868 11748
rect 8812 11694 8814 11746
rect 8814 11694 8866 11746
rect 8866 11694 8868 11746
rect 8812 11692 8868 11694
rect 8972 11746 9028 11748
rect 8972 11694 8974 11746
rect 8974 11694 9026 11746
rect 9026 11694 9028 11746
rect 8972 11692 9028 11694
rect 9292 11746 9348 11748
rect 9292 11694 9294 11746
rect 9294 11694 9346 11746
rect 9346 11694 9348 11746
rect 9292 11692 9348 11694
rect 9452 11746 9508 11748
rect 9452 11694 9454 11746
rect 9454 11694 9506 11746
rect 9506 11694 9508 11746
rect 9452 11692 9508 11694
rect 9772 11746 9828 11748
rect 9772 11694 9774 11746
rect 9774 11694 9826 11746
rect 9826 11694 9828 11746
rect 9772 11692 9828 11694
rect 10092 11746 10148 11748
rect 10092 11694 10094 11746
rect 10094 11694 10146 11746
rect 10146 11694 10148 11746
rect 10092 11692 10148 11694
rect 10412 11746 10468 11748
rect 10412 11694 10414 11746
rect 10414 11694 10466 11746
rect 10466 11694 10468 11746
rect 10412 11692 10468 11694
rect 10732 11746 10788 11748
rect 10732 11694 10734 11746
rect 10734 11694 10786 11746
rect 10786 11694 10788 11746
rect 10732 11692 10788 11694
rect 11052 11746 11108 11748
rect 11052 11694 11054 11746
rect 11054 11694 11106 11746
rect 11106 11694 11108 11746
rect 11052 11692 11108 11694
rect 11372 11746 11428 11748
rect 11372 11694 11374 11746
rect 11374 11694 11426 11746
rect 11426 11694 11428 11746
rect 11372 11692 11428 11694
rect 11532 11746 11588 11748
rect 11532 11694 11534 11746
rect 11534 11694 11586 11746
rect 11586 11694 11588 11746
rect 11532 11692 11588 11694
rect 11852 11746 11908 11748
rect 11852 11694 11854 11746
rect 11854 11694 11906 11746
rect 11906 11694 11908 11746
rect 11852 11692 11908 11694
rect 12012 11746 12068 11748
rect 12012 11694 12014 11746
rect 12014 11694 12066 11746
rect 12066 11694 12068 11746
rect 12012 11692 12068 11694
rect 12332 11746 12388 11748
rect 12332 11694 12334 11746
rect 12334 11694 12386 11746
rect 12386 11694 12388 11746
rect 12332 11692 12388 11694
rect 8492 11586 8548 11588
rect 8492 11534 8494 11586
rect 8494 11534 8546 11586
rect 8546 11534 8548 11586
rect 8492 11532 8548 11534
rect 8812 11586 8868 11588
rect 8812 11534 8814 11586
rect 8814 11534 8866 11586
rect 8866 11534 8868 11586
rect 8812 11532 8868 11534
rect 8972 11586 9028 11588
rect 8972 11534 8974 11586
rect 8974 11534 9026 11586
rect 9026 11534 9028 11586
rect 8972 11532 9028 11534
rect 9292 11586 9348 11588
rect 9292 11534 9294 11586
rect 9294 11534 9346 11586
rect 9346 11534 9348 11586
rect 9292 11532 9348 11534
rect 9452 11586 9508 11588
rect 9452 11534 9454 11586
rect 9454 11534 9506 11586
rect 9506 11534 9508 11586
rect 9452 11532 9508 11534
rect 9772 11586 9828 11588
rect 9772 11534 9774 11586
rect 9774 11534 9826 11586
rect 9826 11534 9828 11586
rect 9772 11532 9828 11534
rect 10092 11586 10148 11588
rect 10092 11534 10094 11586
rect 10094 11534 10146 11586
rect 10146 11534 10148 11586
rect 10092 11532 10148 11534
rect 10412 11586 10468 11588
rect 10412 11534 10414 11586
rect 10414 11534 10466 11586
rect 10466 11534 10468 11586
rect 10412 11532 10468 11534
rect 10732 11586 10788 11588
rect 10732 11534 10734 11586
rect 10734 11534 10786 11586
rect 10786 11534 10788 11586
rect 10732 11532 10788 11534
rect 11052 11586 11108 11588
rect 11052 11534 11054 11586
rect 11054 11534 11106 11586
rect 11106 11534 11108 11586
rect 11052 11532 11108 11534
rect 11372 11586 11428 11588
rect 11372 11534 11374 11586
rect 11374 11534 11426 11586
rect 11426 11534 11428 11586
rect 11372 11532 11428 11534
rect 11532 11586 11588 11588
rect 11532 11534 11534 11586
rect 11534 11534 11586 11586
rect 11586 11534 11588 11586
rect 11532 11532 11588 11534
rect 11852 11586 11908 11588
rect 11852 11534 11854 11586
rect 11854 11534 11906 11586
rect 11906 11534 11908 11586
rect 11852 11532 11908 11534
rect 12012 11586 12068 11588
rect 12012 11534 12014 11586
rect 12014 11534 12066 11586
rect 12066 11534 12068 11586
rect 12012 11532 12068 11534
rect 12332 11586 12388 11588
rect 12332 11534 12334 11586
rect 12334 11534 12386 11586
rect 12386 11534 12388 11586
rect 12332 11532 12388 11534
rect 8492 11426 8548 11428
rect 8492 11374 8494 11426
rect 8494 11374 8546 11426
rect 8546 11374 8548 11426
rect 8492 11372 8548 11374
rect 8812 11426 8868 11428
rect 8812 11374 8814 11426
rect 8814 11374 8866 11426
rect 8866 11374 8868 11426
rect 8812 11372 8868 11374
rect 8972 11426 9028 11428
rect 8972 11374 8974 11426
rect 8974 11374 9026 11426
rect 9026 11374 9028 11426
rect 8972 11372 9028 11374
rect 9292 11426 9348 11428
rect 9292 11374 9294 11426
rect 9294 11374 9346 11426
rect 9346 11374 9348 11426
rect 9292 11372 9348 11374
rect 9452 11426 9508 11428
rect 9452 11374 9454 11426
rect 9454 11374 9506 11426
rect 9506 11374 9508 11426
rect 9452 11372 9508 11374
rect 9772 11426 9828 11428
rect 9772 11374 9774 11426
rect 9774 11374 9826 11426
rect 9826 11374 9828 11426
rect 9772 11372 9828 11374
rect 10092 11426 10148 11428
rect 10092 11374 10094 11426
rect 10094 11374 10146 11426
rect 10146 11374 10148 11426
rect 10092 11372 10148 11374
rect 10412 11426 10468 11428
rect 10412 11374 10414 11426
rect 10414 11374 10466 11426
rect 10466 11374 10468 11426
rect 10412 11372 10468 11374
rect 10732 11426 10788 11428
rect 10732 11374 10734 11426
rect 10734 11374 10786 11426
rect 10786 11374 10788 11426
rect 10732 11372 10788 11374
rect 11052 11426 11108 11428
rect 11052 11374 11054 11426
rect 11054 11374 11106 11426
rect 11106 11374 11108 11426
rect 11052 11372 11108 11374
rect 11372 11426 11428 11428
rect 11372 11374 11374 11426
rect 11374 11374 11426 11426
rect 11426 11374 11428 11426
rect 11372 11372 11428 11374
rect 11532 11426 11588 11428
rect 11532 11374 11534 11426
rect 11534 11374 11586 11426
rect 11586 11374 11588 11426
rect 11532 11372 11588 11374
rect 11852 11426 11908 11428
rect 11852 11374 11854 11426
rect 11854 11374 11906 11426
rect 11906 11374 11908 11426
rect 11852 11372 11908 11374
rect 12012 11426 12068 11428
rect 12012 11374 12014 11426
rect 12014 11374 12066 11426
rect 12066 11374 12068 11426
rect 12012 11372 12068 11374
rect 12332 11426 12388 11428
rect 12332 11374 12334 11426
rect 12334 11374 12386 11426
rect 12386 11374 12388 11426
rect 12332 11372 12388 11374
rect 8492 11266 8548 11268
rect 8492 11214 8494 11266
rect 8494 11214 8546 11266
rect 8546 11214 8548 11266
rect 8492 11212 8548 11214
rect 8812 11266 8868 11268
rect 8812 11214 8814 11266
rect 8814 11214 8866 11266
rect 8866 11214 8868 11266
rect 8812 11212 8868 11214
rect 8972 11266 9028 11268
rect 8972 11214 8974 11266
rect 8974 11214 9026 11266
rect 9026 11214 9028 11266
rect 8972 11212 9028 11214
rect 9292 11266 9348 11268
rect 9292 11214 9294 11266
rect 9294 11214 9346 11266
rect 9346 11214 9348 11266
rect 9292 11212 9348 11214
rect 9452 11266 9508 11268
rect 9452 11214 9454 11266
rect 9454 11214 9506 11266
rect 9506 11214 9508 11266
rect 9452 11212 9508 11214
rect 9772 11266 9828 11268
rect 9772 11214 9774 11266
rect 9774 11214 9826 11266
rect 9826 11214 9828 11266
rect 9772 11212 9828 11214
rect 10092 11266 10148 11268
rect 10092 11214 10094 11266
rect 10094 11214 10146 11266
rect 10146 11214 10148 11266
rect 10092 11212 10148 11214
rect 10412 11266 10468 11268
rect 10412 11214 10414 11266
rect 10414 11214 10466 11266
rect 10466 11214 10468 11266
rect 10412 11212 10468 11214
rect 10732 11266 10788 11268
rect 10732 11214 10734 11266
rect 10734 11214 10786 11266
rect 10786 11214 10788 11266
rect 10732 11212 10788 11214
rect 11052 11266 11108 11268
rect 11052 11214 11054 11266
rect 11054 11214 11106 11266
rect 11106 11214 11108 11266
rect 11052 11212 11108 11214
rect 11372 11266 11428 11268
rect 11372 11214 11374 11266
rect 11374 11214 11426 11266
rect 11426 11214 11428 11266
rect 11372 11212 11428 11214
rect 11532 11266 11588 11268
rect 11532 11214 11534 11266
rect 11534 11214 11586 11266
rect 11586 11214 11588 11266
rect 11532 11212 11588 11214
rect 11852 11266 11908 11268
rect 11852 11214 11854 11266
rect 11854 11214 11906 11266
rect 11906 11214 11908 11266
rect 11852 11212 11908 11214
rect 12012 11266 12068 11268
rect 12012 11214 12014 11266
rect 12014 11214 12066 11266
rect 12066 11214 12068 11266
rect 12012 11212 12068 11214
rect 12332 11266 12388 11268
rect 12332 11214 12334 11266
rect 12334 11214 12386 11266
rect 12386 11214 12388 11266
rect 12332 11212 12388 11214
rect 8492 11106 8548 11108
rect 8492 11054 8494 11106
rect 8494 11054 8546 11106
rect 8546 11054 8548 11106
rect 8492 11052 8548 11054
rect 8812 11106 8868 11108
rect 8812 11054 8814 11106
rect 8814 11054 8866 11106
rect 8866 11054 8868 11106
rect 8812 11052 8868 11054
rect 8972 11106 9028 11108
rect 8972 11054 8974 11106
rect 8974 11054 9026 11106
rect 9026 11054 9028 11106
rect 8972 11052 9028 11054
rect 9292 11106 9348 11108
rect 9292 11054 9294 11106
rect 9294 11054 9346 11106
rect 9346 11054 9348 11106
rect 9292 11052 9348 11054
rect 9452 11106 9508 11108
rect 9452 11054 9454 11106
rect 9454 11054 9506 11106
rect 9506 11054 9508 11106
rect 9452 11052 9508 11054
rect 9772 11106 9828 11108
rect 9772 11054 9774 11106
rect 9774 11054 9826 11106
rect 9826 11054 9828 11106
rect 9772 11052 9828 11054
rect 10092 11106 10148 11108
rect 10092 11054 10094 11106
rect 10094 11054 10146 11106
rect 10146 11054 10148 11106
rect 10092 11052 10148 11054
rect 10412 11106 10468 11108
rect 10412 11054 10414 11106
rect 10414 11054 10466 11106
rect 10466 11054 10468 11106
rect 10412 11052 10468 11054
rect 10732 11106 10788 11108
rect 10732 11054 10734 11106
rect 10734 11054 10786 11106
rect 10786 11054 10788 11106
rect 10732 11052 10788 11054
rect 11052 11106 11108 11108
rect 11052 11054 11054 11106
rect 11054 11054 11106 11106
rect 11106 11054 11108 11106
rect 11052 11052 11108 11054
rect 11372 11106 11428 11108
rect 11372 11054 11374 11106
rect 11374 11054 11426 11106
rect 11426 11054 11428 11106
rect 11372 11052 11428 11054
rect 11532 11106 11588 11108
rect 11532 11054 11534 11106
rect 11534 11054 11586 11106
rect 11586 11054 11588 11106
rect 11532 11052 11588 11054
rect 11852 11106 11908 11108
rect 11852 11054 11854 11106
rect 11854 11054 11906 11106
rect 11906 11054 11908 11106
rect 11852 11052 11908 11054
rect 12012 11106 12068 11108
rect 12012 11054 12014 11106
rect 12014 11054 12066 11106
rect 12066 11054 12068 11106
rect 12012 11052 12068 11054
rect 12332 11106 12388 11108
rect 12332 11054 12334 11106
rect 12334 11054 12386 11106
rect 12386 11054 12388 11106
rect 12332 11052 12388 11054
rect 8492 10946 8548 10948
rect 8492 10894 8494 10946
rect 8494 10894 8546 10946
rect 8546 10894 8548 10946
rect 8492 10892 8548 10894
rect 8812 10946 8868 10948
rect 8812 10894 8814 10946
rect 8814 10894 8866 10946
rect 8866 10894 8868 10946
rect 8812 10892 8868 10894
rect 8972 10946 9028 10948
rect 8972 10894 8974 10946
rect 8974 10894 9026 10946
rect 9026 10894 9028 10946
rect 8972 10892 9028 10894
rect 9292 10946 9348 10948
rect 9292 10894 9294 10946
rect 9294 10894 9346 10946
rect 9346 10894 9348 10946
rect 9292 10892 9348 10894
rect 9452 10946 9508 10948
rect 9452 10894 9454 10946
rect 9454 10894 9506 10946
rect 9506 10894 9508 10946
rect 9452 10892 9508 10894
rect 9772 10946 9828 10948
rect 9772 10894 9774 10946
rect 9774 10894 9826 10946
rect 9826 10894 9828 10946
rect 9772 10892 9828 10894
rect 10092 10946 10148 10948
rect 10092 10894 10094 10946
rect 10094 10894 10146 10946
rect 10146 10894 10148 10946
rect 10092 10892 10148 10894
rect 10412 10946 10468 10948
rect 10412 10894 10414 10946
rect 10414 10894 10466 10946
rect 10466 10894 10468 10946
rect 10412 10892 10468 10894
rect 10732 10946 10788 10948
rect 10732 10894 10734 10946
rect 10734 10894 10786 10946
rect 10786 10894 10788 10946
rect 10732 10892 10788 10894
rect 11052 10946 11108 10948
rect 11052 10894 11054 10946
rect 11054 10894 11106 10946
rect 11106 10894 11108 10946
rect 11052 10892 11108 10894
rect 11372 10946 11428 10948
rect 11372 10894 11374 10946
rect 11374 10894 11426 10946
rect 11426 10894 11428 10946
rect 11372 10892 11428 10894
rect 11532 10946 11588 10948
rect 11532 10894 11534 10946
rect 11534 10894 11586 10946
rect 11586 10894 11588 10946
rect 11532 10892 11588 10894
rect 11852 10946 11908 10948
rect 11852 10894 11854 10946
rect 11854 10894 11906 10946
rect 11906 10894 11908 10946
rect 11852 10892 11908 10894
rect 12012 10946 12068 10948
rect 12012 10894 12014 10946
rect 12014 10894 12066 10946
rect 12066 10894 12068 10946
rect 12012 10892 12068 10894
rect 12332 10946 12388 10948
rect 12332 10894 12334 10946
rect 12334 10894 12386 10946
rect 12386 10894 12388 10946
rect 12332 10892 12388 10894
rect 8492 10786 8548 10788
rect 8492 10734 8494 10786
rect 8494 10734 8546 10786
rect 8546 10734 8548 10786
rect 8492 10732 8548 10734
rect 8812 10786 8868 10788
rect 8812 10734 8814 10786
rect 8814 10734 8866 10786
rect 8866 10734 8868 10786
rect 8812 10732 8868 10734
rect 8972 10786 9028 10788
rect 8972 10734 8974 10786
rect 8974 10734 9026 10786
rect 9026 10734 9028 10786
rect 8972 10732 9028 10734
rect 9292 10786 9348 10788
rect 9292 10734 9294 10786
rect 9294 10734 9346 10786
rect 9346 10734 9348 10786
rect 9292 10732 9348 10734
rect 9452 10786 9508 10788
rect 9452 10734 9454 10786
rect 9454 10734 9506 10786
rect 9506 10734 9508 10786
rect 9452 10732 9508 10734
rect 9772 10786 9828 10788
rect 9772 10734 9774 10786
rect 9774 10734 9826 10786
rect 9826 10734 9828 10786
rect 9772 10732 9828 10734
rect 10092 10786 10148 10788
rect 10092 10734 10094 10786
rect 10094 10734 10146 10786
rect 10146 10734 10148 10786
rect 10092 10732 10148 10734
rect 10412 10786 10468 10788
rect 10412 10734 10414 10786
rect 10414 10734 10466 10786
rect 10466 10734 10468 10786
rect 10412 10732 10468 10734
rect 10732 10786 10788 10788
rect 10732 10734 10734 10786
rect 10734 10734 10786 10786
rect 10786 10734 10788 10786
rect 10732 10732 10788 10734
rect 11052 10786 11108 10788
rect 11052 10734 11054 10786
rect 11054 10734 11106 10786
rect 11106 10734 11108 10786
rect 11052 10732 11108 10734
rect 11372 10786 11428 10788
rect 11372 10734 11374 10786
rect 11374 10734 11426 10786
rect 11426 10734 11428 10786
rect 11372 10732 11428 10734
rect 11532 10786 11588 10788
rect 11532 10734 11534 10786
rect 11534 10734 11586 10786
rect 11586 10734 11588 10786
rect 11532 10732 11588 10734
rect 11852 10786 11908 10788
rect 11852 10734 11854 10786
rect 11854 10734 11906 10786
rect 11906 10734 11908 10786
rect 11852 10732 11908 10734
rect 12012 10786 12068 10788
rect 12012 10734 12014 10786
rect 12014 10734 12066 10786
rect 12066 10734 12068 10786
rect 12012 10732 12068 10734
rect 12332 10786 12388 10788
rect 12332 10734 12334 10786
rect 12334 10734 12386 10786
rect 12386 10734 12388 10786
rect 12332 10732 12388 10734
rect 8492 10626 8548 10628
rect 8492 10574 8494 10626
rect 8494 10574 8546 10626
rect 8546 10574 8548 10626
rect 8492 10572 8548 10574
rect 8812 10626 8868 10628
rect 8812 10574 8814 10626
rect 8814 10574 8866 10626
rect 8866 10574 8868 10626
rect 8812 10572 8868 10574
rect 8972 10626 9028 10628
rect 8972 10574 8974 10626
rect 8974 10574 9026 10626
rect 9026 10574 9028 10626
rect 8972 10572 9028 10574
rect 9292 10626 9348 10628
rect 9292 10574 9294 10626
rect 9294 10574 9346 10626
rect 9346 10574 9348 10626
rect 9292 10572 9348 10574
rect 9452 10626 9508 10628
rect 9452 10574 9454 10626
rect 9454 10574 9506 10626
rect 9506 10574 9508 10626
rect 9452 10572 9508 10574
rect 9772 10626 9828 10628
rect 9772 10574 9774 10626
rect 9774 10574 9826 10626
rect 9826 10574 9828 10626
rect 9772 10572 9828 10574
rect 10092 10626 10148 10628
rect 10092 10574 10094 10626
rect 10094 10574 10146 10626
rect 10146 10574 10148 10626
rect 10092 10572 10148 10574
rect 10412 10626 10468 10628
rect 10412 10574 10414 10626
rect 10414 10574 10466 10626
rect 10466 10574 10468 10626
rect 10412 10572 10468 10574
rect 10732 10626 10788 10628
rect 10732 10574 10734 10626
rect 10734 10574 10786 10626
rect 10786 10574 10788 10626
rect 10732 10572 10788 10574
rect 11052 10626 11108 10628
rect 11052 10574 11054 10626
rect 11054 10574 11106 10626
rect 11106 10574 11108 10626
rect 11052 10572 11108 10574
rect 11372 10626 11428 10628
rect 11372 10574 11374 10626
rect 11374 10574 11426 10626
rect 11426 10574 11428 10626
rect 11372 10572 11428 10574
rect 11532 10626 11588 10628
rect 11532 10574 11534 10626
rect 11534 10574 11586 10626
rect 11586 10574 11588 10626
rect 11532 10572 11588 10574
rect 11852 10626 11908 10628
rect 11852 10574 11854 10626
rect 11854 10574 11906 10626
rect 11906 10574 11908 10626
rect 11852 10572 11908 10574
rect 12012 10626 12068 10628
rect 12012 10574 12014 10626
rect 12014 10574 12066 10626
rect 12066 10574 12068 10626
rect 12012 10572 12068 10574
rect 12332 10626 12388 10628
rect 12332 10574 12334 10626
rect 12334 10574 12386 10626
rect 12386 10574 12388 10626
rect 12332 10572 12388 10574
rect 8492 10466 8548 10468
rect 8492 10414 8494 10466
rect 8494 10414 8546 10466
rect 8546 10414 8548 10466
rect 8492 10412 8548 10414
rect 8812 10466 8868 10468
rect 8812 10414 8814 10466
rect 8814 10414 8866 10466
rect 8866 10414 8868 10466
rect 8812 10412 8868 10414
rect 8972 10466 9028 10468
rect 8972 10414 8974 10466
rect 8974 10414 9026 10466
rect 9026 10414 9028 10466
rect 8972 10412 9028 10414
rect 9292 10466 9348 10468
rect 9292 10414 9294 10466
rect 9294 10414 9346 10466
rect 9346 10414 9348 10466
rect 9292 10412 9348 10414
rect 9452 10466 9508 10468
rect 9452 10414 9454 10466
rect 9454 10414 9506 10466
rect 9506 10414 9508 10466
rect 9452 10412 9508 10414
rect 9772 10466 9828 10468
rect 9772 10414 9774 10466
rect 9774 10414 9826 10466
rect 9826 10414 9828 10466
rect 9772 10412 9828 10414
rect 10092 10466 10148 10468
rect 10092 10414 10094 10466
rect 10094 10414 10146 10466
rect 10146 10414 10148 10466
rect 10092 10412 10148 10414
rect 10412 10466 10468 10468
rect 10412 10414 10414 10466
rect 10414 10414 10466 10466
rect 10466 10414 10468 10466
rect 10412 10412 10468 10414
rect 10732 10466 10788 10468
rect 10732 10414 10734 10466
rect 10734 10414 10786 10466
rect 10786 10414 10788 10466
rect 10732 10412 10788 10414
rect 11052 10466 11108 10468
rect 11052 10414 11054 10466
rect 11054 10414 11106 10466
rect 11106 10414 11108 10466
rect 11052 10412 11108 10414
rect 11372 10466 11428 10468
rect 11372 10414 11374 10466
rect 11374 10414 11426 10466
rect 11426 10414 11428 10466
rect 11372 10412 11428 10414
rect 11532 10466 11588 10468
rect 11532 10414 11534 10466
rect 11534 10414 11586 10466
rect 11586 10414 11588 10466
rect 11532 10412 11588 10414
rect 11852 10466 11908 10468
rect 11852 10414 11854 10466
rect 11854 10414 11906 10466
rect 11906 10414 11908 10466
rect 11852 10412 11908 10414
rect 12012 10466 12068 10468
rect 12012 10414 12014 10466
rect 12014 10414 12066 10466
rect 12066 10414 12068 10466
rect 12012 10412 12068 10414
rect 12332 10466 12388 10468
rect 12332 10414 12334 10466
rect 12334 10414 12386 10466
rect 12386 10414 12388 10466
rect 12332 10412 12388 10414
rect 8492 10306 8548 10308
rect 8492 10254 8494 10306
rect 8494 10254 8546 10306
rect 8546 10254 8548 10306
rect 8492 10252 8548 10254
rect 8812 10306 8868 10308
rect 8812 10254 8814 10306
rect 8814 10254 8866 10306
rect 8866 10254 8868 10306
rect 8812 10252 8868 10254
rect 8972 10306 9028 10308
rect 8972 10254 8974 10306
rect 8974 10254 9026 10306
rect 9026 10254 9028 10306
rect 8972 10252 9028 10254
rect 9292 10306 9348 10308
rect 9292 10254 9294 10306
rect 9294 10254 9346 10306
rect 9346 10254 9348 10306
rect 9292 10252 9348 10254
rect 9452 10306 9508 10308
rect 9452 10254 9454 10306
rect 9454 10254 9506 10306
rect 9506 10254 9508 10306
rect 9452 10252 9508 10254
rect 9772 10306 9828 10308
rect 9772 10254 9774 10306
rect 9774 10254 9826 10306
rect 9826 10254 9828 10306
rect 9772 10252 9828 10254
rect 10092 10306 10148 10308
rect 10092 10254 10094 10306
rect 10094 10254 10146 10306
rect 10146 10254 10148 10306
rect 10092 10252 10148 10254
rect 10412 10306 10468 10308
rect 10412 10254 10414 10306
rect 10414 10254 10466 10306
rect 10466 10254 10468 10306
rect 10412 10252 10468 10254
rect 10732 10306 10788 10308
rect 10732 10254 10734 10306
rect 10734 10254 10786 10306
rect 10786 10254 10788 10306
rect 10732 10252 10788 10254
rect 11052 10306 11108 10308
rect 11052 10254 11054 10306
rect 11054 10254 11106 10306
rect 11106 10254 11108 10306
rect 11052 10252 11108 10254
rect 11372 10306 11428 10308
rect 11372 10254 11374 10306
rect 11374 10254 11426 10306
rect 11426 10254 11428 10306
rect 11372 10252 11428 10254
rect 11532 10306 11588 10308
rect 11532 10254 11534 10306
rect 11534 10254 11586 10306
rect 11586 10254 11588 10306
rect 11532 10252 11588 10254
rect 11852 10306 11908 10308
rect 11852 10254 11854 10306
rect 11854 10254 11906 10306
rect 11906 10254 11908 10306
rect 11852 10252 11908 10254
rect 12012 10306 12068 10308
rect 12012 10254 12014 10306
rect 12014 10254 12066 10306
rect 12066 10254 12068 10306
rect 12012 10252 12068 10254
rect 12332 10306 12388 10308
rect 12332 10254 12334 10306
rect 12334 10254 12386 10306
rect 12386 10254 12388 10306
rect 12332 10252 12388 10254
rect 8492 10146 8548 10148
rect 8492 10094 8494 10146
rect 8494 10094 8546 10146
rect 8546 10094 8548 10146
rect 8492 10092 8548 10094
rect 8812 10146 8868 10148
rect 8812 10094 8814 10146
rect 8814 10094 8866 10146
rect 8866 10094 8868 10146
rect 8812 10092 8868 10094
rect 8972 10146 9028 10148
rect 8972 10094 8974 10146
rect 8974 10094 9026 10146
rect 9026 10094 9028 10146
rect 8972 10092 9028 10094
rect 9292 10146 9348 10148
rect 9292 10094 9294 10146
rect 9294 10094 9346 10146
rect 9346 10094 9348 10146
rect 9292 10092 9348 10094
rect 9452 10146 9508 10148
rect 9452 10094 9454 10146
rect 9454 10094 9506 10146
rect 9506 10094 9508 10146
rect 9452 10092 9508 10094
rect 9772 10146 9828 10148
rect 9772 10094 9774 10146
rect 9774 10094 9826 10146
rect 9826 10094 9828 10146
rect 9772 10092 9828 10094
rect 10092 10146 10148 10148
rect 10092 10094 10094 10146
rect 10094 10094 10146 10146
rect 10146 10094 10148 10146
rect 10092 10092 10148 10094
rect 10412 10146 10468 10148
rect 10412 10094 10414 10146
rect 10414 10094 10466 10146
rect 10466 10094 10468 10146
rect 10412 10092 10468 10094
rect 10732 10146 10788 10148
rect 10732 10094 10734 10146
rect 10734 10094 10786 10146
rect 10786 10094 10788 10146
rect 10732 10092 10788 10094
rect 11052 10146 11108 10148
rect 11052 10094 11054 10146
rect 11054 10094 11106 10146
rect 11106 10094 11108 10146
rect 11052 10092 11108 10094
rect 11372 10146 11428 10148
rect 11372 10094 11374 10146
rect 11374 10094 11426 10146
rect 11426 10094 11428 10146
rect 11372 10092 11428 10094
rect 11532 10146 11588 10148
rect 11532 10094 11534 10146
rect 11534 10094 11586 10146
rect 11586 10094 11588 10146
rect 11532 10092 11588 10094
rect 11852 10146 11908 10148
rect 11852 10094 11854 10146
rect 11854 10094 11906 10146
rect 11906 10094 11908 10146
rect 11852 10092 11908 10094
rect 12012 10146 12068 10148
rect 12012 10094 12014 10146
rect 12014 10094 12066 10146
rect 12066 10094 12068 10146
rect 12012 10092 12068 10094
rect 12332 10146 12388 10148
rect 12332 10094 12334 10146
rect 12334 10094 12386 10146
rect 12386 10094 12388 10146
rect 12332 10092 12388 10094
rect 8492 9986 8548 9988
rect 8492 9934 8494 9986
rect 8494 9934 8546 9986
rect 8546 9934 8548 9986
rect 8492 9932 8548 9934
rect 8812 9986 8868 9988
rect 8812 9934 8814 9986
rect 8814 9934 8866 9986
rect 8866 9934 8868 9986
rect 8812 9932 8868 9934
rect 8972 9986 9028 9988
rect 8972 9934 8974 9986
rect 8974 9934 9026 9986
rect 9026 9934 9028 9986
rect 8972 9932 9028 9934
rect 9292 9986 9348 9988
rect 9292 9934 9294 9986
rect 9294 9934 9346 9986
rect 9346 9934 9348 9986
rect 9292 9932 9348 9934
rect 9452 9986 9508 9988
rect 9452 9934 9454 9986
rect 9454 9934 9506 9986
rect 9506 9934 9508 9986
rect 9452 9932 9508 9934
rect 9772 9986 9828 9988
rect 9772 9934 9774 9986
rect 9774 9934 9826 9986
rect 9826 9934 9828 9986
rect 9772 9932 9828 9934
rect 10092 9986 10148 9988
rect 10092 9934 10094 9986
rect 10094 9934 10146 9986
rect 10146 9934 10148 9986
rect 10092 9932 10148 9934
rect 10412 9986 10468 9988
rect 10412 9934 10414 9986
rect 10414 9934 10466 9986
rect 10466 9934 10468 9986
rect 10412 9932 10468 9934
rect 10732 9986 10788 9988
rect 10732 9934 10734 9986
rect 10734 9934 10786 9986
rect 10786 9934 10788 9986
rect 10732 9932 10788 9934
rect 11052 9986 11108 9988
rect 11052 9934 11054 9986
rect 11054 9934 11106 9986
rect 11106 9934 11108 9986
rect 11052 9932 11108 9934
rect 11372 9986 11428 9988
rect 11372 9934 11374 9986
rect 11374 9934 11426 9986
rect 11426 9934 11428 9986
rect 11372 9932 11428 9934
rect 11532 9986 11588 9988
rect 11532 9934 11534 9986
rect 11534 9934 11586 9986
rect 11586 9934 11588 9986
rect 11532 9932 11588 9934
rect 11852 9986 11908 9988
rect 11852 9934 11854 9986
rect 11854 9934 11906 9986
rect 11906 9934 11908 9986
rect 11852 9932 11908 9934
rect 12012 9986 12068 9988
rect 12012 9934 12014 9986
rect 12014 9934 12066 9986
rect 12066 9934 12068 9986
rect 12012 9932 12068 9934
rect 12332 9986 12388 9988
rect 12332 9934 12334 9986
rect 12334 9934 12386 9986
rect 12386 9934 12388 9986
rect 12332 9932 12388 9934
rect 8492 9826 8548 9828
rect 8492 9774 8494 9826
rect 8494 9774 8546 9826
rect 8546 9774 8548 9826
rect 8492 9772 8548 9774
rect 8812 9826 8868 9828
rect 8812 9774 8814 9826
rect 8814 9774 8866 9826
rect 8866 9774 8868 9826
rect 8812 9772 8868 9774
rect 8972 9826 9028 9828
rect 8972 9774 8974 9826
rect 8974 9774 9026 9826
rect 9026 9774 9028 9826
rect 8972 9772 9028 9774
rect 9292 9826 9348 9828
rect 9292 9774 9294 9826
rect 9294 9774 9346 9826
rect 9346 9774 9348 9826
rect 9292 9772 9348 9774
rect 9452 9826 9508 9828
rect 9452 9774 9454 9826
rect 9454 9774 9506 9826
rect 9506 9774 9508 9826
rect 9452 9772 9508 9774
rect 9772 9826 9828 9828
rect 9772 9774 9774 9826
rect 9774 9774 9826 9826
rect 9826 9774 9828 9826
rect 9772 9772 9828 9774
rect 10092 9826 10148 9828
rect 10092 9774 10094 9826
rect 10094 9774 10146 9826
rect 10146 9774 10148 9826
rect 10092 9772 10148 9774
rect 10412 9826 10468 9828
rect 10412 9774 10414 9826
rect 10414 9774 10466 9826
rect 10466 9774 10468 9826
rect 10412 9772 10468 9774
rect 10732 9826 10788 9828
rect 10732 9774 10734 9826
rect 10734 9774 10786 9826
rect 10786 9774 10788 9826
rect 10732 9772 10788 9774
rect 11052 9826 11108 9828
rect 11052 9774 11054 9826
rect 11054 9774 11106 9826
rect 11106 9774 11108 9826
rect 11052 9772 11108 9774
rect 11372 9826 11428 9828
rect 11372 9774 11374 9826
rect 11374 9774 11426 9826
rect 11426 9774 11428 9826
rect 11372 9772 11428 9774
rect 11532 9826 11588 9828
rect 11532 9774 11534 9826
rect 11534 9774 11586 9826
rect 11586 9774 11588 9826
rect 11532 9772 11588 9774
rect 11852 9826 11908 9828
rect 11852 9774 11854 9826
rect 11854 9774 11906 9826
rect 11906 9774 11908 9826
rect 11852 9772 11908 9774
rect 12012 9826 12068 9828
rect 12012 9774 12014 9826
rect 12014 9774 12066 9826
rect 12066 9774 12068 9826
rect 12012 9772 12068 9774
rect 12332 9826 12388 9828
rect 12332 9774 12334 9826
rect 12334 9774 12386 9826
rect 12386 9774 12388 9826
rect 12332 9772 12388 9774
rect 11692 9612 11748 9668
rect 8492 9506 8548 9508
rect 8492 9454 8494 9506
rect 8494 9454 8546 9506
rect 8546 9454 8548 9506
rect 8492 9452 8548 9454
rect 8812 9506 8868 9508
rect 8812 9454 8814 9506
rect 8814 9454 8866 9506
rect 8866 9454 8868 9506
rect 8812 9452 8868 9454
rect 8972 9506 9028 9508
rect 8972 9454 8974 9506
rect 8974 9454 9026 9506
rect 9026 9454 9028 9506
rect 8972 9452 9028 9454
rect 9292 9506 9348 9508
rect 9292 9454 9294 9506
rect 9294 9454 9346 9506
rect 9346 9454 9348 9506
rect 9292 9452 9348 9454
rect 9452 9506 9508 9508
rect 9452 9454 9454 9506
rect 9454 9454 9506 9506
rect 9506 9454 9508 9506
rect 9452 9452 9508 9454
rect 9772 9506 9828 9508
rect 9772 9454 9774 9506
rect 9774 9454 9826 9506
rect 9826 9454 9828 9506
rect 9772 9452 9828 9454
rect 10092 9506 10148 9508
rect 10092 9454 10094 9506
rect 10094 9454 10146 9506
rect 10146 9454 10148 9506
rect 10092 9452 10148 9454
rect 10412 9506 10468 9508
rect 10412 9454 10414 9506
rect 10414 9454 10466 9506
rect 10466 9454 10468 9506
rect 10412 9452 10468 9454
rect 10732 9506 10788 9508
rect 10732 9454 10734 9506
rect 10734 9454 10786 9506
rect 10786 9454 10788 9506
rect 10732 9452 10788 9454
rect 11052 9506 11108 9508
rect 11052 9454 11054 9506
rect 11054 9454 11106 9506
rect 11106 9454 11108 9506
rect 11052 9452 11108 9454
rect 11372 9506 11428 9508
rect 11372 9454 11374 9506
rect 11374 9454 11426 9506
rect 11426 9454 11428 9506
rect 11372 9452 11428 9454
rect 11532 9506 11588 9508
rect 11532 9454 11534 9506
rect 11534 9454 11586 9506
rect 11586 9454 11588 9506
rect 11532 9452 11588 9454
rect 11852 9506 11908 9508
rect 11852 9454 11854 9506
rect 11854 9454 11906 9506
rect 11906 9454 11908 9506
rect 11852 9452 11908 9454
rect 12012 9506 12068 9508
rect 12012 9454 12014 9506
rect 12014 9454 12066 9506
rect 12066 9454 12068 9506
rect 12012 9452 12068 9454
rect 12332 9506 12388 9508
rect 12332 9454 12334 9506
rect 12334 9454 12386 9506
rect 12386 9454 12388 9506
rect 12332 9452 12388 9454
rect 8492 9346 8548 9348
rect 8492 9294 8494 9346
rect 8494 9294 8546 9346
rect 8546 9294 8548 9346
rect 8492 9292 8548 9294
rect 8812 9346 8868 9348
rect 8812 9294 8814 9346
rect 8814 9294 8866 9346
rect 8866 9294 8868 9346
rect 8812 9292 8868 9294
rect 8972 9346 9028 9348
rect 8972 9294 8974 9346
rect 8974 9294 9026 9346
rect 9026 9294 9028 9346
rect 8972 9292 9028 9294
rect 9292 9346 9348 9348
rect 9292 9294 9294 9346
rect 9294 9294 9346 9346
rect 9346 9294 9348 9346
rect 9292 9292 9348 9294
rect 9452 9346 9508 9348
rect 9452 9294 9454 9346
rect 9454 9294 9506 9346
rect 9506 9294 9508 9346
rect 9452 9292 9508 9294
rect 9772 9346 9828 9348
rect 9772 9294 9774 9346
rect 9774 9294 9826 9346
rect 9826 9294 9828 9346
rect 9772 9292 9828 9294
rect 10092 9346 10148 9348
rect 10092 9294 10094 9346
rect 10094 9294 10146 9346
rect 10146 9294 10148 9346
rect 10092 9292 10148 9294
rect 10412 9346 10468 9348
rect 10412 9294 10414 9346
rect 10414 9294 10466 9346
rect 10466 9294 10468 9346
rect 10412 9292 10468 9294
rect 10732 9346 10788 9348
rect 10732 9294 10734 9346
rect 10734 9294 10786 9346
rect 10786 9294 10788 9346
rect 10732 9292 10788 9294
rect 11052 9346 11108 9348
rect 11052 9294 11054 9346
rect 11054 9294 11106 9346
rect 11106 9294 11108 9346
rect 11052 9292 11108 9294
rect 11372 9346 11428 9348
rect 11372 9294 11374 9346
rect 11374 9294 11426 9346
rect 11426 9294 11428 9346
rect 11372 9292 11428 9294
rect 11532 9346 11588 9348
rect 11532 9294 11534 9346
rect 11534 9294 11586 9346
rect 11586 9294 11588 9346
rect 11532 9292 11588 9294
rect 11852 9346 11908 9348
rect 11852 9294 11854 9346
rect 11854 9294 11906 9346
rect 11906 9294 11908 9346
rect 11852 9292 11908 9294
rect 12012 9346 12068 9348
rect 12012 9294 12014 9346
rect 12014 9294 12066 9346
rect 12066 9294 12068 9346
rect 12012 9292 12068 9294
rect 12332 9346 12388 9348
rect 12332 9294 12334 9346
rect 12334 9294 12386 9346
rect 12386 9294 12388 9346
rect 12332 9292 12388 9294
rect 12172 9132 12228 9188
rect 8492 9026 8548 9028
rect 8492 8974 8494 9026
rect 8494 8974 8546 9026
rect 8546 8974 8548 9026
rect 8492 8972 8548 8974
rect 8812 9026 8868 9028
rect 8812 8974 8814 9026
rect 8814 8974 8866 9026
rect 8866 8974 8868 9026
rect 8812 8972 8868 8974
rect 8972 9026 9028 9028
rect 8972 8974 8974 9026
rect 8974 8974 9026 9026
rect 9026 8974 9028 9026
rect 8972 8972 9028 8974
rect 9292 9026 9348 9028
rect 9292 8974 9294 9026
rect 9294 8974 9346 9026
rect 9346 8974 9348 9026
rect 9292 8972 9348 8974
rect 9452 9026 9508 9028
rect 9452 8974 9454 9026
rect 9454 8974 9506 9026
rect 9506 8974 9508 9026
rect 9452 8972 9508 8974
rect 9772 9026 9828 9028
rect 9772 8974 9774 9026
rect 9774 8974 9826 9026
rect 9826 8974 9828 9026
rect 9772 8972 9828 8974
rect 10092 9026 10148 9028
rect 10092 8974 10094 9026
rect 10094 8974 10146 9026
rect 10146 8974 10148 9026
rect 10092 8972 10148 8974
rect 10412 9026 10468 9028
rect 10412 8974 10414 9026
rect 10414 8974 10466 9026
rect 10466 8974 10468 9026
rect 10412 8972 10468 8974
rect 10732 9026 10788 9028
rect 10732 8974 10734 9026
rect 10734 8974 10786 9026
rect 10786 8974 10788 9026
rect 10732 8972 10788 8974
rect 11052 9026 11108 9028
rect 11052 8974 11054 9026
rect 11054 8974 11106 9026
rect 11106 8974 11108 9026
rect 11052 8972 11108 8974
rect 11372 9026 11428 9028
rect 11372 8974 11374 9026
rect 11374 8974 11426 9026
rect 11426 8974 11428 9026
rect 11372 8972 11428 8974
rect 11532 9026 11588 9028
rect 11532 8974 11534 9026
rect 11534 8974 11586 9026
rect 11586 8974 11588 9026
rect 11532 8972 11588 8974
rect 11852 9026 11908 9028
rect 11852 8974 11854 9026
rect 11854 8974 11906 9026
rect 11906 8974 11908 9026
rect 11852 8972 11908 8974
rect 12012 9026 12068 9028
rect 12012 8974 12014 9026
rect 12014 8974 12066 9026
rect 12066 8974 12068 9026
rect 12012 8972 12068 8974
rect 12332 9026 12388 9028
rect 12332 8974 12334 9026
rect 12334 8974 12386 9026
rect 12386 8974 12388 9026
rect 12332 8972 12388 8974
rect 8492 8866 8548 8868
rect 8492 8814 8494 8866
rect 8494 8814 8546 8866
rect 8546 8814 8548 8866
rect 8492 8812 8548 8814
rect 8812 8866 8868 8868
rect 8812 8814 8814 8866
rect 8814 8814 8866 8866
rect 8866 8814 8868 8866
rect 8812 8812 8868 8814
rect 8972 8866 9028 8868
rect 8972 8814 8974 8866
rect 8974 8814 9026 8866
rect 9026 8814 9028 8866
rect 8972 8812 9028 8814
rect 9292 8866 9348 8868
rect 9292 8814 9294 8866
rect 9294 8814 9346 8866
rect 9346 8814 9348 8866
rect 9292 8812 9348 8814
rect 9452 8866 9508 8868
rect 9452 8814 9454 8866
rect 9454 8814 9506 8866
rect 9506 8814 9508 8866
rect 9452 8812 9508 8814
rect 9772 8866 9828 8868
rect 9772 8814 9774 8866
rect 9774 8814 9826 8866
rect 9826 8814 9828 8866
rect 9772 8812 9828 8814
rect 10092 8866 10148 8868
rect 10092 8814 10094 8866
rect 10094 8814 10146 8866
rect 10146 8814 10148 8866
rect 10092 8812 10148 8814
rect 10412 8866 10468 8868
rect 10412 8814 10414 8866
rect 10414 8814 10466 8866
rect 10466 8814 10468 8866
rect 10412 8812 10468 8814
rect 10732 8866 10788 8868
rect 10732 8814 10734 8866
rect 10734 8814 10786 8866
rect 10786 8814 10788 8866
rect 10732 8812 10788 8814
rect 11052 8866 11108 8868
rect 11052 8814 11054 8866
rect 11054 8814 11106 8866
rect 11106 8814 11108 8866
rect 11052 8812 11108 8814
rect 11372 8866 11428 8868
rect 11372 8814 11374 8866
rect 11374 8814 11426 8866
rect 11426 8814 11428 8866
rect 11372 8812 11428 8814
rect 11532 8866 11588 8868
rect 11532 8814 11534 8866
rect 11534 8814 11586 8866
rect 11586 8814 11588 8866
rect 11532 8812 11588 8814
rect 11852 8866 11908 8868
rect 11852 8814 11854 8866
rect 11854 8814 11906 8866
rect 11906 8814 11908 8866
rect 11852 8812 11908 8814
rect 12012 8866 12068 8868
rect 12012 8814 12014 8866
rect 12014 8814 12066 8866
rect 12066 8814 12068 8866
rect 12012 8812 12068 8814
rect 12332 8866 12388 8868
rect 12332 8814 12334 8866
rect 12334 8814 12386 8866
rect 12386 8814 12388 8866
rect 12332 8812 12388 8814
rect 8492 8706 8548 8708
rect 8492 8654 8494 8706
rect 8494 8654 8546 8706
rect 8546 8654 8548 8706
rect 8492 8652 8548 8654
rect 8812 8706 8868 8708
rect 8812 8654 8814 8706
rect 8814 8654 8866 8706
rect 8866 8654 8868 8706
rect 8812 8652 8868 8654
rect 8972 8706 9028 8708
rect 8972 8654 8974 8706
rect 8974 8654 9026 8706
rect 9026 8654 9028 8706
rect 8972 8652 9028 8654
rect 9292 8706 9348 8708
rect 9292 8654 9294 8706
rect 9294 8654 9346 8706
rect 9346 8654 9348 8706
rect 9292 8652 9348 8654
rect 9452 8706 9508 8708
rect 9452 8654 9454 8706
rect 9454 8654 9506 8706
rect 9506 8654 9508 8706
rect 9452 8652 9508 8654
rect 9772 8706 9828 8708
rect 9772 8654 9774 8706
rect 9774 8654 9826 8706
rect 9826 8654 9828 8706
rect 9772 8652 9828 8654
rect 10092 8706 10148 8708
rect 10092 8654 10094 8706
rect 10094 8654 10146 8706
rect 10146 8654 10148 8706
rect 10092 8652 10148 8654
rect 10412 8706 10468 8708
rect 10412 8654 10414 8706
rect 10414 8654 10466 8706
rect 10466 8654 10468 8706
rect 10412 8652 10468 8654
rect 10732 8706 10788 8708
rect 10732 8654 10734 8706
rect 10734 8654 10786 8706
rect 10786 8654 10788 8706
rect 10732 8652 10788 8654
rect 11052 8706 11108 8708
rect 11052 8654 11054 8706
rect 11054 8654 11106 8706
rect 11106 8654 11108 8706
rect 11052 8652 11108 8654
rect 11372 8706 11428 8708
rect 11372 8654 11374 8706
rect 11374 8654 11426 8706
rect 11426 8654 11428 8706
rect 11372 8652 11428 8654
rect 11532 8706 11588 8708
rect 11532 8654 11534 8706
rect 11534 8654 11586 8706
rect 11586 8654 11588 8706
rect 11532 8652 11588 8654
rect 11852 8706 11908 8708
rect 11852 8654 11854 8706
rect 11854 8654 11906 8706
rect 11906 8654 11908 8706
rect 11852 8652 11908 8654
rect 12012 8706 12068 8708
rect 12012 8654 12014 8706
rect 12014 8654 12066 8706
rect 12066 8654 12068 8706
rect 12012 8652 12068 8654
rect 12332 8706 12388 8708
rect 12332 8654 12334 8706
rect 12334 8654 12386 8706
rect 12386 8654 12388 8706
rect 12332 8652 12388 8654
rect 8492 8546 8548 8548
rect 8492 8494 8494 8546
rect 8494 8494 8546 8546
rect 8546 8494 8548 8546
rect 8492 8492 8548 8494
rect 8812 8546 8868 8548
rect 8812 8494 8814 8546
rect 8814 8494 8866 8546
rect 8866 8494 8868 8546
rect 8812 8492 8868 8494
rect 8972 8546 9028 8548
rect 8972 8494 8974 8546
rect 8974 8494 9026 8546
rect 9026 8494 9028 8546
rect 8972 8492 9028 8494
rect 9292 8546 9348 8548
rect 9292 8494 9294 8546
rect 9294 8494 9346 8546
rect 9346 8494 9348 8546
rect 9292 8492 9348 8494
rect 9452 8546 9508 8548
rect 9452 8494 9454 8546
rect 9454 8494 9506 8546
rect 9506 8494 9508 8546
rect 9452 8492 9508 8494
rect 9772 8546 9828 8548
rect 9772 8494 9774 8546
rect 9774 8494 9826 8546
rect 9826 8494 9828 8546
rect 9772 8492 9828 8494
rect 10092 8546 10148 8548
rect 10092 8494 10094 8546
rect 10094 8494 10146 8546
rect 10146 8494 10148 8546
rect 10092 8492 10148 8494
rect 10412 8546 10468 8548
rect 10412 8494 10414 8546
rect 10414 8494 10466 8546
rect 10466 8494 10468 8546
rect 10412 8492 10468 8494
rect 10732 8546 10788 8548
rect 10732 8494 10734 8546
rect 10734 8494 10786 8546
rect 10786 8494 10788 8546
rect 10732 8492 10788 8494
rect 11052 8546 11108 8548
rect 11052 8494 11054 8546
rect 11054 8494 11106 8546
rect 11106 8494 11108 8546
rect 11052 8492 11108 8494
rect 11372 8546 11428 8548
rect 11372 8494 11374 8546
rect 11374 8494 11426 8546
rect 11426 8494 11428 8546
rect 11372 8492 11428 8494
rect 11532 8546 11588 8548
rect 11532 8494 11534 8546
rect 11534 8494 11586 8546
rect 11586 8494 11588 8546
rect 11532 8492 11588 8494
rect 11852 8546 11908 8548
rect 11852 8494 11854 8546
rect 11854 8494 11906 8546
rect 11906 8494 11908 8546
rect 11852 8492 11908 8494
rect 12012 8546 12068 8548
rect 12012 8494 12014 8546
rect 12014 8494 12066 8546
rect 12066 8494 12068 8546
rect 12012 8492 12068 8494
rect 12332 8546 12388 8548
rect 12332 8494 12334 8546
rect 12334 8494 12386 8546
rect 12386 8494 12388 8546
rect 12332 8492 12388 8494
rect 8492 8386 8548 8388
rect 8492 8334 8494 8386
rect 8494 8334 8546 8386
rect 8546 8334 8548 8386
rect 8492 8332 8548 8334
rect 8812 8386 8868 8388
rect 8812 8334 8814 8386
rect 8814 8334 8866 8386
rect 8866 8334 8868 8386
rect 8812 8332 8868 8334
rect 8972 8386 9028 8388
rect 8972 8334 8974 8386
rect 8974 8334 9026 8386
rect 9026 8334 9028 8386
rect 8972 8332 9028 8334
rect 9292 8386 9348 8388
rect 9292 8334 9294 8386
rect 9294 8334 9346 8386
rect 9346 8334 9348 8386
rect 9292 8332 9348 8334
rect 9452 8386 9508 8388
rect 9452 8334 9454 8386
rect 9454 8334 9506 8386
rect 9506 8334 9508 8386
rect 9452 8332 9508 8334
rect 9772 8386 9828 8388
rect 9772 8334 9774 8386
rect 9774 8334 9826 8386
rect 9826 8334 9828 8386
rect 9772 8332 9828 8334
rect 10092 8386 10148 8388
rect 10092 8334 10094 8386
rect 10094 8334 10146 8386
rect 10146 8334 10148 8386
rect 10092 8332 10148 8334
rect 10412 8386 10468 8388
rect 10412 8334 10414 8386
rect 10414 8334 10466 8386
rect 10466 8334 10468 8386
rect 10412 8332 10468 8334
rect 10732 8386 10788 8388
rect 10732 8334 10734 8386
rect 10734 8334 10786 8386
rect 10786 8334 10788 8386
rect 10732 8332 10788 8334
rect 11052 8386 11108 8388
rect 11052 8334 11054 8386
rect 11054 8334 11106 8386
rect 11106 8334 11108 8386
rect 11052 8332 11108 8334
rect 11372 8386 11428 8388
rect 11372 8334 11374 8386
rect 11374 8334 11426 8386
rect 11426 8334 11428 8386
rect 11372 8332 11428 8334
rect 11532 8386 11588 8388
rect 11532 8334 11534 8386
rect 11534 8334 11586 8386
rect 11586 8334 11588 8386
rect 11532 8332 11588 8334
rect 11852 8386 11908 8388
rect 11852 8334 11854 8386
rect 11854 8334 11906 8386
rect 11906 8334 11908 8386
rect 11852 8332 11908 8334
rect 12012 8386 12068 8388
rect 12012 8334 12014 8386
rect 12014 8334 12066 8386
rect 12066 8334 12068 8386
rect 12012 8332 12068 8334
rect 12332 8386 12388 8388
rect 12332 8334 12334 8386
rect 12334 8334 12386 8386
rect 12386 8334 12388 8386
rect 12332 8332 12388 8334
rect 8492 8226 8548 8228
rect 8492 8174 8494 8226
rect 8494 8174 8546 8226
rect 8546 8174 8548 8226
rect 8492 8172 8548 8174
rect 8812 8226 8868 8228
rect 8812 8174 8814 8226
rect 8814 8174 8866 8226
rect 8866 8174 8868 8226
rect 8812 8172 8868 8174
rect 8972 8226 9028 8228
rect 8972 8174 8974 8226
rect 8974 8174 9026 8226
rect 9026 8174 9028 8226
rect 8972 8172 9028 8174
rect 9292 8226 9348 8228
rect 9292 8174 9294 8226
rect 9294 8174 9346 8226
rect 9346 8174 9348 8226
rect 9292 8172 9348 8174
rect 9452 8226 9508 8228
rect 9452 8174 9454 8226
rect 9454 8174 9506 8226
rect 9506 8174 9508 8226
rect 9452 8172 9508 8174
rect 9772 8226 9828 8228
rect 9772 8174 9774 8226
rect 9774 8174 9826 8226
rect 9826 8174 9828 8226
rect 9772 8172 9828 8174
rect 10092 8226 10148 8228
rect 10092 8174 10094 8226
rect 10094 8174 10146 8226
rect 10146 8174 10148 8226
rect 10092 8172 10148 8174
rect 10412 8226 10468 8228
rect 10412 8174 10414 8226
rect 10414 8174 10466 8226
rect 10466 8174 10468 8226
rect 10412 8172 10468 8174
rect 10732 8226 10788 8228
rect 10732 8174 10734 8226
rect 10734 8174 10786 8226
rect 10786 8174 10788 8226
rect 10732 8172 10788 8174
rect 11052 8226 11108 8228
rect 11052 8174 11054 8226
rect 11054 8174 11106 8226
rect 11106 8174 11108 8226
rect 11052 8172 11108 8174
rect 11372 8226 11428 8228
rect 11372 8174 11374 8226
rect 11374 8174 11426 8226
rect 11426 8174 11428 8226
rect 11372 8172 11428 8174
rect 11532 8226 11588 8228
rect 11532 8174 11534 8226
rect 11534 8174 11586 8226
rect 11586 8174 11588 8226
rect 11532 8172 11588 8174
rect 11852 8226 11908 8228
rect 11852 8174 11854 8226
rect 11854 8174 11906 8226
rect 11906 8174 11908 8226
rect 11852 8172 11908 8174
rect 12012 8226 12068 8228
rect 12012 8174 12014 8226
rect 12014 8174 12066 8226
rect 12066 8174 12068 8226
rect 12012 8172 12068 8174
rect 12332 8226 12388 8228
rect 12332 8174 12334 8226
rect 12334 8174 12386 8226
rect 12386 8174 12388 8226
rect 12332 8172 12388 8174
rect 8492 8066 8548 8068
rect 8492 8014 8494 8066
rect 8494 8014 8546 8066
rect 8546 8014 8548 8066
rect 8492 8012 8548 8014
rect 8812 8066 8868 8068
rect 8812 8014 8814 8066
rect 8814 8014 8866 8066
rect 8866 8014 8868 8066
rect 8812 8012 8868 8014
rect 8972 8066 9028 8068
rect 8972 8014 8974 8066
rect 8974 8014 9026 8066
rect 9026 8014 9028 8066
rect 8972 8012 9028 8014
rect 9292 8066 9348 8068
rect 9292 8014 9294 8066
rect 9294 8014 9346 8066
rect 9346 8014 9348 8066
rect 9292 8012 9348 8014
rect 9452 8066 9508 8068
rect 9452 8014 9454 8066
rect 9454 8014 9506 8066
rect 9506 8014 9508 8066
rect 9452 8012 9508 8014
rect 9772 8066 9828 8068
rect 9772 8014 9774 8066
rect 9774 8014 9826 8066
rect 9826 8014 9828 8066
rect 9772 8012 9828 8014
rect 10092 8066 10148 8068
rect 10092 8014 10094 8066
rect 10094 8014 10146 8066
rect 10146 8014 10148 8066
rect 10092 8012 10148 8014
rect 10412 8066 10468 8068
rect 10412 8014 10414 8066
rect 10414 8014 10466 8066
rect 10466 8014 10468 8066
rect 10412 8012 10468 8014
rect 10732 8066 10788 8068
rect 10732 8014 10734 8066
rect 10734 8014 10786 8066
rect 10786 8014 10788 8066
rect 10732 8012 10788 8014
rect 11052 8066 11108 8068
rect 11052 8014 11054 8066
rect 11054 8014 11106 8066
rect 11106 8014 11108 8066
rect 11052 8012 11108 8014
rect 11372 8066 11428 8068
rect 11372 8014 11374 8066
rect 11374 8014 11426 8066
rect 11426 8014 11428 8066
rect 11372 8012 11428 8014
rect 11532 8066 11588 8068
rect 11532 8014 11534 8066
rect 11534 8014 11586 8066
rect 11586 8014 11588 8066
rect 11532 8012 11588 8014
rect 11852 8066 11908 8068
rect 11852 8014 11854 8066
rect 11854 8014 11906 8066
rect 11906 8014 11908 8066
rect 11852 8012 11908 8014
rect 12012 8066 12068 8068
rect 12012 8014 12014 8066
rect 12014 8014 12066 8066
rect 12066 8014 12068 8066
rect 12012 8012 12068 8014
rect 12332 8066 12388 8068
rect 12332 8014 12334 8066
rect 12334 8014 12386 8066
rect 12386 8014 12388 8066
rect 12332 8012 12388 8014
rect 8492 7906 8548 7908
rect 8492 7854 8494 7906
rect 8494 7854 8546 7906
rect 8546 7854 8548 7906
rect 8492 7852 8548 7854
rect 8812 7906 8868 7908
rect 8812 7854 8814 7906
rect 8814 7854 8866 7906
rect 8866 7854 8868 7906
rect 8812 7852 8868 7854
rect 8972 7906 9028 7908
rect 8972 7854 8974 7906
rect 8974 7854 9026 7906
rect 9026 7854 9028 7906
rect 8972 7852 9028 7854
rect 9292 7906 9348 7908
rect 9292 7854 9294 7906
rect 9294 7854 9346 7906
rect 9346 7854 9348 7906
rect 9292 7852 9348 7854
rect 9452 7906 9508 7908
rect 9452 7854 9454 7906
rect 9454 7854 9506 7906
rect 9506 7854 9508 7906
rect 9452 7852 9508 7854
rect 9772 7906 9828 7908
rect 9772 7854 9774 7906
rect 9774 7854 9826 7906
rect 9826 7854 9828 7906
rect 9772 7852 9828 7854
rect 10092 7906 10148 7908
rect 10092 7854 10094 7906
rect 10094 7854 10146 7906
rect 10146 7854 10148 7906
rect 10092 7852 10148 7854
rect 10412 7906 10468 7908
rect 10412 7854 10414 7906
rect 10414 7854 10466 7906
rect 10466 7854 10468 7906
rect 10412 7852 10468 7854
rect 10732 7906 10788 7908
rect 10732 7854 10734 7906
rect 10734 7854 10786 7906
rect 10786 7854 10788 7906
rect 10732 7852 10788 7854
rect 11052 7906 11108 7908
rect 11052 7854 11054 7906
rect 11054 7854 11106 7906
rect 11106 7854 11108 7906
rect 11052 7852 11108 7854
rect 11372 7906 11428 7908
rect 11372 7854 11374 7906
rect 11374 7854 11426 7906
rect 11426 7854 11428 7906
rect 11372 7852 11428 7854
rect 11532 7906 11588 7908
rect 11532 7854 11534 7906
rect 11534 7854 11586 7906
rect 11586 7854 11588 7906
rect 11532 7852 11588 7854
rect 11852 7906 11908 7908
rect 11852 7854 11854 7906
rect 11854 7854 11906 7906
rect 11906 7854 11908 7906
rect 11852 7852 11908 7854
rect 12012 7906 12068 7908
rect 12012 7854 12014 7906
rect 12014 7854 12066 7906
rect 12066 7854 12068 7906
rect 12012 7852 12068 7854
rect 12332 7906 12388 7908
rect 12332 7854 12334 7906
rect 12334 7854 12386 7906
rect 12386 7854 12388 7906
rect 12332 7852 12388 7854
rect 8492 7746 8548 7748
rect 8492 7694 8494 7746
rect 8494 7694 8546 7746
rect 8546 7694 8548 7746
rect 8492 7692 8548 7694
rect 8812 7746 8868 7748
rect 8812 7694 8814 7746
rect 8814 7694 8866 7746
rect 8866 7694 8868 7746
rect 8812 7692 8868 7694
rect 8972 7746 9028 7748
rect 8972 7694 8974 7746
rect 8974 7694 9026 7746
rect 9026 7694 9028 7746
rect 8972 7692 9028 7694
rect 9292 7746 9348 7748
rect 9292 7694 9294 7746
rect 9294 7694 9346 7746
rect 9346 7694 9348 7746
rect 9292 7692 9348 7694
rect 9452 7746 9508 7748
rect 9452 7694 9454 7746
rect 9454 7694 9506 7746
rect 9506 7694 9508 7746
rect 9452 7692 9508 7694
rect 9772 7746 9828 7748
rect 9772 7694 9774 7746
rect 9774 7694 9826 7746
rect 9826 7694 9828 7746
rect 9772 7692 9828 7694
rect 10092 7746 10148 7748
rect 10092 7694 10094 7746
rect 10094 7694 10146 7746
rect 10146 7694 10148 7746
rect 10092 7692 10148 7694
rect 10412 7746 10468 7748
rect 10412 7694 10414 7746
rect 10414 7694 10466 7746
rect 10466 7694 10468 7746
rect 10412 7692 10468 7694
rect 10732 7746 10788 7748
rect 10732 7694 10734 7746
rect 10734 7694 10786 7746
rect 10786 7694 10788 7746
rect 10732 7692 10788 7694
rect 11052 7746 11108 7748
rect 11052 7694 11054 7746
rect 11054 7694 11106 7746
rect 11106 7694 11108 7746
rect 11052 7692 11108 7694
rect 11372 7746 11428 7748
rect 11372 7694 11374 7746
rect 11374 7694 11426 7746
rect 11426 7694 11428 7746
rect 11372 7692 11428 7694
rect 11532 7746 11588 7748
rect 11532 7694 11534 7746
rect 11534 7694 11586 7746
rect 11586 7694 11588 7746
rect 11532 7692 11588 7694
rect 11852 7746 11908 7748
rect 11852 7694 11854 7746
rect 11854 7694 11906 7746
rect 11906 7694 11908 7746
rect 11852 7692 11908 7694
rect 12012 7746 12068 7748
rect 12012 7694 12014 7746
rect 12014 7694 12066 7746
rect 12066 7694 12068 7746
rect 12012 7692 12068 7694
rect 12332 7746 12388 7748
rect 12332 7694 12334 7746
rect 12334 7694 12386 7746
rect 12386 7694 12388 7746
rect 12332 7692 12388 7694
rect 8652 7532 8708 7588
rect 8492 7426 8548 7428
rect 8492 7374 8494 7426
rect 8494 7374 8546 7426
rect 8546 7374 8548 7426
rect 8492 7372 8548 7374
rect 8812 7426 8868 7428
rect 8812 7374 8814 7426
rect 8814 7374 8866 7426
rect 8866 7374 8868 7426
rect 8812 7372 8868 7374
rect 8972 7426 9028 7428
rect 8972 7374 8974 7426
rect 8974 7374 9026 7426
rect 9026 7374 9028 7426
rect 8972 7372 9028 7374
rect 9292 7426 9348 7428
rect 9292 7374 9294 7426
rect 9294 7374 9346 7426
rect 9346 7374 9348 7426
rect 9292 7372 9348 7374
rect 9452 7426 9508 7428
rect 9452 7374 9454 7426
rect 9454 7374 9506 7426
rect 9506 7374 9508 7426
rect 9452 7372 9508 7374
rect 9772 7426 9828 7428
rect 9772 7374 9774 7426
rect 9774 7374 9826 7426
rect 9826 7374 9828 7426
rect 9772 7372 9828 7374
rect 10092 7426 10148 7428
rect 10092 7374 10094 7426
rect 10094 7374 10146 7426
rect 10146 7374 10148 7426
rect 10092 7372 10148 7374
rect 10412 7426 10468 7428
rect 10412 7374 10414 7426
rect 10414 7374 10466 7426
rect 10466 7374 10468 7426
rect 10412 7372 10468 7374
rect 10732 7426 10788 7428
rect 10732 7374 10734 7426
rect 10734 7374 10786 7426
rect 10786 7374 10788 7426
rect 10732 7372 10788 7374
rect 11052 7426 11108 7428
rect 11052 7374 11054 7426
rect 11054 7374 11106 7426
rect 11106 7374 11108 7426
rect 11052 7372 11108 7374
rect 11372 7426 11428 7428
rect 11372 7374 11374 7426
rect 11374 7374 11426 7426
rect 11426 7374 11428 7426
rect 11372 7372 11428 7374
rect 11532 7426 11588 7428
rect 11532 7374 11534 7426
rect 11534 7374 11586 7426
rect 11586 7374 11588 7426
rect 11532 7372 11588 7374
rect 11852 7426 11908 7428
rect 11852 7374 11854 7426
rect 11854 7374 11906 7426
rect 11906 7374 11908 7426
rect 11852 7372 11908 7374
rect 12012 7426 12068 7428
rect 12012 7374 12014 7426
rect 12014 7374 12066 7426
rect 12066 7374 12068 7426
rect 12012 7372 12068 7374
rect 12332 7426 12388 7428
rect 12332 7374 12334 7426
rect 12334 7374 12386 7426
rect 12386 7374 12388 7426
rect 12332 7372 12388 7374
rect 8492 7266 8548 7268
rect 8492 7214 8494 7266
rect 8494 7214 8546 7266
rect 8546 7214 8548 7266
rect 8492 7212 8548 7214
rect 8812 7266 8868 7268
rect 8812 7214 8814 7266
rect 8814 7214 8866 7266
rect 8866 7214 8868 7266
rect 8812 7212 8868 7214
rect 8972 7266 9028 7268
rect 8972 7214 8974 7266
rect 8974 7214 9026 7266
rect 9026 7214 9028 7266
rect 8972 7212 9028 7214
rect 9292 7266 9348 7268
rect 9292 7214 9294 7266
rect 9294 7214 9346 7266
rect 9346 7214 9348 7266
rect 9292 7212 9348 7214
rect 9452 7266 9508 7268
rect 9452 7214 9454 7266
rect 9454 7214 9506 7266
rect 9506 7214 9508 7266
rect 9452 7212 9508 7214
rect 9772 7266 9828 7268
rect 9772 7214 9774 7266
rect 9774 7214 9826 7266
rect 9826 7214 9828 7266
rect 9772 7212 9828 7214
rect 10092 7266 10148 7268
rect 10092 7214 10094 7266
rect 10094 7214 10146 7266
rect 10146 7214 10148 7266
rect 10092 7212 10148 7214
rect 10412 7266 10468 7268
rect 10412 7214 10414 7266
rect 10414 7214 10466 7266
rect 10466 7214 10468 7266
rect 10412 7212 10468 7214
rect 10732 7266 10788 7268
rect 10732 7214 10734 7266
rect 10734 7214 10786 7266
rect 10786 7214 10788 7266
rect 10732 7212 10788 7214
rect 11052 7266 11108 7268
rect 11052 7214 11054 7266
rect 11054 7214 11106 7266
rect 11106 7214 11108 7266
rect 11052 7212 11108 7214
rect 11372 7266 11428 7268
rect 11372 7214 11374 7266
rect 11374 7214 11426 7266
rect 11426 7214 11428 7266
rect 11372 7212 11428 7214
rect 11532 7266 11588 7268
rect 11532 7214 11534 7266
rect 11534 7214 11586 7266
rect 11586 7214 11588 7266
rect 11532 7212 11588 7214
rect 11852 7266 11908 7268
rect 11852 7214 11854 7266
rect 11854 7214 11906 7266
rect 11906 7214 11908 7266
rect 11852 7212 11908 7214
rect 12012 7266 12068 7268
rect 12012 7214 12014 7266
rect 12014 7214 12066 7266
rect 12066 7214 12068 7266
rect 12012 7212 12068 7214
rect 12332 7266 12388 7268
rect 12332 7214 12334 7266
rect 12334 7214 12386 7266
rect 12386 7214 12388 7266
rect 12332 7212 12388 7214
rect 9132 7052 9188 7108
rect 8492 6946 8548 6948
rect 8492 6894 8494 6946
rect 8494 6894 8546 6946
rect 8546 6894 8548 6946
rect 8492 6892 8548 6894
rect 8812 6946 8868 6948
rect 8812 6894 8814 6946
rect 8814 6894 8866 6946
rect 8866 6894 8868 6946
rect 8812 6892 8868 6894
rect 8972 6946 9028 6948
rect 8972 6894 8974 6946
rect 8974 6894 9026 6946
rect 9026 6894 9028 6946
rect 8972 6892 9028 6894
rect 9292 6946 9348 6948
rect 9292 6894 9294 6946
rect 9294 6894 9346 6946
rect 9346 6894 9348 6946
rect 9292 6892 9348 6894
rect 9452 6946 9508 6948
rect 9452 6894 9454 6946
rect 9454 6894 9506 6946
rect 9506 6894 9508 6946
rect 9452 6892 9508 6894
rect 9772 6946 9828 6948
rect 9772 6894 9774 6946
rect 9774 6894 9826 6946
rect 9826 6894 9828 6946
rect 9772 6892 9828 6894
rect 10092 6946 10148 6948
rect 10092 6894 10094 6946
rect 10094 6894 10146 6946
rect 10146 6894 10148 6946
rect 10092 6892 10148 6894
rect 10412 6946 10468 6948
rect 10412 6894 10414 6946
rect 10414 6894 10466 6946
rect 10466 6894 10468 6946
rect 10412 6892 10468 6894
rect 10732 6946 10788 6948
rect 10732 6894 10734 6946
rect 10734 6894 10786 6946
rect 10786 6894 10788 6946
rect 10732 6892 10788 6894
rect 11052 6946 11108 6948
rect 11052 6894 11054 6946
rect 11054 6894 11106 6946
rect 11106 6894 11108 6946
rect 11052 6892 11108 6894
rect 11372 6946 11428 6948
rect 11372 6894 11374 6946
rect 11374 6894 11426 6946
rect 11426 6894 11428 6946
rect 11372 6892 11428 6894
rect 11532 6946 11588 6948
rect 11532 6894 11534 6946
rect 11534 6894 11586 6946
rect 11586 6894 11588 6946
rect 11532 6892 11588 6894
rect 11852 6946 11908 6948
rect 11852 6894 11854 6946
rect 11854 6894 11906 6946
rect 11906 6894 11908 6946
rect 11852 6892 11908 6894
rect 12012 6946 12068 6948
rect 12012 6894 12014 6946
rect 12014 6894 12066 6946
rect 12066 6894 12068 6946
rect 12012 6892 12068 6894
rect 12332 6946 12388 6948
rect 12332 6894 12334 6946
rect 12334 6894 12386 6946
rect 12386 6894 12388 6946
rect 12332 6892 12388 6894
rect 8492 6786 8548 6788
rect 8492 6734 8494 6786
rect 8494 6734 8546 6786
rect 8546 6734 8548 6786
rect 8492 6732 8548 6734
rect 8812 6786 8868 6788
rect 8812 6734 8814 6786
rect 8814 6734 8866 6786
rect 8866 6734 8868 6786
rect 8812 6732 8868 6734
rect 8972 6786 9028 6788
rect 8972 6734 8974 6786
rect 8974 6734 9026 6786
rect 9026 6734 9028 6786
rect 8972 6732 9028 6734
rect 9292 6786 9348 6788
rect 9292 6734 9294 6786
rect 9294 6734 9346 6786
rect 9346 6734 9348 6786
rect 9292 6732 9348 6734
rect 9452 6786 9508 6788
rect 9452 6734 9454 6786
rect 9454 6734 9506 6786
rect 9506 6734 9508 6786
rect 9452 6732 9508 6734
rect 9772 6786 9828 6788
rect 9772 6734 9774 6786
rect 9774 6734 9826 6786
rect 9826 6734 9828 6786
rect 9772 6732 9828 6734
rect 10092 6786 10148 6788
rect 10092 6734 10094 6786
rect 10094 6734 10146 6786
rect 10146 6734 10148 6786
rect 10092 6732 10148 6734
rect 10412 6786 10468 6788
rect 10412 6734 10414 6786
rect 10414 6734 10466 6786
rect 10466 6734 10468 6786
rect 10412 6732 10468 6734
rect 10732 6786 10788 6788
rect 10732 6734 10734 6786
rect 10734 6734 10786 6786
rect 10786 6734 10788 6786
rect 10732 6732 10788 6734
rect 11052 6786 11108 6788
rect 11052 6734 11054 6786
rect 11054 6734 11106 6786
rect 11106 6734 11108 6786
rect 11052 6732 11108 6734
rect 11372 6786 11428 6788
rect 11372 6734 11374 6786
rect 11374 6734 11426 6786
rect 11426 6734 11428 6786
rect 11372 6732 11428 6734
rect 11532 6786 11588 6788
rect 11532 6734 11534 6786
rect 11534 6734 11586 6786
rect 11586 6734 11588 6786
rect 11532 6732 11588 6734
rect 11852 6786 11908 6788
rect 11852 6734 11854 6786
rect 11854 6734 11906 6786
rect 11906 6734 11908 6786
rect 11852 6732 11908 6734
rect 12012 6786 12068 6788
rect 12012 6734 12014 6786
rect 12014 6734 12066 6786
rect 12066 6734 12068 6786
rect 12012 6732 12068 6734
rect 12332 6786 12388 6788
rect 12332 6734 12334 6786
rect 12334 6734 12386 6786
rect 12386 6734 12388 6786
rect 12332 6732 12388 6734
rect 11692 6572 11748 6628
rect 8492 6466 8548 6468
rect 8492 6414 8494 6466
rect 8494 6414 8546 6466
rect 8546 6414 8548 6466
rect 8492 6412 8548 6414
rect 8812 6466 8868 6468
rect 8812 6414 8814 6466
rect 8814 6414 8866 6466
rect 8866 6414 8868 6466
rect 8812 6412 8868 6414
rect 8972 6466 9028 6468
rect 8972 6414 8974 6466
rect 8974 6414 9026 6466
rect 9026 6414 9028 6466
rect 8972 6412 9028 6414
rect 9292 6466 9348 6468
rect 9292 6414 9294 6466
rect 9294 6414 9346 6466
rect 9346 6414 9348 6466
rect 9292 6412 9348 6414
rect 9452 6466 9508 6468
rect 9452 6414 9454 6466
rect 9454 6414 9506 6466
rect 9506 6414 9508 6466
rect 9452 6412 9508 6414
rect 9772 6466 9828 6468
rect 9772 6414 9774 6466
rect 9774 6414 9826 6466
rect 9826 6414 9828 6466
rect 9772 6412 9828 6414
rect 10092 6466 10148 6468
rect 10092 6414 10094 6466
rect 10094 6414 10146 6466
rect 10146 6414 10148 6466
rect 10092 6412 10148 6414
rect 10412 6466 10468 6468
rect 10412 6414 10414 6466
rect 10414 6414 10466 6466
rect 10466 6414 10468 6466
rect 10412 6412 10468 6414
rect 10732 6466 10788 6468
rect 10732 6414 10734 6466
rect 10734 6414 10786 6466
rect 10786 6414 10788 6466
rect 10732 6412 10788 6414
rect 11052 6466 11108 6468
rect 11052 6414 11054 6466
rect 11054 6414 11106 6466
rect 11106 6414 11108 6466
rect 11052 6412 11108 6414
rect 11372 6466 11428 6468
rect 11372 6414 11374 6466
rect 11374 6414 11426 6466
rect 11426 6414 11428 6466
rect 11372 6412 11428 6414
rect 11532 6466 11588 6468
rect 11532 6414 11534 6466
rect 11534 6414 11586 6466
rect 11586 6414 11588 6466
rect 11532 6412 11588 6414
rect 11852 6466 11908 6468
rect 11852 6414 11854 6466
rect 11854 6414 11906 6466
rect 11906 6414 11908 6466
rect 11852 6412 11908 6414
rect 12012 6466 12068 6468
rect 12012 6414 12014 6466
rect 12014 6414 12066 6466
rect 12066 6414 12068 6466
rect 12012 6412 12068 6414
rect 12332 6466 12388 6468
rect 12332 6414 12334 6466
rect 12334 6414 12386 6466
rect 12386 6414 12388 6466
rect 12332 6412 12388 6414
rect 8492 6306 8548 6308
rect 8492 6254 8494 6306
rect 8494 6254 8546 6306
rect 8546 6254 8548 6306
rect 8492 6252 8548 6254
rect 8812 6306 8868 6308
rect 8812 6254 8814 6306
rect 8814 6254 8866 6306
rect 8866 6254 8868 6306
rect 8812 6252 8868 6254
rect 8972 6306 9028 6308
rect 8972 6254 8974 6306
rect 8974 6254 9026 6306
rect 9026 6254 9028 6306
rect 8972 6252 9028 6254
rect 9292 6306 9348 6308
rect 9292 6254 9294 6306
rect 9294 6254 9346 6306
rect 9346 6254 9348 6306
rect 9292 6252 9348 6254
rect 9452 6306 9508 6308
rect 9452 6254 9454 6306
rect 9454 6254 9506 6306
rect 9506 6254 9508 6306
rect 9452 6252 9508 6254
rect 9772 6306 9828 6308
rect 9772 6254 9774 6306
rect 9774 6254 9826 6306
rect 9826 6254 9828 6306
rect 9772 6252 9828 6254
rect 10092 6306 10148 6308
rect 10092 6254 10094 6306
rect 10094 6254 10146 6306
rect 10146 6254 10148 6306
rect 10092 6252 10148 6254
rect 10412 6306 10468 6308
rect 10412 6254 10414 6306
rect 10414 6254 10466 6306
rect 10466 6254 10468 6306
rect 10412 6252 10468 6254
rect 10732 6306 10788 6308
rect 10732 6254 10734 6306
rect 10734 6254 10786 6306
rect 10786 6254 10788 6306
rect 10732 6252 10788 6254
rect 11052 6306 11108 6308
rect 11052 6254 11054 6306
rect 11054 6254 11106 6306
rect 11106 6254 11108 6306
rect 11052 6252 11108 6254
rect 11372 6306 11428 6308
rect 11372 6254 11374 6306
rect 11374 6254 11426 6306
rect 11426 6254 11428 6306
rect 11372 6252 11428 6254
rect 11532 6306 11588 6308
rect 11532 6254 11534 6306
rect 11534 6254 11586 6306
rect 11586 6254 11588 6306
rect 11532 6252 11588 6254
rect 11852 6306 11908 6308
rect 11852 6254 11854 6306
rect 11854 6254 11906 6306
rect 11906 6254 11908 6306
rect 11852 6252 11908 6254
rect 12012 6306 12068 6308
rect 12012 6254 12014 6306
rect 12014 6254 12066 6306
rect 12066 6254 12068 6306
rect 12012 6252 12068 6254
rect 12332 6306 12388 6308
rect 12332 6254 12334 6306
rect 12334 6254 12386 6306
rect 12386 6254 12388 6306
rect 12332 6252 12388 6254
rect 8492 6146 8548 6148
rect 8492 6094 8494 6146
rect 8494 6094 8546 6146
rect 8546 6094 8548 6146
rect 8492 6092 8548 6094
rect 8812 6146 8868 6148
rect 8812 6094 8814 6146
rect 8814 6094 8866 6146
rect 8866 6094 8868 6146
rect 8812 6092 8868 6094
rect 8972 6146 9028 6148
rect 8972 6094 8974 6146
rect 8974 6094 9026 6146
rect 9026 6094 9028 6146
rect 8972 6092 9028 6094
rect 9292 6146 9348 6148
rect 9292 6094 9294 6146
rect 9294 6094 9346 6146
rect 9346 6094 9348 6146
rect 9292 6092 9348 6094
rect 9452 6146 9508 6148
rect 9452 6094 9454 6146
rect 9454 6094 9506 6146
rect 9506 6094 9508 6146
rect 9452 6092 9508 6094
rect 9772 6146 9828 6148
rect 9772 6094 9774 6146
rect 9774 6094 9826 6146
rect 9826 6094 9828 6146
rect 9772 6092 9828 6094
rect 10092 6146 10148 6148
rect 10092 6094 10094 6146
rect 10094 6094 10146 6146
rect 10146 6094 10148 6146
rect 10092 6092 10148 6094
rect 10412 6146 10468 6148
rect 10412 6094 10414 6146
rect 10414 6094 10466 6146
rect 10466 6094 10468 6146
rect 10412 6092 10468 6094
rect 10732 6146 10788 6148
rect 10732 6094 10734 6146
rect 10734 6094 10786 6146
rect 10786 6094 10788 6146
rect 10732 6092 10788 6094
rect 11052 6146 11108 6148
rect 11052 6094 11054 6146
rect 11054 6094 11106 6146
rect 11106 6094 11108 6146
rect 11052 6092 11108 6094
rect 11372 6146 11428 6148
rect 11372 6094 11374 6146
rect 11374 6094 11426 6146
rect 11426 6094 11428 6146
rect 11372 6092 11428 6094
rect 11532 6146 11588 6148
rect 11532 6094 11534 6146
rect 11534 6094 11586 6146
rect 11586 6094 11588 6146
rect 11532 6092 11588 6094
rect 11852 6146 11908 6148
rect 11852 6094 11854 6146
rect 11854 6094 11906 6146
rect 11906 6094 11908 6146
rect 11852 6092 11908 6094
rect 12012 6146 12068 6148
rect 12012 6094 12014 6146
rect 12014 6094 12066 6146
rect 12066 6094 12068 6146
rect 12012 6092 12068 6094
rect 12332 6146 12388 6148
rect 12332 6094 12334 6146
rect 12334 6094 12386 6146
rect 12386 6094 12388 6146
rect 12332 6092 12388 6094
rect 8492 5986 8548 5988
rect 8492 5934 8494 5986
rect 8494 5934 8546 5986
rect 8546 5934 8548 5986
rect 8492 5932 8548 5934
rect 8812 5986 8868 5988
rect 8812 5934 8814 5986
rect 8814 5934 8866 5986
rect 8866 5934 8868 5986
rect 8812 5932 8868 5934
rect 8972 5986 9028 5988
rect 8972 5934 8974 5986
rect 8974 5934 9026 5986
rect 9026 5934 9028 5986
rect 8972 5932 9028 5934
rect 9292 5986 9348 5988
rect 9292 5934 9294 5986
rect 9294 5934 9346 5986
rect 9346 5934 9348 5986
rect 9292 5932 9348 5934
rect 9452 5986 9508 5988
rect 9452 5934 9454 5986
rect 9454 5934 9506 5986
rect 9506 5934 9508 5986
rect 9452 5932 9508 5934
rect 9772 5986 9828 5988
rect 9772 5934 9774 5986
rect 9774 5934 9826 5986
rect 9826 5934 9828 5986
rect 9772 5932 9828 5934
rect 10092 5986 10148 5988
rect 10092 5934 10094 5986
rect 10094 5934 10146 5986
rect 10146 5934 10148 5986
rect 10092 5932 10148 5934
rect 10412 5986 10468 5988
rect 10412 5934 10414 5986
rect 10414 5934 10466 5986
rect 10466 5934 10468 5986
rect 10412 5932 10468 5934
rect 10732 5986 10788 5988
rect 10732 5934 10734 5986
rect 10734 5934 10786 5986
rect 10786 5934 10788 5986
rect 10732 5932 10788 5934
rect 11052 5986 11108 5988
rect 11052 5934 11054 5986
rect 11054 5934 11106 5986
rect 11106 5934 11108 5986
rect 11052 5932 11108 5934
rect 11372 5986 11428 5988
rect 11372 5934 11374 5986
rect 11374 5934 11426 5986
rect 11426 5934 11428 5986
rect 11372 5932 11428 5934
rect 11532 5986 11588 5988
rect 11532 5934 11534 5986
rect 11534 5934 11586 5986
rect 11586 5934 11588 5986
rect 11532 5932 11588 5934
rect 11852 5986 11908 5988
rect 11852 5934 11854 5986
rect 11854 5934 11906 5986
rect 11906 5934 11908 5986
rect 11852 5932 11908 5934
rect 12012 5986 12068 5988
rect 12012 5934 12014 5986
rect 12014 5934 12066 5986
rect 12066 5934 12068 5986
rect 12012 5932 12068 5934
rect 12332 5986 12388 5988
rect 12332 5934 12334 5986
rect 12334 5934 12386 5986
rect 12386 5934 12388 5986
rect 12332 5932 12388 5934
rect 8492 5826 8548 5828
rect 8492 5774 8494 5826
rect 8494 5774 8546 5826
rect 8546 5774 8548 5826
rect 8492 5772 8548 5774
rect 8812 5826 8868 5828
rect 8812 5774 8814 5826
rect 8814 5774 8866 5826
rect 8866 5774 8868 5826
rect 8812 5772 8868 5774
rect 8972 5826 9028 5828
rect 8972 5774 8974 5826
rect 8974 5774 9026 5826
rect 9026 5774 9028 5826
rect 8972 5772 9028 5774
rect 9292 5826 9348 5828
rect 9292 5774 9294 5826
rect 9294 5774 9346 5826
rect 9346 5774 9348 5826
rect 9292 5772 9348 5774
rect 9452 5826 9508 5828
rect 9452 5774 9454 5826
rect 9454 5774 9506 5826
rect 9506 5774 9508 5826
rect 9452 5772 9508 5774
rect 9772 5826 9828 5828
rect 9772 5774 9774 5826
rect 9774 5774 9826 5826
rect 9826 5774 9828 5826
rect 9772 5772 9828 5774
rect 10092 5826 10148 5828
rect 10092 5774 10094 5826
rect 10094 5774 10146 5826
rect 10146 5774 10148 5826
rect 10092 5772 10148 5774
rect 10412 5826 10468 5828
rect 10412 5774 10414 5826
rect 10414 5774 10466 5826
rect 10466 5774 10468 5826
rect 10412 5772 10468 5774
rect 10732 5826 10788 5828
rect 10732 5774 10734 5826
rect 10734 5774 10786 5826
rect 10786 5774 10788 5826
rect 10732 5772 10788 5774
rect 11052 5826 11108 5828
rect 11052 5774 11054 5826
rect 11054 5774 11106 5826
rect 11106 5774 11108 5826
rect 11052 5772 11108 5774
rect 11372 5826 11428 5828
rect 11372 5774 11374 5826
rect 11374 5774 11426 5826
rect 11426 5774 11428 5826
rect 11372 5772 11428 5774
rect 11532 5826 11588 5828
rect 11532 5774 11534 5826
rect 11534 5774 11586 5826
rect 11586 5774 11588 5826
rect 11532 5772 11588 5774
rect 11852 5826 11908 5828
rect 11852 5774 11854 5826
rect 11854 5774 11906 5826
rect 11906 5774 11908 5826
rect 11852 5772 11908 5774
rect 12012 5826 12068 5828
rect 12012 5774 12014 5826
rect 12014 5774 12066 5826
rect 12066 5774 12068 5826
rect 12012 5772 12068 5774
rect 12332 5826 12388 5828
rect 12332 5774 12334 5826
rect 12334 5774 12386 5826
rect 12386 5774 12388 5826
rect 12332 5772 12388 5774
rect 8492 5666 8548 5668
rect 8492 5614 8494 5666
rect 8494 5614 8546 5666
rect 8546 5614 8548 5666
rect 8492 5612 8548 5614
rect 8812 5666 8868 5668
rect 8812 5614 8814 5666
rect 8814 5614 8866 5666
rect 8866 5614 8868 5666
rect 8812 5612 8868 5614
rect 8972 5666 9028 5668
rect 8972 5614 8974 5666
rect 8974 5614 9026 5666
rect 9026 5614 9028 5666
rect 8972 5612 9028 5614
rect 9292 5666 9348 5668
rect 9292 5614 9294 5666
rect 9294 5614 9346 5666
rect 9346 5614 9348 5666
rect 9292 5612 9348 5614
rect 9452 5666 9508 5668
rect 9452 5614 9454 5666
rect 9454 5614 9506 5666
rect 9506 5614 9508 5666
rect 9452 5612 9508 5614
rect 9772 5666 9828 5668
rect 9772 5614 9774 5666
rect 9774 5614 9826 5666
rect 9826 5614 9828 5666
rect 9772 5612 9828 5614
rect 10092 5666 10148 5668
rect 10092 5614 10094 5666
rect 10094 5614 10146 5666
rect 10146 5614 10148 5666
rect 10092 5612 10148 5614
rect 10412 5666 10468 5668
rect 10412 5614 10414 5666
rect 10414 5614 10466 5666
rect 10466 5614 10468 5666
rect 10412 5612 10468 5614
rect 10732 5666 10788 5668
rect 10732 5614 10734 5666
rect 10734 5614 10786 5666
rect 10786 5614 10788 5666
rect 10732 5612 10788 5614
rect 11052 5666 11108 5668
rect 11052 5614 11054 5666
rect 11054 5614 11106 5666
rect 11106 5614 11108 5666
rect 11052 5612 11108 5614
rect 11372 5666 11428 5668
rect 11372 5614 11374 5666
rect 11374 5614 11426 5666
rect 11426 5614 11428 5666
rect 11372 5612 11428 5614
rect 11532 5666 11588 5668
rect 11532 5614 11534 5666
rect 11534 5614 11586 5666
rect 11586 5614 11588 5666
rect 11532 5612 11588 5614
rect 11852 5666 11908 5668
rect 11852 5614 11854 5666
rect 11854 5614 11906 5666
rect 11906 5614 11908 5666
rect 11852 5612 11908 5614
rect 12012 5666 12068 5668
rect 12012 5614 12014 5666
rect 12014 5614 12066 5666
rect 12066 5614 12068 5666
rect 12012 5612 12068 5614
rect 12332 5666 12388 5668
rect 12332 5614 12334 5666
rect 12334 5614 12386 5666
rect 12386 5614 12388 5666
rect 12332 5612 12388 5614
rect 8492 5506 8548 5508
rect 8492 5454 8494 5506
rect 8494 5454 8546 5506
rect 8546 5454 8548 5506
rect 8492 5452 8548 5454
rect 8812 5506 8868 5508
rect 8812 5454 8814 5506
rect 8814 5454 8866 5506
rect 8866 5454 8868 5506
rect 8812 5452 8868 5454
rect 8972 5506 9028 5508
rect 8972 5454 8974 5506
rect 8974 5454 9026 5506
rect 9026 5454 9028 5506
rect 8972 5452 9028 5454
rect 9292 5506 9348 5508
rect 9292 5454 9294 5506
rect 9294 5454 9346 5506
rect 9346 5454 9348 5506
rect 9292 5452 9348 5454
rect 9452 5506 9508 5508
rect 9452 5454 9454 5506
rect 9454 5454 9506 5506
rect 9506 5454 9508 5506
rect 9452 5452 9508 5454
rect 9772 5506 9828 5508
rect 9772 5454 9774 5506
rect 9774 5454 9826 5506
rect 9826 5454 9828 5506
rect 9772 5452 9828 5454
rect 10092 5506 10148 5508
rect 10092 5454 10094 5506
rect 10094 5454 10146 5506
rect 10146 5454 10148 5506
rect 10092 5452 10148 5454
rect 10412 5506 10468 5508
rect 10412 5454 10414 5506
rect 10414 5454 10466 5506
rect 10466 5454 10468 5506
rect 10412 5452 10468 5454
rect 10732 5506 10788 5508
rect 10732 5454 10734 5506
rect 10734 5454 10786 5506
rect 10786 5454 10788 5506
rect 10732 5452 10788 5454
rect 11052 5506 11108 5508
rect 11052 5454 11054 5506
rect 11054 5454 11106 5506
rect 11106 5454 11108 5506
rect 11052 5452 11108 5454
rect 11372 5506 11428 5508
rect 11372 5454 11374 5506
rect 11374 5454 11426 5506
rect 11426 5454 11428 5506
rect 11372 5452 11428 5454
rect 11532 5506 11588 5508
rect 11532 5454 11534 5506
rect 11534 5454 11586 5506
rect 11586 5454 11588 5506
rect 11532 5452 11588 5454
rect 11852 5506 11908 5508
rect 11852 5454 11854 5506
rect 11854 5454 11906 5506
rect 11906 5454 11908 5506
rect 11852 5452 11908 5454
rect 12012 5506 12068 5508
rect 12012 5454 12014 5506
rect 12014 5454 12066 5506
rect 12066 5454 12068 5506
rect 12012 5452 12068 5454
rect 12332 5506 12388 5508
rect 12332 5454 12334 5506
rect 12334 5454 12386 5506
rect 12386 5454 12388 5506
rect 12332 5452 12388 5454
rect 8492 5346 8548 5348
rect 8492 5294 8494 5346
rect 8494 5294 8546 5346
rect 8546 5294 8548 5346
rect 8492 5292 8548 5294
rect 8812 5346 8868 5348
rect 8812 5294 8814 5346
rect 8814 5294 8866 5346
rect 8866 5294 8868 5346
rect 8812 5292 8868 5294
rect 8972 5346 9028 5348
rect 8972 5294 8974 5346
rect 8974 5294 9026 5346
rect 9026 5294 9028 5346
rect 8972 5292 9028 5294
rect 9292 5346 9348 5348
rect 9292 5294 9294 5346
rect 9294 5294 9346 5346
rect 9346 5294 9348 5346
rect 9292 5292 9348 5294
rect 9452 5346 9508 5348
rect 9452 5294 9454 5346
rect 9454 5294 9506 5346
rect 9506 5294 9508 5346
rect 9452 5292 9508 5294
rect 9772 5346 9828 5348
rect 9772 5294 9774 5346
rect 9774 5294 9826 5346
rect 9826 5294 9828 5346
rect 9772 5292 9828 5294
rect 10092 5346 10148 5348
rect 10092 5294 10094 5346
rect 10094 5294 10146 5346
rect 10146 5294 10148 5346
rect 10092 5292 10148 5294
rect 10412 5346 10468 5348
rect 10412 5294 10414 5346
rect 10414 5294 10466 5346
rect 10466 5294 10468 5346
rect 10412 5292 10468 5294
rect 10732 5346 10788 5348
rect 10732 5294 10734 5346
rect 10734 5294 10786 5346
rect 10786 5294 10788 5346
rect 10732 5292 10788 5294
rect 11052 5346 11108 5348
rect 11052 5294 11054 5346
rect 11054 5294 11106 5346
rect 11106 5294 11108 5346
rect 11052 5292 11108 5294
rect 11372 5346 11428 5348
rect 11372 5294 11374 5346
rect 11374 5294 11426 5346
rect 11426 5294 11428 5346
rect 11372 5292 11428 5294
rect 11532 5346 11588 5348
rect 11532 5294 11534 5346
rect 11534 5294 11586 5346
rect 11586 5294 11588 5346
rect 11532 5292 11588 5294
rect 11852 5346 11908 5348
rect 11852 5294 11854 5346
rect 11854 5294 11906 5346
rect 11906 5294 11908 5346
rect 11852 5292 11908 5294
rect 12012 5346 12068 5348
rect 12012 5294 12014 5346
rect 12014 5294 12066 5346
rect 12066 5294 12068 5346
rect 12012 5292 12068 5294
rect 12332 5346 12388 5348
rect 12332 5294 12334 5346
rect 12334 5294 12386 5346
rect 12386 5294 12388 5346
rect 12332 5292 12388 5294
rect 8492 5186 8548 5188
rect 8492 5134 8494 5186
rect 8494 5134 8546 5186
rect 8546 5134 8548 5186
rect 8492 5132 8548 5134
rect 8812 5186 8868 5188
rect 8812 5134 8814 5186
rect 8814 5134 8866 5186
rect 8866 5134 8868 5186
rect 8812 5132 8868 5134
rect 8972 5186 9028 5188
rect 8972 5134 8974 5186
rect 8974 5134 9026 5186
rect 9026 5134 9028 5186
rect 8972 5132 9028 5134
rect 9292 5186 9348 5188
rect 9292 5134 9294 5186
rect 9294 5134 9346 5186
rect 9346 5134 9348 5186
rect 9292 5132 9348 5134
rect 9452 5186 9508 5188
rect 9452 5134 9454 5186
rect 9454 5134 9506 5186
rect 9506 5134 9508 5186
rect 9452 5132 9508 5134
rect 9772 5186 9828 5188
rect 9772 5134 9774 5186
rect 9774 5134 9826 5186
rect 9826 5134 9828 5186
rect 9772 5132 9828 5134
rect 10092 5186 10148 5188
rect 10092 5134 10094 5186
rect 10094 5134 10146 5186
rect 10146 5134 10148 5186
rect 10092 5132 10148 5134
rect 10412 5186 10468 5188
rect 10412 5134 10414 5186
rect 10414 5134 10466 5186
rect 10466 5134 10468 5186
rect 10412 5132 10468 5134
rect 10732 5186 10788 5188
rect 10732 5134 10734 5186
rect 10734 5134 10786 5186
rect 10786 5134 10788 5186
rect 10732 5132 10788 5134
rect 11052 5186 11108 5188
rect 11052 5134 11054 5186
rect 11054 5134 11106 5186
rect 11106 5134 11108 5186
rect 11052 5132 11108 5134
rect 11372 5186 11428 5188
rect 11372 5134 11374 5186
rect 11374 5134 11426 5186
rect 11426 5134 11428 5186
rect 11372 5132 11428 5134
rect 11532 5186 11588 5188
rect 11532 5134 11534 5186
rect 11534 5134 11586 5186
rect 11586 5134 11588 5186
rect 11532 5132 11588 5134
rect 11852 5186 11908 5188
rect 11852 5134 11854 5186
rect 11854 5134 11906 5186
rect 11906 5134 11908 5186
rect 11852 5132 11908 5134
rect 12012 5186 12068 5188
rect 12012 5134 12014 5186
rect 12014 5134 12066 5186
rect 12066 5134 12068 5186
rect 12012 5132 12068 5134
rect 12332 5186 12388 5188
rect 12332 5134 12334 5186
rect 12334 5134 12386 5186
rect 12386 5134 12388 5186
rect 12332 5132 12388 5134
rect 8492 5026 8548 5028
rect 8492 4974 8494 5026
rect 8494 4974 8546 5026
rect 8546 4974 8548 5026
rect 8492 4972 8548 4974
rect 8812 5026 8868 5028
rect 8812 4974 8814 5026
rect 8814 4974 8866 5026
rect 8866 4974 8868 5026
rect 8812 4972 8868 4974
rect 8972 5026 9028 5028
rect 8972 4974 8974 5026
rect 8974 4974 9026 5026
rect 9026 4974 9028 5026
rect 8972 4972 9028 4974
rect 9292 5026 9348 5028
rect 9292 4974 9294 5026
rect 9294 4974 9346 5026
rect 9346 4974 9348 5026
rect 9292 4972 9348 4974
rect 9452 5026 9508 5028
rect 9452 4974 9454 5026
rect 9454 4974 9506 5026
rect 9506 4974 9508 5026
rect 9452 4972 9508 4974
rect 9772 5026 9828 5028
rect 9772 4974 9774 5026
rect 9774 4974 9826 5026
rect 9826 4974 9828 5026
rect 9772 4972 9828 4974
rect 10092 5026 10148 5028
rect 10092 4974 10094 5026
rect 10094 4974 10146 5026
rect 10146 4974 10148 5026
rect 10092 4972 10148 4974
rect 10412 5026 10468 5028
rect 10412 4974 10414 5026
rect 10414 4974 10466 5026
rect 10466 4974 10468 5026
rect 10412 4972 10468 4974
rect 10732 5026 10788 5028
rect 10732 4974 10734 5026
rect 10734 4974 10786 5026
rect 10786 4974 10788 5026
rect 10732 4972 10788 4974
rect 11052 5026 11108 5028
rect 11052 4974 11054 5026
rect 11054 4974 11106 5026
rect 11106 4974 11108 5026
rect 11052 4972 11108 4974
rect 11372 5026 11428 5028
rect 11372 4974 11374 5026
rect 11374 4974 11426 5026
rect 11426 4974 11428 5026
rect 11372 4972 11428 4974
rect 11532 5026 11588 5028
rect 11532 4974 11534 5026
rect 11534 4974 11586 5026
rect 11586 4974 11588 5026
rect 11532 4972 11588 4974
rect 11852 5026 11908 5028
rect 11852 4974 11854 5026
rect 11854 4974 11906 5026
rect 11906 4974 11908 5026
rect 11852 4972 11908 4974
rect 12012 5026 12068 5028
rect 12012 4974 12014 5026
rect 12014 4974 12066 5026
rect 12066 4974 12068 5026
rect 12012 4972 12068 4974
rect 12332 5026 12388 5028
rect 12332 4974 12334 5026
rect 12334 4974 12386 5026
rect 12386 4974 12388 5026
rect 12332 4972 12388 4974
rect 8492 4866 8548 4868
rect 8492 4814 8494 4866
rect 8494 4814 8546 4866
rect 8546 4814 8548 4866
rect 8492 4812 8548 4814
rect 8812 4866 8868 4868
rect 8812 4814 8814 4866
rect 8814 4814 8866 4866
rect 8866 4814 8868 4866
rect 8812 4812 8868 4814
rect 8972 4866 9028 4868
rect 8972 4814 8974 4866
rect 8974 4814 9026 4866
rect 9026 4814 9028 4866
rect 8972 4812 9028 4814
rect 9292 4866 9348 4868
rect 9292 4814 9294 4866
rect 9294 4814 9346 4866
rect 9346 4814 9348 4866
rect 9292 4812 9348 4814
rect 9452 4866 9508 4868
rect 9452 4814 9454 4866
rect 9454 4814 9506 4866
rect 9506 4814 9508 4866
rect 9452 4812 9508 4814
rect 9772 4866 9828 4868
rect 9772 4814 9774 4866
rect 9774 4814 9826 4866
rect 9826 4814 9828 4866
rect 9772 4812 9828 4814
rect 10092 4866 10148 4868
rect 10092 4814 10094 4866
rect 10094 4814 10146 4866
rect 10146 4814 10148 4866
rect 10092 4812 10148 4814
rect 10412 4866 10468 4868
rect 10412 4814 10414 4866
rect 10414 4814 10466 4866
rect 10466 4814 10468 4866
rect 10412 4812 10468 4814
rect 10732 4866 10788 4868
rect 10732 4814 10734 4866
rect 10734 4814 10786 4866
rect 10786 4814 10788 4866
rect 10732 4812 10788 4814
rect 11052 4866 11108 4868
rect 11052 4814 11054 4866
rect 11054 4814 11106 4866
rect 11106 4814 11108 4866
rect 11052 4812 11108 4814
rect 11372 4866 11428 4868
rect 11372 4814 11374 4866
rect 11374 4814 11426 4866
rect 11426 4814 11428 4866
rect 11372 4812 11428 4814
rect 11532 4866 11588 4868
rect 11532 4814 11534 4866
rect 11534 4814 11586 4866
rect 11586 4814 11588 4866
rect 11532 4812 11588 4814
rect 11852 4866 11908 4868
rect 11852 4814 11854 4866
rect 11854 4814 11906 4866
rect 11906 4814 11908 4866
rect 11852 4812 11908 4814
rect 12012 4866 12068 4868
rect 12012 4814 12014 4866
rect 12014 4814 12066 4866
rect 12066 4814 12068 4866
rect 12012 4812 12068 4814
rect 12332 4866 12388 4868
rect 12332 4814 12334 4866
rect 12334 4814 12386 4866
rect 12386 4814 12388 4866
rect 12332 4812 12388 4814
rect 8492 4706 8548 4708
rect 8492 4654 8494 4706
rect 8494 4654 8546 4706
rect 8546 4654 8548 4706
rect 8492 4652 8548 4654
rect 8812 4706 8868 4708
rect 8812 4654 8814 4706
rect 8814 4654 8866 4706
rect 8866 4654 8868 4706
rect 8812 4652 8868 4654
rect 8972 4706 9028 4708
rect 8972 4654 8974 4706
rect 8974 4654 9026 4706
rect 9026 4654 9028 4706
rect 8972 4652 9028 4654
rect 9292 4706 9348 4708
rect 9292 4654 9294 4706
rect 9294 4654 9346 4706
rect 9346 4654 9348 4706
rect 9292 4652 9348 4654
rect 9452 4706 9508 4708
rect 9452 4654 9454 4706
rect 9454 4654 9506 4706
rect 9506 4654 9508 4706
rect 9452 4652 9508 4654
rect 9772 4706 9828 4708
rect 9772 4654 9774 4706
rect 9774 4654 9826 4706
rect 9826 4654 9828 4706
rect 9772 4652 9828 4654
rect 10092 4706 10148 4708
rect 10092 4654 10094 4706
rect 10094 4654 10146 4706
rect 10146 4654 10148 4706
rect 10092 4652 10148 4654
rect 10412 4706 10468 4708
rect 10412 4654 10414 4706
rect 10414 4654 10466 4706
rect 10466 4654 10468 4706
rect 10412 4652 10468 4654
rect 10732 4706 10788 4708
rect 10732 4654 10734 4706
rect 10734 4654 10786 4706
rect 10786 4654 10788 4706
rect 10732 4652 10788 4654
rect 11052 4706 11108 4708
rect 11052 4654 11054 4706
rect 11054 4654 11106 4706
rect 11106 4654 11108 4706
rect 11052 4652 11108 4654
rect 11372 4706 11428 4708
rect 11372 4654 11374 4706
rect 11374 4654 11426 4706
rect 11426 4654 11428 4706
rect 11372 4652 11428 4654
rect 11532 4706 11588 4708
rect 11532 4654 11534 4706
rect 11534 4654 11586 4706
rect 11586 4654 11588 4706
rect 11532 4652 11588 4654
rect 11852 4706 11908 4708
rect 11852 4654 11854 4706
rect 11854 4654 11906 4706
rect 11906 4654 11908 4706
rect 11852 4652 11908 4654
rect 12012 4706 12068 4708
rect 12012 4654 12014 4706
rect 12014 4654 12066 4706
rect 12066 4654 12068 4706
rect 12012 4652 12068 4654
rect 12332 4706 12388 4708
rect 12332 4654 12334 4706
rect 12334 4654 12386 4706
rect 12386 4654 12388 4706
rect 12332 4652 12388 4654
rect 8492 4546 8548 4548
rect 8492 4494 8494 4546
rect 8494 4494 8546 4546
rect 8546 4494 8548 4546
rect 8492 4492 8548 4494
rect 8812 4546 8868 4548
rect 8812 4494 8814 4546
rect 8814 4494 8866 4546
rect 8866 4494 8868 4546
rect 8812 4492 8868 4494
rect 8972 4546 9028 4548
rect 8972 4494 8974 4546
rect 8974 4494 9026 4546
rect 9026 4494 9028 4546
rect 8972 4492 9028 4494
rect 9292 4546 9348 4548
rect 9292 4494 9294 4546
rect 9294 4494 9346 4546
rect 9346 4494 9348 4546
rect 9292 4492 9348 4494
rect 9452 4546 9508 4548
rect 9452 4494 9454 4546
rect 9454 4494 9506 4546
rect 9506 4494 9508 4546
rect 9452 4492 9508 4494
rect 9772 4546 9828 4548
rect 9772 4494 9774 4546
rect 9774 4494 9826 4546
rect 9826 4494 9828 4546
rect 9772 4492 9828 4494
rect 10092 4546 10148 4548
rect 10092 4494 10094 4546
rect 10094 4494 10146 4546
rect 10146 4494 10148 4546
rect 10092 4492 10148 4494
rect 10412 4546 10468 4548
rect 10412 4494 10414 4546
rect 10414 4494 10466 4546
rect 10466 4494 10468 4546
rect 10412 4492 10468 4494
rect 10732 4546 10788 4548
rect 10732 4494 10734 4546
rect 10734 4494 10786 4546
rect 10786 4494 10788 4546
rect 10732 4492 10788 4494
rect 11052 4546 11108 4548
rect 11052 4494 11054 4546
rect 11054 4494 11106 4546
rect 11106 4494 11108 4546
rect 11052 4492 11108 4494
rect 11372 4546 11428 4548
rect 11372 4494 11374 4546
rect 11374 4494 11426 4546
rect 11426 4494 11428 4546
rect 11372 4492 11428 4494
rect 11532 4546 11588 4548
rect 11532 4494 11534 4546
rect 11534 4494 11586 4546
rect 11586 4494 11588 4546
rect 11532 4492 11588 4494
rect 11852 4546 11908 4548
rect 11852 4494 11854 4546
rect 11854 4494 11906 4546
rect 11906 4494 11908 4546
rect 11852 4492 11908 4494
rect 12012 4546 12068 4548
rect 12012 4494 12014 4546
rect 12014 4494 12066 4546
rect 12066 4494 12068 4546
rect 12012 4492 12068 4494
rect 12332 4546 12388 4548
rect 12332 4494 12334 4546
rect 12334 4494 12386 4546
rect 12386 4494 12388 4546
rect 12332 4492 12388 4494
rect 8492 4386 8548 4388
rect 8492 4334 8494 4386
rect 8494 4334 8546 4386
rect 8546 4334 8548 4386
rect 8492 4332 8548 4334
rect 8812 4386 8868 4388
rect 8812 4334 8814 4386
rect 8814 4334 8866 4386
rect 8866 4334 8868 4386
rect 8812 4332 8868 4334
rect 8972 4386 9028 4388
rect 8972 4334 8974 4386
rect 8974 4334 9026 4386
rect 9026 4334 9028 4386
rect 8972 4332 9028 4334
rect 9292 4386 9348 4388
rect 9292 4334 9294 4386
rect 9294 4334 9346 4386
rect 9346 4334 9348 4386
rect 9292 4332 9348 4334
rect 9452 4386 9508 4388
rect 9452 4334 9454 4386
rect 9454 4334 9506 4386
rect 9506 4334 9508 4386
rect 9452 4332 9508 4334
rect 9772 4386 9828 4388
rect 9772 4334 9774 4386
rect 9774 4334 9826 4386
rect 9826 4334 9828 4386
rect 9772 4332 9828 4334
rect 10092 4386 10148 4388
rect 10092 4334 10094 4386
rect 10094 4334 10146 4386
rect 10146 4334 10148 4386
rect 10092 4332 10148 4334
rect 10412 4386 10468 4388
rect 10412 4334 10414 4386
rect 10414 4334 10466 4386
rect 10466 4334 10468 4386
rect 10412 4332 10468 4334
rect 10732 4386 10788 4388
rect 10732 4334 10734 4386
rect 10734 4334 10786 4386
rect 10786 4334 10788 4386
rect 10732 4332 10788 4334
rect 11052 4386 11108 4388
rect 11052 4334 11054 4386
rect 11054 4334 11106 4386
rect 11106 4334 11108 4386
rect 11052 4332 11108 4334
rect 11372 4386 11428 4388
rect 11372 4334 11374 4386
rect 11374 4334 11426 4386
rect 11426 4334 11428 4386
rect 11372 4332 11428 4334
rect 11532 4386 11588 4388
rect 11532 4334 11534 4386
rect 11534 4334 11586 4386
rect 11586 4334 11588 4386
rect 11532 4332 11588 4334
rect 11852 4386 11908 4388
rect 11852 4334 11854 4386
rect 11854 4334 11906 4386
rect 11906 4334 11908 4386
rect 11852 4332 11908 4334
rect 12012 4386 12068 4388
rect 12012 4334 12014 4386
rect 12014 4334 12066 4386
rect 12066 4334 12068 4386
rect 12012 4332 12068 4334
rect 12332 4386 12388 4388
rect 12332 4334 12334 4386
rect 12334 4334 12386 4386
rect 12386 4334 12388 4386
rect 12332 4332 12388 4334
rect 8492 4226 8548 4228
rect 8492 4174 8494 4226
rect 8494 4174 8546 4226
rect 8546 4174 8548 4226
rect 8492 4172 8548 4174
rect 8812 4226 8868 4228
rect 8812 4174 8814 4226
rect 8814 4174 8866 4226
rect 8866 4174 8868 4226
rect 8812 4172 8868 4174
rect 8972 4226 9028 4228
rect 8972 4174 8974 4226
rect 8974 4174 9026 4226
rect 9026 4174 9028 4226
rect 8972 4172 9028 4174
rect 9292 4226 9348 4228
rect 9292 4174 9294 4226
rect 9294 4174 9346 4226
rect 9346 4174 9348 4226
rect 9292 4172 9348 4174
rect 9452 4226 9508 4228
rect 9452 4174 9454 4226
rect 9454 4174 9506 4226
rect 9506 4174 9508 4226
rect 9452 4172 9508 4174
rect 9772 4226 9828 4228
rect 9772 4174 9774 4226
rect 9774 4174 9826 4226
rect 9826 4174 9828 4226
rect 9772 4172 9828 4174
rect 10092 4226 10148 4228
rect 10092 4174 10094 4226
rect 10094 4174 10146 4226
rect 10146 4174 10148 4226
rect 10092 4172 10148 4174
rect 10412 4226 10468 4228
rect 10412 4174 10414 4226
rect 10414 4174 10466 4226
rect 10466 4174 10468 4226
rect 10412 4172 10468 4174
rect 10732 4226 10788 4228
rect 10732 4174 10734 4226
rect 10734 4174 10786 4226
rect 10786 4174 10788 4226
rect 10732 4172 10788 4174
rect 11052 4226 11108 4228
rect 11052 4174 11054 4226
rect 11054 4174 11106 4226
rect 11106 4174 11108 4226
rect 11052 4172 11108 4174
rect 11372 4226 11428 4228
rect 11372 4174 11374 4226
rect 11374 4174 11426 4226
rect 11426 4174 11428 4226
rect 11372 4172 11428 4174
rect 11532 4226 11588 4228
rect 11532 4174 11534 4226
rect 11534 4174 11586 4226
rect 11586 4174 11588 4226
rect 11532 4172 11588 4174
rect 11852 4226 11908 4228
rect 11852 4174 11854 4226
rect 11854 4174 11906 4226
rect 11906 4174 11908 4226
rect 11852 4172 11908 4174
rect 12012 4226 12068 4228
rect 12012 4174 12014 4226
rect 12014 4174 12066 4226
rect 12066 4174 12068 4226
rect 12012 4172 12068 4174
rect 12332 4226 12388 4228
rect 12332 4174 12334 4226
rect 12334 4174 12386 4226
rect 12386 4174 12388 4226
rect 12332 4172 12388 4174
rect 8492 4066 8548 4068
rect 8492 4014 8494 4066
rect 8494 4014 8546 4066
rect 8546 4014 8548 4066
rect 8492 4012 8548 4014
rect 8812 4066 8868 4068
rect 8812 4014 8814 4066
rect 8814 4014 8866 4066
rect 8866 4014 8868 4066
rect 8812 4012 8868 4014
rect 8972 4066 9028 4068
rect 8972 4014 8974 4066
rect 8974 4014 9026 4066
rect 9026 4014 9028 4066
rect 8972 4012 9028 4014
rect 9292 4066 9348 4068
rect 9292 4014 9294 4066
rect 9294 4014 9346 4066
rect 9346 4014 9348 4066
rect 9292 4012 9348 4014
rect 9452 4066 9508 4068
rect 9452 4014 9454 4066
rect 9454 4014 9506 4066
rect 9506 4014 9508 4066
rect 9452 4012 9508 4014
rect 9772 4066 9828 4068
rect 9772 4014 9774 4066
rect 9774 4014 9826 4066
rect 9826 4014 9828 4066
rect 9772 4012 9828 4014
rect 10092 4066 10148 4068
rect 10092 4014 10094 4066
rect 10094 4014 10146 4066
rect 10146 4014 10148 4066
rect 10092 4012 10148 4014
rect 10412 4066 10468 4068
rect 10412 4014 10414 4066
rect 10414 4014 10466 4066
rect 10466 4014 10468 4066
rect 10412 4012 10468 4014
rect 10732 4066 10788 4068
rect 10732 4014 10734 4066
rect 10734 4014 10786 4066
rect 10786 4014 10788 4066
rect 10732 4012 10788 4014
rect 11052 4066 11108 4068
rect 11052 4014 11054 4066
rect 11054 4014 11106 4066
rect 11106 4014 11108 4066
rect 11052 4012 11108 4014
rect 11372 4066 11428 4068
rect 11372 4014 11374 4066
rect 11374 4014 11426 4066
rect 11426 4014 11428 4066
rect 11372 4012 11428 4014
rect 11532 4066 11588 4068
rect 11532 4014 11534 4066
rect 11534 4014 11586 4066
rect 11586 4014 11588 4066
rect 11532 4012 11588 4014
rect 11852 4066 11908 4068
rect 11852 4014 11854 4066
rect 11854 4014 11906 4066
rect 11906 4014 11908 4066
rect 11852 4012 11908 4014
rect 12012 4066 12068 4068
rect 12012 4014 12014 4066
rect 12014 4014 12066 4066
rect 12066 4014 12068 4066
rect 12012 4012 12068 4014
rect 12332 4066 12388 4068
rect 12332 4014 12334 4066
rect 12334 4014 12386 4066
rect 12386 4014 12388 4066
rect 12332 4012 12388 4014
rect 8492 3906 8548 3908
rect 8492 3854 8494 3906
rect 8494 3854 8546 3906
rect 8546 3854 8548 3906
rect 8492 3852 8548 3854
rect 8812 3906 8868 3908
rect 8812 3854 8814 3906
rect 8814 3854 8866 3906
rect 8866 3854 8868 3906
rect 8812 3852 8868 3854
rect 8972 3906 9028 3908
rect 8972 3854 8974 3906
rect 8974 3854 9026 3906
rect 9026 3854 9028 3906
rect 8972 3852 9028 3854
rect 9292 3906 9348 3908
rect 9292 3854 9294 3906
rect 9294 3854 9346 3906
rect 9346 3854 9348 3906
rect 9292 3852 9348 3854
rect 9452 3906 9508 3908
rect 9452 3854 9454 3906
rect 9454 3854 9506 3906
rect 9506 3854 9508 3906
rect 9452 3852 9508 3854
rect 9772 3906 9828 3908
rect 9772 3854 9774 3906
rect 9774 3854 9826 3906
rect 9826 3854 9828 3906
rect 9772 3852 9828 3854
rect 10092 3906 10148 3908
rect 10092 3854 10094 3906
rect 10094 3854 10146 3906
rect 10146 3854 10148 3906
rect 10092 3852 10148 3854
rect 10412 3906 10468 3908
rect 10412 3854 10414 3906
rect 10414 3854 10466 3906
rect 10466 3854 10468 3906
rect 10412 3852 10468 3854
rect 10732 3906 10788 3908
rect 10732 3854 10734 3906
rect 10734 3854 10786 3906
rect 10786 3854 10788 3906
rect 10732 3852 10788 3854
rect 11052 3906 11108 3908
rect 11052 3854 11054 3906
rect 11054 3854 11106 3906
rect 11106 3854 11108 3906
rect 11052 3852 11108 3854
rect 11372 3906 11428 3908
rect 11372 3854 11374 3906
rect 11374 3854 11426 3906
rect 11426 3854 11428 3906
rect 11372 3852 11428 3854
rect 11532 3906 11588 3908
rect 11532 3854 11534 3906
rect 11534 3854 11586 3906
rect 11586 3854 11588 3906
rect 11532 3852 11588 3854
rect 11852 3906 11908 3908
rect 11852 3854 11854 3906
rect 11854 3854 11906 3906
rect 11906 3854 11908 3906
rect 11852 3852 11908 3854
rect 12012 3906 12068 3908
rect 12012 3854 12014 3906
rect 12014 3854 12066 3906
rect 12066 3854 12068 3906
rect 12012 3852 12068 3854
rect 12332 3906 12388 3908
rect 12332 3854 12334 3906
rect 12334 3854 12386 3906
rect 12386 3854 12388 3906
rect 12332 3852 12388 3854
rect 9132 3612 9188 3668
rect 8492 3426 8548 3428
rect 8492 3374 8494 3426
rect 8494 3374 8546 3426
rect 8546 3374 8548 3426
rect 8492 3372 8548 3374
rect 8812 3426 8868 3428
rect 8812 3374 8814 3426
rect 8814 3374 8866 3426
rect 8866 3374 8868 3426
rect 8812 3372 8868 3374
rect 8972 3426 9028 3428
rect 8972 3374 8974 3426
rect 8974 3374 9026 3426
rect 9026 3374 9028 3426
rect 8972 3372 9028 3374
rect 9292 3426 9348 3428
rect 9292 3374 9294 3426
rect 9294 3374 9346 3426
rect 9346 3374 9348 3426
rect 9292 3372 9348 3374
rect 9452 3426 9508 3428
rect 9452 3374 9454 3426
rect 9454 3374 9506 3426
rect 9506 3374 9508 3426
rect 9452 3372 9508 3374
rect 9772 3426 9828 3428
rect 9772 3374 9774 3426
rect 9774 3374 9826 3426
rect 9826 3374 9828 3426
rect 9772 3372 9828 3374
rect 10092 3426 10148 3428
rect 10092 3374 10094 3426
rect 10094 3374 10146 3426
rect 10146 3374 10148 3426
rect 10092 3372 10148 3374
rect 10412 3426 10468 3428
rect 10412 3374 10414 3426
rect 10414 3374 10466 3426
rect 10466 3374 10468 3426
rect 10412 3372 10468 3374
rect 10732 3426 10788 3428
rect 10732 3374 10734 3426
rect 10734 3374 10786 3426
rect 10786 3374 10788 3426
rect 10732 3372 10788 3374
rect 11052 3426 11108 3428
rect 11052 3374 11054 3426
rect 11054 3374 11106 3426
rect 11106 3374 11108 3426
rect 11052 3372 11108 3374
rect 11372 3426 11428 3428
rect 11372 3374 11374 3426
rect 11374 3374 11426 3426
rect 11426 3374 11428 3426
rect 11372 3372 11428 3374
rect 11532 3426 11588 3428
rect 11532 3374 11534 3426
rect 11534 3374 11586 3426
rect 11586 3374 11588 3426
rect 11532 3372 11588 3374
rect 11852 3426 11908 3428
rect 11852 3374 11854 3426
rect 11854 3374 11906 3426
rect 11906 3374 11908 3426
rect 11852 3372 11908 3374
rect 12012 3426 12068 3428
rect 12012 3374 12014 3426
rect 12014 3374 12066 3426
rect 12066 3374 12068 3426
rect 12012 3372 12068 3374
rect 12332 3426 12388 3428
rect 12332 3374 12334 3426
rect 12334 3374 12386 3426
rect 12386 3374 12388 3426
rect 12332 3372 12388 3374
rect 8492 3266 8548 3268
rect 8492 3214 8494 3266
rect 8494 3214 8546 3266
rect 8546 3214 8548 3266
rect 8492 3212 8548 3214
rect 8812 3266 8868 3268
rect 8812 3214 8814 3266
rect 8814 3214 8866 3266
rect 8866 3214 8868 3266
rect 8812 3212 8868 3214
rect 8972 3266 9028 3268
rect 8972 3214 8974 3266
rect 8974 3214 9026 3266
rect 9026 3214 9028 3266
rect 8972 3212 9028 3214
rect 9292 3266 9348 3268
rect 9292 3214 9294 3266
rect 9294 3214 9346 3266
rect 9346 3214 9348 3266
rect 9292 3212 9348 3214
rect 9452 3266 9508 3268
rect 9452 3214 9454 3266
rect 9454 3214 9506 3266
rect 9506 3214 9508 3266
rect 9452 3212 9508 3214
rect 9772 3266 9828 3268
rect 9772 3214 9774 3266
rect 9774 3214 9826 3266
rect 9826 3214 9828 3266
rect 9772 3212 9828 3214
rect 10092 3266 10148 3268
rect 10092 3214 10094 3266
rect 10094 3214 10146 3266
rect 10146 3214 10148 3266
rect 10092 3212 10148 3214
rect 10412 3266 10468 3268
rect 10412 3214 10414 3266
rect 10414 3214 10466 3266
rect 10466 3214 10468 3266
rect 10412 3212 10468 3214
rect 10732 3266 10788 3268
rect 10732 3214 10734 3266
rect 10734 3214 10786 3266
rect 10786 3214 10788 3266
rect 10732 3212 10788 3214
rect 11052 3266 11108 3268
rect 11052 3214 11054 3266
rect 11054 3214 11106 3266
rect 11106 3214 11108 3266
rect 11052 3212 11108 3214
rect 11372 3266 11428 3268
rect 11372 3214 11374 3266
rect 11374 3214 11426 3266
rect 11426 3214 11428 3266
rect 11372 3212 11428 3214
rect 11532 3266 11588 3268
rect 11532 3214 11534 3266
rect 11534 3214 11586 3266
rect 11586 3214 11588 3266
rect 11532 3212 11588 3214
rect 11852 3266 11908 3268
rect 11852 3214 11854 3266
rect 11854 3214 11906 3266
rect 11906 3214 11908 3266
rect 11852 3212 11908 3214
rect 12012 3266 12068 3268
rect 12012 3214 12014 3266
rect 12014 3214 12066 3266
rect 12066 3214 12068 3266
rect 12012 3212 12068 3214
rect 12332 3266 12388 3268
rect 12332 3214 12334 3266
rect 12334 3214 12386 3266
rect 12386 3214 12388 3266
rect 12332 3212 12388 3214
rect 8492 3106 8548 3108
rect 8492 3054 8494 3106
rect 8494 3054 8546 3106
rect 8546 3054 8548 3106
rect 8492 3052 8548 3054
rect 8812 3106 8868 3108
rect 8812 3054 8814 3106
rect 8814 3054 8866 3106
rect 8866 3054 8868 3106
rect 8812 3052 8868 3054
rect 8972 3106 9028 3108
rect 8972 3054 8974 3106
rect 8974 3054 9026 3106
rect 9026 3054 9028 3106
rect 8972 3052 9028 3054
rect 9292 3106 9348 3108
rect 9292 3054 9294 3106
rect 9294 3054 9346 3106
rect 9346 3054 9348 3106
rect 9292 3052 9348 3054
rect 9452 3106 9508 3108
rect 9452 3054 9454 3106
rect 9454 3054 9506 3106
rect 9506 3054 9508 3106
rect 9452 3052 9508 3054
rect 9772 3106 9828 3108
rect 9772 3054 9774 3106
rect 9774 3054 9826 3106
rect 9826 3054 9828 3106
rect 9772 3052 9828 3054
rect 10092 3106 10148 3108
rect 10092 3054 10094 3106
rect 10094 3054 10146 3106
rect 10146 3054 10148 3106
rect 10092 3052 10148 3054
rect 10412 3106 10468 3108
rect 10412 3054 10414 3106
rect 10414 3054 10466 3106
rect 10466 3054 10468 3106
rect 10412 3052 10468 3054
rect 10732 3106 10788 3108
rect 10732 3054 10734 3106
rect 10734 3054 10786 3106
rect 10786 3054 10788 3106
rect 10732 3052 10788 3054
rect 11052 3106 11108 3108
rect 11052 3054 11054 3106
rect 11054 3054 11106 3106
rect 11106 3054 11108 3106
rect 11052 3052 11108 3054
rect 11372 3106 11428 3108
rect 11372 3054 11374 3106
rect 11374 3054 11426 3106
rect 11426 3054 11428 3106
rect 11372 3052 11428 3054
rect 11532 3106 11588 3108
rect 11532 3054 11534 3106
rect 11534 3054 11586 3106
rect 11586 3054 11588 3106
rect 11532 3052 11588 3054
rect 11852 3106 11908 3108
rect 11852 3054 11854 3106
rect 11854 3054 11906 3106
rect 11906 3054 11908 3106
rect 11852 3052 11908 3054
rect 12012 3106 12068 3108
rect 12012 3054 12014 3106
rect 12014 3054 12066 3106
rect 12066 3054 12068 3106
rect 12012 3052 12068 3054
rect 12332 3106 12388 3108
rect 12332 3054 12334 3106
rect 12334 3054 12386 3106
rect 12386 3054 12388 3106
rect 12332 3052 12388 3054
rect 8492 2946 8548 2948
rect 8492 2894 8494 2946
rect 8494 2894 8546 2946
rect 8546 2894 8548 2946
rect 8492 2892 8548 2894
rect 8812 2946 8868 2948
rect 8812 2894 8814 2946
rect 8814 2894 8866 2946
rect 8866 2894 8868 2946
rect 8812 2892 8868 2894
rect 8972 2946 9028 2948
rect 8972 2894 8974 2946
rect 8974 2894 9026 2946
rect 9026 2894 9028 2946
rect 8972 2892 9028 2894
rect 9292 2946 9348 2948
rect 9292 2894 9294 2946
rect 9294 2894 9346 2946
rect 9346 2894 9348 2946
rect 9292 2892 9348 2894
rect 9452 2946 9508 2948
rect 9452 2894 9454 2946
rect 9454 2894 9506 2946
rect 9506 2894 9508 2946
rect 9452 2892 9508 2894
rect 9772 2946 9828 2948
rect 9772 2894 9774 2946
rect 9774 2894 9826 2946
rect 9826 2894 9828 2946
rect 9772 2892 9828 2894
rect 10092 2946 10148 2948
rect 10092 2894 10094 2946
rect 10094 2894 10146 2946
rect 10146 2894 10148 2946
rect 10092 2892 10148 2894
rect 10412 2946 10468 2948
rect 10412 2894 10414 2946
rect 10414 2894 10466 2946
rect 10466 2894 10468 2946
rect 10412 2892 10468 2894
rect 10732 2946 10788 2948
rect 10732 2894 10734 2946
rect 10734 2894 10786 2946
rect 10786 2894 10788 2946
rect 10732 2892 10788 2894
rect 11052 2946 11108 2948
rect 11052 2894 11054 2946
rect 11054 2894 11106 2946
rect 11106 2894 11108 2946
rect 11052 2892 11108 2894
rect 11372 2946 11428 2948
rect 11372 2894 11374 2946
rect 11374 2894 11426 2946
rect 11426 2894 11428 2946
rect 11372 2892 11428 2894
rect 11532 2946 11588 2948
rect 11532 2894 11534 2946
rect 11534 2894 11586 2946
rect 11586 2894 11588 2946
rect 11532 2892 11588 2894
rect 11852 2946 11908 2948
rect 11852 2894 11854 2946
rect 11854 2894 11906 2946
rect 11906 2894 11908 2946
rect 11852 2892 11908 2894
rect 12012 2946 12068 2948
rect 12012 2894 12014 2946
rect 12014 2894 12066 2946
rect 12066 2894 12068 2946
rect 12012 2892 12068 2894
rect 12332 2946 12388 2948
rect 12332 2894 12334 2946
rect 12334 2894 12386 2946
rect 12386 2894 12388 2946
rect 12332 2892 12388 2894
rect 8492 2786 8548 2788
rect 8492 2734 8494 2786
rect 8494 2734 8546 2786
rect 8546 2734 8548 2786
rect 8492 2732 8548 2734
rect 8812 2786 8868 2788
rect 8812 2734 8814 2786
rect 8814 2734 8866 2786
rect 8866 2734 8868 2786
rect 8812 2732 8868 2734
rect 8972 2786 9028 2788
rect 8972 2734 8974 2786
rect 8974 2734 9026 2786
rect 9026 2734 9028 2786
rect 8972 2732 9028 2734
rect 9292 2786 9348 2788
rect 9292 2734 9294 2786
rect 9294 2734 9346 2786
rect 9346 2734 9348 2786
rect 9292 2732 9348 2734
rect 9452 2786 9508 2788
rect 9452 2734 9454 2786
rect 9454 2734 9506 2786
rect 9506 2734 9508 2786
rect 9452 2732 9508 2734
rect 9772 2786 9828 2788
rect 9772 2734 9774 2786
rect 9774 2734 9826 2786
rect 9826 2734 9828 2786
rect 9772 2732 9828 2734
rect 10092 2786 10148 2788
rect 10092 2734 10094 2786
rect 10094 2734 10146 2786
rect 10146 2734 10148 2786
rect 10092 2732 10148 2734
rect 10412 2786 10468 2788
rect 10412 2734 10414 2786
rect 10414 2734 10466 2786
rect 10466 2734 10468 2786
rect 10412 2732 10468 2734
rect 10732 2786 10788 2788
rect 10732 2734 10734 2786
rect 10734 2734 10786 2786
rect 10786 2734 10788 2786
rect 10732 2732 10788 2734
rect 11052 2786 11108 2788
rect 11052 2734 11054 2786
rect 11054 2734 11106 2786
rect 11106 2734 11108 2786
rect 11052 2732 11108 2734
rect 11372 2786 11428 2788
rect 11372 2734 11374 2786
rect 11374 2734 11426 2786
rect 11426 2734 11428 2786
rect 11372 2732 11428 2734
rect 11532 2786 11588 2788
rect 11532 2734 11534 2786
rect 11534 2734 11586 2786
rect 11586 2734 11588 2786
rect 11532 2732 11588 2734
rect 11852 2786 11908 2788
rect 11852 2734 11854 2786
rect 11854 2734 11906 2786
rect 11906 2734 11908 2786
rect 11852 2732 11908 2734
rect 12012 2786 12068 2788
rect 12012 2734 12014 2786
rect 12014 2734 12066 2786
rect 12066 2734 12068 2786
rect 12012 2732 12068 2734
rect 12332 2786 12388 2788
rect 12332 2734 12334 2786
rect 12334 2734 12386 2786
rect 12386 2734 12388 2786
rect 12332 2732 12388 2734
rect 8492 2626 8548 2628
rect 8492 2574 8494 2626
rect 8494 2574 8546 2626
rect 8546 2574 8548 2626
rect 8492 2572 8548 2574
rect 8812 2626 8868 2628
rect 8812 2574 8814 2626
rect 8814 2574 8866 2626
rect 8866 2574 8868 2626
rect 8812 2572 8868 2574
rect 8972 2626 9028 2628
rect 8972 2574 8974 2626
rect 8974 2574 9026 2626
rect 9026 2574 9028 2626
rect 8972 2572 9028 2574
rect 9292 2626 9348 2628
rect 9292 2574 9294 2626
rect 9294 2574 9346 2626
rect 9346 2574 9348 2626
rect 9292 2572 9348 2574
rect 9452 2626 9508 2628
rect 9452 2574 9454 2626
rect 9454 2574 9506 2626
rect 9506 2574 9508 2626
rect 9452 2572 9508 2574
rect 9772 2626 9828 2628
rect 9772 2574 9774 2626
rect 9774 2574 9826 2626
rect 9826 2574 9828 2626
rect 9772 2572 9828 2574
rect 10092 2626 10148 2628
rect 10092 2574 10094 2626
rect 10094 2574 10146 2626
rect 10146 2574 10148 2626
rect 10092 2572 10148 2574
rect 10412 2626 10468 2628
rect 10412 2574 10414 2626
rect 10414 2574 10466 2626
rect 10466 2574 10468 2626
rect 10412 2572 10468 2574
rect 10732 2626 10788 2628
rect 10732 2574 10734 2626
rect 10734 2574 10786 2626
rect 10786 2574 10788 2626
rect 10732 2572 10788 2574
rect 11052 2626 11108 2628
rect 11052 2574 11054 2626
rect 11054 2574 11106 2626
rect 11106 2574 11108 2626
rect 11052 2572 11108 2574
rect 11372 2626 11428 2628
rect 11372 2574 11374 2626
rect 11374 2574 11426 2626
rect 11426 2574 11428 2626
rect 11372 2572 11428 2574
rect 11532 2626 11588 2628
rect 11532 2574 11534 2626
rect 11534 2574 11586 2626
rect 11586 2574 11588 2626
rect 11532 2572 11588 2574
rect 11852 2626 11908 2628
rect 11852 2574 11854 2626
rect 11854 2574 11906 2626
rect 11906 2574 11908 2626
rect 11852 2572 11908 2574
rect 12012 2626 12068 2628
rect 12012 2574 12014 2626
rect 12014 2574 12066 2626
rect 12066 2574 12068 2626
rect 12012 2572 12068 2574
rect 12332 2626 12388 2628
rect 12332 2574 12334 2626
rect 12334 2574 12386 2626
rect 12386 2574 12388 2626
rect 12332 2572 12388 2574
rect 8492 2466 8548 2468
rect 8492 2414 8494 2466
rect 8494 2414 8546 2466
rect 8546 2414 8548 2466
rect 8492 2412 8548 2414
rect 8812 2466 8868 2468
rect 8812 2414 8814 2466
rect 8814 2414 8866 2466
rect 8866 2414 8868 2466
rect 8812 2412 8868 2414
rect 8972 2466 9028 2468
rect 8972 2414 8974 2466
rect 8974 2414 9026 2466
rect 9026 2414 9028 2466
rect 8972 2412 9028 2414
rect 9292 2466 9348 2468
rect 9292 2414 9294 2466
rect 9294 2414 9346 2466
rect 9346 2414 9348 2466
rect 9292 2412 9348 2414
rect 9452 2466 9508 2468
rect 9452 2414 9454 2466
rect 9454 2414 9506 2466
rect 9506 2414 9508 2466
rect 9452 2412 9508 2414
rect 9772 2466 9828 2468
rect 9772 2414 9774 2466
rect 9774 2414 9826 2466
rect 9826 2414 9828 2466
rect 9772 2412 9828 2414
rect 10092 2466 10148 2468
rect 10092 2414 10094 2466
rect 10094 2414 10146 2466
rect 10146 2414 10148 2466
rect 10092 2412 10148 2414
rect 10412 2466 10468 2468
rect 10412 2414 10414 2466
rect 10414 2414 10466 2466
rect 10466 2414 10468 2466
rect 10412 2412 10468 2414
rect 10732 2466 10788 2468
rect 10732 2414 10734 2466
rect 10734 2414 10786 2466
rect 10786 2414 10788 2466
rect 10732 2412 10788 2414
rect 11052 2466 11108 2468
rect 11052 2414 11054 2466
rect 11054 2414 11106 2466
rect 11106 2414 11108 2466
rect 11052 2412 11108 2414
rect 11372 2466 11428 2468
rect 11372 2414 11374 2466
rect 11374 2414 11426 2466
rect 11426 2414 11428 2466
rect 11372 2412 11428 2414
rect 11532 2466 11588 2468
rect 11532 2414 11534 2466
rect 11534 2414 11586 2466
rect 11586 2414 11588 2466
rect 11532 2412 11588 2414
rect 11852 2466 11908 2468
rect 11852 2414 11854 2466
rect 11854 2414 11906 2466
rect 11906 2414 11908 2466
rect 11852 2412 11908 2414
rect 12012 2466 12068 2468
rect 12012 2414 12014 2466
rect 12014 2414 12066 2466
rect 12066 2414 12068 2466
rect 12012 2412 12068 2414
rect 12332 2466 12388 2468
rect 12332 2414 12334 2466
rect 12334 2414 12386 2466
rect 12386 2414 12388 2466
rect 12332 2412 12388 2414
rect 8492 2306 8548 2308
rect 8492 2254 8494 2306
rect 8494 2254 8546 2306
rect 8546 2254 8548 2306
rect 8492 2252 8548 2254
rect 8812 2306 8868 2308
rect 8812 2254 8814 2306
rect 8814 2254 8866 2306
rect 8866 2254 8868 2306
rect 8812 2252 8868 2254
rect 8972 2306 9028 2308
rect 8972 2254 8974 2306
rect 8974 2254 9026 2306
rect 9026 2254 9028 2306
rect 8972 2252 9028 2254
rect 9292 2306 9348 2308
rect 9292 2254 9294 2306
rect 9294 2254 9346 2306
rect 9346 2254 9348 2306
rect 9292 2252 9348 2254
rect 9452 2306 9508 2308
rect 9452 2254 9454 2306
rect 9454 2254 9506 2306
rect 9506 2254 9508 2306
rect 9452 2252 9508 2254
rect 9772 2306 9828 2308
rect 9772 2254 9774 2306
rect 9774 2254 9826 2306
rect 9826 2254 9828 2306
rect 9772 2252 9828 2254
rect 10092 2306 10148 2308
rect 10092 2254 10094 2306
rect 10094 2254 10146 2306
rect 10146 2254 10148 2306
rect 10092 2252 10148 2254
rect 10412 2306 10468 2308
rect 10412 2254 10414 2306
rect 10414 2254 10466 2306
rect 10466 2254 10468 2306
rect 10412 2252 10468 2254
rect 10732 2306 10788 2308
rect 10732 2254 10734 2306
rect 10734 2254 10786 2306
rect 10786 2254 10788 2306
rect 10732 2252 10788 2254
rect 11052 2306 11108 2308
rect 11052 2254 11054 2306
rect 11054 2254 11106 2306
rect 11106 2254 11108 2306
rect 11052 2252 11108 2254
rect 11372 2306 11428 2308
rect 11372 2254 11374 2306
rect 11374 2254 11426 2306
rect 11426 2254 11428 2306
rect 11372 2252 11428 2254
rect 11532 2306 11588 2308
rect 11532 2254 11534 2306
rect 11534 2254 11586 2306
rect 11586 2254 11588 2306
rect 11532 2252 11588 2254
rect 11852 2306 11908 2308
rect 11852 2254 11854 2306
rect 11854 2254 11906 2306
rect 11906 2254 11908 2306
rect 11852 2252 11908 2254
rect 12012 2306 12068 2308
rect 12012 2254 12014 2306
rect 12014 2254 12066 2306
rect 12066 2254 12068 2306
rect 12012 2252 12068 2254
rect 12332 2306 12388 2308
rect 12332 2254 12334 2306
rect 12334 2254 12386 2306
rect 12386 2254 12388 2306
rect 12332 2252 12388 2254
rect 8492 2146 8548 2148
rect 8492 2094 8494 2146
rect 8494 2094 8546 2146
rect 8546 2094 8548 2146
rect 8492 2092 8548 2094
rect 8812 2146 8868 2148
rect 8812 2094 8814 2146
rect 8814 2094 8866 2146
rect 8866 2094 8868 2146
rect 8812 2092 8868 2094
rect 8972 2146 9028 2148
rect 8972 2094 8974 2146
rect 8974 2094 9026 2146
rect 9026 2094 9028 2146
rect 8972 2092 9028 2094
rect 9292 2146 9348 2148
rect 9292 2094 9294 2146
rect 9294 2094 9346 2146
rect 9346 2094 9348 2146
rect 9292 2092 9348 2094
rect 9452 2146 9508 2148
rect 9452 2094 9454 2146
rect 9454 2094 9506 2146
rect 9506 2094 9508 2146
rect 9452 2092 9508 2094
rect 9772 2146 9828 2148
rect 9772 2094 9774 2146
rect 9774 2094 9826 2146
rect 9826 2094 9828 2146
rect 9772 2092 9828 2094
rect 10092 2146 10148 2148
rect 10092 2094 10094 2146
rect 10094 2094 10146 2146
rect 10146 2094 10148 2146
rect 10092 2092 10148 2094
rect 10412 2146 10468 2148
rect 10412 2094 10414 2146
rect 10414 2094 10466 2146
rect 10466 2094 10468 2146
rect 10412 2092 10468 2094
rect 10732 2146 10788 2148
rect 10732 2094 10734 2146
rect 10734 2094 10786 2146
rect 10786 2094 10788 2146
rect 10732 2092 10788 2094
rect 11052 2146 11108 2148
rect 11052 2094 11054 2146
rect 11054 2094 11106 2146
rect 11106 2094 11108 2146
rect 11052 2092 11108 2094
rect 11372 2146 11428 2148
rect 11372 2094 11374 2146
rect 11374 2094 11426 2146
rect 11426 2094 11428 2146
rect 11372 2092 11428 2094
rect 11532 2146 11588 2148
rect 11532 2094 11534 2146
rect 11534 2094 11586 2146
rect 11586 2094 11588 2146
rect 11532 2092 11588 2094
rect 11852 2146 11908 2148
rect 11852 2094 11854 2146
rect 11854 2094 11906 2146
rect 11906 2094 11908 2146
rect 11852 2092 11908 2094
rect 12012 2146 12068 2148
rect 12012 2094 12014 2146
rect 12014 2094 12066 2146
rect 12066 2094 12068 2146
rect 12012 2092 12068 2094
rect 12332 2146 12388 2148
rect 12332 2094 12334 2146
rect 12334 2094 12386 2146
rect 12386 2094 12388 2146
rect 12332 2092 12388 2094
rect 8492 1986 8548 1988
rect 8492 1934 8494 1986
rect 8494 1934 8546 1986
rect 8546 1934 8548 1986
rect 8492 1932 8548 1934
rect 8812 1986 8868 1988
rect 8812 1934 8814 1986
rect 8814 1934 8866 1986
rect 8866 1934 8868 1986
rect 8812 1932 8868 1934
rect 8972 1986 9028 1988
rect 8972 1934 8974 1986
rect 8974 1934 9026 1986
rect 9026 1934 9028 1986
rect 8972 1932 9028 1934
rect 9292 1986 9348 1988
rect 9292 1934 9294 1986
rect 9294 1934 9346 1986
rect 9346 1934 9348 1986
rect 9292 1932 9348 1934
rect 9452 1986 9508 1988
rect 9452 1934 9454 1986
rect 9454 1934 9506 1986
rect 9506 1934 9508 1986
rect 9452 1932 9508 1934
rect 9772 1986 9828 1988
rect 9772 1934 9774 1986
rect 9774 1934 9826 1986
rect 9826 1934 9828 1986
rect 9772 1932 9828 1934
rect 10092 1986 10148 1988
rect 10092 1934 10094 1986
rect 10094 1934 10146 1986
rect 10146 1934 10148 1986
rect 10092 1932 10148 1934
rect 10412 1986 10468 1988
rect 10412 1934 10414 1986
rect 10414 1934 10466 1986
rect 10466 1934 10468 1986
rect 10412 1932 10468 1934
rect 10732 1986 10788 1988
rect 10732 1934 10734 1986
rect 10734 1934 10786 1986
rect 10786 1934 10788 1986
rect 10732 1932 10788 1934
rect 11052 1986 11108 1988
rect 11052 1934 11054 1986
rect 11054 1934 11106 1986
rect 11106 1934 11108 1986
rect 11052 1932 11108 1934
rect 11372 1986 11428 1988
rect 11372 1934 11374 1986
rect 11374 1934 11426 1986
rect 11426 1934 11428 1986
rect 11372 1932 11428 1934
rect 11532 1986 11588 1988
rect 11532 1934 11534 1986
rect 11534 1934 11586 1986
rect 11586 1934 11588 1986
rect 11532 1932 11588 1934
rect 11852 1986 11908 1988
rect 11852 1934 11854 1986
rect 11854 1934 11906 1986
rect 11906 1934 11908 1986
rect 11852 1932 11908 1934
rect 12012 1986 12068 1988
rect 12012 1934 12014 1986
rect 12014 1934 12066 1986
rect 12066 1934 12068 1986
rect 12012 1932 12068 1934
rect 12332 1986 12388 1988
rect 12332 1934 12334 1986
rect 12334 1934 12386 1986
rect 12386 1934 12388 1986
rect 12332 1932 12388 1934
rect 12172 1772 12228 1828
rect 8492 1666 8548 1668
rect 8492 1614 8494 1666
rect 8494 1614 8546 1666
rect 8546 1614 8548 1666
rect 8492 1612 8548 1614
rect 8812 1666 8868 1668
rect 8812 1614 8814 1666
rect 8814 1614 8866 1666
rect 8866 1614 8868 1666
rect 8812 1612 8868 1614
rect 8972 1666 9028 1668
rect 8972 1614 8974 1666
rect 8974 1614 9026 1666
rect 9026 1614 9028 1666
rect 8972 1612 9028 1614
rect 9292 1666 9348 1668
rect 9292 1614 9294 1666
rect 9294 1614 9346 1666
rect 9346 1614 9348 1666
rect 9292 1612 9348 1614
rect 9452 1666 9508 1668
rect 9452 1614 9454 1666
rect 9454 1614 9506 1666
rect 9506 1614 9508 1666
rect 9452 1612 9508 1614
rect 9772 1666 9828 1668
rect 9772 1614 9774 1666
rect 9774 1614 9826 1666
rect 9826 1614 9828 1666
rect 9772 1612 9828 1614
rect 10092 1666 10148 1668
rect 10092 1614 10094 1666
rect 10094 1614 10146 1666
rect 10146 1614 10148 1666
rect 10092 1612 10148 1614
rect 10412 1666 10468 1668
rect 10412 1614 10414 1666
rect 10414 1614 10466 1666
rect 10466 1614 10468 1666
rect 10412 1612 10468 1614
rect 10732 1666 10788 1668
rect 10732 1614 10734 1666
rect 10734 1614 10786 1666
rect 10786 1614 10788 1666
rect 10732 1612 10788 1614
rect 11052 1666 11108 1668
rect 11052 1614 11054 1666
rect 11054 1614 11106 1666
rect 11106 1614 11108 1666
rect 11052 1612 11108 1614
rect 11372 1666 11428 1668
rect 11372 1614 11374 1666
rect 11374 1614 11426 1666
rect 11426 1614 11428 1666
rect 11372 1612 11428 1614
rect 11532 1666 11588 1668
rect 11532 1614 11534 1666
rect 11534 1614 11586 1666
rect 11586 1614 11588 1666
rect 11532 1612 11588 1614
rect 11852 1666 11908 1668
rect 11852 1614 11854 1666
rect 11854 1614 11906 1666
rect 11906 1614 11908 1666
rect 11852 1612 11908 1614
rect 12012 1666 12068 1668
rect 12012 1614 12014 1666
rect 12014 1614 12066 1666
rect 12066 1614 12068 1666
rect 12012 1612 12068 1614
rect 12332 1666 12388 1668
rect 12332 1614 12334 1666
rect 12334 1614 12386 1666
rect 12386 1614 12388 1666
rect 12332 1612 12388 1614
rect 8492 1506 8548 1508
rect 8492 1454 8494 1506
rect 8494 1454 8546 1506
rect 8546 1454 8548 1506
rect 8492 1452 8548 1454
rect 8812 1506 8868 1508
rect 8812 1454 8814 1506
rect 8814 1454 8866 1506
rect 8866 1454 8868 1506
rect 8812 1452 8868 1454
rect 8972 1506 9028 1508
rect 8972 1454 8974 1506
rect 8974 1454 9026 1506
rect 9026 1454 9028 1506
rect 8972 1452 9028 1454
rect 9292 1506 9348 1508
rect 9292 1454 9294 1506
rect 9294 1454 9346 1506
rect 9346 1454 9348 1506
rect 9292 1452 9348 1454
rect 9452 1506 9508 1508
rect 9452 1454 9454 1506
rect 9454 1454 9506 1506
rect 9506 1454 9508 1506
rect 9452 1452 9508 1454
rect 9772 1506 9828 1508
rect 9772 1454 9774 1506
rect 9774 1454 9826 1506
rect 9826 1454 9828 1506
rect 9772 1452 9828 1454
rect 10092 1506 10148 1508
rect 10092 1454 10094 1506
rect 10094 1454 10146 1506
rect 10146 1454 10148 1506
rect 10092 1452 10148 1454
rect 10412 1506 10468 1508
rect 10412 1454 10414 1506
rect 10414 1454 10466 1506
rect 10466 1454 10468 1506
rect 10412 1452 10468 1454
rect 10732 1506 10788 1508
rect 10732 1454 10734 1506
rect 10734 1454 10786 1506
rect 10786 1454 10788 1506
rect 10732 1452 10788 1454
rect 11052 1506 11108 1508
rect 11052 1454 11054 1506
rect 11054 1454 11106 1506
rect 11106 1454 11108 1506
rect 11052 1452 11108 1454
rect 11372 1506 11428 1508
rect 11372 1454 11374 1506
rect 11374 1454 11426 1506
rect 11426 1454 11428 1506
rect 11372 1452 11428 1454
rect 11532 1506 11588 1508
rect 11532 1454 11534 1506
rect 11534 1454 11586 1506
rect 11586 1454 11588 1506
rect 11532 1452 11588 1454
rect 11852 1506 11908 1508
rect 11852 1454 11854 1506
rect 11854 1454 11906 1506
rect 11906 1454 11908 1506
rect 11852 1452 11908 1454
rect 12012 1506 12068 1508
rect 12012 1454 12014 1506
rect 12014 1454 12066 1506
rect 12066 1454 12068 1506
rect 12012 1452 12068 1454
rect 12332 1506 12388 1508
rect 12332 1454 12334 1506
rect 12334 1454 12386 1506
rect 12386 1454 12388 1506
rect 12332 1452 12388 1454
rect 8492 1346 8548 1348
rect 8492 1294 8494 1346
rect 8494 1294 8546 1346
rect 8546 1294 8548 1346
rect 8492 1292 8548 1294
rect 8812 1346 8868 1348
rect 8812 1294 8814 1346
rect 8814 1294 8866 1346
rect 8866 1294 8868 1346
rect 8812 1292 8868 1294
rect 8972 1346 9028 1348
rect 8972 1294 8974 1346
rect 8974 1294 9026 1346
rect 9026 1294 9028 1346
rect 8972 1292 9028 1294
rect 9292 1346 9348 1348
rect 9292 1294 9294 1346
rect 9294 1294 9346 1346
rect 9346 1294 9348 1346
rect 9292 1292 9348 1294
rect 9452 1346 9508 1348
rect 9452 1294 9454 1346
rect 9454 1294 9506 1346
rect 9506 1294 9508 1346
rect 9452 1292 9508 1294
rect 9772 1346 9828 1348
rect 9772 1294 9774 1346
rect 9774 1294 9826 1346
rect 9826 1294 9828 1346
rect 9772 1292 9828 1294
rect 10092 1346 10148 1348
rect 10092 1294 10094 1346
rect 10094 1294 10146 1346
rect 10146 1294 10148 1346
rect 10092 1292 10148 1294
rect 10412 1346 10468 1348
rect 10412 1294 10414 1346
rect 10414 1294 10466 1346
rect 10466 1294 10468 1346
rect 10412 1292 10468 1294
rect 10732 1346 10788 1348
rect 10732 1294 10734 1346
rect 10734 1294 10786 1346
rect 10786 1294 10788 1346
rect 10732 1292 10788 1294
rect 11052 1346 11108 1348
rect 11052 1294 11054 1346
rect 11054 1294 11106 1346
rect 11106 1294 11108 1346
rect 11052 1292 11108 1294
rect 11372 1346 11428 1348
rect 11372 1294 11374 1346
rect 11374 1294 11426 1346
rect 11426 1294 11428 1346
rect 11372 1292 11428 1294
rect 11532 1346 11588 1348
rect 11532 1294 11534 1346
rect 11534 1294 11586 1346
rect 11586 1294 11588 1346
rect 11532 1292 11588 1294
rect 11852 1346 11908 1348
rect 11852 1294 11854 1346
rect 11854 1294 11906 1346
rect 11906 1294 11908 1346
rect 11852 1292 11908 1294
rect 12012 1346 12068 1348
rect 12012 1294 12014 1346
rect 12014 1294 12066 1346
rect 12066 1294 12068 1346
rect 12012 1292 12068 1294
rect 12332 1346 12388 1348
rect 12332 1294 12334 1346
rect 12334 1294 12386 1346
rect 12386 1294 12388 1346
rect 12332 1292 12388 1294
rect 8492 1186 8548 1188
rect 8492 1134 8494 1186
rect 8494 1134 8546 1186
rect 8546 1134 8548 1186
rect 8492 1132 8548 1134
rect 8812 1186 8868 1188
rect 8812 1134 8814 1186
rect 8814 1134 8866 1186
rect 8866 1134 8868 1186
rect 8812 1132 8868 1134
rect 8972 1186 9028 1188
rect 8972 1134 8974 1186
rect 8974 1134 9026 1186
rect 9026 1134 9028 1186
rect 8972 1132 9028 1134
rect 9292 1186 9348 1188
rect 9292 1134 9294 1186
rect 9294 1134 9346 1186
rect 9346 1134 9348 1186
rect 9292 1132 9348 1134
rect 9452 1186 9508 1188
rect 9452 1134 9454 1186
rect 9454 1134 9506 1186
rect 9506 1134 9508 1186
rect 9452 1132 9508 1134
rect 9772 1186 9828 1188
rect 9772 1134 9774 1186
rect 9774 1134 9826 1186
rect 9826 1134 9828 1186
rect 9772 1132 9828 1134
rect 10092 1186 10148 1188
rect 10092 1134 10094 1186
rect 10094 1134 10146 1186
rect 10146 1134 10148 1186
rect 10092 1132 10148 1134
rect 10412 1186 10468 1188
rect 10412 1134 10414 1186
rect 10414 1134 10466 1186
rect 10466 1134 10468 1186
rect 10412 1132 10468 1134
rect 10732 1186 10788 1188
rect 10732 1134 10734 1186
rect 10734 1134 10786 1186
rect 10786 1134 10788 1186
rect 10732 1132 10788 1134
rect 11052 1186 11108 1188
rect 11052 1134 11054 1186
rect 11054 1134 11106 1186
rect 11106 1134 11108 1186
rect 11052 1132 11108 1134
rect 11372 1186 11428 1188
rect 11372 1134 11374 1186
rect 11374 1134 11426 1186
rect 11426 1134 11428 1186
rect 11372 1132 11428 1134
rect 11532 1186 11588 1188
rect 11532 1134 11534 1186
rect 11534 1134 11586 1186
rect 11586 1134 11588 1186
rect 11532 1132 11588 1134
rect 11852 1186 11908 1188
rect 11852 1134 11854 1186
rect 11854 1134 11906 1186
rect 11906 1134 11908 1186
rect 11852 1132 11908 1134
rect 12012 1186 12068 1188
rect 12012 1134 12014 1186
rect 12014 1134 12066 1186
rect 12066 1134 12068 1186
rect 12012 1132 12068 1134
rect 12332 1186 12388 1188
rect 12332 1134 12334 1186
rect 12334 1134 12386 1186
rect 12386 1134 12388 1186
rect 12332 1132 12388 1134
rect 8492 1026 8548 1028
rect 8492 974 8494 1026
rect 8494 974 8546 1026
rect 8546 974 8548 1026
rect 8492 972 8548 974
rect 8812 1026 8868 1028
rect 8812 974 8814 1026
rect 8814 974 8866 1026
rect 8866 974 8868 1026
rect 8812 972 8868 974
rect 8972 1026 9028 1028
rect 8972 974 8974 1026
rect 8974 974 9026 1026
rect 9026 974 9028 1026
rect 8972 972 9028 974
rect 9292 1026 9348 1028
rect 9292 974 9294 1026
rect 9294 974 9346 1026
rect 9346 974 9348 1026
rect 9292 972 9348 974
rect 9452 1026 9508 1028
rect 9452 974 9454 1026
rect 9454 974 9506 1026
rect 9506 974 9508 1026
rect 9452 972 9508 974
rect 9772 1026 9828 1028
rect 9772 974 9774 1026
rect 9774 974 9826 1026
rect 9826 974 9828 1026
rect 9772 972 9828 974
rect 10092 1026 10148 1028
rect 10092 974 10094 1026
rect 10094 974 10146 1026
rect 10146 974 10148 1026
rect 10092 972 10148 974
rect 10412 1026 10468 1028
rect 10412 974 10414 1026
rect 10414 974 10466 1026
rect 10466 974 10468 1026
rect 10412 972 10468 974
rect 10732 1026 10788 1028
rect 10732 974 10734 1026
rect 10734 974 10786 1026
rect 10786 974 10788 1026
rect 10732 972 10788 974
rect 11052 1026 11108 1028
rect 11052 974 11054 1026
rect 11054 974 11106 1026
rect 11106 974 11108 1026
rect 11052 972 11108 974
rect 11372 1026 11428 1028
rect 11372 974 11374 1026
rect 11374 974 11426 1026
rect 11426 974 11428 1026
rect 11372 972 11428 974
rect 11532 1026 11588 1028
rect 11532 974 11534 1026
rect 11534 974 11586 1026
rect 11586 974 11588 1026
rect 11532 972 11588 974
rect 11852 1026 11908 1028
rect 11852 974 11854 1026
rect 11854 974 11906 1026
rect 11906 974 11908 1026
rect 11852 972 11908 974
rect 12012 1026 12068 1028
rect 12012 974 12014 1026
rect 12014 974 12066 1026
rect 12066 974 12068 1026
rect 12012 972 12068 974
rect 12332 1026 12388 1028
rect 12332 974 12334 1026
rect 12334 974 12386 1026
rect 12386 974 12388 1026
rect 12332 972 12388 974
rect 8652 732 8708 788
rect 8492 546 8548 548
rect 8492 494 8494 546
rect 8494 494 8546 546
rect 8546 494 8548 546
rect 8492 492 8548 494
rect 8812 546 8868 548
rect 8812 494 8814 546
rect 8814 494 8866 546
rect 8866 494 8868 546
rect 8812 492 8868 494
rect 8972 546 9028 548
rect 8972 494 8974 546
rect 8974 494 9026 546
rect 9026 494 9028 546
rect 8972 492 9028 494
rect 9292 546 9348 548
rect 9292 494 9294 546
rect 9294 494 9346 546
rect 9346 494 9348 546
rect 9292 492 9348 494
rect 9452 546 9508 548
rect 9452 494 9454 546
rect 9454 494 9506 546
rect 9506 494 9508 546
rect 9452 492 9508 494
rect 9772 546 9828 548
rect 9772 494 9774 546
rect 9774 494 9826 546
rect 9826 494 9828 546
rect 9772 492 9828 494
rect 10092 546 10148 548
rect 10092 494 10094 546
rect 10094 494 10146 546
rect 10146 494 10148 546
rect 10092 492 10148 494
rect 10412 546 10468 548
rect 10412 494 10414 546
rect 10414 494 10466 546
rect 10466 494 10468 546
rect 10412 492 10468 494
rect 10732 546 10788 548
rect 10732 494 10734 546
rect 10734 494 10786 546
rect 10786 494 10788 546
rect 10732 492 10788 494
rect 11052 546 11108 548
rect 11052 494 11054 546
rect 11054 494 11106 546
rect 11106 494 11108 546
rect 11052 492 11108 494
rect 11372 546 11428 548
rect 11372 494 11374 546
rect 11374 494 11426 546
rect 11426 494 11428 546
rect 11372 492 11428 494
rect 11532 546 11588 548
rect 11532 494 11534 546
rect 11534 494 11586 546
rect 11586 494 11588 546
rect 11532 492 11588 494
rect 11852 546 11908 548
rect 11852 494 11854 546
rect 11854 494 11906 546
rect 11906 494 11908 546
rect 11852 492 11908 494
rect 12012 546 12068 548
rect 12012 494 12014 546
rect 12014 494 12066 546
rect 12066 494 12068 546
rect 12012 492 12068 494
rect 12332 546 12388 548
rect 12332 494 12334 546
rect 12334 494 12386 546
rect 12386 494 12388 546
rect 12332 492 12388 494
rect 8492 386 8548 388
rect 8492 334 8494 386
rect 8494 334 8546 386
rect 8546 334 8548 386
rect 8492 332 8548 334
rect 8812 386 8868 388
rect 8812 334 8814 386
rect 8814 334 8866 386
rect 8866 334 8868 386
rect 8812 332 8868 334
rect 8972 386 9028 388
rect 8972 334 8974 386
rect 8974 334 9026 386
rect 9026 334 9028 386
rect 8972 332 9028 334
rect 9292 386 9348 388
rect 9292 334 9294 386
rect 9294 334 9346 386
rect 9346 334 9348 386
rect 9292 332 9348 334
rect 9452 386 9508 388
rect 9452 334 9454 386
rect 9454 334 9506 386
rect 9506 334 9508 386
rect 9452 332 9508 334
rect 9772 386 9828 388
rect 9772 334 9774 386
rect 9774 334 9826 386
rect 9826 334 9828 386
rect 9772 332 9828 334
rect 10092 386 10148 388
rect 10092 334 10094 386
rect 10094 334 10146 386
rect 10146 334 10148 386
rect 10092 332 10148 334
rect 10412 386 10468 388
rect 10412 334 10414 386
rect 10414 334 10466 386
rect 10466 334 10468 386
rect 10412 332 10468 334
rect 10732 386 10788 388
rect 10732 334 10734 386
rect 10734 334 10786 386
rect 10786 334 10788 386
rect 10732 332 10788 334
rect 11052 386 11108 388
rect 11052 334 11054 386
rect 11054 334 11106 386
rect 11106 334 11108 386
rect 11052 332 11108 334
rect 11372 386 11428 388
rect 11372 334 11374 386
rect 11374 334 11426 386
rect 11426 334 11428 386
rect 11372 332 11428 334
rect 11532 386 11588 388
rect 11532 334 11534 386
rect 11534 334 11586 386
rect 11586 334 11588 386
rect 11532 332 11588 334
rect 11852 386 11908 388
rect 11852 334 11854 386
rect 11854 334 11906 386
rect 11906 334 11908 386
rect 11852 332 11908 334
rect 12012 386 12068 388
rect 12012 334 12014 386
rect 12014 334 12066 386
rect 12066 334 12068 386
rect 12012 332 12068 334
rect 12332 386 12388 388
rect 12332 334 12334 386
rect 12334 334 12386 386
rect 12386 334 12388 386
rect 12332 332 12388 334
rect 8492 226 8548 228
rect 8492 174 8494 226
rect 8494 174 8546 226
rect 8546 174 8548 226
rect 8492 172 8548 174
rect 8812 226 8868 228
rect 8812 174 8814 226
rect 8814 174 8866 226
rect 8866 174 8868 226
rect 8812 172 8868 174
rect 8972 226 9028 228
rect 8972 174 8974 226
rect 8974 174 9026 226
rect 9026 174 9028 226
rect 8972 172 9028 174
rect 9292 226 9348 228
rect 9292 174 9294 226
rect 9294 174 9346 226
rect 9346 174 9348 226
rect 9292 172 9348 174
rect 9452 226 9508 228
rect 9452 174 9454 226
rect 9454 174 9506 226
rect 9506 174 9508 226
rect 9452 172 9508 174
rect 9772 226 9828 228
rect 9772 174 9774 226
rect 9774 174 9826 226
rect 9826 174 9828 226
rect 9772 172 9828 174
rect 10092 226 10148 228
rect 10092 174 10094 226
rect 10094 174 10146 226
rect 10146 174 10148 226
rect 10092 172 10148 174
rect 10412 226 10468 228
rect 10412 174 10414 226
rect 10414 174 10466 226
rect 10466 174 10468 226
rect 10412 172 10468 174
rect 10732 226 10788 228
rect 10732 174 10734 226
rect 10734 174 10786 226
rect 10786 174 10788 226
rect 10732 172 10788 174
rect 11052 226 11108 228
rect 11052 174 11054 226
rect 11054 174 11106 226
rect 11106 174 11108 226
rect 11052 172 11108 174
rect 11372 226 11428 228
rect 11372 174 11374 226
rect 11374 174 11426 226
rect 11426 174 11428 226
rect 11372 172 11428 174
rect 11532 226 11588 228
rect 11532 174 11534 226
rect 11534 174 11586 226
rect 11586 174 11588 226
rect 11532 172 11588 174
rect 11852 226 11908 228
rect 11852 174 11854 226
rect 11854 174 11906 226
rect 11906 174 11908 226
rect 11852 172 11908 174
rect 12012 226 12068 228
rect 12012 174 12014 226
rect 12014 174 12066 226
rect 12066 174 12068 226
rect 12012 172 12068 174
rect 12332 226 12388 228
rect 12332 174 12334 226
rect 12334 174 12386 226
rect 12386 174 12388 226
rect 12332 172 12388 174
rect 8492 66 8548 68
rect 8492 14 8494 66
rect 8494 14 8546 66
rect 8546 14 8548 66
rect 8492 12 8548 14
rect 8812 66 8868 68
rect 8812 14 8814 66
rect 8814 14 8866 66
rect 8866 14 8868 66
rect 8812 12 8868 14
rect 8972 66 9028 68
rect 8972 14 8974 66
rect 8974 14 9026 66
rect 9026 14 9028 66
rect 8972 12 9028 14
rect 9292 66 9348 68
rect 9292 14 9294 66
rect 9294 14 9346 66
rect 9346 14 9348 66
rect 9292 12 9348 14
rect 9452 66 9508 68
rect 9452 14 9454 66
rect 9454 14 9506 66
rect 9506 14 9508 66
rect 9452 12 9508 14
rect 9772 66 9828 68
rect 9772 14 9774 66
rect 9774 14 9826 66
rect 9826 14 9828 66
rect 9772 12 9828 14
rect 10092 66 10148 68
rect 10092 14 10094 66
rect 10094 14 10146 66
rect 10146 14 10148 66
rect 10092 12 10148 14
rect 10412 66 10468 68
rect 10412 14 10414 66
rect 10414 14 10466 66
rect 10466 14 10468 66
rect 10412 12 10468 14
rect 10732 66 10788 68
rect 10732 14 10734 66
rect 10734 14 10786 66
rect 10786 14 10788 66
rect 10732 12 10788 14
rect 11052 66 11108 68
rect 11052 14 11054 66
rect 11054 14 11106 66
rect 11106 14 11108 66
rect 11052 12 11108 14
rect 11372 66 11428 68
rect 11372 14 11374 66
rect 11374 14 11426 66
rect 11426 14 11428 66
rect 11372 12 11428 14
rect 11532 66 11588 68
rect 11532 14 11534 66
rect 11534 14 11586 66
rect 11586 14 11588 66
rect 11532 12 11588 14
rect 11852 66 11908 68
rect 11852 14 11854 66
rect 11854 14 11906 66
rect 11906 14 11908 66
rect 11852 12 11908 14
rect 12012 66 12068 68
rect 12012 14 12014 66
rect 12014 14 12066 66
rect 12066 14 12068 66
rect 12012 12 12068 14
rect 12332 66 12388 68
rect 12332 14 12334 66
rect 12334 14 12386 66
rect 12386 14 12388 66
rect 12332 12 12388 14
<< metal3 >>
rect 8480 31432 8560 31520
rect 8480 31368 8488 31432
rect 8552 31368 8560 31432
rect 8480 31272 8560 31368
rect 8480 31208 8488 31272
rect 8552 31208 8560 31272
rect 8480 31112 8560 31208
rect 8480 31048 8488 31112
rect 8552 31048 8560 31112
rect 8480 30952 8560 31048
rect 8480 30888 8488 30952
rect 8552 30888 8560 30952
rect 8480 30792 8560 30888
rect 8480 30728 8488 30792
rect 8552 30728 8560 30792
rect 8480 30632 8560 30728
rect 8480 30568 8488 30632
rect 8552 30568 8560 30632
rect 8480 30472 8560 30568
rect 8480 30408 8488 30472
rect 8552 30408 8560 30472
rect 8480 30312 8560 30408
rect 8480 30248 8488 30312
rect 8552 30248 8560 30312
rect 8480 30152 8560 30248
rect 8480 30088 8488 30152
rect 8552 30088 8560 30152
rect 8480 29992 8560 30088
rect 8480 29928 8488 29992
rect 8552 29928 8560 29992
rect 8480 29832 8560 29928
rect 8480 29768 8488 29832
rect 8552 29768 8560 29832
rect 8480 29672 8560 29768
rect 8480 29608 8488 29672
rect 8552 29608 8560 29672
rect 8480 29512 8560 29608
rect 8480 29448 8488 29512
rect 8552 29448 8560 29512
rect 8480 29352 8560 29448
rect 8480 29288 8488 29352
rect 8552 29288 8560 29352
rect 8480 29192 8560 29288
rect 8480 29128 8488 29192
rect 8552 29128 8560 29192
rect 8480 29032 8560 29128
rect 8480 28968 8488 29032
rect 8552 28968 8560 29032
rect 8480 28872 8560 28968
rect 8480 28808 8488 28872
rect 8552 28808 8560 28872
rect 8480 28712 8560 28808
rect 8480 28648 8488 28712
rect 8552 28648 8560 28712
rect 8480 28552 8560 28648
rect 8480 28488 8488 28552
rect 8552 28488 8560 28552
rect 8480 28392 8560 28488
rect 8480 28328 8488 28392
rect 8552 28328 8560 28392
rect 8480 28232 8560 28328
rect 8480 28168 8488 28232
rect 8552 28168 8560 28232
rect 8480 28072 8560 28168
rect 8480 28008 8488 28072
rect 8552 28008 8560 28072
rect 8480 27912 8560 28008
rect 8480 27848 8488 27912
rect 8552 27848 8560 27912
rect 8480 27752 8560 27848
rect 8480 27688 8488 27752
rect 8552 27688 8560 27752
rect 8480 27592 8560 27688
rect 8480 27528 8488 27592
rect 8552 27528 8560 27592
rect 8480 27432 8560 27528
rect 8480 27368 8488 27432
rect 8552 27368 8560 27432
rect 8480 27272 8560 27368
rect 8480 27208 8488 27272
rect 8552 27208 8560 27272
rect 8480 27112 8560 27208
rect 8480 27048 8488 27112
rect 8552 27048 8560 27112
rect 8480 26952 8560 27048
rect 8480 26888 8488 26952
rect 8552 26888 8560 26952
rect 8480 26792 8560 26888
rect 8480 26728 8488 26792
rect 8552 26728 8560 26792
rect 8480 26632 8560 26728
rect 8480 26568 8488 26632
rect 8552 26568 8560 26632
rect 8480 26472 8560 26568
rect 8480 26408 8488 26472
rect 8552 26408 8560 26472
rect 8480 26312 8560 26408
rect 8480 26248 8488 26312
rect 8552 26248 8560 26312
rect 8480 26152 8560 26248
rect 8480 26088 8488 26152
rect 8552 26088 8560 26152
rect 8480 25992 8560 26088
rect 8480 25928 8488 25992
rect 8552 25928 8560 25992
rect 8480 25832 8560 25928
rect 8480 25768 8488 25832
rect 8552 25768 8560 25832
rect 8480 25672 8560 25768
rect 8480 25608 8488 25672
rect 8552 25608 8560 25672
rect 8480 25512 8560 25608
rect 8480 25448 8488 25512
rect 8552 25448 8560 25512
rect 8480 25352 8560 25448
rect 8480 25288 8488 25352
rect 8552 25288 8560 25352
rect 8480 25192 8560 25288
rect 8480 25128 8488 25192
rect 8552 25128 8560 25192
rect 8480 25032 8560 25128
rect 8480 24968 8488 25032
rect 8552 24968 8560 25032
rect 8480 24872 8560 24968
rect 8480 24808 8488 24872
rect 8552 24808 8560 24872
rect 8480 24712 8560 24808
rect 8480 24648 8488 24712
rect 8552 24648 8560 24712
rect 8480 24552 8560 24648
rect 8480 24488 8488 24552
rect 8552 24488 8560 24552
rect 8480 24392 8560 24488
rect 8480 24328 8488 24392
rect 8552 24328 8560 24392
rect 8480 24232 8560 24328
rect 8480 24168 8488 24232
rect 8552 24168 8560 24232
rect 8480 24072 8560 24168
rect 8480 24008 8488 24072
rect 8552 24008 8560 24072
rect 8480 23912 8560 24008
rect 8480 23848 8488 23912
rect 8552 23848 8560 23912
rect 8480 23752 8560 23848
rect 8480 23688 8488 23752
rect 8552 23688 8560 23752
rect 8480 23592 8560 23688
rect 8480 23528 8488 23592
rect 8552 23528 8560 23592
rect 8480 23432 8560 23528
rect 8480 23368 8488 23432
rect 8552 23368 8560 23432
rect 8480 23272 8560 23368
rect 8480 23208 8488 23272
rect 8552 23208 8560 23272
rect 8480 23112 8560 23208
rect 8480 23048 8488 23112
rect 8552 23048 8560 23112
rect 8480 22952 8560 23048
rect 8480 22888 8488 22952
rect 8552 22888 8560 22952
rect 8480 22792 8560 22888
rect 8480 22728 8488 22792
rect 8552 22728 8560 22792
rect 8480 22632 8560 22728
rect 8480 22568 8488 22632
rect 8552 22568 8560 22632
rect 8480 22472 8560 22568
rect 8480 22408 8488 22472
rect 8552 22408 8560 22472
rect 8480 22312 8560 22408
rect 8480 22248 8488 22312
rect 8552 22248 8560 22312
rect 8480 22152 8560 22248
rect 8480 22088 8488 22152
rect 8552 22088 8560 22152
rect 8480 21992 8560 22088
rect 8480 21928 8488 21992
rect 8552 21928 8560 21992
rect 8480 21832 8560 21928
rect 8480 21768 8488 21832
rect 8552 21768 8560 21832
rect 8480 21672 8560 21768
rect 8480 21608 8488 21672
rect 8552 21608 8560 21672
rect 8480 21512 8560 21608
rect 8480 21448 8488 21512
rect 8552 21448 8560 21512
rect 8480 21352 8560 21448
rect 8480 21288 8488 21352
rect 8552 21288 8560 21352
rect 8480 21192 8560 21288
rect 8480 21128 8488 21192
rect 8552 21128 8560 21192
rect 8480 21032 8560 21128
rect 8480 20968 8488 21032
rect 8552 20968 8560 21032
rect 8480 20872 8560 20968
rect 8480 20808 8488 20872
rect 8552 20808 8560 20872
rect 8480 20712 8560 20808
rect 8480 20648 8488 20712
rect 8552 20648 8560 20712
rect 8480 20552 8560 20648
rect 8480 20488 8488 20552
rect 8552 20488 8560 20552
rect 8480 20392 8560 20488
rect 8480 20328 8488 20392
rect 8552 20328 8560 20392
rect 8480 20232 8560 20328
rect 8480 20168 8488 20232
rect 8552 20168 8560 20232
rect 8480 20072 8560 20168
rect 8480 20008 8488 20072
rect 8552 20008 8560 20072
rect 8480 19912 8560 20008
rect 8480 19848 8488 19912
rect 8552 19848 8560 19912
rect 8480 19752 8560 19848
rect 8480 19688 8488 19752
rect 8552 19688 8560 19752
rect 8480 19592 8560 19688
rect 8480 19528 8488 19592
rect 8552 19528 8560 19592
rect 8480 19432 8560 19528
rect 8480 19368 8488 19432
rect 8552 19368 8560 19432
rect 8480 19272 8560 19368
rect 8480 19208 8488 19272
rect 8552 19208 8560 19272
rect 8480 19112 8560 19208
rect 8480 19048 8488 19112
rect 8552 19048 8560 19112
rect 8480 18952 8560 19048
rect 8480 18888 8488 18952
rect 8552 18888 8560 18952
rect 8480 18792 8560 18888
rect 8480 18728 8488 18792
rect 8552 18728 8560 18792
rect 8480 18632 8560 18728
rect 8480 18568 8488 18632
rect 8552 18568 8560 18632
rect 8480 18472 8560 18568
rect 8480 18408 8488 18472
rect 8552 18408 8560 18472
rect 8480 18312 8560 18408
rect 8480 18248 8488 18312
rect 8552 18248 8560 18312
rect 8480 18152 8560 18248
rect 8480 18088 8488 18152
rect 8552 18088 8560 18152
rect 8480 17992 8560 18088
rect 8480 17928 8488 17992
rect 8552 17928 8560 17992
rect 8480 17832 8560 17928
rect 8480 17768 8488 17832
rect 8552 17768 8560 17832
rect 8480 17672 8560 17768
rect 8480 17608 8488 17672
rect 8552 17608 8560 17672
rect 8480 17512 8560 17608
rect 8480 17448 8488 17512
rect 8552 17448 8560 17512
rect 8480 17352 8560 17448
rect 8480 17288 8488 17352
rect 8552 17288 8560 17352
rect 8480 17192 8560 17288
rect 8480 17128 8488 17192
rect 8552 17128 8560 17192
rect 8480 17032 8560 17128
rect 8480 16968 8488 17032
rect 8552 16968 8560 17032
rect 8480 16872 8560 16968
rect 8480 16808 8488 16872
rect 8552 16808 8560 16872
rect 8480 16712 8560 16808
rect 8480 16648 8488 16712
rect 8552 16648 8560 16712
rect 8480 16552 8560 16648
rect 8480 16488 8488 16552
rect 8552 16488 8560 16552
rect 8480 16392 8560 16488
rect 8480 16328 8488 16392
rect 8552 16328 8560 16392
rect 8480 16232 8560 16328
rect 8480 16168 8488 16232
rect 8552 16168 8560 16232
rect 8480 16072 8560 16168
rect 8480 16008 8488 16072
rect 8552 16008 8560 16072
rect 8480 15912 8560 16008
rect 8480 15848 8488 15912
rect 8552 15848 8560 15912
rect 8480 15752 8560 15848
rect 8480 15688 8488 15752
rect 8552 15688 8560 15752
rect 8480 15592 8560 15688
rect 8480 15528 8488 15592
rect 8552 15528 8560 15592
rect 8480 15432 8560 15528
rect 8480 15368 8488 15432
rect 8552 15368 8560 15432
rect 8480 15272 8560 15368
rect 8480 15208 8488 15272
rect 8552 15208 8560 15272
rect 8480 15112 8560 15208
rect 8480 15048 8488 15112
rect 8552 15048 8560 15112
rect 8480 14952 8560 15048
rect 8480 14888 8488 14952
rect 8552 14888 8560 14952
rect 8480 14792 8560 14888
rect 8480 14728 8488 14792
rect 8552 14728 8560 14792
rect 8480 14632 8560 14728
rect 8480 14568 8488 14632
rect 8552 14568 8560 14632
rect 8480 14472 8560 14568
rect 8480 14408 8488 14472
rect 8552 14408 8560 14472
rect 8480 14312 8560 14408
rect 8480 14248 8488 14312
rect 8552 14248 8560 14312
rect 8480 14152 8560 14248
rect 8480 14088 8488 14152
rect 8552 14088 8560 14152
rect 8480 13992 8560 14088
rect 8480 13928 8488 13992
rect 8552 13928 8560 13992
rect 8480 13832 8560 13928
rect 8480 13768 8488 13832
rect 8552 13768 8560 13832
rect 8480 13672 8560 13768
rect 8480 13608 8488 13672
rect 8552 13608 8560 13672
rect 8480 13512 8560 13608
rect 8480 13448 8488 13512
rect 8552 13448 8560 13512
rect 8480 13352 8560 13448
rect 8480 13288 8488 13352
rect 8552 13288 8560 13352
rect 8480 13192 8560 13288
rect 8480 13128 8488 13192
rect 8552 13128 8560 13192
rect 8480 13032 8560 13128
rect 8480 12968 8488 13032
rect 8552 12968 8560 13032
rect 8480 12872 8560 12968
rect 8480 12808 8488 12872
rect 8552 12808 8560 12872
rect 8480 12712 8560 12808
rect 8480 12648 8488 12712
rect 8552 12648 8560 12712
rect 8480 12552 8560 12648
rect 8480 12488 8488 12552
rect 8552 12488 8560 12552
rect 8480 12392 8560 12488
rect 8480 12328 8488 12392
rect 8552 12328 8560 12392
rect 8480 12232 8560 12328
rect 8480 12168 8488 12232
rect 8552 12168 8560 12232
rect 8480 12072 8560 12168
rect 8480 12008 8488 12072
rect 8552 12008 8560 12072
rect 8480 11912 8560 12008
rect 8480 11848 8488 11912
rect 8552 11848 8560 11912
rect 8480 11752 8560 11848
rect 8480 11688 8488 11752
rect 8552 11688 8560 11752
rect 8480 11592 8560 11688
rect 8480 11528 8488 11592
rect 8552 11528 8560 11592
rect 8480 11432 8560 11528
rect 8480 11368 8488 11432
rect 8552 11368 8560 11432
rect 8480 11272 8560 11368
rect 8480 11208 8488 11272
rect 8552 11208 8560 11272
rect 8480 11112 8560 11208
rect 8480 11048 8488 11112
rect 8552 11048 8560 11112
rect 8480 10952 8560 11048
rect 8480 10888 8488 10952
rect 8552 10888 8560 10952
rect 8480 10792 8560 10888
rect 8480 10728 8488 10792
rect 8552 10728 8560 10792
rect 8480 10632 8560 10728
rect 8480 10568 8488 10632
rect 8552 10568 8560 10632
rect 8480 10472 8560 10568
rect 8480 10408 8488 10472
rect 8552 10408 8560 10472
rect 8480 10312 8560 10408
rect 8480 10248 8488 10312
rect 8552 10248 8560 10312
rect 8480 10152 8560 10248
rect 8480 10088 8488 10152
rect 8552 10088 8560 10152
rect 8480 9992 8560 10088
rect 8480 9928 8488 9992
rect 8552 9928 8560 9992
rect 8480 9832 8560 9928
rect 8480 9768 8488 9832
rect 8552 9768 8560 9832
rect 8480 9672 8560 9768
rect 8480 9608 8488 9672
rect 8552 9608 8560 9672
rect 8480 9512 8560 9608
rect 8480 9448 8488 9512
rect 8552 9448 8560 9512
rect 8480 9352 8560 9448
rect 8480 9288 8488 9352
rect 8552 9288 8560 9352
rect 8480 9192 8560 9288
rect 8480 9128 8488 9192
rect 8552 9128 8560 9192
rect 8480 9032 8560 9128
rect 8480 8968 8488 9032
rect 8552 8968 8560 9032
rect 8480 8872 8560 8968
rect 8480 8808 8488 8872
rect 8552 8808 8560 8872
rect 8480 8712 8560 8808
rect 8480 8648 8488 8712
rect 8552 8648 8560 8712
rect 8480 8552 8560 8648
rect 8480 8488 8488 8552
rect 8552 8488 8560 8552
rect 8480 8392 8560 8488
rect 8480 8328 8488 8392
rect 8552 8328 8560 8392
rect 8480 8232 8560 8328
rect 8480 8168 8488 8232
rect 8552 8168 8560 8232
rect 8480 8072 8560 8168
rect 8480 8008 8488 8072
rect 8552 8008 8560 8072
rect 8480 7912 8560 8008
rect 8480 7848 8488 7912
rect 8552 7848 8560 7912
rect 8480 7752 8560 7848
rect 8480 7688 8488 7752
rect 8552 7688 8560 7752
rect 8480 7592 8560 7688
rect 8480 7528 8488 7592
rect 8552 7528 8560 7592
rect 8480 7432 8560 7528
rect 8480 7368 8488 7432
rect 8552 7368 8560 7432
rect 8480 7272 8560 7368
rect 8480 7208 8488 7272
rect 8552 7208 8560 7272
rect 8480 7112 8560 7208
rect 8480 7048 8488 7112
rect 8552 7048 8560 7112
rect 8480 6952 8560 7048
rect 8480 6888 8488 6952
rect 8552 6888 8560 6952
rect 8480 6792 8560 6888
rect 8480 6728 8488 6792
rect 8552 6728 8560 6792
rect 8480 6632 8560 6728
rect 8480 6568 8488 6632
rect 8552 6568 8560 6632
rect 8480 6472 8560 6568
rect 8480 6408 8488 6472
rect 8552 6408 8560 6472
rect 8480 6312 8560 6408
rect 8480 6248 8488 6312
rect 8552 6248 8560 6312
rect 8480 6152 8560 6248
rect 8480 6088 8488 6152
rect 8552 6088 8560 6152
rect 8480 5992 8560 6088
rect 8480 5928 8488 5992
rect 8552 5928 8560 5992
rect 8480 5832 8560 5928
rect 8480 5768 8488 5832
rect 8552 5768 8560 5832
rect 8480 5672 8560 5768
rect 8480 5608 8488 5672
rect 8552 5608 8560 5672
rect 8480 5512 8560 5608
rect 8480 5448 8488 5512
rect 8552 5448 8560 5512
rect 8480 5352 8560 5448
rect 8480 5288 8488 5352
rect 8552 5288 8560 5352
rect 8480 5192 8560 5288
rect 8480 5128 8488 5192
rect 8552 5128 8560 5192
rect 8480 5032 8560 5128
rect 8480 4968 8488 5032
rect 8552 4968 8560 5032
rect 8480 4872 8560 4968
rect 8480 4808 8488 4872
rect 8552 4808 8560 4872
rect 8480 4712 8560 4808
rect 8480 4648 8488 4712
rect 8552 4648 8560 4712
rect 8480 4552 8560 4648
rect 8480 4488 8488 4552
rect 8552 4488 8560 4552
rect 8480 4392 8560 4488
rect 8480 4328 8488 4392
rect 8552 4328 8560 4392
rect 8480 4232 8560 4328
rect 8480 4168 8488 4232
rect 8552 4168 8560 4232
rect 8480 4072 8560 4168
rect 8480 4008 8488 4072
rect 8552 4008 8560 4072
rect 8480 3912 8560 4008
rect 8480 3848 8488 3912
rect 8552 3848 8560 3912
rect 8480 3752 8560 3848
rect 8480 3688 8488 3752
rect 8552 3688 8560 3752
rect 8480 3592 8560 3688
rect 8480 3528 8488 3592
rect 8552 3528 8560 3592
rect 8480 3432 8560 3528
rect 8480 3368 8488 3432
rect 8552 3368 8560 3432
rect 8480 3272 8560 3368
rect 8480 3208 8488 3272
rect 8552 3208 8560 3272
rect 8480 3112 8560 3208
rect 8480 3048 8488 3112
rect 8552 3048 8560 3112
rect 8480 2952 8560 3048
rect 8480 2888 8488 2952
rect 8552 2888 8560 2952
rect 8480 2792 8560 2888
rect 8480 2728 8488 2792
rect 8552 2728 8560 2792
rect 8480 2632 8560 2728
rect 8480 2568 8488 2632
rect 8552 2568 8560 2632
rect 8480 2472 8560 2568
rect 8480 2408 8488 2472
rect 8552 2408 8560 2472
rect 8480 2312 8560 2408
rect 8480 2248 8488 2312
rect 8552 2248 8560 2312
rect 8480 2152 8560 2248
rect 8480 2088 8488 2152
rect 8552 2088 8560 2152
rect 8480 1992 8560 2088
rect 8480 1928 8488 1992
rect 8552 1928 8560 1992
rect 8480 1832 8560 1928
rect 8480 1768 8488 1832
rect 8552 1768 8560 1832
rect 8480 1672 8560 1768
rect 8480 1608 8488 1672
rect 8552 1608 8560 1672
rect 8480 1512 8560 1608
rect 8480 1448 8488 1512
rect 8552 1448 8560 1512
rect 8480 1352 8560 1448
rect 8480 1288 8488 1352
rect 8552 1288 8560 1352
rect 8480 1192 8560 1288
rect 8480 1128 8488 1192
rect 8552 1128 8560 1192
rect 8480 1032 8560 1128
rect 8480 968 8488 1032
rect 8552 968 8560 1032
rect 8480 872 8560 968
rect 8480 808 8488 872
rect 8552 808 8560 872
rect 8480 712 8560 808
rect 8480 648 8488 712
rect 8552 648 8560 712
rect 8480 552 8560 648
rect 8480 488 8488 552
rect 8552 488 8560 552
rect 8480 392 8560 488
rect 8480 328 8488 392
rect 8552 328 8560 392
rect 8480 232 8560 328
rect 8480 168 8488 232
rect 8552 168 8560 232
rect 8480 72 8560 168
rect 8480 8 8488 72
rect 8552 8 8560 72
rect 8480 -1528 8560 8
rect 8640 7588 8720 31520
rect 8640 7532 8652 7588
rect 8708 7532 8720 7588
rect 8640 788 8720 7532
rect 8640 732 8652 788
rect 8708 732 8720 788
rect 8640 0 8720 732
rect 8800 31432 8880 31520
rect 8800 31368 8808 31432
rect 8872 31368 8880 31432
rect 8800 31272 8880 31368
rect 8800 31208 8808 31272
rect 8872 31208 8880 31272
rect 8800 31112 8880 31208
rect 8800 31048 8808 31112
rect 8872 31048 8880 31112
rect 8800 30952 8880 31048
rect 8800 30888 8808 30952
rect 8872 30888 8880 30952
rect 8800 30792 8880 30888
rect 8800 30728 8808 30792
rect 8872 30728 8880 30792
rect 8800 30632 8880 30728
rect 8800 30568 8808 30632
rect 8872 30568 8880 30632
rect 8800 30472 8880 30568
rect 8800 30408 8808 30472
rect 8872 30408 8880 30472
rect 8800 30312 8880 30408
rect 8800 30248 8808 30312
rect 8872 30248 8880 30312
rect 8800 30152 8880 30248
rect 8800 30088 8808 30152
rect 8872 30088 8880 30152
rect 8800 29992 8880 30088
rect 8800 29928 8808 29992
rect 8872 29928 8880 29992
rect 8800 29832 8880 29928
rect 8800 29768 8808 29832
rect 8872 29768 8880 29832
rect 8800 29672 8880 29768
rect 8800 29608 8808 29672
rect 8872 29608 8880 29672
rect 8800 29512 8880 29608
rect 8800 29448 8808 29512
rect 8872 29448 8880 29512
rect 8800 29352 8880 29448
rect 8800 29288 8808 29352
rect 8872 29288 8880 29352
rect 8800 29192 8880 29288
rect 8800 29128 8808 29192
rect 8872 29128 8880 29192
rect 8800 29032 8880 29128
rect 8800 28968 8808 29032
rect 8872 28968 8880 29032
rect 8800 28872 8880 28968
rect 8800 28808 8808 28872
rect 8872 28808 8880 28872
rect 8800 28712 8880 28808
rect 8800 28648 8808 28712
rect 8872 28648 8880 28712
rect 8800 28552 8880 28648
rect 8800 28488 8808 28552
rect 8872 28488 8880 28552
rect 8800 28392 8880 28488
rect 8800 28328 8808 28392
rect 8872 28328 8880 28392
rect 8800 28232 8880 28328
rect 8800 28168 8808 28232
rect 8872 28168 8880 28232
rect 8800 28072 8880 28168
rect 8800 28008 8808 28072
rect 8872 28008 8880 28072
rect 8800 27912 8880 28008
rect 8800 27848 8808 27912
rect 8872 27848 8880 27912
rect 8800 27752 8880 27848
rect 8800 27688 8808 27752
rect 8872 27688 8880 27752
rect 8800 27592 8880 27688
rect 8800 27528 8808 27592
rect 8872 27528 8880 27592
rect 8800 27432 8880 27528
rect 8800 27368 8808 27432
rect 8872 27368 8880 27432
rect 8800 27272 8880 27368
rect 8800 27208 8808 27272
rect 8872 27208 8880 27272
rect 8800 27112 8880 27208
rect 8800 27048 8808 27112
rect 8872 27048 8880 27112
rect 8800 26952 8880 27048
rect 8800 26888 8808 26952
rect 8872 26888 8880 26952
rect 8800 26792 8880 26888
rect 8800 26728 8808 26792
rect 8872 26728 8880 26792
rect 8800 26632 8880 26728
rect 8800 26568 8808 26632
rect 8872 26568 8880 26632
rect 8800 26472 8880 26568
rect 8800 26408 8808 26472
rect 8872 26408 8880 26472
rect 8800 26312 8880 26408
rect 8800 26248 8808 26312
rect 8872 26248 8880 26312
rect 8800 26152 8880 26248
rect 8800 26088 8808 26152
rect 8872 26088 8880 26152
rect 8800 25992 8880 26088
rect 8800 25928 8808 25992
rect 8872 25928 8880 25992
rect 8800 25832 8880 25928
rect 8800 25768 8808 25832
rect 8872 25768 8880 25832
rect 8800 25672 8880 25768
rect 8800 25608 8808 25672
rect 8872 25608 8880 25672
rect 8800 25512 8880 25608
rect 8800 25448 8808 25512
rect 8872 25448 8880 25512
rect 8800 25352 8880 25448
rect 8800 25288 8808 25352
rect 8872 25288 8880 25352
rect 8800 25192 8880 25288
rect 8800 25128 8808 25192
rect 8872 25128 8880 25192
rect 8800 25032 8880 25128
rect 8800 24968 8808 25032
rect 8872 24968 8880 25032
rect 8800 24872 8880 24968
rect 8800 24808 8808 24872
rect 8872 24808 8880 24872
rect 8800 24712 8880 24808
rect 8800 24648 8808 24712
rect 8872 24648 8880 24712
rect 8800 24552 8880 24648
rect 8800 24488 8808 24552
rect 8872 24488 8880 24552
rect 8800 24392 8880 24488
rect 8800 24328 8808 24392
rect 8872 24328 8880 24392
rect 8800 24232 8880 24328
rect 8800 24168 8808 24232
rect 8872 24168 8880 24232
rect 8800 24072 8880 24168
rect 8800 24008 8808 24072
rect 8872 24008 8880 24072
rect 8800 23912 8880 24008
rect 8800 23848 8808 23912
rect 8872 23848 8880 23912
rect 8800 23752 8880 23848
rect 8800 23688 8808 23752
rect 8872 23688 8880 23752
rect 8800 23592 8880 23688
rect 8800 23528 8808 23592
rect 8872 23528 8880 23592
rect 8800 23432 8880 23528
rect 8800 23368 8808 23432
rect 8872 23368 8880 23432
rect 8800 23272 8880 23368
rect 8800 23208 8808 23272
rect 8872 23208 8880 23272
rect 8800 23112 8880 23208
rect 8800 23048 8808 23112
rect 8872 23048 8880 23112
rect 8800 22952 8880 23048
rect 8800 22888 8808 22952
rect 8872 22888 8880 22952
rect 8800 22792 8880 22888
rect 8800 22728 8808 22792
rect 8872 22728 8880 22792
rect 8800 22632 8880 22728
rect 8800 22568 8808 22632
rect 8872 22568 8880 22632
rect 8800 22472 8880 22568
rect 8800 22408 8808 22472
rect 8872 22408 8880 22472
rect 8800 22312 8880 22408
rect 8800 22248 8808 22312
rect 8872 22248 8880 22312
rect 8800 22152 8880 22248
rect 8800 22088 8808 22152
rect 8872 22088 8880 22152
rect 8800 21992 8880 22088
rect 8800 21928 8808 21992
rect 8872 21928 8880 21992
rect 8800 21832 8880 21928
rect 8800 21768 8808 21832
rect 8872 21768 8880 21832
rect 8800 21672 8880 21768
rect 8800 21608 8808 21672
rect 8872 21608 8880 21672
rect 8800 21512 8880 21608
rect 8800 21448 8808 21512
rect 8872 21448 8880 21512
rect 8800 21352 8880 21448
rect 8800 21288 8808 21352
rect 8872 21288 8880 21352
rect 8800 21192 8880 21288
rect 8800 21128 8808 21192
rect 8872 21128 8880 21192
rect 8800 21032 8880 21128
rect 8800 20968 8808 21032
rect 8872 20968 8880 21032
rect 8800 20872 8880 20968
rect 8800 20808 8808 20872
rect 8872 20808 8880 20872
rect 8800 20712 8880 20808
rect 8800 20648 8808 20712
rect 8872 20648 8880 20712
rect 8800 20552 8880 20648
rect 8800 20488 8808 20552
rect 8872 20488 8880 20552
rect 8800 20392 8880 20488
rect 8800 20328 8808 20392
rect 8872 20328 8880 20392
rect 8800 20232 8880 20328
rect 8800 20168 8808 20232
rect 8872 20168 8880 20232
rect 8800 20072 8880 20168
rect 8800 20008 8808 20072
rect 8872 20008 8880 20072
rect 8800 19912 8880 20008
rect 8800 19848 8808 19912
rect 8872 19848 8880 19912
rect 8800 19752 8880 19848
rect 8800 19688 8808 19752
rect 8872 19688 8880 19752
rect 8800 19592 8880 19688
rect 8800 19528 8808 19592
rect 8872 19528 8880 19592
rect 8800 19432 8880 19528
rect 8800 19368 8808 19432
rect 8872 19368 8880 19432
rect 8800 19272 8880 19368
rect 8800 19208 8808 19272
rect 8872 19208 8880 19272
rect 8800 19112 8880 19208
rect 8800 19048 8808 19112
rect 8872 19048 8880 19112
rect 8800 18952 8880 19048
rect 8800 18888 8808 18952
rect 8872 18888 8880 18952
rect 8800 18792 8880 18888
rect 8800 18728 8808 18792
rect 8872 18728 8880 18792
rect 8800 18632 8880 18728
rect 8800 18568 8808 18632
rect 8872 18568 8880 18632
rect 8800 18472 8880 18568
rect 8800 18408 8808 18472
rect 8872 18408 8880 18472
rect 8800 18312 8880 18408
rect 8800 18248 8808 18312
rect 8872 18248 8880 18312
rect 8800 18152 8880 18248
rect 8800 18088 8808 18152
rect 8872 18088 8880 18152
rect 8800 17992 8880 18088
rect 8800 17928 8808 17992
rect 8872 17928 8880 17992
rect 8800 17832 8880 17928
rect 8800 17768 8808 17832
rect 8872 17768 8880 17832
rect 8800 17672 8880 17768
rect 8800 17608 8808 17672
rect 8872 17608 8880 17672
rect 8800 17512 8880 17608
rect 8800 17448 8808 17512
rect 8872 17448 8880 17512
rect 8800 17352 8880 17448
rect 8800 17288 8808 17352
rect 8872 17288 8880 17352
rect 8800 17192 8880 17288
rect 8800 17128 8808 17192
rect 8872 17128 8880 17192
rect 8800 17032 8880 17128
rect 8800 16968 8808 17032
rect 8872 16968 8880 17032
rect 8800 16872 8880 16968
rect 8800 16808 8808 16872
rect 8872 16808 8880 16872
rect 8800 16712 8880 16808
rect 8800 16648 8808 16712
rect 8872 16648 8880 16712
rect 8800 16552 8880 16648
rect 8800 16488 8808 16552
rect 8872 16488 8880 16552
rect 8800 16392 8880 16488
rect 8800 16328 8808 16392
rect 8872 16328 8880 16392
rect 8800 16232 8880 16328
rect 8800 16168 8808 16232
rect 8872 16168 8880 16232
rect 8800 16072 8880 16168
rect 8800 16008 8808 16072
rect 8872 16008 8880 16072
rect 8800 15912 8880 16008
rect 8800 15848 8808 15912
rect 8872 15848 8880 15912
rect 8800 15752 8880 15848
rect 8800 15688 8808 15752
rect 8872 15688 8880 15752
rect 8800 15592 8880 15688
rect 8800 15528 8808 15592
rect 8872 15528 8880 15592
rect 8800 15432 8880 15528
rect 8800 15368 8808 15432
rect 8872 15368 8880 15432
rect 8800 15272 8880 15368
rect 8800 15208 8808 15272
rect 8872 15208 8880 15272
rect 8800 15112 8880 15208
rect 8800 15048 8808 15112
rect 8872 15048 8880 15112
rect 8800 14952 8880 15048
rect 8800 14888 8808 14952
rect 8872 14888 8880 14952
rect 8800 14792 8880 14888
rect 8800 14728 8808 14792
rect 8872 14728 8880 14792
rect 8800 14632 8880 14728
rect 8800 14568 8808 14632
rect 8872 14568 8880 14632
rect 8800 14472 8880 14568
rect 8800 14408 8808 14472
rect 8872 14408 8880 14472
rect 8800 14312 8880 14408
rect 8800 14248 8808 14312
rect 8872 14248 8880 14312
rect 8800 14152 8880 14248
rect 8800 14088 8808 14152
rect 8872 14088 8880 14152
rect 8800 13992 8880 14088
rect 8800 13928 8808 13992
rect 8872 13928 8880 13992
rect 8800 13832 8880 13928
rect 8800 13768 8808 13832
rect 8872 13768 8880 13832
rect 8800 13672 8880 13768
rect 8800 13608 8808 13672
rect 8872 13608 8880 13672
rect 8800 13512 8880 13608
rect 8800 13448 8808 13512
rect 8872 13448 8880 13512
rect 8800 13352 8880 13448
rect 8800 13288 8808 13352
rect 8872 13288 8880 13352
rect 8800 13192 8880 13288
rect 8800 13128 8808 13192
rect 8872 13128 8880 13192
rect 8800 13032 8880 13128
rect 8800 12968 8808 13032
rect 8872 12968 8880 13032
rect 8800 12872 8880 12968
rect 8800 12808 8808 12872
rect 8872 12808 8880 12872
rect 8800 12712 8880 12808
rect 8800 12648 8808 12712
rect 8872 12648 8880 12712
rect 8800 12552 8880 12648
rect 8800 12488 8808 12552
rect 8872 12488 8880 12552
rect 8800 12392 8880 12488
rect 8800 12328 8808 12392
rect 8872 12328 8880 12392
rect 8800 12232 8880 12328
rect 8800 12168 8808 12232
rect 8872 12168 8880 12232
rect 8800 12072 8880 12168
rect 8800 12008 8808 12072
rect 8872 12008 8880 12072
rect 8800 11912 8880 12008
rect 8800 11848 8808 11912
rect 8872 11848 8880 11912
rect 8800 11752 8880 11848
rect 8800 11688 8808 11752
rect 8872 11688 8880 11752
rect 8800 11592 8880 11688
rect 8800 11528 8808 11592
rect 8872 11528 8880 11592
rect 8800 11432 8880 11528
rect 8800 11368 8808 11432
rect 8872 11368 8880 11432
rect 8800 11272 8880 11368
rect 8800 11208 8808 11272
rect 8872 11208 8880 11272
rect 8800 11112 8880 11208
rect 8800 11048 8808 11112
rect 8872 11048 8880 11112
rect 8800 10952 8880 11048
rect 8800 10888 8808 10952
rect 8872 10888 8880 10952
rect 8800 10792 8880 10888
rect 8800 10728 8808 10792
rect 8872 10728 8880 10792
rect 8800 10632 8880 10728
rect 8800 10568 8808 10632
rect 8872 10568 8880 10632
rect 8800 10472 8880 10568
rect 8800 10408 8808 10472
rect 8872 10408 8880 10472
rect 8800 10312 8880 10408
rect 8800 10248 8808 10312
rect 8872 10248 8880 10312
rect 8800 10152 8880 10248
rect 8800 10088 8808 10152
rect 8872 10088 8880 10152
rect 8800 9992 8880 10088
rect 8800 9928 8808 9992
rect 8872 9928 8880 9992
rect 8800 9832 8880 9928
rect 8800 9768 8808 9832
rect 8872 9768 8880 9832
rect 8800 9672 8880 9768
rect 8800 9608 8808 9672
rect 8872 9608 8880 9672
rect 8800 9512 8880 9608
rect 8800 9448 8808 9512
rect 8872 9448 8880 9512
rect 8800 9352 8880 9448
rect 8800 9288 8808 9352
rect 8872 9288 8880 9352
rect 8800 9192 8880 9288
rect 8800 9128 8808 9192
rect 8872 9128 8880 9192
rect 8800 9032 8880 9128
rect 8800 8968 8808 9032
rect 8872 8968 8880 9032
rect 8800 8872 8880 8968
rect 8800 8808 8808 8872
rect 8872 8808 8880 8872
rect 8800 8712 8880 8808
rect 8800 8648 8808 8712
rect 8872 8648 8880 8712
rect 8800 8552 8880 8648
rect 8800 8488 8808 8552
rect 8872 8488 8880 8552
rect 8800 8392 8880 8488
rect 8800 8328 8808 8392
rect 8872 8328 8880 8392
rect 8800 8232 8880 8328
rect 8800 8168 8808 8232
rect 8872 8168 8880 8232
rect 8800 8072 8880 8168
rect 8800 8008 8808 8072
rect 8872 8008 8880 8072
rect 8800 7912 8880 8008
rect 8800 7848 8808 7912
rect 8872 7848 8880 7912
rect 8800 7752 8880 7848
rect 8800 7688 8808 7752
rect 8872 7688 8880 7752
rect 8800 7592 8880 7688
rect 8800 7528 8808 7592
rect 8872 7528 8880 7592
rect 8800 7432 8880 7528
rect 8800 7368 8808 7432
rect 8872 7368 8880 7432
rect 8800 7272 8880 7368
rect 8800 7208 8808 7272
rect 8872 7208 8880 7272
rect 8800 7112 8880 7208
rect 8800 7048 8808 7112
rect 8872 7048 8880 7112
rect 8800 6952 8880 7048
rect 8800 6888 8808 6952
rect 8872 6888 8880 6952
rect 8800 6792 8880 6888
rect 8800 6728 8808 6792
rect 8872 6728 8880 6792
rect 8800 6632 8880 6728
rect 8800 6568 8808 6632
rect 8872 6568 8880 6632
rect 8800 6472 8880 6568
rect 8800 6408 8808 6472
rect 8872 6408 8880 6472
rect 8800 6312 8880 6408
rect 8800 6248 8808 6312
rect 8872 6248 8880 6312
rect 8800 6152 8880 6248
rect 8800 6088 8808 6152
rect 8872 6088 8880 6152
rect 8800 5992 8880 6088
rect 8800 5928 8808 5992
rect 8872 5928 8880 5992
rect 8800 5832 8880 5928
rect 8800 5768 8808 5832
rect 8872 5768 8880 5832
rect 8800 5672 8880 5768
rect 8800 5608 8808 5672
rect 8872 5608 8880 5672
rect 8800 5512 8880 5608
rect 8800 5448 8808 5512
rect 8872 5448 8880 5512
rect 8800 5352 8880 5448
rect 8800 5288 8808 5352
rect 8872 5288 8880 5352
rect 8800 5192 8880 5288
rect 8800 5128 8808 5192
rect 8872 5128 8880 5192
rect 8800 5032 8880 5128
rect 8800 4968 8808 5032
rect 8872 4968 8880 5032
rect 8800 4872 8880 4968
rect 8800 4808 8808 4872
rect 8872 4808 8880 4872
rect 8800 4712 8880 4808
rect 8800 4648 8808 4712
rect 8872 4648 8880 4712
rect 8800 4552 8880 4648
rect 8800 4488 8808 4552
rect 8872 4488 8880 4552
rect 8800 4392 8880 4488
rect 8800 4328 8808 4392
rect 8872 4328 8880 4392
rect 8800 4232 8880 4328
rect 8800 4168 8808 4232
rect 8872 4168 8880 4232
rect 8800 4072 8880 4168
rect 8800 4008 8808 4072
rect 8872 4008 8880 4072
rect 8800 3912 8880 4008
rect 8800 3848 8808 3912
rect 8872 3848 8880 3912
rect 8800 3752 8880 3848
rect 8800 3688 8808 3752
rect 8872 3688 8880 3752
rect 8800 3592 8880 3688
rect 8800 3528 8808 3592
rect 8872 3528 8880 3592
rect 8800 3432 8880 3528
rect 8800 3368 8808 3432
rect 8872 3368 8880 3432
rect 8800 3272 8880 3368
rect 8800 3208 8808 3272
rect 8872 3208 8880 3272
rect 8800 3112 8880 3208
rect 8800 3048 8808 3112
rect 8872 3048 8880 3112
rect 8800 2952 8880 3048
rect 8800 2888 8808 2952
rect 8872 2888 8880 2952
rect 8800 2792 8880 2888
rect 8800 2728 8808 2792
rect 8872 2728 8880 2792
rect 8800 2632 8880 2728
rect 8800 2568 8808 2632
rect 8872 2568 8880 2632
rect 8800 2472 8880 2568
rect 8800 2408 8808 2472
rect 8872 2408 8880 2472
rect 8800 2312 8880 2408
rect 8800 2248 8808 2312
rect 8872 2248 8880 2312
rect 8800 2152 8880 2248
rect 8800 2088 8808 2152
rect 8872 2088 8880 2152
rect 8800 1992 8880 2088
rect 8800 1928 8808 1992
rect 8872 1928 8880 1992
rect 8800 1832 8880 1928
rect 8800 1768 8808 1832
rect 8872 1768 8880 1832
rect 8800 1672 8880 1768
rect 8800 1608 8808 1672
rect 8872 1608 8880 1672
rect 8800 1512 8880 1608
rect 8800 1448 8808 1512
rect 8872 1448 8880 1512
rect 8800 1352 8880 1448
rect 8800 1288 8808 1352
rect 8872 1288 8880 1352
rect 8800 1192 8880 1288
rect 8800 1128 8808 1192
rect 8872 1128 8880 1192
rect 8800 1032 8880 1128
rect 8800 968 8808 1032
rect 8872 968 8880 1032
rect 8800 872 8880 968
rect 8800 808 8808 872
rect 8872 808 8880 872
rect 8800 712 8880 808
rect 8800 648 8808 712
rect 8872 648 8880 712
rect 8800 552 8880 648
rect 8800 488 8808 552
rect 8872 488 8880 552
rect 8800 392 8880 488
rect 8800 328 8808 392
rect 8872 328 8880 392
rect 8800 232 8880 328
rect 8800 168 8808 232
rect 8872 168 8880 232
rect 8800 72 8880 168
rect 8800 8 8808 72
rect 8872 8 8880 72
rect 8480 -1592 8488 -1528
rect 8552 -1592 8560 -1528
rect 8480 -1608 8560 -1592
rect 8480 -1672 8488 -1608
rect 8552 -1672 8560 -1608
rect 8480 -1688 8560 -1672
rect 8480 -1752 8488 -1688
rect 8552 -1752 8560 -1688
rect 8480 -1768 8560 -1752
rect 8480 -1832 8488 -1768
rect 8552 -1832 8560 -1768
rect 8480 -1848 8560 -1832
rect 8480 -1912 8488 -1848
rect 8552 -1912 8560 -1848
rect 8480 -1920 8560 -1912
rect 8800 -1528 8880 8
rect 8800 -1592 8808 -1528
rect 8872 -1592 8880 -1528
rect 8800 -1608 8880 -1592
rect 8800 -1672 8808 -1608
rect 8872 -1672 8880 -1608
rect 8800 -1688 8880 -1672
rect 8800 -1752 8808 -1688
rect 8872 -1752 8880 -1688
rect 8800 -1768 8880 -1752
rect 8800 -1832 8808 -1768
rect 8872 -1832 8880 -1768
rect 8800 -1848 8880 -1832
rect 8800 -1912 8808 -1848
rect 8872 -1912 8880 -1848
rect 8800 -1920 8880 -1912
rect 8960 31432 9040 31520
rect 8960 31368 8968 31432
rect 9032 31368 9040 31432
rect 8960 31272 9040 31368
rect 8960 31208 8968 31272
rect 9032 31208 9040 31272
rect 8960 31112 9040 31208
rect 8960 31048 8968 31112
rect 9032 31048 9040 31112
rect 8960 30952 9040 31048
rect 8960 30888 8968 30952
rect 9032 30888 9040 30952
rect 8960 30792 9040 30888
rect 8960 30728 8968 30792
rect 9032 30728 9040 30792
rect 8960 30632 9040 30728
rect 8960 30568 8968 30632
rect 9032 30568 9040 30632
rect 8960 30472 9040 30568
rect 8960 30408 8968 30472
rect 9032 30408 9040 30472
rect 8960 30312 9040 30408
rect 8960 30248 8968 30312
rect 9032 30248 9040 30312
rect 8960 30152 9040 30248
rect 8960 30088 8968 30152
rect 9032 30088 9040 30152
rect 8960 29992 9040 30088
rect 8960 29928 8968 29992
rect 9032 29928 9040 29992
rect 8960 29832 9040 29928
rect 8960 29768 8968 29832
rect 9032 29768 9040 29832
rect 8960 29672 9040 29768
rect 8960 29608 8968 29672
rect 9032 29608 9040 29672
rect 8960 29512 9040 29608
rect 8960 29448 8968 29512
rect 9032 29448 9040 29512
rect 8960 29352 9040 29448
rect 8960 29288 8968 29352
rect 9032 29288 9040 29352
rect 8960 29192 9040 29288
rect 8960 29128 8968 29192
rect 9032 29128 9040 29192
rect 8960 29032 9040 29128
rect 8960 28968 8968 29032
rect 9032 28968 9040 29032
rect 8960 28872 9040 28968
rect 8960 28808 8968 28872
rect 9032 28808 9040 28872
rect 8960 28712 9040 28808
rect 8960 28648 8968 28712
rect 9032 28648 9040 28712
rect 8960 28552 9040 28648
rect 8960 28488 8968 28552
rect 9032 28488 9040 28552
rect 8960 28392 9040 28488
rect 8960 28328 8968 28392
rect 9032 28328 9040 28392
rect 8960 28232 9040 28328
rect 8960 28168 8968 28232
rect 9032 28168 9040 28232
rect 8960 28072 9040 28168
rect 8960 28008 8968 28072
rect 9032 28008 9040 28072
rect 8960 27912 9040 28008
rect 8960 27848 8968 27912
rect 9032 27848 9040 27912
rect 8960 27752 9040 27848
rect 8960 27688 8968 27752
rect 9032 27688 9040 27752
rect 8960 27592 9040 27688
rect 8960 27528 8968 27592
rect 9032 27528 9040 27592
rect 8960 27432 9040 27528
rect 8960 27368 8968 27432
rect 9032 27368 9040 27432
rect 8960 27272 9040 27368
rect 8960 27208 8968 27272
rect 9032 27208 9040 27272
rect 8960 27112 9040 27208
rect 8960 27048 8968 27112
rect 9032 27048 9040 27112
rect 8960 26952 9040 27048
rect 8960 26888 8968 26952
rect 9032 26888 9040 26952
rect 8960 26792 9040 26888
rect 8960 26728 8968 26792
rect 9032 26728 9040 26792
rect 8960 26632 9040 26728
rect 8960 26568 8968 26632
rect 9032 26568 9040 26632
rect 8960 26472 9040 26568
rect 8960 26408 8968 26472
rect 9032 26408 9040 26472
rect 8960 26312 9040 26408
rect 8960 26248 8968 26312
rect 9032 26248 9040 26312
rect 8960 26152 9040 26248
rect 8960 26088 8968 26152
rect 9032 26088 9040 26152
rect 8960 25992 9040 26088
rect 8960 25928 8968 25992
rect 9032 25928 9040 25992
rect 8960 25832 9040 25928
rect 8960 25768 8968 25832
rect 9032 25768 9040 25832
rect 8960 25672 9040 25768
rect 8960 25608 8968 25672
rect 9032 25608 9040 25672
rect 8960 25512 9040 25608
rect 8960 25448 8968 25512
rect 9032 25448 9040 25512
rect 8960 25352 9040 25448
rect 8960 25288 8968 25352
rect 9032 25288 9040 25352
rect 8960 25192 9040 25288
rect 8960 25128 8968 25192
rect 9032 25128 9040 25192
rect 8960 25032 9040 25128
rect 8960 24968 8968 25032
rect 9032 24968 9040 25032
rect 8960 24872 9040 24968
rect 8960 24808 8968 24872
rect 9032 24808 9040 24872
rect 8960 24712 9040 24808
rect 8960 24648 8968 24712
rect 9032 24648 9040 24712
rect 8960 24552 9040 24648
rect 8960 24488 8968 24552
rect 9032 24488 9040 24552
rect 8960 24392 9040 24488
rect 8960 24328 8968 24392
rect 9032 24328 9040 24392
rect 8960 24232 9040 24328
rect 8960 24168 8968 24232
rect 9032 24168 9040 24232
rect 8960 24072 9040 24168
rect 8960 24008 8968 24072
rect 9032 24008 9040 24072
rect 8960 23912 9040 24008
rect 8960 23848 8968 23912
rect 9032 23848 9040 23912
rect 8960 23752 9040 23848
rect 8960 23688 8968 23752
rect 9032 23688 9040 23752
rect 8960 23592 9040 23688
rect 8960 23528 8968 23592
rect 9032 23528 9040 23592
rect 8960 23432 9040 23528
rect 8960 23368 8968 23432
rect 9032 23368 9040 23432
rect 8960 23272 9040 23368
rect 8960 23208 8968 23272
rect 9032 23208 9040 23272
rect 8960 23112 9040 23208
rect 8960 23048 8968 23112
rect 9032 23048 9040 23112
rect 8960 22952 9040 23048
rect 8960 22888 8968 22952
rect 9032 22888 9040 22952
rect 8960 22792 9040 22888
rect 8960 22728 8968 22792
rect 9032 22728 9040 22792
rect 8960 22632 9040 22728
rect 8960 22568 8968 22632
rect 9032 22568 9040 22632
rect 8960 22472 9040 22568
rect 8960 22408 8968 22472
rect 9032 22408 9040 22472
rect 8960 22312 9040 22408
rect 8960 22248 8968 22312
rect 9032 22248 9040 22312
rect 8960 22152 9040 22248
rect 8960 22088 8968 22152
rect 9032 22088 9040 22152
rect 8960 21992 9040 22088
rect 8960 21928 8968 21992
rect 9032 21928 9040 21992
rect 8960 21832 9040 21928
rect 8960 21768 8968 21832
rect 9032 21768 9040 21832
rect 8960 21672 9040 21768
rect 8960 21608 8968 21672
rect 9032 21608 9040 21672
rect 8960 21512 9040 21608
rect 8960 21448 8968 21512
rect 9032 21448 9040 21512
rect 8960 21352 9040 21448
rect 8960 21288 8968 21352
rect 9032 21288 9040 21352
rect 8960 21192 9040 21288
rect 8960 21128 8968 21192
rect 9032 21128 9040 21192
rect 8960 21032 9040 21128
rect 8960 20968 8968 21032
rect 9032 20968 9040 21032
rect 8960 20872 9040 20968
rect 8960 20808 8968 20872
rect 9032 20808 9040 20872
rect 8960 20712 9040 20808
rect 8960 20648 8968 20712
rect 9032 20648 9040 20712
rect 8960 20552 9040 20648
rect 8960 20488 8968 20552
rect 9032 20488 9040 20552
rect 8960 20392 9040 20488
rect 8960 20328 8968 20392
rect 9032 20328 9040 20392
rect 8960 20232 9040 20328
rect 8960 20168 8968 20232
rect 9032 20168 9040 20232
rect 8960 20072 9040 20168
rect 8960 20008 8968 20072
rect 9032 20008 9040 20072
rect 8960 19912 9040 20008
rect 8960 19848 8968 19912
rect 9032 19848 9040 19912
rect 8960 19752 9040 19848
rect 8960 19688 8968 19752
rect 9032 19688 9040 19752
rect 8960 19592 9040 19688
rect 8960 19528 8968 19592
rect 9032 19528 9040 19592
rect 8960 19432 9040 19528
rect 8960 19368 8968 19432
rect 9032 19368 9040 19432
rect 8960 19272 9040 19368
rect 8960 19208 8968 19272
rect 9032 19208 9040 19272
rect 8960 19112 9040 19208
rect 8960 19048 8968 19112
rect 9032 19048 9040 19112
rect 8960 18952 9040 19048
rect 8960 18888 8968 18952
rect 9032 18888 9040 18952
rect 8960 18792 9040 18888
rect 8960 18728 8968 18792
rect 9032 18728 9040 18792
rect 8960 18632 9040 18728
rect 8960 18568 8968 18632
rect 9032 18568 9040 18632
rect 8960 18472 9040 18568
rect 8960 18408 8968 18472
rect 9032 18408 9040 18472
rect 8960 18312 9040 18408
rect 8960 18248 8968 18312
rect 9032 18248 9040 18312
rect 8960 18152 9040 18248
rect 8960 18088 8968 18152
rect 9032 18088 9040 18152
rect 8960 17992 9040 18088
rect 8960 17928 8968 17992
rect 9032 17928 9040 17992
rect 8960 17832 9040 17928
rect 8960 17768 8968 17832
rect 9032 17768 9040 17832
rect 8960 17672 9040 17768
rect 8960 17608 8968 17672
rect 9032 17608 9040 17672
rect 8960 17512 9040 17608
rect 8960 17448 8968 17512
rect 9032 17448 9040 17512
rect 8960 17352 9040 17448
rect 8960 17288 8968 17352
rect 9032 17288 9040 17352
rect 8960 17192 9040 17288
rect 8960 17128 8968 17192
rect 9032 17128 9040 17192
rect 8960 17032 9040 17128
rect 8960 16968 8968 17032
rect 9032 16968 9040 17032
rect 8960 16872 9040 16968
rect 8960 16808 8968 16872
rect 9032 16808 9040 16872
rect 8960 16712 9040 16808
rect 8960 16648 8968 16712
rect 9032 16648 9040 16712
rect 8960 16552 9040 16648
rect 8960 16488 8968 16552
rect 9032 16488 9040 16552
rect 8960 16392 9040 16488
rect 8960 16328 8968 16392
rect 9032 16328 9040 16392
rect 8960 16232 9040 16328
rect 8960 16168 8968 16232
rect 9032 16168 9040 16232
rect 8960 16072 9040 16168
rect 8960 16008 8968 16072
rect 9032 16008 9040 16072
rect 8960 15912 9040 16008
rect 8960 15848 8968 15912
rect 9032 15848 9040 15912
rect 8960 15752 9040 15848
rect 8960 15688 8968 15752
rect 9032 15688 9040 15752
rect 8960 15592 9040 15688
rect 8960 15528 8968 15592
rect 9032 15528 9040 15592
rect 8960 15432 9040 15528
rect 8960 15368 8968 15432
rect 9032 15368 9040 15432
rect 8960 15272 9040 15368
rect 8960 15208 8968 15272
rect 9032 15208 9040 15272
rect 8960 15112 9040 15208
rect 8960 15048 8968 15112
rect 9032 15048 9040 15112
rect 8960 14952 9040 15048
rect 8960 14888 8968 14952
rect 9032 14888 9040 14952
rect 8960 14792 9040 14888
rect 8960 14728 8968 14792
rect 9032 14728 9040 14792
rect 8960 14632 9040 14728
rect 8960 14568 8968 14632
rect 9032 14568 9040 14632
rect 8960 14472 9040 14568
rect 8960 14408 8968 14472
rect 9032 14408 9040 14472
rect 8960 14312 9040 14408
rect 8960 14248 8968 14312
rect 9032 14248 9040 14312
rect 8960 14152 9040 14248
rect 8960 14088 8968 14152
rect 9032 14088 9040 14152
rect 8960 13992 9040 14088
rect 8960 13928 8968 13992
rect 9032 13928 9040 13992
rect 8960 13832 9040 13928
rect 8960 13768 8968 13832
rect 9032 13768 9040 13832
rect 8960 13672 9040 13768
rect 8960 13608 8968 13672
rect 9032 13608 9040 13672
rect 8960 13512 9040 13608
rect 8960 13448 8968 13512
rect 9032 13448 9040 13512
rect 8960 13352 9040 13448
rect 8960 13288 8968 13352
rect 9032 13288 9040 13352
rect 8960 13192 9040 13288
rect 8960 13128 8968 13192
rect 9032 13128 9040 13192
rect 8960 13032 9040 13128
rect 8960 12968 8968 13032
rect 9032 12968 9040 13032
rect 8960 12872 9040 12968
rect 8960 12808 8968 12872
rect 9032 12808 9040 12872
rect 8960 12712 9040 12808
rect 8960 12648 8968 12712
rect 9032 12648 9040 12712
rect 8960 12552 9040 12648
rect 8960 12488 8968 12552
rect 9032 12488 9040 12552
rect 8960 12392 9040 12488
rect 8960 12328 8968 12392
rect 9032 12328 9040 12392
rect 8960 12232 9040 12328
rect 8960 12168 8968 12232
rect 9032 12168 9040 12232
rect 8960 12072 9040 12168
rect 8960 12008 8968 12072
rect 9032 12008 9040 12072
rect 8960 11912 9040 12008
rect 8960 11848 8968 11912
rect 9032 11848 9040 11912
rect 8960 11752 9040 11848
rect 8960 11688 8968 11752
rect 9032 11688 9040 11752
rect 8960 11592 9040 11688
rect 8960 11528 8968 11592
rect 9032 11528 9040 11592
rect 8960 11432 9040 11528
rect 8960 11368 8968 11432
rect 9032 11368 9040 11432
rect 8960 11272 9040 11368
rect 8960 11208 8968 11272
rect 9032 11208 9040 11272
rect 8960 11112 9040 11208
rect 8960 11048 8968 11112
rect 9032 11048 9040 11112
rect 8960 10952 9040 11048
rect 8960 10888 8968 10952
rect 9032 10888 9040 10952
rect 8960 10792 9040 10888
rect 8960 10728 8968 10792
rect 9032 10728 9040 10792
rect 8960 10632 9040 10728
rect 8960 10568 8968 10632
rect 9032 10568 9040 10632
rect 8960 10472 9040 10568
rect 8960 10408 8968 10472
rect 9032 10408 9040 10472
rect 8960 10312 9040 10408
rect 8960 10248 8968 10312
rect 9032 10248 9040 10312
rect 8960 10152 9040 10248
rect 8960 10088 8968 10152
rect 9032 10088 9040 10152
rect 8960 9992 9040 10088
rect 8960 9928 8968 9992
rect 9032 9928 9040 9992
rect 8960 9832 9040 9928
rect 8960 9768 8968 9832
rect 9032 9768 9040 9832
rect 8960 9672 9040 9768
rect 8960 9608 8968 9672
rect 9032 9608 9040 9672
rect 8960 9512 9040 9608
rect 8960 9448 8968 9512
rect 9032 9448 9040 9512
rect 8960 9352 9040 9448
rect 8960 9288 8968 9352
rect 9032 9288 9040 9352
rect 8960 9192 9040 9288
rect 8960 9128 8968 9192
rect 9032 9128 9040 9192
rect 8960 9032 9040 9128
rect 8960 8968 8968 9032
rect 9032 8968 9040 9032
rect 8960 8872 9040 8968
rect 8960 8808 8968 8872
rect 9032 8808 9040 8872
rect 8960 8712 9040 8808
rect 8960 8648 8968 8712
rect 9032 8648 9040 8712
rect 8960 8552 9040 8648
rect 8960 8488 8968 8552
rect 9032 8488 9040 8552
rect 8960 8392 9040 8488
rect 8960 8328 8968 8392
rect 9032 8328 9040 8392
rect 8960 8232 9040 8328
rect 8960 8168 8968 8232
rect 9032 8168 9040 8232
rect 8960 8072 9040 8168
rect 8960 8008 8968 8072
rect 9032 8008 9040 8072
rect 8960 7912 9040 8008
rect 8960 7848 8968 7912
rect 9032 7848 9040 7912
rect 8960 7752 9040 7848
rect 8960 7688 8968 7752
rect 9032 7688 9040 7752
rect 8960 7592 9040 7688
rect 8960 7528 8968 7592
rect 9032 7528 9040 7592
rect 8960 7432 9040 7528
rect 8960 7368 8968 7432
rect 9032 7368 9040 7432
rect 8960 7272 9040 7368
rect 8960 7208 8968 7272
rect 9032 7208 9040 7272
rect 8960 7112 9040 7208
rect 8960 7048 8968 7112
rect 9032 7048 9040 7112
rect 8960 6952 9040 7048
rect 8960 6888 8968 6952
rect 9032 6888 9040 6952
rect 8960 6792 9040 6888
rect 8960 6728 8968 6792
rect 9032 6728 9040 6792
rect 8960 6632 9040 6728
rect 8960 6568 8968 6632
rect 9032 6568 9040 6632
rect 8960 6472 9040 6568
rect 8960 6408 8968 6472
rect 9032 6408 9040 6472
rect 8960 6312 9040 6408
rect 8960 6248 8968 6312
rect 9032 6248 9040 6312
rect 8960 6152 9040 6248
rect 8960 6088 8968 6152
rect 9032 6088 9040 6152
rect 8960 5992 9040 6088
rect 8960 5928 8968 5992
rect 9032 5928 9040 5992
rect 8960 5832 9040 5928
rect 8960 5768 8968 5832
rect 9032 5768 9040 5832
rect 8960 5672 9040 5768
rect 8960 5608 8968 5672
rect 9032 5608 9040 5672
rect 8960 5512 9040 5608
rect 8960 5448 8968 5512
rect 9032 5448 9040 5512
rect 8960 5352 9040 5448
rect 8960 5288 8968 5352
rect 9032 5288 9040 5352
rect 8960 5192 9040 5288
rect 8960 5128 8968 5192
rect 9032 5128 9040 5192
rect 8960 5032 9040 5128
rect 8960 4968 8968 5032
rect 9032 4968 9040 5032
rect 8960 4872 9040 4968
rect 8960 4808 8968 4872
rect 9032 4808 9040 4872
rect 8960 4712 9040 4808
rect 8960 4648 8968 4712
rect 9032 4648 9040 4712
rect 8960 4552 9040 4648
rect 8960 4488 8968 4552
rect 9032 4488 9040 4552
rect 8960 4392 9040 4488
rect 8960 4328 8968 4392
rect 9032 4328 9040 4392
rect 8960 4232 9040 4328
rect 8960 4168 8968 4232
rect 9032 4168 9040 4232
rect 8960 4072 9040 4168
rect 8960 4008 8968 4072
rect 9032 4008 9040 4072
rect 8960 3912 9040 4008
rect 8960 3848 8968 3912
rect 9032 3848 9040 3912
rect 8960 3752 9040 3848
rect 8960 3688 8968 3752
rect 9032 3688 9040 3752
rect 8960 3592 9040 3688
rect 8960 3528 8968 3592
rect 9032 3528 9040 3592
rect 8960 3432 9040 3528
rect 8960 3368 8968 3432
rect 9032 3368 9040 3432
rect 8960 3272 9040 3368
rect 8960 3208 8968 3272
rect 9032 3208 9040 3272
rect 8960 3112 9040 3208
rect 8960 3048 8968 3112
rect 9032 3048 9040 3112
rect 8960 2952 9040 3048
rect 8960 2888 8968 2952
rect 9032 2888 9040 2952
rect 8960 2792 9040 2888
rect 8960 2728 8968 2792
rect 9032 2728 9040 2792
rect 8960 2632 9040 2728
rect 8960 2568 8968 2632
rect 9032 2568 9040 2632
rect 8960 2472 9040 2568
rect 8960 2408 8968 2472
rect 9032 2408 9040 2472
rect 8960 2312 9040 2408
rect 8960 2248 8968 2312
rect 9032 2248 9040 2312
rect 8960 2152 9040 2248
rect 8960 2088 8968 2152
rect 9032 2088 9040 2152
rect 8960 1992 9040 2088
rect 8960 1928 8968 1992
rect 9032 1928 9040 1992
rect 8960 1832 9040 1928
rect 8960 1768 8968 1832
rect 9032 1768 9040 1832
rect 8960 1672 9040 1768
rect 8960 1608 8968 1672
rect 9032 1608 9040 1672
rect 8960 1512 9040 1608
rect 8960 1448 8968 1512
rect 9032 1448 9040 1512
rect 8960 1352 9040 1448
rect 8960 1288 8968 1352
rect 9032 1288 9040 1352
rect 8960 1192 9040 1288
rect 8960 1128 8968 1192
rect 9032 1128 9040 1192
rect 8960 1032 9040 1128
rect 8960 968 8968 1032
rect 9032 968 9040 1032
rect 8960 872 9040 968
rect 8960 808 8968 872
rect 9032 808 9040 872
rect 8960 712 9040 808
rect 8960 648 8968 712
rect 9032 648 9040 712
rect 8960 552 9040 648
rect 8960 488 8968 552
rect 9032 488 9040 552
rect 8960 392 9040 488
rect 8960 328 8968 392
rect 9032 328 9040 392
rect 8960 232 9040 328
rect 8960 168 8968 232
rect 9032 168 9040 232
rect 8960 72 9040 168
rect 8960 8 8968 72
rect 9032 8 9040 72
rect 8960 -568 9040 8
rect 8960 -632 8968 -568
rect 9032 -632 9040 -568
rect 8960 -648 9040 -632
rect 8960 -712 8968 -648
rect 9032 -712 9040 -648
rect 8960 -728 9040 -712
rect 8960 -792 8968 -728
rect 9032 -792 9040 -728
rect 8960 -808 9040 -792
rect 8960 -872 8968 -808
rect 9032 -872 9040 -808
rect 8960 -888 9040 -872
rect 8960 -952 8968 -888
rect 9032 -952 9040 -888
rect 240 -2008 320 -2000
rect 240 -2072 248 -2008
rect 312 -2072 320 -2008
rect 240 -4568 320 -2072
rect 8960 -2008 9040 -952
rect 8960 -2072 8968 -2008
rect 9032 -2072 9040 -2008
rect 8960 -2080 9040 -2072
rect 9120 30148 9200 31520
rect 9120 30092 9132 30148
rect 9188 30092 9200 30148
rect 9120 24868 9200 30092
rect 9120 24812 9132 24868
rect 9188 24812 9200 24868
rect 9120 21988 9200 24812
rect 9120 21932 9132 21988
rect 9188 21932 9200 21988
rect 9120 16708 9200 21932
rect 9120 16652 9132 16708
rect 9188 16652 9200 16708
rect 9120 13828 9200 16652
rect 9120 13772 9132 13828
rect 9188 13772 9200 13828
rect 9120 7108 9200 13772
rect 9120 7052 9132 7108
rect 9188 7052 9200 7108
rect 9120 3668 9200 7052
rect 9120 3612 9132 3668
rect 9188 3612 9200 3668
rect 9120 -2160 9200 3612
rect 9280 31432 9360 31520
rect 9280 31368 9288 31432
rect 9352 31368 9360 31432
rect 9280 31272 9360 31368
rect 9280 31208 9288 31272
rect 9352 31208 9360 31272
rect 9280 31112 9360 31208
rect 9280 31048 9288 31112
rect 9352 31048 9360 31112
rect 9280 30952 9360 31048
rect 9280 30888 9288 30952
rect 9352 30888 9360 30952
rect 9280 30792 9360 30888
rect 9280 30728 9288 30792
rect 9352 30728 9360 30792
rect 9280 30632 9360 30728
rect 9280 30568 9288 30632
rect 9352 30568 9360 30632
rect 9280 30472 9360 30568
rect 9280 30408 9288 30472
rect 9352 30408 9360 30472
rect 9280 30312 9360 30408
rect 9280 30248 9288 30312
rect 9352 30248 9360 30312
rect 9280 30152 9360 30248
rect 9280 30088 9288 30152
rect 9352 30088 9360 30152
rect 9280 29992 9360 30088
rect 9280 29928 9288 29992
rect 9352 29928 9360 29992
rect 9280 29832 9360 29928
rect 9280 29768 9288 29832
rect 9352 29768 9360 29832
rect 9280 29672 9360 29768
rect 9280 29608 9288 29672
rect 9352 29608 9360 29672
rect 9280 29512 9360 29608
rect 9280 29448 9288 29512
rect 9352 29448 9360 29512
rect 9280 29352 9360 29448
rect 9280 29288 9288 29352
rect 9352 29288 9360 29352
rect 9280 29192 9360 29288
rect 9280 29128 9288 29192
rect 9352 29128 9360 29192
rect 9280 29032 9360 29128
rect 9280 28968 9288 29032
rect 9352 28968 9360 29032
rect 9280 28872 9360 28968
rect 9280 28808 9288 28872
rect 9352 28808 9360 28872
rect 9280 28712 9360 28808
rect 9280 28648 9288 28712
rect 9352 28648 9360 28712
rect 9280 28552 9360 28648
rect 9280 28488 9288 28552
rect 9352 28488 9360 28552
rect 9280 28392 9360 28488
rect 9280 28328 9288 28392
rect 9352 28328 9360 28392
rect 9280 28232 9360 28328
rect 9280 28168 9288 28232
rect 9352 28168 9360 28232
rect 9280 28072 9360 28168
rect 9280 28008 9288 28072
rect 9352 28008 9360 28072
rect 9280 27912 9360 28008
rect 9280 27848 9288 27912
rect 9352 27848 9360 27912
rect 9280 27752 9360 27848
rect 9280 27688 9288 27752
rect 9352 27688 9360 27752
rect 9280 27592 9360 27688
rect 9280 27528 9288 27592
rect 9352 27528 9360 27592
rect 9280 27432 9360 27528
rect 9280 27368 9288 27432
rect 9352 27368 9360 27432
rect 9280 27272 9360 27368
rect 9280 27208 9288 27272
rect 9352 27208 9360 27272
rect 9280 27112 9360 27208
rect 9280 27048 9288 27112
rect 9352 27048 9360 27112
rect 9280 26952 9360 27048
rect 9280 26888 9288 26952
rect 9352 26888 9360 26952
rect 9280 26792 9360 26888
rect 9280 26728 9288 26792
rect 9352 26728 9360 26792
rect 9280 26632 9360 26728
rect 9280 26568 9288 26632
rect 9352 26568 9360 26632
rect 9280 26472 9360 26568
rect 9280 26408 9288 26472
rect 9352 26408 9360 26472
rect 9280 26312 9360 26408
rect 9280 26248 9288 26312
rect 9352 26248 9360 26312
rect 9280 26152 9360 26248
rect 9280 26088 9288 26152
rect 9352 26088 9360 26152
rect 9280 25992 9360 26088
rect 9280 25928 9288 25992
rect 9352 25928 9360 25992
rect 9280 25832 9360 25928
rect 9280 25768 9288 25832
rect 9352 25768 9360 25832
rect 9280 25672 9360 25768
rect 9280 25608 9288 25672
rect 9352 25608 9360 25672
rect 9280 25512 9360 25608
rect 9280 25448 9288 25512
rect 9352 25448 9360 25512
rect 9280 25352 9360 25448
rect 9280 25288 9288 25352
rect 9352 25288 9360 25352
rect 9280 25192 9360 25288
rect 9280 25128 9288 25192
rect 9352 25128 9360 25192
rect 9280 25032 9360 25128
rect 9280 24968 9288 25032
rect 9352 24968 9360 25032
rect 9280 24872 9360 24968
rect 9280 24808 9288 24872
rect 9352 24808 9360 24872
rect 9280 24712 9360 24808
rect 9280 24648 9288 24712
rect 9352 24648 9360 24712
rect 9280 24552 9360 24648
rect 9280 24488 9288 24552
rect 9352 24488 9360 24552
rect 9280 24392 9360 24488
rect 9280 24328 9288 24392
rect 9352 24328 9360 24392
rect 9280 24232 9360 24328
rect 9280 24168 9288 24232
rect 9352 24168 9360 24232
rect 9280 24072 9360 24168
rect 9280 24008 9288 24072
rect 9352 24008 9360 24072
rect 9280 23912 9360 24008
rect 9280 23848 9288 23912
rect 9352 23848 9360 23912
rect 9280 23752 9360 23848
rect 9280 23688 9288 23752
rect 9352 23688 9360 23752
rect 9280 23592 9360 23688
rect 9280 23528 9288 23592
rect 9352 23528 9360 23592
rect 9280 23432 9360 23528
rect 9280 23368 9288 23432
rect 9352 23368 9360 23432
rect 9280 23272 9360 23368
rect 9280 23208 9288 23272
rect 9352 23208 9360 23272
rect 9280 23112 9360 23208
rect 9280 23048 9288 23112
rect 9352 23048 9360 23112
rect 9280 22952 9360 23048
rect 9280 22888 9288 22952
rect 9352 22888 9360 22952
rect 9280 22792 9360 22888
rect 9280 22728 9288 22792
rect 9352 22728 9360 22792
rect 9280 22632 9360 22728
rect 9280 22568 9288 22632
rect 9352 22568 9360 22632
rect 9280 22472 9360 22568
rect 9280 22408 9288 22472
rect 9352 22408 9360 22472
rect 9280 22312 9360 22408
rect 9280 22248 9288 22312
rect 9352 22248 9360 22312
rect 9280 22152 9360 22248
rect 9280 22088 9288 22152
rect 9352 22088 9360 22152
rect 9280 21992 9360 22088
rect 9280 21928 9288 21992
rect 9352 21928 9360 21992
rect 9280 21832 9360 21928
rect 9280 21768 9288 21832
rect 9352 21768 9360 21832
rect 9280 21672 9360 21768
rect 9280 21608 9288 21672
rect 9352 21608 9360 21672
rect 9280 21512 9360 21608
rect 9280 21448 9288 21512
rect 9352 21448 9360 21512
rect 9280 21352 9360 21448
rect 9280 21288 9288 21352
rect 9352 21288 9360 21352
rect 9280 21192 9360 21288
rect 9280 21128 9288 21192
rect 9352 21128 9360 21192
rect 9280 21032 9360 21128
rect 9280 20968 9288 21032
rect 9352 20968 9360 21032
rect 9280 20872 9360 20968
rect 9280 20808 9288 20872
rect 9352 20808 9360 20872
rect 9280 20712 9360 20808
rect 9280 20648 9288 20712
rect 9352 20648 9360 20712
rect 9280 20552 9360 20648
rect 9280 20488 9288 20552
rect 9352 20488 9360 20552
rect 9280 20392 9360 20488
rect 9280 20328 9288 20392
rect 9352 20328 9360 20392
rect 9280 20232 9360 20328
rect 9280 20168 9288 20232
rect 9352 20168 9360 20232
rect 9280 20072 9360 20168
rect 9280 20008 9288 20072
rect 9352 20008 9360 20072
rect 9280 19912 9360 20008
rect 9280 19848 9288 19912
rect 9352 19848 9360 19912
rect 9280 19752 9360 19848
rect 9280 19688 9288 19752
rect 9352 19688 9360 19752
rect 9280 19592 9360 19688
rect 9280 19528 9288 19592
rect 9352 19528 9360 19592
rect 9280 19432 9360 19528
rect 9280 19368 9288 19432
rect 9352 19368 9360 19432
rect 9280 19272 9360 19368
rect 9280 19208 9288 19272
rect 9352 19208 9360 19272
rect 9280 19112 9360 19208
rect 9280 19048 9288 19112
rect 9352 19048 9360 19112
rect 9280 18952 9360 19048
rect 9280 18888 9288 18952
rect 9352 18888 9360 18952
rect 9280 18792 9360 18888
rect 9280 18728 9288 18792
rect 9352 18728 9360 18792
rect 9280 18632 9360 18728
rect 9280 18568 9288 18632
rect 9352 18568 9360 18632
rect 9280 18472 9360 18568
rect 9280 18408 9288 18472
rect 9352 18408 9360 18472
rect 9280 18312 9360 18408
rect 9280 18248 9288 18312
rect 9352 18248 9360 18312
rect 9280 18152 9360 18248
rect 9280 18088 9288 18152
rect 9352 18088 9360 18152
rect 9280 17992 9360 18088
rect 9280 17928 9288 17992
rect 9352 17928 9360 17992
rect 9280 17832 9360 17928
rect 9280 17768 9288 17832
rect 9352 17768 9360 17832
rect 9280 17672 9360 17768
rect 9280 17608 9288 17672
rect 9352 17608 9360 17672
rect 9280 17512 9360 17608
rect 9280 17448 9288 17512
rect 9352 17448 9360 17512
rect 9280 17352 9360 17448
rect 9280 17288 9288 17352
rect 9352 17288 9360 17352
rect 9280 17192 9360 17288
rect 9280 17128 9288 17192
rect 9352 17128 9360 17192
rect 9280 17032 9360 17128
rect 9280 16968 9288 17032
rect 9352 16968 9360 17032
rect 9280 16872 9360 16968
rect 9280 16808 9288 16872
rect 9352 16808 9360 16872
rect 9280 16712 9360 16808
rect 9280 16648 9288 16712
rect 9352 16648 9360 16712
rect 9280 16552 9360 16648
rect 9280 16488 9288 16552
rect 9352 16488 9360 16552
rect 9280 16392 9360 16488
rect 9280 16328 9288 16392
rect 9352 16328 9360 16392
rect 9280 16232 9360 16328
rect 9280 16168 9288 16232
rect 9352 16168 9360 16232
rect 9280 16072 9360 16168
rect 9280 16008 9288 16072
rect 9352 16008 9360 16072
rect 9280 15912 9360 16008
rect 9280 15848 9288 15912
rect 9352 15848 9360 15912
rect 9280 15752 9360 15848
rect 9280 15688 9288 15752
rect 9352 15688 9360 15752
rect 9280 15592 9360 15688
rect 9280 15528 9288 15592
rect 9352 15528 9360 15592
rect 9280 15432 9360 15528
rect 9280 15368 9288 15432
rect 9352 15368 9360 15432
rect 9280 15272 9360 15368
rect 9280 15208 9288 15272
rect 9352 15208 9360 15272
rect 9280 15112 9360 15208
rect 9280 15048 9288 15112
rect 9352 15048 9360 15112
rect 9280 14952 9360 15048
rect 9280 14888 9288 14952
rect 9352 14888 9360 14952
rect 9280 14792 9360 14888
rect 9280 14728 9288 14792
rect 9352 14728 9360 14792
rect 9280 14632 9360 14728
rect 9280 14568 9288 14632
rect 9352 14568 9360 14632
rect 9280 14472 9360 14568
rect 9280 14408 9288 14472
rect 9352 14408 9360 14472
rect 9280 14312 9360 14408
rect 9280 14248 9288 14312
rect 9352 14248 9360 14312
rect 9280 14152 9360 14248
rect 9280 14088 9288 14152
rect 9352 14088 9360 14152
rect 9280 13992 9360 14088
rect 9280 13928 9288 13992
rect 9352 13928 9360 13992
rect 9280 13832 9360 13928
rect 9280 13768 9288 13832
rect 9352 13768 9360 13832
rect 9280 13672 9360 13768
rect 9280 13608 9288 13672
rect 9352 13608 9360 13672
rect 9280 13512 9360 13608
rect 9280 13448 9288 13512
rect 9352 13448 9360 13512
rect 9280 13352 9360 13448
rect 9280 13288 9288 13352
rect 9352 13288 9360 13352
rect 9280 13192 9360 13288
rect 9280 13128 9288 13192
rect 9352 13128 9360 13192
rect 9280 13032 9360 13128
rect 9280 12968 9288 13032
rect 9352 12968 9360 13032
rect 9280 12872 9360 12968
rect 9280 12808 9288 12872
rect 9352 12808 9360 12872
rect 9280 12712 9360 12808
rect 9280 12648 9288 12712
rect 9352 12648 9360 12712
rect 9280 12552 9360 12648
rect 9280 12488 9288 12552
rect 9352 12488 9360 12552
rect 9280 12392 9360 12488
rect 9280 12328 9288 12392
rect 9352 12328 9360 12392
rect 9280 12232 9360 12328
rect 9280 12168 9288 12232
rect 9352 12168 9360 12232
rect 9280 12072 9360 12168
rect 9280 12008 9288 12072
rect 9352 12008 9360 12072
rect 9280 11912 9360 12008
rect 9280 11848 9288 11912
rect 9352 11848 9360 11912
rect 9280 11752 9360 11848
rect 9280 11688 9288 11752
rect 9352 11688 9360 11752
rect 9280 11592 9360 11688
rect 9280 11528 9288 11592
rect 9352 11528 9360 11592
rect 9280 11432 9360 11528
rect 9280 11368 9288 11432
rect 9352 11368 9360 11432
rect 9280 11272 9360 11368
rect 9280 11208 9288 11272
rect 9352 11208 9360 11272
rect 9280 11112 9360 11208
rect 9280 11048 9288 11112
rect 9352 11048 9360 11112
rect 9280 10952 9360 11048
rect 9280 10888 9288 10952
rect 9352 10888 9360 10952
rect 9280 10792 9360 10888
rect 9280 10728 9288 10792
rect 9352 10728 9360 10792
rect 9280 10632 9360 10728
rect 9280 10568 9288 10632
rect 9352 10568 9360 10632
rect 9280 10472 9360 10568
rect 9280 10408 9288 10472
rect 9352 10408 9360 10472
rect 9280 10312 9360 10408
rect 9280 10248 9288 10312
rect 9352 10248 9360 10312
rect 9280 10152 9360 10248
rect 9280 10088 9288 10152
rect 9352 10088 9360 10152
rect 9280 9992 9360 10088
rect 9280 9928 9288 9992
rect 9352 9928 9360 9992
rect 9280 9832 9360 9928
rect 9280 9768 9288 9832
rect 9352 9768 9360 9832
rect 9280 9672 9360 9768
rect 9280 9608 9288 9672
rect 9352 9608 9360 9672
rect 9280 9512 9360 9608
rect 9280 9448 9288 9512
rect 9352 9448 9360 9512
rect 9280 9352 9360 9448
rect 9280 9288 9288 9352
rect 9352 9288 9360 9352
rect 9280 9192 9360 9288
rect 9280 9128 9288 9192
rect 9352 9128 9360 9192
rect 9280 9032 9360 9128
rect 9280 8968 9288 9032
rect 9352 8968 9360 9032
rect 9280 8872 9360 8968
rect 9280 8808 9288 8872
rect 9352 8808 9360 8872
rect 9280 8712 9360 8808
rect 9280 8648 9288 8712
rect 9352 8648 9360 8712
rect 9280 8552 9360 8648
rect 9280 8488 9288 8552
rect 9352 8488 9360 8552
rect 9280 8392 9360 8488
rect 9280 8328 9288 8392
rect 9352 8328 9360 8392
rect 9280 8232 9360 8328
rect 9280 8168 9288 8232
rect 9352 8168 9360 8232
rect 9280 8072 9360 8168
rect 9280 8008 9288 8072
rect 9352 8008 9360 8072
rect 9280 7912 9360 8008
rect 9280 7848 9288 7912
rect 9352 7848 9360 7912
rect 9280 7752 9360 7848
rect 9280 7688 9288 7752
rect 9352 7688 9360 7752
rect 9280 7592 9360 7688
rect 9280 7528 9288 7592
rect 9352 7528 9360 7592
rect 9280 7432 9360 7528
rect 9280 7368 9288 7432
rect 9352 7368 9360 7432
rect 9280 7272 9360 7368
rect 9280 7208 9288 7272
rect 9352 7208 9360 7272
rect 9280 7112 9360 7208
rect 9280 7048 9288 7112
rect 9352 7048 9360 7112
rect 9280 6952 9360 7048
rect 9280 6888 9288 6952
rect 9352 6888 9360 6952
rect 9280 6792 9360 6888
rect 9280 6728 9288 6792
rect 9352 6728 9360 6792
rect 9280 6632 9360 6728
rect 9280 6568 9288 6632
rect 9352 6568 9360 6632
rect 9280 6472 9360 6568
rect 9280 6408 9288 6472
rect 9352 6408 9360 6472
rect 9280 6312 9360 6408
rect 9280 6248 9288 6312
rect 9352 6248 9360 6312
rect 9280 6152 9360 6248
rect 9280 6088 9288 6152
rect 9352 6088 9360 6152
rect 9280 5992 9360 6088
rect 9280 5928 9288 5992
rect 9352 5928 9360 5992
rect 9280 5832 9360 5928
rect 9280 5768 9288 5832
rect 9352 5768 9360 5832
rect 9280 5672 9360 5768
rect 9280 5608 9288 5672
rect 9352 5608 9360 5672
rect 9280 5512 9360 5608
rect 9280 5448 9288 5512
rect 9352 5448 9360 5512
rect 9280 5352 9360 5448
rect 9280 5288 9288 5352
rect 9352 5288 9360 5352
rect 9280 5192 9360 5288
rect 9280 5128 9288 5192
rect 9352 5128 9360 5192
rect 9280 5032 9360 5128
rect 9280 4968 9288 5032
rect 9352 4968 9360 5032
rect 9280 4872 9360 4968
rect 9280 4808 9288 4872
rect 9352 4808 9360 4872
rect 9280 4712 9360 4808
rect 9280 4648 9288 4712
rect 9352 4648 9360 4712
rect 9280 4552 9360 4648
rect 9280 4488 9288 4552
rect 9352 4488 9360 4552
rect 9280 4392 9360 4488
rect 9280 4328 9288 4392
rect 9352 4328 9360 4392
rect 9280 4232 9360 4328
rect 9280 4168 9288 4232
rect 9352 4168 9360 4232
rect 9280 4072 9360 4168
rect 9280 4008 9288 4072
rect 9352 4008 9360 4072
rect 9280 3912 9360 4008
rect 9280 3848 9288 3912
rect 9352 3848 9360 3912
rect 9280 3752 9360 3848
rect 9280 3688 9288 3752
rect 9352 3688 9360 3752
rect 9280 3592 9360 3688
rect 9280 3528 9288 3592
rect 9352 3528 9360 3592
rect 9280 3432 9360 3528
rect 9280 3368 9288 3432
rect 9352 3368 9360 3432
rect 9280 3272 9360 3368
rect 9280 3208 9288 3272
rect 9352 3208 9360 3272
rect 9280 3112 9360 3208
rect 9280 3048 9288 3112
rect 9352 3048 9360 3112
rect 9280 2952 9360 3048
rect 9280 2888 9288 2952
rect 9352 2888 9360 2952
rect 9280 2792 9360 2888
rect 9280 2728 9288 2792
rect 9352 2728 9360 2792
rect 9280 2632 9360 2728
rect 9280 2568 9288 2632
rect 9352 2568 9360 2632
rect 9280 2472 9360 2568
rect 9280 2408 9288 2472
rect 9352 2408 9360 2472
rect 9280 2312 9360 2408
rect 9280 2248 9288 2312
rect 9352 2248 9360 2312
rect 9280 2152 9360 2248
rect 9280 2088 9288 2152
rect 9352 2088 9360 2152
rect 9280 1992 9360 2088
rect 9280 1928 9288 1992
rect 9352 1928 9360 1992
rect 9280 1832 9360 1928
rect 9280 1768 9288 1832
rect 9352 1768 9360 1832
rect 9280 1672 9360 1768
rect 9280 1608 9288 1672
rect 9352 1608 9360 1672
rect 9280 1512 9360 1608
rect 9280 1448 9288 1512
rect 9352 1448 9360 1512
rect 9280 1352 9360 1448
rect 9280 1288 9288 1352
rect 9352 1288 9360 1352
rect 9280 1192 9360 1288
rect 9280 1128 9288 1192
rect 9352 1128 9360 1192
rect 9280 1032 9360 1128
rect 9280 968 9288 1032
rect 9352 968 9360 1032
rect 9280 872 9360 968
rect 9280 808 9288 872
rect 9352 808 9360 872
rect 9280 712 9360 808
rect 9280 648 9288 712
rect 9352 648 9360 712
rect 9280 552 9360 648
rect 9280 488 9288 552
rect 9352 488 9360 552
rect 9280 392 9360 488
rect 9280 328 9288 392
rect 9352 328 9360 392
rect 9280 232 9360 328
rect 9280 168 9288 232
rect 9352 168 9360 232
rect 9280 72 9360 168
rect 9280 8 9288 72
rect 9352 8 9360 72
rect 9280 -568 9360 8
rect 9280 -632 9288 -568
rect 9352 -632 9360 -568
rect 9280 -648 9360 -632
rect 9280 -712 9288 -648
rect 9352 -712 9360 -648
rect 9280 -728 9360 -712
rect 9280 -792 9288 -728
rect 9352 -792 9360 -728
rect 9280 -808 9360 -792
rect 9280 -872 9288 -808
rect 9352 -872 9360 -808
rect 9280 -888 9360 -872
rect 9280 -952 9288 -888
rect 9352 -952 9360 -888
rect 9280 -2008 9360 -952
rect 9440 31432 9520 31520
rect 9440 31368 9448 31432
rect 9512 31368 9520 31432
rect 9440 31272 9520 31368
rect 9440 31208 9448 31272
rect 9512 31208 9520 31272
rect 9440 31112 9520 31208
rect 9440 31048 9448 31112
rect 9512 31048 9520 31112
rect 9440 30952 9520 31048
rect 9440 30888 9448 30952
rect 9512 30888 9520 30952
rect 9440 30792 9520 30888
rect 9440 30728 9448 30792
rect 9512 30728 9520 30792
rect 9440 30632 9520 30728
rect 9440 30568 9448 30632
rect 9512 30568 9520 30632
rect 9440 30472 9520 30568
rect 9440 30408 9448 30472
rect 9512 30408 9520 30472
rect 9440 30312 9520 30408
rect 9440 30248 9448 30312
rect 9512 30248 9520 30312
rect 9440 30152 9520 30248
rect 9440 30088 9448 30152
rect 9512 30088 9520 30152
rect 9440 29992 9520 30088
rect 9440 29928 9448 29992
rect 9512 29928 9520 29992
rect 9440 29832 9520 29928
rect 9440 29768 9448 29832
rect 9512 29768 9520 29832
rect 9440 29672 9520 29768
rect 9440 29608 9448 29672
rect 9512 29608 9520 29672
rect 9440 29512 9520 29608
rect 9440 29448 9448 29512
rect 9512 29448 9520 29512
rect 9440 29352 9520 29448
rect 9440 29288 9448 29352
rect 9512 29288 9520 29352
rect 9440 29192 9520 29288
rect 9440 29128 9448 29192
rect 9512 29128 9520 29192
rect 9440 29032 9520 29128
rect 9440 28968 9448 29032
rect 9512 28968 9520 29032
rect 9440 28872 9520 28968
rect 9440 28808 9448 28872
rect 9512 28808 9520 28872
rect 9440 28712 9520 28808
rect 9440 28648 9448 28712
rect 9512 28648 9520 28712
rect 9440 28552 9520 28648
rect 9440 28488 9448 28552
rect 9512 28488 9520 28552
rect 9440 28392 9520 28488
rect 9440 28328 9448 28392
rect 9512 28328 9520 28392
rect 9440 28232 9520 28328
rect 9440 28168 9448 28232
rect 9512 28168 9520 28232
rect 9440 28072 9520 28168
rect 9440 28008 9448 28072
rect 9512 28008 9520 28072
rect 9440 27912 9520 28008
rect 9440 27848 9448 27912
rect 9512 27848 9520 27912
rect 9440 27752 9520 27848
rect 9440 27688 9448 27752
rect 9512 27688 9520 27752
rect 9440 27592 9520 27688
rect 9440 27528 9448 27592
rect 9512 27528 9520 27592
rect 9440 27432 9520 27528
rect 9440 27368 9448 27432
rect 9512 27368 9520 27432
rect 9440 27272 9520 27368
rect 9440 27208 9448 27272
rect 9512 27208 9520 27272
rect 9440 27112 9520 27208
rect 9440 27048 9448 27112
rect 9512 27048 9520 27112
rect 9440 26952 9520 27048
rect 9440 26888 9448 26952
rect 9512 26888 9520 26952
rect 9440 26792 9520 26888
rect 9440 26728 9448 26792
rect 9512 26728 9520 26792
rect 9440 26632 9520 26728
rect 9440 26568 9448 26632
rect 9512 26568 9520 26632
rect 9440 26472 9520 26568
rect 9440 26408 9448 26472
rect 9512 26408 9520 26472
rect 9440 26312 9520 26408
rect 9440 26248 9448 26312
rect 9512 26248 9520 26312
rect 9440 26152 9520 26248
rect 9440 26088 9448 26152
rect 9512 26088 9520 26152
rect 9440 25992 9520 26088
rect 9440 25928 9448 25992
rect 9512 25928 9520 25992
rect 9440 25832 9520 25928
rect 9440 25768 9448 25832
rect 9512 25768 9520 25832
rect 9440 25672 9520 25768
rect 9440 25608 9448 25672
rect 9512 25608 9520 25672
rect 9440 25512 9520 25608
rect 9440 25448 9448 25512
rect 9512 25448 9520 25512
rect 9440 25352 9520 25448
rect 9440 25288 9448 25352
rect 9512 25288 9520 25352
rect 9440 25192 9520 25288
rect 9440 25128 9448 25192
rect 9512 25128 9520 25192
rect 9440 25032 9520 25128
rect 9440 24968 9448 25032
rect 9512 24968 9520 25032
rect 9440 24872 9520 24968
rect 9440 24808 9448 24872
rect 9512 24808 9520 24872
rect 9440 24712 9520 24808
rect 9440 24648 9448 24712
rect 9512 24648 9520 24712
rect 9440 24552 9520 24648
rect 9440 24488 9448 24552
rect 9512 24488 9520 24552
rect 9440 24392 9520 24488
rect 9440 24328 9448 24392
rect 9512 24328 9520 24392
rect 9440 24232 9520 24328
rect 9440 24168 9448 24232
rect 9512 24168 9520 24232
rect 9440 24072 9520 24168
rect 9440 24008 9448 24072
rect 9512 24008 9520 24072
rect 9440 23912 9520 24008
rect 9440 23848 9448 23912
rect 9512 23848 9520 23912
rect 9440 23752 9520 23848
rect 9440 23688 9448 23752
rect 9512 23688 9520 23752
rect 9440 23592 9520 23688
rect 9440 23528 9448 23592
rect 9512 23528 9520 23592
rect 9440 23432 9520 23528
rect 9440 23368 9448 23432
rect 9512 23368 9520 23432
rect 9440 23272 9520 23368
rect 9440 23208 9448 23272
rect 9512 23208 9520 23272
rect 9440 23112 9520 23208
rect 9440 23048 9448 23112
rect 9512 23048 9520 23112
rect 9440 22952 9520 23048
rect 9440 22888 9448 22952
rect 9512 22888 9520 22952
rect 9440 22792 9520 22888
rect 9440 22728 9448 22792
rect 9512 22728 9520 22792
rect 9440 22632 9520 22728
rect 9440 22568 9448 22632
rect 9512 22568 9520 22632
rect 9440 22472 9520 22568
rect 9440 22408 9448 22472
rect 9512 22408 9520 22472
rect 9440 22312 9520 22408
rect 9440 22248 9448 22312
rect 9512 22248 9520 22312
rect 9440 22152 9520 22248
rect 9440 22088 9448 22152
rect 9512 22088 9520 22152
rect 9440 21992 9520 22088
rect 9440 21928 9448 21992
rect 9512 21928 9520 21992
rect 9440 21832 9520 21928
rect 9440 21768 9448 21832
rect 9512 21768 9520 21832
rect 9440 21672 9520 21768
rect 9440 21608 9448 21672
rect 9512 21608 9520 21672
rect 9440 21512 9520 21608
rect 9440 21448 9448 21512
rect 9512 21448 9520 21512
rect 9440 21352 9520 21448
rect 9440 21288 9448 21352
rect 9512 21288 9520 21352
rect 9440 21192 9520 21288
rect 9440 21128 9448 21192
rect 9512 21128 9520 21192
rect 9440 21032 9520 21128
rect 9440 20968 9448 21032
rect 9512 20968 9520 21032
rect 9440 20872 9520 20968
rect 9440 20808 9448 20872
rect 9512 20808 9520 20872
rect 9440 20712 9520 20808
rect 9440 20648 9448 20712
rect 9512 20648 9520 20712
rect 9440 20552 9520 20648
rect 9440 20488 9448 20552
rect 9512 20488 9520 20552
rect 9440 20392 9520 20488
rect 9440 20328 9448 20392
rect 9512 20328 9520 20392
rect 9440 20232 9520 20328
rect 9440 20168 9448 20232
rect 9512 20168 9520 20232
rect 9440 20072 9520 20168
rect 9440 20008 9448 20072
rect 9512 20008 9520 20072
rect 9440 19912 9520 20008
rect 9440 19848 9448 19912
rect 9512 19848 9520 19912
rect 9440 19752 9520 19848
rect 9440 19688 9448 19752
rect 9512 19688 9520 19752
rect 9440 19592 9520 19688
rect 9440 19528 9448 19592
rect 9512 19528 9520 19592
rect 9440 19432 9520 19528
rect 9440 19368 9448 19432
rect 9512 19368 9520 19432
rect 9440 19272 9520 19368
rect 9440 19208 9448 19272
rect 9512 19208 9520 19272
rect 9440 19112 9520 19208
rect 9440 19048 9448 19112
rect 9512 19048 9520 19112
rect 9440 18952 9520 19048
rect 9440 18888 9448 18952
rect 9512 18888 9520 18952
rect 9440 18792 9520 18888
rect 9440 18728 9448 18792
rect 9512 18728 9520 18792
rect 9440 18632 9520 18728
rect 9440 18568 9448 18632
rect 9512 18568 9520 18632
rect 9440 18472 9520 18568
rect 9440 18408 9448 18472
rect 9512 18408 9520 18472
rect 9440 18312 9520 18408
rect 9440 18248 9448 18312
rect 9512 18248 9520 18312
rect 9440 18152 9520 18248
rect 9440 18088 9448 18152
rect 9512 18088 9520 18152
rect 9440 17992 9520 18088
rect 9440 17928 9448 17992
rect 9512 17928 9520 17992
rect 9440 17832 9520 17928
rect 9440 17768 9448 17832
rect 9512 17768 9520 17832
rect 9440 17672 9520 17768
rect 9440 17608 9448 17672
rect 9512 17608 9520 17672
rect 9440 17512 9520 17608
rect 9440 17448 9448 17512
rect 9512 17448 9520 17512
rect 9440 17352 9520 17448
rect 9440 17288 9448 17352
rect 9512 17288 9520 17352
rect 9440 17192 9520 17288
rect 9440 17128 9448 17192
rect 9512 17128 9520 17192
rect 9440 17032 9520 17128
rect 9440 16968 9448 17032
rect 9512 16968 9520 17032
rect 9440 16872 9520 16968
rect 9440 16808 9448 16872
rect 9512 16808 9520 16872
rect 9440 16712 9520 16808
rect 9440 16648 9448 16712
rect 9512 16648 9520 16712
rect 9440 16552 9520 16648
rect 9440 16488 9448 16552
rect 9512 16488 9520 16552
rect 9440 16392 9520 16488
rect 9440 16328 9448 16392
rect 9512 16328 9520 16392
rect 9440 16232 9520 16328
rect 9440 16168 9448 16232
rect 9512 16168 9520 16232
rect 9440 16072 9520 16168
rect 9440 16008 9448 16072
rect 9512 16008 9520 16072
rect 9440 15912 9520 16008
rect 9440 15848 9448 15912
rect 9512 15848 9520 15912
rect 9440 15752 9520 15848
rect 9440 15688 9448 15752
rect 9512 15688 9520 15752
rect 9440 15592 9520 15688
rect 9440 15528 9448 15592
rect 9512 15528 9520 15592
rect 9440 15432 9520 15528
rect 9440 15368 9448 15432
rect 9512 15368 9520 15432
rect 9440 15272 9520 15368
rect 9440 15208 9448 15272
rect 9512 15208 9520 15272
rect 9440 15112 9520 15208
rect 9440 15048 9448 15112
rect 9512 15048 9520 15112
rect 9440 14952 9520 15048
rect 9440 14888 9448 14952
rect 9512 14888 9520 14952
rect 9440 14792 9520 14888
rect 9440 14728 9448 14792
rect 9512 14728 9520 14792
rect 9440 14632 9520 14728
rect 9440 14568 9448 14632
rect 9512 14568 9520 14632
rect 9440 14472 9520 14568
rect 9440 14408 9448 14472
rect 9512 14408 9520 14472
rect 9440 14312 9520 14408
rect 9440 14248 9448 14312
rect 9512 14248 9520 14312
rect 9440 14152 9520 14248
rect 9440 14088 9448 14152
rect 9512 14088 9520 14152
rect 9440 13992 9520 14088
rect 9440 13928 9448 13992
rect 9512 13928 9520 13992
rect 9440 13832 9520 13928
rect 9440 13768 9448 13832
rect 9512 13768 9520 13832
rect 9440 13672 9520 13768
rect 9440 13608 9448 13672
rect 9512 13608 9520 13672
rect 9440 13512 9520 13608
rect 9440 13448 9448 13512
rect 9512 13448 9520 13512
rect 9440 13352 9520 13448
rect 9440 13288 9448 13352
rect 9512 13288 9520 13352
rect 9440 13192 9520 13288
rect 9440 13128 9448 13192
rect 9512 13128 9520 13192
rect 9440 13032 9520 13128
rect 9440 12968 9448 13032
rect 9512 12968 9520 13032
rect 9440 12872 9520 12968
rect 9440 12808 9448 12872
rect 9512 12808 9520 12872
rect 9440 12712 9520 12808
rect 9440 12648 9448 12712
rect 9512 12648 9520 12712
rect 9440 12552 9520 12648
rect 9440 12488 9448 12552
rect 9512 12488 9520 12552
rect 9440 12392 9520 12488
rect 9440 12328 9448 12392
rect 9512 12328 9520 12392
rect 9440 12232 9520 12328
rect 9440 12168 9448 12232
rect 9512 12168 9520 12232
rect 9440 12072 9520 12168
rect 9440 12008 9448 12072
rect 9512 12008 9520 12072
rect 9440 11912 9520 12008
rect 9440 11848 9448 11912
rect 9512 11848 9520 11912
rect 9440 11752 9520 11848
rect 9440 11688 9448 11752
rect 9512 11688 9520 11752
rect 9440 11592 9520 11688
rect 9440 11528 9448 11592
rect 9512 11528 9520 11592
rect 9440 11432 9520 11528
rect 9440 11368 9448 11432
rect 9512 11368 9520 11432
rect 9440 11272 9520 11368
rect 9440 11208 9448 11272
rect 9512 11208 9520 11272
rect 9440 11112 9520 11208
rect 9440 11048 9448 11112
rect 9512 11048 9520 11112
rect 9440 10952 9520 11048
rect 9440 10888 9448 10952
rect 9512 10888 9520 10952
rect 9440 10792 9520 10888
rect 9440 10728 9448 10792
rect 9512 10728 9520 10792
rect 9440 10632 9520 10728
rect 9440 10568 9448 10632
rect 9512 10568 9520 10632
rect 9440 10472 9520 10568
rect 9440 10408 9448 10472
rect 9512 10408 9520 10472
rect 9440 10312 9520 10408
rect 9440 10248 9448 10312
rect 9512 10248 9520 10312
rect 9440 10152 9520 10248
rect 9440 10088 9448 10152
rect 9512 10088 9520 10152
rect 9440 9992 9520 10088
rect 9440 9928 9448 9992
rect 9512 9928 9520 9992
rect 9440 9832 9520 9928
rect 9440 9768 9448 9832
rect 9512 9768 9520 9832
rect 9440 9672 9520 9768
rect 9440 9608 9448 9672
rect 9512 9608 9520 9672
rect 9440 9512 9520 9608
rect 9440 9448 9448 9512
rect 9512 9448 9520 9512
rect 9440 9352 9520 9448
rect 9440 9288 9448 9352
rect 9512 9288 9520 9352
rect 9440 9192 9520 9288
rect 9440 9128 9448 9192
rect 9512 9128 9520 9192
rect 9440 9032 9520 9128
rect 9440 8968 9448 9032
rect 9512 8968 9520 9032
rect 9440 8872 9520 8968
rect 9440 8808 9448 8872
rect 9512 8808 9520 8872
rect 9440 8712 9520 8808
rect 9440 8648 9448 8712
rect 9512 8648 9520 8712
rect 9440 8552 9520 8648
rect 9440 8488 9448 8552
rect 9512 8488 9520 8552
rect 9440 8392 9520 8488
rect 9440 8328 9448 8392
rect 9512 8328 9520 8392
rect 9440 8232 9520 8328
rect 9440 8168 9448 8232
rect 9512 8168 9520 8232
rect 9440 8072 9520 8168
rect 9440 8008 9448 8072
rect 9512 8008 9520 8072
rect 9440 7912 9520 8008
rect 9440 7848 9448 7912
rect 9512 7848 9520 7912
rect 9440 7752 9520 7848
rect 9440 7688 9448 7752
rect 9512 7688 9520 7752
rect 9440 7592 9520 7688
rect 9440 7528 9448 7592
rect 9512 7528 9520 7592
rect 9440 7432 9520 7528
rect 9440 7368 9448 7432
rect 9512 7368 9520 7432
rect 9440 7272 9520 7368
rect 9440 7208 9448 7272
rect 9512 7208 9520 7272
rect 9440 7112 9520 7208
rect 9440 7048 9448 7112
rect 9512 7048 9520 7112
rect 9440 6952 9520 7048
rect 9440 6888 9448 6952
rect 9512 6888 9520 6952
rect 9440 6792 9520 6888
rect 9440 6728 9448 6792
rect 9512 6728 9520 6792
rect 9440 6632 9520 6728
rect 9440 6568 9448 6632
rect 9512 6568 9520 6632
rect 9440 6472 9520 6568
rect 9440 6408 9448 6472
rect 9512 6408 9520 6472
rect 9440 6312 9520 6408
rect 9440 6248 9448 6312
rect 9512 6248 9520 6312
rect 9440 6152 9520 6248
rect 9440 6088 9448 6152
rect 9512 6088 9520 6152
rect 9440 5992 9520 6088
rect 9440 5928 9448 5992
rect 9512 5928 9520 5992
rect 9440 5832 9520 5928
rect 9440 5768 9448 5832
rect 9512 5768 9520 5832
rect 9440 5672 9520 5768
rect 9440 5608 9448 5672
rect 9512 5608 9520 5672
rect 9440 5512 9520 5608
rect 9440 5448 9448 5512
rect 9512 5448 9520 5512
rect 9440 5352 9520 5448
rect 9440 5288 9448 5352
rect 9512 5288 9520 5352
rect 9440 5192 9520 5288
rect 9440 5128 9448 5192
rect 9512 5128 9520 5192
rect 9440 5032 9520 5128
rect 9440 4968 9448 5032
rect 9512 4968 9520 5032
rect 9440 4872 9520 4968
rect 9440 4808 9448 4872
rect 9512 4808 9520 4872
rect 9440 4712 9520 4808
rect 9440 4648 9448 4712
rect 9512 4648 9520 4712
rect 9440 4552 9520 4648
rect 9440 4488 9448 4552
rect 9512 4488 9520 4552
rect 9440 4392 9520 4488
rect 9440 4328 9448 4392
rect 9512 4328 9520 4392
rect 9440 4232 9520 4328
rect 9440 4168 9448 4232
rect 9512 4168 9520 4232
rect 9440 4072 9520 4168
rect 9440 4008 9448 4072
rect 9512 4008 9520 4072
rect 9440 3912 9520 4008
rect 9440 3848 9448 3912
rect 9512 3848 9520 3912
rect 9440 3752 9520 3848
rect 9440 3688 9448 3752
rect 9512 3688 9520 3752
rect 9440 3592 9520 3688
rect 9440 3528 9448 3592
rect 9512 3528 9520 3592
rect 9440 3432 9520 3528
rect 9440 3368 9448 3432
rect 9512 3368 9520 3432
rect 9440 3272 9520 3368
rect 9440 3208 9448 3272
rect 9512 3208 9520 3272
rect 9440 3112 9520 3208
rect 9440 3048 9448 3112
rect 9512 3048 9520 3112
rect 9440 2952 9520 3048
rect 9440 2888 9448 2952
rect 9512 2888 9520 2952
rect 9440 2792 9520 2888
rect 9440 2728 9448 2792
rect 9512 2728 9520 2792
rect 9440 2632 9520 2728
rect 9440 2568 9448 2632
rect 9512 2568 9520 2632
rect 9440 2472 9520 2568
rect 9440 2408 9448 2472
rect 9512 2408 9520 2472
rect 9440 2312 9520 2408
rect 9440 2248 9448 2312
rect 9512 2248 9520 2312
rect 9440 2152 9520 2248
rect 9440 2088 9448 2152
rect 9512 2088 9520 2152
rect 9440 1992 9520 2088
rect 9440 1928 9448 1992
rect 9512 1928 9520 1992
rect 9440 1832 9520 1928
rect 9440 1768 9448 1832
rect 9512 1768 9520 1832
rect 9440 1672 9520 1768
rect 9440 1608 9448 1672
rect 9512 1608 9520 1672
rect 9440 1512 9520 1608
rect 9440 1448 9448 1512
rect 9512 1448 9520 1512
rect 9440 1352 9520 1448
rect 9440 1288 9448 1352
rect 9512 1288 9520 1352
rect 9440 1192 9520 1288
rect 9440 1128 9448 1192
rect 9512 1128 9520 1192
rect 9440 1032 9520 1128
rect 9440 968 9448 1032
rect 9512 968 9520 1032
rect 9440 872 9520 968
rect 9440 808 9448 872
rect 9512 808 9520 872
rect 9440 712 9520 808
rect 9440 648 9448 712
rect 9512 648 9520 712
rect 9440 552 9520 648
rect 9440 488 9448 552
rect 9512 488 9520 552
rect 9440 392 9520 488
rect 9440 328 9448 392
rect 9512 328 9520 392
rect 9440 232 9520 328
rect 9440 168 9448 232
rect 9512 168 9520 232
rect 9440 72 9520 168
rect 9440 8 9448 72
rect 9512 8 9520 72
rect 9440 -1048 9520 8
rect 9600 12308 9680 31520
rect 9600 12252 9612 12308
rect 9668 12252 9680 12308
rect 9600 0 9680 12252
rect 9760 31432 9840 31520
rect 9760 31368 9768 31432
rect 9832 31368 9840 31432
rect 9760 31272 9840 31368
rect 9760 31208 9768 31272
rect 9832 31208 9840 31272
rect 9760 31112 9840 31208
rect 9760 31048 9768 31112
rect 9832 31048 9840 31112
rect 9760 30952 9840 31048
rect 9760 30888 9768 30952
rect 9832 30888 9840 30952
rect 9760 30792 9840 30888
rect 9760 30728 9768 30792
rect 9832 30728 9840 30792
rect 9760 30632 9840 30728
rect 9760 30568 9768 30632
rect 9832 30568 9840 30632
rect 9760 30472 9840 30568
rect 9760 30408 9768 30472
rect 9832 30408 9840 30472
rect 9760 30312 9840 30408
rect 9760 30248 9768 30312
rect 9832 30248 9840 30312
rect 9760 30152 9840 30248
rect 9760 30088 9768 30152
rect 9832 30088 9840 30152
rect 9760 29992 9840 30088
rect 9760 29928 9768 29992
rect 9832 29928 9840 29992
rect 9760 29832 9840 29928
rect 9760 29768 9768 29832
rect 9832 29768 9840 29832
rect 9760 29672 9840 29768
rect 9760 29608 9768 29672
rect 9832 29608 9840 29672
rect 9760 29512 9840 29608
rect 9760 29448 9768 29512
rect 9832 29448 9840 29512
rect 9760 29352 9840 29448
rect 9760 29288 9768 29352
rect 9832 29288 9840 29352
rect 9760 29192 9840 29288
rect 9760 29128 9768 29192
rect 9832 29128 9840 29192
rect 9760 29032 9840 29128
rect 9760 28968 9768 29032
rect 9832 28968 9840 29032
rect 9760 28872 9840 28968
rect 9760 28808 9768 28872
rect 9832 28808 9840 28872
rect 9760 28712 9840 28808
rect 9760 28648 9768 28712
rect 9832 28648 9840 28712
rect 9760 28552 9840 28648
rect 9760 28488 9768 28552
rect 9832 28488 9840 28552
rect 9760 28392 9840 28488
rect 9760 28328 9768 28392
rect 9832 28328 9840 28392
rect 9760 28232 9840 28328
rect 9760 28168 9768 28232
rect 9832 28168 9840 28232
rect 9760 28072 9840 28168
rect 9760 28008 9768 28072
rect 9832 28008 9840 28072
rect 9760 27912 9840 28008
rect 9760 27848 9768 27912
rect 9832 27848 9840 27912
rect 9760 27752 9840 27848
rect 9760 27688 9768 27752
rect 9832 27688 9840 27752
rect 9760 27592 9840 27688
rect 9760 27528 9768 27592
rect 9832 27528 9840 27592
rect 9760 27432 9840 27528
rect 9760 27368 9768 27432
rect 9832 27368 9840 27432
rect 9760 27272 9840 27368
rect 9760 27208 9768 27272
rect 9832 27208 9840 27272
rect 9760 27112 9840 27208
rect 9760 27048 9768 27112
rect 9832 27048 9840 27112
rect 9760 26952 9840 27048
rect 9760 26888 9768 26952
rect 9832 26888 9840 26952
rect 9760 26792 9840 26888
rect 9760 26728 9768 26792
rect 9832 26728 9840 26792
rect 9760 26632 9840 26728
rect 9760 26568 9768 26632
rect 9832 26568 9840 26632
rect 9760 26472 9840 26568
rect 9760 26408 9768 26472
rect 9832 26408 9840 26472
rect 9760 26312 9840 26408
rect 9760 26248 9768 26312
rect 9832 26248 9840 26312
rect 9760 26152 9840 26248
rect 9760 26088 9768 26152
rect 9832 26088 9840 26152
rect 9760 25992 9840 26088
rect 9760 25928 9768 25992
rect 9832 25928 9840 25992
rect 9760 25832 9840 25928
rect 9760 25768 9768 25832
rect 9832 25768 9840 25832
rect 9760 25672 9840 25768
rect 9760 25608 9768 25672
rect 9832 25608 9840 25672
rect 9760 25512 9840 25608
rect 9760 25448 9768 25512
rect 9832 25448 9840 25512
rect 9760 25352 9840 25448
rect 9760 25288 9768 25352
rect 9832 25288 9840 25352
rect 9760 25192 9840 25288
rect 9760 25128 9768 25192
rect 9832 25128 9840 25192
rect 9760 25032 9840 25128
rect 9760 24968 9768 25032
rect 9832 24968 9840 25032
rect 9760 24872 9840 24968
rect 9760 24808 9768 24872
rect 9832 24808 9840 24872
rect 9760 24712 9840 24808
rect 9760 24648 9768 24712
rect 9832 24648 9840 24712
rect 9760 24552 9840 24648
rect 9760 24488 9768 24552
rect 9832 24488 9840 24552
rect 9760 24392 9840 24488
rect 9760 24328 9768 24392
rect 9832 24328 9840 24392
rect 9760 24232 9840 24328
rect 9760 24168 9768 24232
rect 9832 24168 9840 24232
rect 9760 24072 9840 24168
rect 9760 24008 9768 24072
rect 9832 24008 9840 24072
rect 9760 23912 9840 24008
rect 9760 23848 9768 23912
rect 9832 23848 9840 23912
rect 9760 23752 9840 23848
rect 9760 23688 9768 23752
rect 9832 23688 9840 23752
rect 9760 23592 9840 23688
rect 9760 23528 9768 23592
rect 9832 23528 9840 23592
rect 9760 23432 9840 23528
rect 9760 23368 9768 23432
rect 9832 23368 9840 23432
rect 9760 23272 9840 23368
rect 9760 23208 9768 23272
rect 9832 23208 9840 23272
rect 9760 23112 9840 23208
rect 9760 23048 9768 23112
rect 9832 23048 9840 23112
rect 9760 22952 9840 23048
rect 9760 22888 9768 22952
rect 9832 22888 9840 22952
rect 9760 22792 9840 22888
rect 9760 22728 9768 22792
rect 9832 22728 9840 22792
rect 9760 22632 9840 22728
rect 9760 22568 9768 22632
rect 9832 22568 9840 22632
rect 9760 22472 9840 22568
rect 9760 22408 9768 22472
rect 9832 22408 9840 22472
rect 9760 22312 9840 22408
rect 9760 22248 9768 22312
rect 9832 22248 9840 22312
rect 9760 22152 9840 22248
rect 9760 22088 9768 22152
rect 9832 22088 9840 22152
rect 9760 21992 9840 22088
rect 9760 21928 9768 21992
rect 9832 21928 9840 21992
rect 9760 21832 9840 21928
rect 9760 21768 9768 21832
rect 9832 21768 9840 21832
rect 9760 21672 9840 21768
rect 9760 21608 9768 21672
rect 9832 21608 9840 21672
rect 9760 21512 9840 21608
rect 9760 21448 9768 21512
rect 9832 21448 9840 21512
rect 9760 21352 9840 21448
rect 9760 21288 9768 21352
rect 9832 21288 9840 21352
rect 9760 21192 9840 21288
rect 9760 21128 9768 21192
rect 9832 21128 9840 21192
rect 9760 21032 9840 21128
rect 9760 20968 9768 21032
rect 9832 20968 9840 21032
rect 9760 20872 9840 20968
rect 9760 20808 9768 20872
rect 9832 20808 9840 20872
rect 9760 20712 9840 20808
rect 9760 20648 9768 20712
rect 9832 20648 9840 20712
rect 9760 20552 9840 20648
rect 9760 20488 9768 20552
rect 9832 20488 9840 20552
rect 9760 20392 9840 20488
rect 9760 20328 9768 20392
rect 9832 20328 9840 20392
rect 9760 20232 9840 20328
rect 9760 20168 9768 20232
rect 9832 20168 9840 20232
rect 9760 20072 9840 20168
rect 9760 20008 9768 20072
rect 9832 20008 9840 20072
rect 9760 19912 9840 20008
rect 9760 19848 9768 19912
rect 9832 19848 9840 19912
rect 9760 19752 9840 19848
rect 9760 19688 9768 19752
rect 9832 19688 9840 19752
rect 9760 19592 9840 19688
rect 9760 19528 9768 19592
rect 9832 19528 9840 19592
rect 9760 19432 9840 19528
rect 9760 19368 9768 19432
rect 9832 19368 9840 19432
rect 9760 19272 9840 19368
rect 9760 19208 9768 19272
rect 9832 19208 9840 19272
rect 9760 19112 9840 19208
rect 9760 19048 9768 19112
rect 9832 19048 9840 19112
rect 9760 18952 9840 19048
rect 9760 18888 9768 18952
rect 9832 18888 9840 18952
rect 9760 18792 9840 18888
rect 9760 18728 9768 18792
rect 9832 18728 9840 18792
rect 9760 18632 9840 18728
rect 9760 18568 9768 18632
rect 9832 18568 9840 18632
rect 9760 18472 9840 18568
rect 9760 18408 9768 18472
rect 9832 18408 9840 18472
rect 9760 18312 9840 18408
rect 9760 18248 9768 18312
rect 9832 18248 9840 18312
rect 9760 18152 9840 18248
rect 9760 18088 9768 18152
rect 9832 18088 9840 18152
rect 9760 17992 9840 18088
rect 9760 17928 9768 17992
rect 9832 17928 9840 17992
rect 9760 17832 9840 17928
rect 9760 17768 9768 17832
rect 9832 17768 9840 17832
rect 9760 17672 9840 17768
rect 9760 17608 9768 17672
rect 9832 17608 9840 17672
rect 9760 17512 9840 17608
rect 9760 17448 9768 17512
rect 9832 17448 9840 17512
rect 9760 17352 9840 17448
rect 9760 17288 9768 17352
rect 9832 17288 9840 17352
rect 9760 17192 9840 17288
rect 9760 17128 9768 17192
rect 9832 17128 9840 17192
rect 9760 17032 9840 17128
rect 9760 16968 9768 17032
rect 9832 16968 9840 17032
rect 9760 16872 9840 16968
rect 9760 16808 9768 16872
rect 9832 16808 9840 16872
rect 9760 16712 9840 16808
rect 9760 16648 9768 16712
rect 9832 16648 9840 16712
rect 9760 16552 9840 16648
rect 9760 16488 9768 16552
rect 9832 16488 9840 16552
rect 9760 16392 9840 16488
rect 9760 16328 9768 16392
rect 9832 16328 9840 16392
rect 9760 16232 9840 16328
rect 9760 16168 9768 16232
rect 9832 16168 9840 16232
rect 9760 16072 9840 16168
rect 9760 16008 9768 16072
rect 9832 16008 9840 16072
rect 9760 15912 9840 16008
rect 9760 15848 9768 15912
rect 9832 15848 9840 15912
rect 9760 15752 9840 15848
rect 9760 15688 9768 15752
rect 9832 15688 9840 15752
rect 9760 15592 9840 15688
rect 9760 15528 9768 15592
rect 9832 15528 9840 15592
rect 9760 15432 9840 15528
rect 9760 15368 9768 15432
rect 9832 15368 9840 15432
rect 9760 15272 9840 15368
rect 9760 15208 9768 15272
rect 9832 15208 9840 15272
rect 9760 15112 9840 15208
rect 9760 15048 9768 15112
rect 9832 15048 9840 15112
rect 9760 14952 9840 15048
rect 9760 14888 9768 14952
rect 9832 14888 9840 14952
rect 9760 14792 9840 14888
rect 9760 14728 9768 14792
rect 9832 14728 9840 14792
rect 9760 14632 9840 14728
rect 9760 14568 9768 14632
rect 9832 14568 9840 14632
rect 9760 14472 9840 14568
rect 9760 14408 9768 14472
rect 9832 14408 9840 14472
rect 9760 14312 9840 14408
rect 9760 14248 9768 14312
rect 9832 14248 9840 14312
rect 9760 14152 9840 14248
rect 9760 14088 9768 14152
rect 9832 14088 9840 14152
rect 9760 13992 9840 14088
rect 9760 13928 9768 13992
rect 9832 13928 9840 13992
rect 9760 13832 9840 13928
rect 9760 13768 9768 13832
rect 9832 13768 9840 13832
rect 9760 13672 9840 13768
rect 9760 13608 9768 13672
rect 9832 13608 9840 13672
rect 9760 13512 9840 13608
rect 9760 13448 9768 13512
rect 9832 13448 9840 13512
rect 9760 13352 9840 13448
rect 9760 13288 9768 13352
rect 9832 13288 9840 13352
rect 9760 13192 9840 13288
rect 9760 13128 9768 13192
rect 9832 13128 9840 13192
rect 9760 13032 9840 13128
rect 9760 12968 9768 13032
rect 9832 12968 9840 13032
rect 9760 12872 9840 12968
rect 9760 12808 9768 12872
rect 9832 12808 9840 12872
rect 9760 12712 9840 12808
rect 9760 12648 9768 12712
rect 9832 12648 9840 12712
rect 9760 12552 9840 12648
rect 9760 12488 9768 12552
rect 9832 12488 9840 12552
rect 9760 12392 9840 12488
rect 9760 12328 9768 12392
rect 9832 12328 9840 12392
rect 9760 12232 9840 12328
rect 9760 12168 9768 12232
rect 9832 12168 9840 12232
rect 9760 12072 9840 12168
rect 9760 12008 9768 12072
rect 9832 12008 9840 12072
rect 9760 11912 9840 12008
rect 9760 11848 9768 11912
rect 9832 11848 9840 11912
rect 9760 11752 9840 11848
rect 9760 11688 9768 11752
rect 9832 11688 9840 11752
rect 9760 11592 9840 11688
rect 9760 11528 9768 11592
rect 9832 11528 9840 11592
rect 9760 11432 9840 11528
rect 9760 11368 9768 11432
rect 9832 11368 9840 11432
rect 9760 11272 9840 11368
rect 9760 11208 9768 11272
rect 9832 11208 9840 11272
rect 9760 11112 9840 11208
rect 9760 11048 9768 11112
rect 9832 11048 9840 11112
rect 9760 10952 9840 11048
rect 9760 10888 9768 10952
rect 9832 10888 9840 10952
rect 9760 10792 9840 10888
rect 9760 10728 9768 10792
rect 9832 10728 9840 10792
rect 9760 10632 9840 10728
rect 9760 10568 9768 10632
rect 9832 10568 9840 10632
rect 9760 10472 9840 10568
rect 9760 10408 9768 10472
rect 9832 10408 9840 10472
rect 9760 10312 9840 10408
rect 9760 10248 9768 10312
rect 9832 10248 9840 10312
rect 9760 10152 9840 10248
rect 9760 10088 9768 10152
rect 9832 10088 9840 10152
rect 9760 9992 9840 10088
rect 9760 9928 9768 9992
rect 9832 9928 9840 9992
rect 9760 9832 9840 9928
rect 9760 9768 9768 9832
rect 9832 9768 9840 9832
rect 9760 9672 9840 9768
rect 9760 9608 9768 9672
rect 9832 9608 9840 9672
rect 9760 9512 9840 9608
rect 9760 9448 9768 9512
rect 9832 9448 9840 9512
rect 9760 9352 9840 9448
rect 9760 9288 9768 9352
rect 9832 9288 9840 9352
rect 9760 9192 9840 9288
rect 9760 9128 9768 9192
rect 9832 9128 9840 9192
rect 9760 9032 9840 9128
rect 9760 8968 9768 9032
rect 9832 8968 9840 9032
rect 9760 8872 9840 8968
rect 9760 8808 9768 8872
rect 9832 8808 9840 8872
rect 9760 8712 9840 8808
rect 9760 8648 9768 8712
rect 9832 8648 9840 8712
rect 9760 8552 9840 8648
rect 9760 8488 9768 8552
rect 9832 8488 9840 8552
rect 9760 8392 9840 8488
rect 9760 8328 9768 8392
rect 9832 8328 9840 8392
rect 9760 8232 9840 8328
rect 9760 8168 9768 8232
rect 9832 8168 9840 8232
rect 9760 8072 9840 8168
rect 9760 8008 9768 8072
rect 9832 8008 9840 8072
rect 9760 7912 9840 8008
rect 9760 7848 9768 7912
rect 9832 7848 9840 7912
rect 9760 7752 9840 7848
rect 9760 7688 9768 7752
rect 9832 7688 9840 7752
rect 9760 7592 9840 7688
rect 9760 7528 9768 7592
rect 9832 7528 9840 7592
rect 9760 7432 9840 7528
rect 9760 7368 9768 7432
rect 9832 7368 9840 7432
rect 9760 7272 9840 7368
rect 9760 7208 9768 7272
rect 9832 7208 9840 7272
rect 9760 7112 9840 7208
rect 9760 7048 9768 7112
rect 9832 7048 9840 7112
rect 9760 6952 9840 7048
rect 9760 6888 9768 6952
rect 9832 6888 9840 6952
rect 9760 6792 9840 6888
rect 9760 6728 9768 6792
rect 9832 6728 9840 6792
rect 9760 6632 9840 6728
rect 9760 6568 9768 6632
rect 9832 6568 9840 6632
rect 9760 6472 9840 6568
rect 9760 6408 9768 6472
rect 9832 6408 9840 6472
rect 9760 6312 9840 6408
rect 9760 6248 9768 6312
rect 9832 6248 9840 6312
rect 9760 6152 9840 6248
rect 9760 6088 9768 6152
rect 9832 6088 9840 6152
rect 9760 5992 9840 6088
rect 9760 5928 9768 5992
rect 9832 5928 9840 5992
rect 9760 5832 9840 5928
rect 9760 5768 9768 5832
rect 9832 5768 9840 5832
rect 9760 5672 9840 5768
rect 9760 5608 9768 5672
rect 9832 5608 9840 5672
rect 9760 5512 9840 5608
rect 9760 5448 9768 5512
rect 9832 5448 9840 5512
rect 9760 5352 9840 5448
rect 9760 5288 9768 5352
rect 9832 5288 9840 5352
rect 9760 5192 9840 5288
rect 9760 5128 9768 5192
rect 9832 5128 9840 5192
rect 9760 5032 9840 5128
rect 9760 4968 9768 5032
rect 9832 4968 9840 5032
rect 9760 4872 9840 4968
rect 9760 4808 9768 4872
rect 9832 4808 9840 4872
rect 9760 4712 9840 4808
rect 9760 4648 9768 4712
rect 9832 4648 9840 4712
rect 9760 4552 9840 4648
rect 9760 4488 9768 4552
rect 9832 4488 9840 4552
rect 9760 4392 9840 4488
rect 9760 4328 9768 4392
rect 9832 4328 9840 4392
rect 9760 4232 9840 4328
rect 9760 4168 9768 4232
rect 9832 4168 9840 4232
rect 9760 4072 9840 4168
rect 9760 4008 9768 4072
rect 9832 4008 9840 4072
rect 9760 3912 9840 4008
rect 9760 3848 9768 3912
rect 9832 3848 9840 3912
rect 9760 3752 9840 3848
rect 9760 3688 9768 3752
rect 9832 3688 9840 3752
rect 9760 3592 9840 3688
rect 9760 3528 9768 3592
rect 9832 3528 9840 3592
rect 9760 3432 9840 3528
rect 9760 3368 9768 3432
rect 9832 3368 9840 3432
rect 9760 3272 9840 3368
rect 9760 3208 9768 3272
rect 9832 3208 9840 3272
rect 9760 3112 9840 3208
rect 9760 3048 9768 3112
rect 9832 3048 9840 3112
rect 9760 2952 9840 3048
rect 9760 2888 9768 2952
rect 9832 2888 9840 2952
rect 9760 2792 9840 2888
rect 9760 2728 9768 2792
rect 9832 2728 9840 2792
rect 9760 2632 9840 2728
rect 9760 2568 9768 2632
rect 9832 2568 9840 2632
rect 9760 2472 9840 2568
rect 9760 2408 9768 2472
rect 9832 2408 9840 2472
rect 9760 2312 9840 2408
rect 9760 2248 9768 2312
rect 9832 2248 9840 2312
rect 9760 2152 9840 2248
rect 9760 2088 9768 2152
rect 9832 2088 9840 2152
rect 9760 1992 9840 2088
rect 9760 1928 9768 1992
rect 9832 1928 9840 1992
rect 9760 1832 9840 1928
rect 9760 1768 9768 1832
rect 9832 1768 9840 1832
rect 9760 1672 9840 1768
rect 9760 1608 9768 1672
rect 9832 1608 9840 1672
rect 9760 1512 9840 1608
rect 9760 1448 9768 1512
rect 9832 1448 9840 1512
rect 9760 1352 9840 1448
rect 9760 1288 9768 1352
rect 9832 1288 9840 1352
rect 9760 1192 9840 1288
rect 9760 1128 9768 1192
rect 9832 1128 9840 1192
rect 9760 1032 9840 1128
rect 9760 968 9768 1032
rect 9832 968 9840 1032
rect 9760 872 9840 968
rect 9760 808 9768 872
rect 9832 808 9840 872
rect 9760 712 9840 808
rect 9760 648 9768 712
rect 9832 648 9840 712
rect 9760 552 9840 648
rect 9760 488 9768 552
rect 9832 488 9840 552
rect 9760 392 9840 488
rect 9760 328 9768 392
rect 9832 328 9840 392
rect 9760 232 9840 328
rect 9760 168 9768 232
rect 9832 168 9840 232
rect 9760 72 9840 168
rect 9760 8 9768 72
rect 9832 8 9840 72
rect 9440 -1112 9448 -1048
rect 9512 -1112 9520 -1048
rect 9440 -1128 9520 -1112
rect 9440 -1192 9448 -1128
rect 9512 -1192 9520 -1128
rect 9440 -1208 9520 -1192
rect 9440 -1272 9448 -1208
rect 9512 -1272 9520 -1208
rect 9440 -1288 9520 -1272
rect 9440 -1352 9448 -1288
rect 9512 -1352 9520 -1288
rect 9440 -1368 9520 -1352
rect 9440 -1432 9448 -1368
rect 9512 -1432 9520 -1368
rect 9440 -1920 9520 -1432
rect 9760 -1048 9840 8
rect 9920 28308 10000 31520
rect 9920 28252 9932 28308
rect 9988 28252 10000 28308
rect 9920 18228 10000 28252
rect 9920 18172 9932 18228
rect 9988 18172 10000 18228
rect 9920 11988 10000 18172
rect 9920 11932 9932 11988
rect 9988 11932 10000 11988
rect 9920 0 10000 11932
rect 10080 31432 10160 31520
rect 10080 31368 10088 31432
rect 10152 31368 10160 31432
rect 10080 31272 10160 31368
rect 10080 31208 10088 31272
rect 10152 31208 10160 31272
rect 10080 31112 10160 31208
rect 10080 31048 10088 31112
rect 10152 31048 10160 31112
rect 10080 30952 10160 31048
rect 10080 30888 10088 30952
rect 10152 30888 10160 30952
rect 10080 30792 10160 30888
rect 10080 30728 10088 30792
rect 10152 30728 10160 30792
rect 10080 30632 10160 30728
rect 10080 30568 10088 30632
rect 10152 30568 10160 30632
rect 10080 30472 10160 30568
rect 10080 30408 10088 30472
rect 10152 30408 10160 30472
rect 10080 30312 10160 30408
rect 10080 30248 10088 30312
rect 10152 30248 10160 30312
rect 10080 30152 10160 30248
rect 10080 30088 10088 30152
rect 10152 30088 10160 30152
rect 10080 29992 10160 30088
rect 10080 29928 10088 29992
rect 10152 29928 10160 29992
rect 10080 29832 10160 29928
rect 10080 29768 10088 29832
rect 10152 29768 10160 29832
rect 10080 29672 10160 29768
rect 10080 29608 10088 29672
rect 10152 29608 10160 29672
rect 10080 29512 10160 29608
rect 10080 29448 10088 29512
rect 10152 29448 10160 29512
rect 10080 29352 10160 29448
rect 10080 29288 10088 29352
rect 10152 29288 10160 29352
rect 10080 29192 10160 29288
rect 10080 29128 10088 29192
rect 10152 29128 10160 29192
rect 10080 29032 10160 29128
rect 10080 28968 10088 29032
rect 10152 28968 10160 29032
rect 10080 28872 10160 28968
rect 10080 28808 10088 28872
rect 10152 28808 10160 28872
rect 10080 28712 10160 28808
rect 10080 28648 10088 28712
rect 10152 28648 10160 28712
rect 10080 28552 10160 28648
rect 10080 28488 10088 28552
rect 10152 28488 10160 28552
rect 10080 28392 10160 28488
rect 10080 28328 10088 28392
rect 10152 28328 10160 28392
rect 10080 28232 10160 28328
rect 10080 28168 10088 28232
rect 10152 28168 10160 28232
rect 10080 28072 10160 28168
rect 10080 28008 10088 28072
rect 10152 28008 10160 28072
rect 10080 27912 10160 28008
rect 10080 27848 10088 27912
rect 10152 27848 10160 27912
rect 10080 27752 10160 27848
rect 10080 27688 10088 27752
rect 10152 27688 10160 27752
rect 10080 27592 10160 27688
rect 10080 27528 10088 27592
rect 10152 27528 10160 27592
rect 10080 27432 10160 27528
rect 10080 27368 10088 27432
rect 10152 27368 10160 27432
rect 10080 27272 10160 27368
rect 10080 27208 10088 27272
rect 10152 27208 10160 27272
rect 10080 27112 10160 27208
rect 10080 27048 10088 27112
rect 10152 27048 10160 27112
rect 10080 26952 10160 27048
rect 10080 26888 10088 26952
rect 10152 26888 10160 26952
rect 10080 26792 10160 26888
rect 10080 26728 10088 26792
rect 10152 26728 10160 26792
rect 10080 26632 10160 26728
rect 10080 26568 10088 26632
rect 10152 26568 10160 26632
rect 10080 26472 10160 26568
rect 10080 26408 10088 26472
rect 10152 26408 10160 26472
rect 10080 26312 10160 26408
rect 10080 26248 10088 26312
rect 10152 26248 10160 26312
rect 10080 26152 10160 26248
rect 10080 26088 10088 26152
rect 10152 26088 10160 26152
rect 10080 25992 10160 26088
rect 10080 25928 10088 25992
rect 10152 25928 10160 25992
rect 10080 25832 10160 25928
rect 10080 25768 10088 25832
rect 10152 25768 10160 25832
rect 10080 25672 10160 25768
rect 10080 25608 10088 25672
rect 10152 25608 10160 25672
rect 10080 25512 10160 25608
rect 10080 25448 10088 25512
rect 10152 25448 10160 25512
rect 10080 25352 10160 25448
rect 10080 25288 10088 25352
rect 10152 25288 10160 25352
rect 10080 25192 10160 25288
rect 10080 25128 10088 25192
rect 10152 25128 10160 25192
rect 10080 25032 10160 25128
rect 10080 24968 10088 25032
rect 10152 24968 10160 25032
rect 10080 24872 10160 24968
rect 10080 24808 10088 24872
rect 10152 24808 10160 24872
rect 10080 24712 10160 24808
rect 10080 24648 10088 24712
rect 10152 24648 10160 24712
rect 10080 24552 10160 24648
rect 10080 24488 10088 24552
rect 10152 24488 10160 24552
rect 10080 24392 10160 24488
rect 10080 24328 10088 24392
rect 10152 24328 10160 24392
rect 10080 24232 10160 24328
rect 10080 24168 10088 24232
rect 10152 24168 10160 24232
rect 10080 24072 10160 24168
rect 10080 24008 10088 24072
rect 10152 24008 10160 24072
rect 10080 23912 10160 24008
rect 10080 23848 10088 23912
rect 10152 23848 10160 23912
rect 10080 23752 10160 23848
rect 10080 23688 10088 23752
rect 10152 23688 10160 23752
rect 10080 23592 10160 23688
rect 10080 23528 10088 23592
rect 10152 23528 10160 23592
rect 10080 23432 10160 23528
rect 10080 23368 10088 23432
rect 10152 23368 10160 23432
rect 10080 23272 10160 23368
rect 10080 23208 10088 23272
rect 10152 23208 10160 23272
rect 10080 23112 10160 23208
rect 10080 23048 10088 23112
rect 10152 23048 10160 23112
rect 10080 22952 10160 23048
rect 10080 22888 10088 22952
rect 10152 22888 10160 22952
rect 10080 22792 10160 22888
rect 10080 22728 10088 22792
rect 10152 22728 10160 22792
rect 10080 22632 10160 22728
rect 10080 22568 10088 22632
rect 10152 22568 10160 22632
rect 10080 22472 10160 22568
rect 10080 22408 10088 22472
rect 10152 22408 10160 22472
rect 10080 22312 10160 22408
rect 10080 22248 10088 22312
rect 10152 22248 10160 22312
rect 10080 22152 10160 22248
rect 10080 22088 10088 22152
rect 10152 22088 10160 22152
rect 10080 21992 10160 22088
rect 10080 21928 10088 21992
rect 10152 21928 10160 21992
rect 10080 21832 10160 21928
rect 10080 21768 10088 21832
rect 10152 21768 10160 21832
rect 10080 21672 10160 21768
rect 10080 21608 10088 21672
rect 10152 21608 10160 21672
rect 10080 21512 10160 21608
rect 10080 21448 10088 21512
rect 10152 21448 10160 21512
rect 10080 21352 10160 21448
rect 10080 21288 10088 21352
rect 10152 21288 10160 21352
rect 10080 21192 10160 21288
rect 10080 21128 10088 21192
rect 10152 21128 10160 21192
rect 10080 21032 10160 21128
rect 10080 20968 10088 21032
rect 10152 20968 10160 21032
rect 10080 20872 10160 20968
rect 10080 20808 10088 20872
rect 10152 20808 10160 20872
rect 10080 20712 10160 20808
rect 10080 20648 10088 20712
rect 10152 20648 10160 20712
rect 10080 20552 10160 20648
rect 10080 20488 10088 20552
rect 10152 20488 10160 20552
rect 10080 20392 10160 20488
rect 10080 20328 10088 20392
rect 10152 20328 10160 20392
rect 10080 20232 10160 20328
rect 10080 20168 10088 20232
rect 10152 20168 10160 20232
rect 10080 20072 10160 20168
rect 10080 20008 10088 20072
rect 10152 20008 10160 20072
rect 10080 19912 10160 20008
rect 10080 19848 10088 19912
rect 10152 19848 10160 19912
rect 10080 19752 10160 19848
rect 10080 19688 10088 19752
rect 10152 19688 10160 19752
rect 10080 19592 10160 19688
rect 10080 19528 10088 19592
rect 10152 19528 10160 19592
rect 10080 19432 10160 19528
rect 10080 19368 10088 19432
rect 10152 19368 10160 19432
rect 10080 19272 10160 19368
rect 10080 19208 10088 19272
rect 10152 19208 10160 19272
rect 10080 19112 10160 19208
rect 10080 19048 10088 19112
rect 10152 19048 10160 19112
rect 10080 18952 10160 19048
rect 10080 18888 10088 18952
rect 10152 18888 10160 18952
rect 10080 18792 10160 18888
rect 10080 18728 10088 18792
rect 10152 18728 10160 18792
rect 10080 18632 10160 18728
rect 10080 18568 10088 18632
rect 10152 18568 10160 18632
rect 10080 18472 10160 18568
rect 10080 18408 10088 18472
rect 10152 18408 10160 18472
rect 10080 18312 10160 18408
rect 10080 18248 10088 18312
rect 10152 18248 10160 18312
rect 10080 18152 10160 18248
rect 10080 18088 10088 18152
rect 10152 18088 10160 18152
rect 10080 17992 10160 18088
rect 10080 17928 10088 17992
rect 10152 17928 10160 17992
rect 10080 17832 10160 17928
rect 10080 17768 10088 17832
rect 10152 17768 10160 17832
rect 10080 17672 10160 17768
rect 10080 17608 10088 17672
rect 10152 17608 10160 17672
rect 10080 17512 10160 17608
rect 10080 17448 10088 17512
rect 10152 17448 10160 17512
rect 10080 17352 10160 17448
rect 10080 17288 10088 17352
rect 10152 17288 10160 17352
rect 10080 17192 10160 17288
rect 10080 17128 10088 17192
rect 10152 17128 10160 17192
rect 10080 17032 10160 17128
rect 10080 16968 10088 17032
rect 10152 16968 10160 17032
rect 10080 16872 10160 16968
rect 10080 16808 10088 16872
rect 10152 16808 10160 16872
rect 10080 16712 10160 16808
rect 10080 16648 10088 16712
rect 10152 16648 10160 16712
rect 10080 16552 10160 16648
rect 10080 16488 10088 16552
rect 10152 16488 10160 16552
rect 10080 16392 10160 16488
rect 10080 16328 10088 16392
rect 10152 16328 10160 16392
rect 10080 16232 10160 16328
rect 10080 16168 10088 16232
rect 10152 16168 10160 16232
rect 10080 16072 10160 16168
rect 10080 16008 10088 16072
rect 10152 16008 10160 16072
rect 10080 15912 10160 16008
rect 10080 15848 10088 15912
rect 10152 15848 10160 15912
rect 10080 15752 10160 15848
rect 10080 15688 10088 15752
rect 10152 15688 10160 15752
rect 10080 15592 10160 15688
rect 10080 15528 10088 15592
rect 10152 15528 10160 15592
rect 10080 15432 10160 15528
rect 10080 15368 10088 15432
rect 10152 15368 10160 15432
rect 10080 15272 10160 15368
rect 10080 15208 10088 15272
rect 10152 15208 10160 15272
rect 10080 15112 10160 15208
rect 10080 15048 10088 15112
rect 10152 15048 10160 15112
rect 10080 14952 10160 15048
rect 10080 14888 10088 14952
rect 10152 14888 10160 14952
rect 10080 14792 10160 14888
rect 10080 14728 10088 14792
rect 10152 14728 10160 14792
rect 10080 14632 10160 14728
rect 10080 14568 10088 14632
rect 10152 14568 10160 14632
rect 10080 14472 10160 14568
rect 10080 14408 10088 14472
rect 10152 14408 10160 14472
rect 10080 14312 10160 14408
rect 10080 14248 10088 14312
rect 10152 14248 10160 14312
rect 10080 14152 10160 14248
rect 10080 14088 10088 14152
rect 10152 14088 10160 14152
rect 10080 13992 10160 14088
rect 10080 13928 10088 13992
rect 10152 13928 10160 13992
rect 10080 13832 10160 13928
rect 10080 13768 10088 13832
rect 10152 13768 10160 13832
rect 10080 13672 10160 13768
rect 10080 13608 10088 13672
rect 10152 13608 10160 13672
rect 10080 13512 10160 13608
rect 10080 13448 10088 13512
rect 10152 13448 10160 13512
rect 10080 13352 10160 13448
rect 10080 13288 10088 13352
rect 10152 13288 10160 13352
rect 10080 13192 10160 13288
rect 10080 13128 10088 13192
rect 10152 13128 10160 13192
rect 10080 13032 10160 13128
rect 10080 12968 10088 13032
rect 10152 12968 10160 13032
rect 10080 12872 10160 12968
rect 10080 12808 10088 12872
rect 10152 12808 10160 12872
rect 10080 12712 10160 12808
rect 10080 12648 10088 12712
rect 10152 12648 10160 12712
rect 10080 12552 10160 12648
rect 10080 12488 10088 12552
rect 10152 12488 10160 12552
rect 10080 12392 10160 12488
rect 10080 12328 10088 12392
rect 10152 12328 10160 12392
rect 10080 12232 10160 12328
rect 10080 12168 10088 12232
rect 10152 12168 10160 12232
rect 10080 12072 10160 12168
rect 10080 12008 10088 12072
rect 10152 12008 10160 12072
rect 10080 11912 10160 12008
rect 10080 11848 10088 11912
rect 10152 11848 10160 11912
rect 10080 11752 10160 11848
rect 10080 11688 10088 11752
rect 10152 11688 10160 11752
rect 10080 11592 10160 11688
rect 10080 11528 10088 11592
rect 10152 11528 10160 11592
rect 10080 11432 10160 11528
rect 10080 11368 10088 11432
rect 10152 11368 10160 11432
rect 10080 11272 10160 11368
rect 10080 11208 10088 11272
rect 10152 11208 10160 11272
rect 10080 11112 10160 11208
rect 10080 11048 10088 11112
rect 10152 11048 10160 11112
rect 10080 10952 10160 11048
rect 10080 10888 10088 10952
rect 10152 10888 10160 10952
rect 10080 10792 10160 10888
rect 10080 10728 10088 10792
rect 10152 10728 10160 10792
rect 10080 10632 10160 10728
rect 10080 10568 10088 10632
rect 10152 10568 10160 10632
rect 10080 10472 10160 10568
rect 10080 10408 10088 10472
rect 10152 10408 10160 10472
rect 10080 10312 10160 10408
rect 10080 10248 10088 10312
rect 10152 10248 10160 10312
rect 10080 10152 10160 10248
rect 10080 10088 10088 10152
rect 10152 10088 10160 10152
rect 10080 9992 10160 10088
rect 10080 9928 10088 9992
rect 10152 9928 10160 9992
rect 10080 9832 10160 9928
rect 10080 9768 10088 9832
rect 10152 9768 10160 9832
rect 10080 9672 10160 9768
rect 10080 9608 10088 9672
rect 10152 9608 10160 9672
rect 10080 9512 10160 9608
rect 10080 9448 10088 9512
rect 10152 9448 10160 9512
rect 10080 9352 10160 9448
rect 10080 9288 10088 9352
rect 10152 9288 10160 9352
rect 10080 9192 10160 9288
rect 10080 9128 10088 9192
rect 10152 9128 10160 9192
rect 10080 9032 10160 9128
rect 10080 8968 10088 9032
rect 10152 8968 10160 9032
rect 10080 8872 10160 8968
rect 10080 8808 10088 8872
rect 10152 8808 10160 8872
rect 10080 8712 10160 8808
rect 10080 8648 10088 8712
rect 10152 8648 10160 8712
rect 10080 8552 10160 8648
rect 10080 8488 10088 8552
rect 10152 8488 10160 8552
rect 10080 8392 10160 8488
rect 10080 8328 10088 8392
rect 10152 8328 10160 8392
rect 10080 8232 10160 8328
rect 10080 8168 10088 8232
rect 10152 8168 10160 8232
rect 10080 8072 10160 8168
rect 10080 8008 10088 8072
rect 10152 8008 10160 8072
rect 10080 7912 10160 8008
rect 10080 7848 10088 7912
rect 10152 7848 10160 7912
rect 10080 7752 10160 7848
rect 10080 7688 10088 7752
rect 10152 7688 10160 7752
rect 10080 7592 10160 7688
rect 10080 7528 10088 7592
rect 10152 7528 10160 7592
rect 10080 7432 10160 7528
rect 10080 7368 10088 7432
rect 10152 7368 10160 7432
rect 10080 7272 10160 7368
rect 10080 7208 10088 7272
rect 10152 7208 10160 7272
rect 10080 7112 10160 7208
rect 10080 7048 10088 7112
rect 10152 7048 10160 7112
rect 10080 6952 10160 7048
rect 10080 6888 10088 6952
rect 10152 6888 10160 6952
rect 10080 6792 10160 6888
rect 10080 6728 10088 6792
rect 10152 6728 10160 6792
rect 10080 6632 10160 6728
rect 10080 6568 10088 6632
rect 10152 6568 10160 6632
rect 10080 6472 10160 6568
rect 10080 6408 10088 6472
rect 10152 6408 10160 6472
rect 10080 6312 10160 6408
rect 10080 6248 10088 6312
rect 10152 6248 10160 6312
rect 10080 6152 10160 6248
rect 10080 6088 10088 6152
rect 10152 6088 10160 6152
rect 10080 5992 10160 6088
rect 10080 5928 10088 5992
rect 10152 5928 10160 5992
rect 10080 5832 10160 5928
rect 10080 5768 10088 5832
rect 10152 5768 10160 5832
rect 10080 5672 10160 5768
rect 10080 5608 10088 5672
rect 10152 5608 10160 5672
rect 10080 5512 10160 5608
rect 10080 5448 10088 5512
rect 10152 5448 10160 5512
rect 10080 5352 10160 5448
rect 10080 5288 10088 5352
rect 10152 5288 10160 5352
rect 10080 5192 10160 5288
rect 10080 5128 10088 5192
rect 10152 5128 10160 5192
rect 10080 5032 10160 5128
rect 10080 4968 10088 5032
rect 10152 4968 10160 5032
rect 10080 4872 10160 4968
rect 10080 4808 10088 4872
rect 10152 4808 10160 4872
rect 10080 4712 10160 4808
rect 10080 4648 10088 4712
rect 10152 4648 10160 4712
rect 10080 4552 10160 4648
rect 10080 4488 10088 4552
rect 10152 4488 10160 4552
rect 10080 4392 10160 4488
rect 10080 4328 10088 4392
rect 10152 4328 10160 4392
rect 10080 4232 10160 4328
rect 10080 4168 10088 4232
rect 10152 4168 10160 4232
rect 10080 4072 10160 4168
rect 10080 4008 10088 4072
rect 10152 4008 10160 4072
rect 10080 3912 10160 4008
rect 10080 3848 10088 3912
rect 10152 3848 10160 3912
rect 10080 3752 10160 3848
rect 10080 3688 10088 3752
rect 10152 3688 10160 3752
rect 10080 3592 10160 3688
rect 10080 3528 10088 3592
rect 10152 3528 10160 3592
rect 10080 3432 10160 3528
rect 10080 3368 10088 3432
rect 10152 3368 10160 3432
rect 10080 3272 10160 3368
rect 10080 3208 10088 3272
rect 10152 3208 10160 3272
rect 10080 3112 10160 3208
rect 10080 3048 10088 3112
rect 10152 3048 10160 3112
rect 10080 2952 10160 3048
rect 10080 2888 10088 2952
rect 10152 2888 10160 2952
rect 10080 2792 10160 2888
rect 10080 2728 10088 2792
rect 10152 2728 10160 2792
rect 10080 2632 10160 2728
rect 10080 2568 10088 2632
rect 10152 2568 10160 2632
rect 10080 2472 10160 2568
rect 10080 2408 10088 2472
rect 10152 2408 10160 2472
rect 10080 2312 10160 2408
rect 10080 2248 10088 2312
rect 10152 2248 10160 2312
rect 10080 2152 10160 2248
rect 10080 2088 10088 2152
rect 10152 2088 10160 2152
rect 10080 1992 10160 2088
rect 10080 1928 10088 1992
rect 10152 1928 10160 1992
rect 10080 1832 10160 1928
rect 10080 1768 10088 1832
rect 10152 1768 10160 1832
rect 10080 1672 10160 1768
rect 10080 1608 10088 1672
rect 10152 1608 10160 1672
rect 10080 1512 10160 1608
rect 10080 1448 10088 1512
rect 10152 1448 10160 1512
rect 10080 1352 10160 1448
rect 10080 1288 10088 1352
rect 10152 1288 10160 1352
rect 10080 1192 10160 1288
rect 10080 1128 10088 1192
rect 10152 1128 10160 1192
rect 10080 1032 10160 1128
rect 10080 968 10088 1032
rect 10152 968 10160 1032
rect 10080 872 10160 968
rect 10080 808 10088 872
rect 10152 808 10160 872
rect 10080 712 10160 808
rect 10080 648 10088 712
rect 10152 648 10160 712
rect 10080 552 10160 648
rect 10080 488 10088 552
rect 10152 488 10160 552
rect 10080 392 10160 488
rect 10080 328 10088 392
rect 10152 328 10160 392
rect 10080 232 10160 328
rect 10080 168 10088 232
rect 10152 168 10160 232
rect 10080 72 10160 168
rect 10080 8 10088 72
rect 10152 8 10160 72
rect 9760 -1112 9768 -1048
rect 9832 -1112 9840 -1048
rect 9760 -1128 9840 -1112
rect 9760 -1192 9768 -1128
rect 9832 -1192 9840 -1128
rect 9760 -1208 9840 -1192
rect 9760 -1272 9768 -1208
rect 9832 -1272 9840 -1208
rect 9760 -1288 9840 -1272
rect 9760 -1352 9768 -1288
rect 9832 -1352 9840 -1288
rect 9760 -1368 9840 -1352
rect 9760 -1432 9768 -1368
rect 9832 -1432 9840 -1368
rect 9760 -1920 9840 -1432
rect 10080 -1048 10160 8
rect 10240 26388 10320 31520
rect 10240 26332 10252 26388
rect 10308 26332 10320 26388
rect 10240 20468 10320 26332
rect 10240 20412 10252 20468
rect 10308 20412 10320 20468
rect 10240 20148 10320 20412
rect 10240 20092 10252 20148
rect 10308 20092 10320 20148
rect 10240 18548 10320 20092
rect 10240 18492 10252 18548
rect 10308 18492 10320 18548
rect 10240 0 10320 18492
rect 10400 31432 10480 31520
rect 10400 31368 10408 31432
rect 10472 31368 10480 31432
rect 10400 31272 10480 31368
rect 10400 31208 10408 31272
rect 10472 31208 10480 31272
rect 10400 31112 10480 31208
rect 10400 31048 10408 31112
rect 10472 31048 10480 31112
rect 10400 30952 10480 31048
rect 10400 30888 10408 30952
rect 10472 30888 10480 30952
rect 10400 30792 10480 30888
rect 10400 30728 10408 30792
rect 10472 30728 10480 30792
rect 10400 30632 10480 30728
rect 10400 30568 10408 30632
rect 10472 30568 10480 30632
rect 10400 30472 10480 30568
rect 10400 30408 10408 30472
rect 10472 30408 10480 30472
rect 10400 30312 10480 30408
rect 10400 30248 10408 30312
rect 10472 30248 10480 30312
rect 10400 30152 10480 30248
rect 10400 30088 10408 30152
rect 10472 30088 10480 30152
rect 10400 29992 10480 30088
rect 10400 29928 10408 29992
rect 10472 29928 10480 29992
rect 10400 29832 10480 29928
rect 10400 29768 10408 29832
rect 10472 29768 10480 29832
rect 10400 29672 10480 29768
rect 10400 29608 10408 29672
rect 10472 29608 10480 29672
rect 10400 29512 10480 29608
rect 10400 29448 10408 29512
rect 10472 29448 10480 29512
rect 10400 29352 10480 29448
rect 10400 29288 10408 29352
rect 10472 29288 10480 29352
rect 10400 29192 10480 29288
rect 10400 29128 10408 29192
rect 10472 29128 10480 29192
rect 10400 29032 10480 29128
rect 10400 28968 10408 29032
rect 10472 28968 10480 29032
rect 10400 28872 10480 28968
rect 10400 28808 10408 28872
rect 10472 28808 10480 28872
rect 10400 28712 10480 28808
rect 10400 28648 10408 28712
rect 10472 28648 10480 28712
rect 10400 28552 10480 28648
rect 10400 28488 10408 28552
rect 10472 28488 10480 28552
rect 10400 28392 10480 28488
rect 10400 28328 10408 28392
rect 10472 28328 10480 28392
rect 10400 28232 10480 28328
rect 10400 28168 10408 28232
rect 10472 28168 10480 28232
rect 10400 28072 10480 28168
rect 10400 28008 10408 28072
rect 10472 28008 10480 28072
rect 10400 27912 10480 28008
rect 10400 27848 10408 27912
rect 10472 27848 10480 27912
rect 10400 27752 10480 27848
rect 10400 27688 10408 27752
rect 10472 27688 10480 27752
rect 10400 27592 10480 27688
rect 10400 27528 10408 27592
rect 10472 27528 10480 27592
rect 10400 27432 10480 27528
rect 10400 27368 10408 27432
rect 10472 27368 10480 27432
rect 10400 27272 10480 27368
rect 10400 27208 10408 27272
rect 10472 27208 10480 27272
rect 10400 27112 10480 27208
rect 10400 27048 10408 27112
rect 10472 27048 10480 27112
rect 10400 26952 10480 27048
rect 10400 26888 10408 26952
rect 10472 26888 10480 26952
rect 10400 26792 10480 26888
rect 10400 26728 10408 26792
rect 10472 26728 10480 26792
rect 10400 26632 10480 26728
rect 10400 26568 10408 26632
rect 10472 26568 10480 26632
rect 10400 26472 10480 26568
rect 10400 26408 10408 26472
rect 10472 26408 10480 26472
rect 10400 26312 10480 26408
rect 10400 26248 10408 26312
rect 10472 26248 10480 26312
rect 10400 26152 10480 26248
rect 10400 26088 10408 26152
rect 10472 26088 10480 26152
rect 10400 25992 10480 26088
rect 10400 25928 10408 25992
rect 10472 25928 10480 25992
rect 10400 25832 10480 25928
rect 10400 25768 10408 25832
rect 10472 25768 10480 25832
rect 10400 25672 10480 25768
rect 10400 25608 10408 25672
rect 10472 25608 10480 25672
rect 10400 25512 10480 25608
rect 10400 25448 10408 25512
rect 10472 25448 10480 25512
rect 10400 25352 10480 25448
rect 10400 25288 10408 25352
rect 10472 25288 10480 25352
rect 10400 25192 10480 25288
rect 10400 25128 10408 25192
rect 10472 25128 10480 25192
rect 10400 25032 10480 25128
rect 10400 24968 10408 25032
rect 10472 24968 10480 25032
rect 10400 24872 10480 24968
rect 10400 24808 10408 24872
rect 10472 24808 10480 24872
rect 10400 24712 10480 24808
rect 10400 24648 10408 24712
rect 10472 24648 10480 24712
rect 10400 24552 10480 24648
rect 10400 24488 10408 24552
rect 10472 24488 10480 24552
rect 10400 24392 10480 24488
rect 10400 24328 10408 24392
rect 10472 24328 10480 24392
rect 10400 24232 10480 24328
rect 10400 24168 10408 24232
rect 10472 24168 10480 24232
rect 10400 24072 10480 24168
rect 10400 24008 10408 24072
rect 10472 24008 10480 24072
rect 10400 23912 10480 24008
rect 10400 23848 10408 23912
rect 10472 23848 10480 23912
rect 10400 23752 10480 23848
rect 10400 23688 10408 23752
rect 10472 23688 10480 23752
rect 10400 23592 10480 23688
rect 10400 23528 10408 23592
rect 10472 23528 10480 23592
rect 10400 23432 10480 23528
rect 10400 23368 10408 23432
rect 10472 23368 10480 23432
rect 10400 23272 10480 23368
rect 10400 23208 10408 23272
rect 10472 23208 10480 23272
rect 10400 23112 10480 23208
rect 10400 23048 10408 23112
rect 10472 23048 10480 23112
rect 10400 22952 10480 23048
rect 10400 22888 10408 22952
rect 10472 22888 10480 22952
rect 10400 22792 10480 22888
rect 10400 22728 10408 22792
rect 10472 22728 10480 22792
rect 10400 22632 10480 22728
rect 10400 22568 10408 22632
rect 10472 22568 10480 22632
rect 10400 22472 10480 22568
rect 10400 22408 10408 22472
rect 10472 22408 10480 22472
rect 10400 22312 10480 22408
rect 10400 22248 10408 22312
rect 10472 22248 10480 22312
rect 10400 22152 10480 22248
rect 10400 22088 10408 22152
rect 10472 22088 10480 22152
rect 10400 21992 10480 22088
rect 10400 21928 10408 21992
rect 10472 21928 10480 21992
rect 10400 21832 10480 21928
rect 10400 21768 10408 21832
rect 10472 21768 10480 21832
rect 10400 21672 10480 21768
rect 10400 21608 10408 21672
rect 10472 21608 10480 21672
rect 10400 21512 10480 21608
rect 10400 21448 10408 21512
rect 10472 21448 10480 21512
rect 10400 21352 10480 21448
rect 10400 21288 10408 21352
rect 10472 21288 10480 21352
rect 10400 21192 10480 21288
rect 10400 21128 10408 21192
rect 10472 21128 10480 21192
rect 10400 21032 10480 21128
rect 10400 20968 10408 21032
rect 10472 20968 10480 21032
rect 10400 20872 10480 20968
rect 10400 20808 10408 20872
rect 10472 20808 10480 20872
rect 10400 20712 10480 20808
rect 10400 20648 10408 20712
rect 10472 20648 10480 20712
rect 10400 20552 10480 20648
rect 10400 20488 10408 20552
rect 10472 20488 10480 20552
rect 10400 20392 10480 20488
rect 10400 20328 10408 20392
rect 10472 20328 10480 20392
rect 10400 20232 10480 20328
rect 10400 20168 10408 20232
rect 10472 20168 10480 20232
rect 10400 20072 10480 20168
rect 10400 20008 10408 20072
rect 10472 20008 10480 20072
rect 10400 19912 10480 20008
rect 10400 19848 10408 19912
rect 10472 19848 10480 19912
rect 10400 19752 10480 19848
rect 10400 19688 10408 19752
rect 10472 19688 10480 19752
rect 10400 19592 10480 19688
rect 10400 19528 10408 19592
rect 10472 19528 10480 19592
rect 10400 19432 10480 19528
rect 10400 19368 10408 19432
rect 10472 19368 10480 19432
rect 10400 19272 10480 19368
rect 10400 19208 10408 19272
rect 10472 19208 10480 19272
rect 10400 19112 10480 19208
rect 10400 19048 10408 19112
rect 10472 19048 10480 19112
rect 10400 18952 10480 19048
rect 10400 18888 10408 18952
rect 10472 18888 10480 18952
rect 10400 18792 10480 18888
rect 10400 18728 10408 18792
rect 10472 18728 10480 18792
rect 10400 18632 10480 18728
rect 10400 18568 10408 18632
rect 10472 18568 10480 18632
rect 10400 18472 10480 18568
rect 10400 18408 10408 18472
rect 10472 18408 10480 18472
rect 10400 18312 10480 18408
rect 10400 18248 10408 18312
rect 10472 18248 10480 18312
rect 10400 18152 10480 18248
rect 10400 18088 10408 18152
rect 10472 18088 10480 18152
rect 10400 17992 10480 18088
rect 10400 17928 10408 17992
rect 10472 17928 10480 17992
rect 10400 17832 10480 17928
rect 10400 17768 10408 17832
rect 10472 17768 10480 17832
rect 10400 17672 10480 17768
rect 10400 17608 10408 17672
rect 10472 17608 10480 17672
rect 10400 17512 10480 17608
rect 10400 17448 10408 17512
rect 10472 17448 10480 17512
rect 10400 17352 10480 17448
rect 10400 17288 10408 17352
rect 10472 17288 10480 17352
rect 10400 17192 10480 17288
rect 10400 17128 10408 17192
rect 10472 17128 10480 17192
rect 10400 17032 10480 17128
rect 10400 16968 10408 17032
rect 10472 16968 10480 17032
rect 10400 16872 10480 16968
rect 10400 16808 10408 16872
rect 10472 16808 10480 16872
rect 10400 16712 10480 16808
rect 10400 16648 10408 16712
rect 10472 16648 10480 16712
rect 10400 16552 10480 16648
rect 10400 16488 10408 16552
rect 10472 16488 10480 16552
rect 10400 16392 10480 16488
rect 10400 16328 10408 16392
rect 10472 16328 10480 16392
rect 10400 16232 10480 16328
rect 10400 16168 10408 16232
rect 10472 16168 10480 16232
rect 10400 16072 10480 16168
rect 10400 16008 10408 16072
rect 10472 16008 10480 16072
rect 10400 15912 10480 16008
rect 10400 15848 10408 15912
rect 10472 15848 10480 15912
rect 10400 15752 10480 15848
rect 10400 15688 10408 15752
rect 10472 15688 10480 15752
rect 10400 15592 10480 15688
rect 10400 15528 10408 15592
rect 10472 15528 10480 15592
rect 10400 15432 10480 15528
rect 10400 15368 10408 15432
rect 10472 15368 10480 15432
rect 10400 15272 10480 15368
rect 10400 15208 10408 15272
rect 10472 15208 10480 15272
rect 10400 15112 10480 15208
rect 10400 15048 10408 15112
rect 10472 15048 10480 15112
rect 10400 14952 10480 15048
rect 10400 14888 10408 14952
rect 10472 14888 10480 14952
rect 10400 14792 10480 14888
rect 10400 14728 10408 14792
rect 10472 14728 10480 14792
rect 10400 14632 10480 14728
rect 10400 14568 10408 14632
rect 10472 14568 10480 14632
rect 10400 14472 10480 14568
rect 10400 14408 10408 14472
rect 10472 14408 10480 14472
rect 10400 14312 10480 14408
rect 10400 14248 10408 14312
rect 10472 14248 10480 14312
rect 10400 14152 10480 14248
rect 10400 14088 10408 14152
rect 10472 14088 10480 14152
rect 10400 13992 10480 14088
rect 10400 13928 10408 13992
rect 10472 13928 10480 13992
rect 10400 13832 10480 13928
rect 10400 13768 10408 13832
rect 10472 13768 10480 13832
rect 10400 13672 10480 13768
rect 10400 13608 10408 13672
rect 10472 13608 10480 13672
rect 10400 13512 10480 13608
rect 10400 13448 10408 13512
rect 10472 13448 10480 13512
rect 10400 13352 10480 13448
rect 10400 13288 10408 13352
rect 10472 13288 10480 13352
rect 10400 13192 10480 13288
rect 10400 13128 10408 13192
rect 10472 13128 10480 13192
rect 10400 13032 10480 13128
rect 10400 12968 10408 13032
rect 10472 12968 10480 13032
rect 10400 12872 10480 12968
rect 10400 12808 10408 12872
rect 10472 12808 10480 12872
rect 10400 12712 10480 12808
rect 10400 12648 10408 12712
rect 10472 12648 10480 12712
rect 10400 12552 10480 12648
rect 10400 12488 10408 12552
rect 10472 12488 10480 12552
rect 10400 12392 10480 12488
rect 10400 12328 10408 12392
rect 10472 12328 10480 12392
rect 10400 12232 10480 12328
rect 10400 12168 10408 12232
rect 10472 12168 10480 12232
rect 10400 12072 10480 12168
rect 10400 12008 10408 12072
rect 10472 12008 10480 12072
rect 10400 11912 10480 12008
rect 10400 11848 10408 11912
rect 10472 11848 10480 11912
rect 10400 11752 10480 11848
rect 10400 11688 10408 11752
rect 10472 11688 10480 11752
rect 10400 11592 10480 11688
rect 10400 11528 10408 11592
rect 10472 11528 10480 11592
rect 10400 11432 10480 11528
rect 10400 11368 10408 11432
rect 10472 11368 10480 11432
rect 10400 11272 10480 11368
rect 10400 11208 10408 11272
rect 10472 11208 10480 11272
rect 10400 11112 10480 11208
rect 10400 11048 10408 11112
rect 10472 11048 10480 11112
rect 10400 10952 10480 11048
rect 10400 10888 10408 10952
rect 10472 10888 10480 10952
rect 10400 10792 10480 10888
rect 10400 10728 10408 10792
rect 10472 10728 10480 10792
rect 10400 10632 10480 10728
rect 10400 10568 10408 10632
rect 10472 10568 10480 10632
rect 10400 10472 10480 10568
rect 10400 10408 10408 10472
rect 10472 10408 10480 10472
rect 10400 10312 10480 10408
rect 10400 10248 10408 10312
rect 10472 10248 10480 10312
rect 10400 10152 10480 10248
rect 10400 10088 10408 10152
rect 10472 10088 10480 10152
rect 10400 9992 10480 10088
rect 10400 9928 10408 9992
rect 10472 9928 10480 9992
rect 10400 9832 10480 9928
rect 10400 9768 10408 9832
rect 10472 9768 10480 9832
rect 10400 9672 10480 9768
rect 10400 9608 10408 9672
rect 10472 9608 10480 9672
rect 10400 9512 10480 9608
rect 10400 9448 10408 9512
rect 10472 9448 10480 9512
rect 10400 9352 10480 9448
rect 10400 9288 10408 9352
rect 10472 9288 10480 9352
rect 10400 9192 10480 9288
rect 10400 9128 10408 9192
rect 10472 9128 10480 9192
rect 10400 9032 10480 9128
rect 10400 8968 10408 9032
rect 10472 8968 10480 9032
rect 10400 8872 10480 8968
rect 10400 8808 10408 8872
rect 10472 8808 10480 8872
rect 10400 8712 10480 8808
rect 10400 8648 10408 8712
rect 10472 8648 10480 8712
rect 10400 8552 10480 8648
rect 10400 8488 10408 8552
rect 10472 8488 10480 8552
rect 10400 8392 10480 8488
rect 10400 8328 10408 8392
rect 10472 8328 10480 8392
rect 10400 8232 10480 8328
rect 10400 8168 10408 8232
rect 10472 8168 10480 8232
rect 10400 8072 10480 8168
rect 10400 8008 10408 8072
rect 10472 8008 10480 8072
rect 10400 7912 10480 8008
rect 10400 7848 10408 7912
rect 10472 7848 10480 7912
rect 10400 7752 10480 7848
rect 10400 7688 10408 7752
rect 10472 7688 10480 7752
rect 10400 7592 10480 7688
rect 10400 7528 10408 7592
rect 10472 7528 10480 7592
rect 10400 7432 10480 7528
rect 10400 7368 10408 7432
rect 10472 7368 10480 7432
rect 10400 7272 10480 7368
rect 10400 7208 10408 7272
rect 10472 7208 10480 7272
rect 10400 7112 10480 7208
rect 10400 7048 10408 7112
rect 10472 7048 10480 7112
rect 10400 6952 10480 7048
rect 10400 6888 10408 6952
rect 10472 6888 10480 6952
rect 10400 6792 10480 6888
rect 10400 6728 10408 6792
rect 10472 6728 10480 6792
rect 10400 6632 10480 6728
rect 10400 6568 10408 6632
rect 10472 6568 10480 6632
rect 10400 6472 10480 6568
rect 10400 6408 10408 6472
rect 10472 6408 10480 6472
rect 10400 6312 10480 6408
rect 10400 6248 10408 6312
rect 10472 6248 10480 6312
rect 10400 6152 10480 6248
rect 10400 6088 10408 6152
rect 10472 6088 10480 6152
rect 10400 5992 10480 6088
rect 10400 5928 10408 5992
rect 10472 5928 10480 5992
rect 10400 5832 10480 5928
rect 10400 5768 10408 5832
rect 10472 5768 10480 5832
rect 10400 5672 10480 5768
rect 10400 5608 10408 5672
rect 10472 5608 10480 5672
rect 10400 5512 10480 5608
rect 10400 5448 10408 5512
rect 10472 5448 10480 5512
rect 10400 5352 10480 5448
rect 10400 5288 10408 5352
rect 10472 5288 10480 5352
rect 10400 5192 10480 5288
rect 10400 5128 10408 5192
rect 10472 5128 10480 5192
rect 10400 5032 10480 5128
rect 10400 4968 10408 5032
rect 10472 4968 10480 5032
rect 10400 4872 10480 4968
rect 10400 4808 10408 4872
rect 10472 4808 10480 4872
rect 10400 4712 10480 4808
rect 10400 4648 10408 4712
rect 10472 4648 10480 4712
rect 10400 4552 10480 4648
rect 10400 4488 10408 4552
rect 10472 4488 10480 4552
rect 10400 4392 10480 4488
rect 10400 4328 10408 4392
rect 10472 4328 10480 4392
rect 10400 4232 10480 4328
rect 10400 4168 10408 4232
rect 10472 4168 10480 4232
rect 10400 4072 10480 4168
rect 10400 4008 10408 4072
rect 10472 4008 10480 4072
rect 10400 3912 10480 4008
rect 10400 3848 10408 3912
rect 10472 3848 10480 3912
rect 10400 3752 10480 3848
rect 10400 3688 10408 3752
rect 10472 3688 10480 3752
rect 10400 3592 10480 3688
rect 10400 3528 10408 3592
rect 10472 3528 10480 3592
rect 10400 3432 10480 3528
rect 10400 3368 10408 3432
rect 10472 3368 10480 3432
rect 10400 3272 10480 3368
rect 10400 3208 10408 3272
rect 10472 3208 10480 3272
rect 10400 3112 10480 3208
rect 10400 3048 10408 3112
rect 10472 3048 10480 3112
rect 10400 2952 10480 3048
rect 10400 2888 10408 2952
rect 10472 2888 10480 2952
rect 10400 2792 10480 2888
rect 10400 2728 10408 2792
rect 10472 2728 10480 2792
rect 10400 2632 10480 2728
rect 10400 2568 10408 2632
rect 10472 2568 10480 2632
rect 10400 2472 10480 2568
rect 10400 2408 10408 2472
rect 10472 2408 10480 2472
rect 10400 2312 10480 2408
rect 10400 2248 10408 2312
rect 10472 2248 10480 2312
rect 10400 2152 10480 2248
rect 10400 2088 10408 2152
rect 10472 2088 10480 2152
rect 10400 1992 10480 2088
rect 10400 1928 10408 1992
rect 10472 1928 10480 1992
rect 10400 1832 10480 1928
rect 10400 1768 10408 1832
rect 10472 1768 10480 1832
rect 10400 1672 10480 1768
rect 10400 1608 10408 1672
rect 10472 1608 10480 1672
rect 10400 1512 10480 1608
rect 10400 1448 10408 1512
rect 10472 1448 10480 1512
rect 10400 1352 10480 1448
rect 10400 1288 10408 1352
rect 10472 1288 10480 1352
rect 10400 1192 10480 1288
rect 10400 1128 10408 1192
rect 10472 1128 10480 1192
rect 10400 1032 10480 1128
rect 10400 968 10408 1032
rect 10472 968 10480 1032
rect 10400 872 10480 968
rect 10400 808 10408 872
rect 10472 808 10480 872
rect 10400 712 10480 808
rect 10400 648 10408 712
rect 10472 648 10480 712
rect 10400 552 10480 648
rect 10400 488 10408 552
rect 10472 488 10480 552
rect 10400 392 10480 488
rect 10400 328 10408 392
rect 10472 328 10480 392
rect 10400 232 10480 328
rect 10400 168 10408 232
rect 10472 168 10480 232
rect 10400 72 10480 168
rect 10400 8 10408 72
rect 10472 8 10480 72
rect 10080 -1112 10088 -1048
rect 10152 -1112 10160 -1048
rect 10080 -1128 10160 -1112
rect 10080 -1192 10088 -1128
rect 10152 -1192 10160 -1128
rect 10080 -1208 10160 -1192
rect 10080 -1272 10088 -1208
rect 10152 -1272 10160 -1208
rect 10080 -1288 10160 -1272
rect 10080 -1352 10088 -1288
rect 10152 -1352 10160 -1288
rect 10080 -1368 10160 -1352
rect 10080 -1432 10088 -1368
rect 10152 -1432 10160 -1368
rect 10080 -1920 10160 -1432
rect 10400 -1048 10480 8
rect 10560 28628 10640 31520
rect 10560 28572 10572 28628
rect 10628 28572 10640 28628
rect 10560 26708 10640 28572
rect 10560 26652 10572 26708
rect 10628 26652 10640 26708
rect 10560 26388 10640 26652
rect 10560 26332 10572 26388
rect 10628 26332 10640 26388
rect 10560 0 10640 26332
rect 10720 31432 10800 31520
rect 10720 31368 10728 31432
rect 10792 31368 10800 31432
rect 10720 31272 10800 31368
rect 10720 31208 10728 31272
rect 10792 31208 10800 31272
rect 10720 31112 10800 31208
rect 10720 31048 10728 31112
rect 10792 31048 10800 31112
rect 10720 30952 10800 31048
rect 10720 30888 10728 30952
rect 10792 30888 10800 30952
rect 10720 30792 10800 30888
rect 10720 30728 10728 30792
rect 10792 30728 10800 30792
rect 10720 30632 10800 30728
rect 10720 30568 10728 30632
rect 10792 30568 10800 30632
rect 10720 30472 10800 30568
rect 10720 30408 10728 30472
rect 10792 30408 10800 30472
rect 10720 30312 10800 30408
rect 10720 30248 10728 30312
rect 10792 30248 10800 30312
rect 10720 30152 10800 30248
rect 10720 30088 10728 30152
rect 10792 30088 10800 30152
rect 10720 29992 10800 30088
rect 10720 29928 10728 29992
rect 10792 29928 10800 29992
rect 10720 29832 10800 29928
rect 10720 29768 10728 29832
rect 10792 29768 10800 29832
rect 10720 29672 10800 29768
rect 10720 29608 10728 29672
rect 10792 29608 10800 29672
rect 10720 29512 10800 29608
rect 10720 29448 10728 29512
rect 10792 29448 10800 29512
rect 10720 29352 10800 29448
rect 10720 29288 10728 29352
rect 10792 29288 10800 29352
rect 10720 29192 10800 29288
rect 10720 29128 10728 29192
rect 10792 29128 10800 29192
rect 10720 29032 10800 29128
rect 10720 28968 10728 29032
rect 10792 28968 10800 29032
rect 10720 28872 10800 28968
rect 10720 28808 10728 28872
rect 10792 28808 10800 28872
rect 10720 28712 10800 28808
rect 10720 28648 10728 28712
rect 10792 28648 10800 28712
rect 10720 28552 10800 28648
rect 10720 28488 10728 28552
rect 10792 28488 10800 28552
rect 10720 28392 10800 28488
rect 10720 28328 10728 28392
rect 10792 28328 10800 28392
rect 10720 28232 10800 28328
rect 10720 28168 10728 28232
rect 10792 28168 10800 28232
rect 10720 28072 10800 28168
rect 10720 28008 10728 28072
rect 10792 28008 10800 28072
rect 10720 27912 10800 28008
rect 10720 27848 10728 27912
rect 10792 27848 10800 27912
rect 10720 27752 10800 27848
rect 10720 27688 10728 27752
rect 10792 27688 10800 27752
rect 10720 27592 10800 27688
rect 10720 27528 10728 27592
rect 10792 27528 10800 27592
rect 10720 27432 10800 27528
rect 10720 27368 10728 27432
rect 10792 27368 10800 27432
rect 10720 27272 10800 27368
rect 10720 27208 10728 27272
rect 10792 27208 10800 27272
rect 10720 27112 10800 27208
rect 10720 27048 10728 27112
rect 10792 27048 10800 27112
rect 10720 26952 10800 27048
rect 10720 26888 10728 26952
rect 10792 26888 10800 26952
rect 10720 26792 10800 26888
rect 10720 26728 10728 26792
rect 10792 26728 10800 26792
rect 10720 26632 10800 26728
rect 10720 26568 10728 26632
rect 10792 26568 10800 26632
rect 10720 26472 10800 26568
rect 10720 26408 10728 26472
rect 10792 26408 10800 26472
rect 10720 26312 10800 26408
rect 10720 26248 10728 26312
rect 10792 26248 10800 26312
rect 10720 26152 10800 26248
rect 10720 26088 10728 26152
rect 10792 26088 10800 26152
rect 10720 25992 10800 26088
rect 10720 25928 10728 25992
rect 10792 25928 10800 25992
rect 10720 25832 10800 25928
rect 10720 25768 10728 25832
rect 10792 25768 10800 25832
rect 10720 25672 10800 25768
rect 10720 25608 10728 25672
rect 10792 25608 10800 25672
rect 10720 25512 10800 25608
rect 10720 25448 10728 25512
rect 10792 25448 10800 25512
rect 10720 25352 10800 25448
rect 10720 25288 10728 25352
rect 10792 25288 10800 25352
rect 10720 25192 10800 25288
rect 10720 25128 10728 25192
rect 10792 25128 10800 25192
rect 10720 25032 10800 25128
rect 10720 24968 10728 25032
rect 10792 24968 10800 25032
rect 10720 24872 10800 24968
rect 10720 24808 10728 24872
rect 10792 24808 10800 24872
rect 10720 24712 10800 24808
rect 10720 24648 10728 24712
rect 10792 24648 10800 24712
rect 10720 24552 10800 24648
rect 10720 24488 10728 24552
rect 10792 24488 10800 24552
rect 10720 24392 10800 24488
rect 10720 24328 10728 24392
rect 10792 24328 10800 24392
rect 10720 24232 10800 24328
rect 10720 24168 10728 24232
rect 10792 24168 10800 24232
rect 10720 24072 10800 24168
rect 10720 24008 10728 24072
rect 10792 24008 10800 24072
rect 10720 23912 10800 24008
rect 10720 23848 10728 23912
rect 10792 23848 10800 23912
rect 10720 23752 10800 23848
rect 10720 23688 10728 23752
rect 10792 23688 10800 23752
rect 10720 23592 10800 23688
rect 10720 23528 10728 23592
rect 10792 23528 10800 23592
rect 10720 23432 10800 23528
rect 10720 23368 10728 23432
rect 10792 23368 10800 23432
rect 10720 23272 10800 23368
rect 10720 23208 10728 23272
rect 10792 23208 10800 23272
rect 10720 23112 10800 23208
rect 10720 23048 10728 23112
rect 10792 23048 10800 23112
rect 10720 22952 10800 23048
rect 10720 22888 10728 22952
rect 10792 22888 10800 22952
rect 10720 22792 10800 22888
rect 10720 22728 10728 22792
rect 10792 22728 10800 22792
rect 10720 22632 10800 22728
rect 10720 22568 10728 22632
rect 10792 22568 10800 22632
rect 10720 22472 10800 22568
rect 10720 22408 10728 22472
rect 10792 22408 10800 22472
rect 10720 22312 10800 22408
rect 10720 22248 10728 22312
rect 10792 22248 10800 22312
rect 10720 22152 10800 22248
rect 10720 22088 10728 22152
rect 10792 22088 10800 22152
rect 10720 21992 10800 22088
rect 10720 21928 10728 21992
rect 10792 21928 10800 21992
rect 10720 21832 10800 21928
rect 10720 21768 10728 21832
rect 10792 21768 10800 21832
rect 10720 21672 10800 21768
rect 10720 21608 10728 21672
rect 10792 21608 10800 21672
rect 10720 21512 10800 21608
rect 10720 21448 10728 21512
rect 10792 21448 10800 21512
rect 10720 21352 10800 21448
rect 10720 21288 10728 21352
rect 10792 21288 10800 21352
rect 10720 21192 10800 21288
rect 10720 21128 10728 21192
rect 10792 21128 10800 21192
rect 10720 21032 10800 21128
rect 10720 20968 10728 21032
rect 10792 20968 10800 21032
rect 10720 20872 10800 20968
rect 10720 20808 10728 20872
rect 10792 20808 10800 20872
rect 10720 20712 10800 20808
rect 10720 20648 10728 20712
rect 10792 20648 10800 20712
rect 10720 20552 10800 20648
rect 10720 20488 10728 20552
rect 10792 20488 10800 20552
rect 10720 20392 10800 20488
rect 10720 20328 10728 20392
rect 10792 20328 10800 20392
rect 10720 20232 10800 20328
rect 10720 20168 10728 20232
rect 10792 20168 10800 20232
rect 10720 20072 10800 20168
rect 10720 20008 10728 20072
rect 10792 20008 10800 20072
rect 10720 19912 10800 20008
rect 10720 19848 10728 19912
rect 10792 19848 10800 19912
rect 10720 19752 10800 19848
rect 10720 19688 10728 19752
rect 10792 19688 10800 19752
rect 10720 19592 10800 19688
rect 10720 19528 10728 19592
rect 10792 19528 10800 19592
rect 10720 19432 10800 19528
rect 10720 19368 10728 19432
rect 10792 19368 10800 19432
rect 10720 19272 10800 19368
rect 10720 19208 10728 19272
rect 10792 19208 10800 19272
rect 10720 19112 10800 19208
rect 10720 19048 10728 19112
rect 10792 19048 10800 19112
rect 10720 18952 10800 19048
rect 10720 18888 10728 18952
rect 10792 18888 10800 18952
rect 10720 18792 10800 18888
rect 10720 18728 10728 18792
rect 10792 18728 10800 18792
rect 10720 18632 10800 18728
rect 10720 18568 10728 18632
rect 10792 18568 10800 18632
rect 10720 18472 10800 18568
rect 10720 18408 10728 18472
rect 10792 18408 10800 18472
rect 10720 18312 10800 18408
rect 10720 18248 10728 18312
rect 10792 18248 10800 18312
rect 10720 18152 10800 18248
rect 10720 18088 10728 18152
rect 10792 18088 10800 18152
rect 10720 17992 10800 18088
rect 10720 17928 10728 17992
rect 10792 17928 10800 17992
rect 10720 17832 10800 17928
rect 10720 17768 10728 17832
rect 10792 17768 10800 17832
rect 10720 17672 10800 17768
rect 10720 17608 10728 17672
rect 10792 17608 10800 17672
rect 10720 17512 10800 17608
rect 10720 17448 10728 17512
rect 10792 17448 10800 17512
rect 10720 17352 10800 17448
rect 10720 17288 10728 17352
rect 10792 17288 10800 17352
rect 10720 17192 10800 17288
rect 10720 17128 10728 17192
rect 10792 17128 10800 17192
rect 10720 17032 10800 17128
rect 10720 16968 10728 17032
rect 10792 16968 10800 17032
rect 10720 16872 10800 16968
rect 10720 16808 10728 16872
rect 10792 16808 10800 16872
rect 10720 16712 10800 16808
rect 10720 16648 10728 16712
rect 10792 16648 10800 16712
rect 10720 16552 10800 16648
rect 10720 16488 10728 16552
rect 10792 16488 10800 16552
rect 10720 16392 10800 16488
rect 10720 16328 10728 16392
rect 10792 16328 10800 16392
rect 10720 16232 10800 16328
rect 10720 16168 10728 16232
rect 10792 16168 10800 16232
rect 10720 16072 10800 16168
rect 10720 16008 10728 16072
rect 10792 16008 10800 16072
rect 10720 15912 10800 16008
rect 10720 15848 10728 15912
rect 10792 15848 10800 15912
rect 10720 15752 10800 15848
rect 10720 15688 10728 15752
rect 10792 15688 10800 15752
rect 10720 15592 10800 15688
rect 10720 15528 10728 15592
rect 10792 15528 10800 15592
rect 10720 15432 10800 15528
rect 10720 15368 10728 15432
rect 10792 15368 10800 15432
rect 10720 15272 10800 15368
rect 10720 15208 10728 15272
rect 10792 15208 10800 15272
rect 10720 15112 10800 15208
rect 10720 15048 10728 15112
rect 10792 15048 10800 15112
rect 10720 14952 10800 15048
rect 10720 14888 10728 14952
rect 10792 14888 10800 14952
rect 10720 14792 10800 14888
rect 10720 14728 10728 14792
rect 10792 14728 10800 14792
rect 10720 14632 10800 14728
rect 10720 14568 10728 14632
rect 10792 14568 10800 14632
rect 10720 14472 10800 14568
rect 10720 14408 10728 14472
rect 10792 14408 10800 14472
rect 10720 14312 10800 14408
rect 10720 14248 10728 14312
rect 10792 14248 10800 14312
rect 10720 14152 10800 14248
rect 10720 14088 10728 14152
rect 10792 14088 10800 14152
rect 10720 13992 10800 14088
rect 10720 13928 10728 13992
rect 10792 13928 10800 13992
rect 10720 13832 10800 13928
rect 10720 13768 10728 13832
rect 10792 13768 10800 13832
rect 10720 13672 10800 13768
rect 10720 13608 10728 13672
rect 10792 13608 10800 13672
rect 10720 13512 10800 13608
rect 10720 13448 10728 13512
rect 10792 13448 10800 13512
rect 10720 13352 10800 13448
rect 10720 13288 10728 13352
rect 10792 13288 10800 13352
rect 10720 13192 10800 13288
rect 10720 13128 10728 13192
rect 10792 13128 10800 13192
rect 10720 13032 10800 13128
rect 10720 12968 10728 13032
rect 10792 12968 10800 13032
rect 10720 12872 10800 12968
rect 10720 12808 10728 12872
rect 10792 12808 10800 12872
rect 10720 12712 10800 12808
rect 10720 12648 10728 12712
rect 10792 12648 10800 12712
rect 10720 12552 10800 12648
rect 10720 12488 10728 12552
rect 10792 12488 10800 12552
rect 10720 12392 10800 12488
rect 10720 12328 10728 12392
rect 10792 12328 10800 12392
rect 10720 12232 10800 12328
rect 10720 12168 10728 12232
rect 10792 12168 10800 12232
rect 10720 12072 10800 12168
rect 10720 12008 10728 12072
rect 10792 12008 10800 12072
rect 10720 11912 10800 12008
rect 10720 11848 10728 11912
rect 10792 11848 10800 11912
rect 10720 11752 10800 11848
rect 10720 11688 10728 11752
rect 10792 11688 10800 11752
rect 10720 11592 10800 11688
rect 10720 11528 10728 11592
rect 10792 11528 10800 11592
rect 10720 11432 10800 11528
rect 10720 11368 10728 11432
rect 10792 11368 10800 11432
rect 10720 11272 10800 11368
rect 10720 11208 10728 11272
rect 10792 11208 10800 11272
rect 10720 11112 10800 11208
rect 10720 11048 10728 11112
rect 10792 11048 10800 11112
rect 10720 10952 10800 11048
rect 10720 10888 10728 10952
rect 10792 10888 10800 10952
rect 10720 10792 10800 10888
rect 10720 10728 10728 10792
rect 10792 10728 10800 10792
rect 10720 10632 10800 10728
rect 10720 10568 10728 10632
rect 10792 10568 10800 10632
rect 10720 10472 10800 10568
rect 10720 10408 10728 10472
rect 10792 10408 10800 10472
rect 10720 10312 10800 10408
rect 10720 10248 10728 10312
rect 10792 10248 10800 10312
rect 10720 10152 10800 10248
rect 10720 10088 10728 10152
rect 10792 10088 10800 10152
rect 10720 9992 10800 10088
rect 10720 9928 10728 9992
rect 10792 9928 10800 9992
rect 10720 9832 10800 9928
rect 10720 9768 10728 9832
rect 10792 9768 10800 9832
rect 10720 9672 10800 9768
rect 10720 9608 10728 9672
rect 10792 9608 10800 9672
rect 10720 9512 10800 9608
rect 10720 9448 10728 9512
rect 10792 9448 10800 9512
rect 10720 9352 10800 9448
rect 10720 9288 10728 9352
rect 10792 9288 10800 9352
rect 10720 9192 10800 9288
rect 10720 9128 10728 9192
rect 10792 9128 10800 9192
rect 10720 9032 10800 9128
rect 10720 8968 10728 9032
rect 10792 8968 10800 9032
rect 10720 8872 10800 8968
rect 10720 8808 10728 8872
rect 10792 8808 10800 8872
rect 10720 8712 10800 8808
rect 10720 8648 10728 8712
rect 10792 8648 10800 8712
rect 10720 8552 10800 8648
rect 10720 8488 10728 8552
rect 10792 8488 10800 8552
rect 10720 8392 10800 8488
rect 10720 8328 10728 8392
rect 10792 8328 10800 8392
rect 10720 8232 10800 8328
rect 10720 8168 10728 8232
rect 10792 8168 10800 8232
rect 10720 8072 10800 8168
rect 10720 8008 10728 8072
rect 10792 8008 10800 8072
rect 10720 7912 10800 8008
rect 10720 7848 10728 7912
rect 10792 7848 10800 7912
rect 10720 7752 10800 7848
rect 10720 7688 10728 7752
rect 10792 7688 10800 7752
rect 10720 7592 10800 7688
rect 10720 7528 10728 7592
rect 10792 7528 10800 7592
rect 10720 7432 10800 7528
rect 10720 7368 10728 7432
rect 10792 7368 10800 7432
rect 10720 7272 10800 7368
rect 10720 7208 10728 7272
rect 10792 7208 10800 7272
rect 10720 7112 10800 7208
rect 10720 7048 10728 7112
rect 10792 7048 10800 7112
rect 10720 6952 10800 7048
rect 10720 6888 10728 6952
rect 10792 6888 10800 6952
rect 10720 6792 10800 6888
rect 10720 6728 10728 6792
rect 10792 6728 10800 6792
rect 10720 6632 10800 6728
rect 10720 6568 10728 6632
rect 10792 6568 10800 6632
rect 10720 6472 10800 6568
rect 10720 6408 10728 6472
rect 10792 6408 10800 6472
rect 10720 6312 10800 6408
rect 10720 6248 10728 6312
rect 10792 6248 10800 6312
rect 10720 6152 10800 6248
rect 10720 6088 10728 6152
rect 10792 6088 10800 6152
rect 10720 5992 10800 6088
rect 10720 5928 10728 5992
rect 10792 5928 10800 5992
rect 10720 5832 10800 5928
rect 10720 5768 10728 5832
rect 10792 5768 10800 5832
rect 10720 5672 10800 5768
rect 10720 5608 10728 5672
rect 10792 5608 10800 5672
rect 10720 5512 10800 5608
rect 10720 5448 10728 5512
rect 10792 5448 10800 5512
rect 10720 5352 10800 5448
rect 10720 5288 10728 5352
rect 10792 5288 10800 5352
rect 10720 5192 10800 5288
rect 10720 5128 10728 5192
rect 10792 5128 10800 5192
rect 10720 5032 10800 5128
rect 10720 4968 10728 5032
rect 10792 4968 10800 5032
rect 10720 4872 10800 4968
rect 10720 4808 10728 4872
rect 10792 4808 10800 4872
rect 10720 4712 10800 4808
rect 10720 4648 10728 4712
rect 10792 4648 10800 4712
rect 10720 4552 10800 4648
rect 10720 4488 10728 4552
rect 10792 4488 10800 4552
rect 10720 4392 10800 4488
rect 10720 4328 10728 4392
rect 10792 4328 10800 4392
rect 10720 4232 10800 4328
rect 10720 4168 10728 4232
rect 10792 4168 10800 4232
rect 10720 4072 10800 4168
rect 10720 4008 10728 4072
rect 10792 4008 10800 4072
rect 10720 3912 10800 4008
rect 10720 3848 10728 3912
rect 10792 3848 10800 3912
rect 10720 3752 10800 3848
rect 10720 3688 10728 3752
rect 10792 3688 10800 3752
rect 10720 3592 10800 3688
rect 10720 3528 10728 3592
rect 10792 3528 10800 3592
rect 10720 3432 10800 3528
rect 10720 3368 10728 3432
rect 10792 3368 10800 3432
rect 10720 3272 10800 3368
rect 10720 3208 10728 3272
rect 10792 3208 10800 3272
rect 10720 3112 10800 3208
rect 10720 3048 10728 3112
rect 10792 3048 10800 3112
rect 10720 2952 10800 3048
rect 10720 2888 10728 2952
rect 10792 2888 10800 2952
rect 10720 2792 10800 2888
rect 10720 2728 10728 2792
rect 10792 2728 10800 2792
rect 10720 2632 10800 2728
rect 10720 2568 10728 2632
rect 10792 2568 10800 2632
rect 10720 2472 10800 2568
rect 10720 2408 10728 2472
rect 10792 2408 10800 2472
rect 10720 2312 10800 2408
rect 10720 2248 10728 2312
rect 10792 2248 10800 2312
rect 10720 2152 10800 2248
rect 10720 2088 10728 2152
rect 10792 2088 10800 2152
rect 10720 1992 10800 2088
rect 10720 1928 10728 1992
rect 10792 1928 10800 1992
rect 10720 1832 10800 1928
rect 10720 1768 10728 1832
rect 10792 1768 10800 1832
rect 10720 1672 10800 1768
rect 10720 1608 10728 1672
rect 10792 1608 10800 1672
rect 10720 1512 10800 1608
rect 10720 1448 10728 1512
rect 10792 1448 10800 1512
rect 10720 1352 10800 1448
rect 10720 1288 10728 1352
rect 10792 1288 10800 1352
rect 10720 1192 10800 1288
rect 10720 1128 10728 1192
rect 10792 1128 10800 1192
rect 10720 1032 10800 1128
rect 10720 968 10728 1032
rect 10792 968 10800 1032
rect 10720 872 10800 968
rect 10720 808 10728 872
rect 10792 808 10800 872
rect 10720 712 10800 808
rect 10720 648 10728 712
rect 10792 648 10800 712
rect 10720 552 10800 648
rect 10720 488 10728 552
rect 10792 488 10800 552
rect 10720 392 10800 488
rect 10720 328 10728 392
rect 10792 328 10800 392
rect 10720 232 10800 328
rect 10720 168 10728 232
rect 10792 168 10800 232
rect 10720 72 10800 168
rect 10720 8 10728 72
rect 10792 8 10800 72
rect 10400 -1112 10408 -1048
rect 10472 -1112 10480 -1048
rect 10400 -1128 10480 -1112
rect 10400 -1192 10408 -1128
rect 10472 -1192 10480 -1128
rect 10400 -1208 10480 -1192
rect 10400 -1272 10408 -1208
rect 10472 -1272 10480 -1208
rect 10400 -1288 10480 -1272
rect 10400 -1352 10408 -1288
rect 10472 -1352 10480 -1288
rect 10400 -1368 10480 -1352
rect 10400 -1432 10408 -1368
rect 10472 -1432 10480 -1368
rect 10400 -1920 10480 -1432
rect 10720 -1048 10800 8
rect 10880 28308 10960 31520
rect 10880 28252 10892 28308
rect 10948 28252 10960 28308
rect 10880 18228 10960 28252
rect 10880 18172 10892 18228
rect 10948 18172 10960 18228
rect 10880 11988 10960 18172
rect 10880 11932 10892 11988
rect 10948 11932 10960 11988
rect 10880 0 10960 11932
rect 11040 31432 11120 31520
rect 11040 31368 11048 31432
rect 11112 31368 11120 31432
rect 11040 31272 11120 31368
rect 11040 31208 11048 31272
rect 11112 31208 11120 31272
rect 11040 31112 11120 31208
rect 11040 31048 11048 31112
rect 11112 31048 11120 31112
rect 11040 30952 11120 31048
rect 11040 30888 11048 30952
rect 11112 30888 11120 30952
rect 11040 30792 11120 30888
rect 11040 30728 11048 30792
rect 11112 30728 11120 30792
rect 11040 30632 11120 30728
rect 11040 30568 11048 30632
rect 11112 30568 11120 30632
rect 11040 30472 11120 30568
rect 11040 30408 11048 30472
rect 11112 30408 11120 30472
rect 11040 30312 11120 30408
rect 11040 30248 11048 30312
rect 11112 30248 11120 30312
rect 11040 30152 11120 30248
rect 11040 30088 11048 30152
rect 11112 30088 11120 30152
rect 11040 29992 11120 30088
rect 11040 29928 11048 29992
rect 11112 29928 11120 29992
rect 11040 29832 11120 29928
rect 11040 29768 11048 29832
rect 11112 29768 11120 29832
rect 11040 29672 11120 29768
rect 11040 29608 11048 29672
rect 11112 29608 11120 29672
rect 11040 29512 11120 29608
rect 11040 29448 11048 29512
rect 11112 29448 11120 29512
rect 11040 29352 11120 29448
rect 11040 29288 11048 29352
rect 11112 29288 11120 29352
rect 11040 29192 11120 29288
rect 11040 29128 11048 29192
rect 11112 29128 11120 29192
rect 11040 29032 11120 29128
rect 11040 28968 11048 29032
rect 11112 28968 11120 29032
rect 11040 28872 11120 28968
rect 11040 28808 11048 28872
rect 11112 28808 11120 28872
rect 11040 28712 11120 28808
rect 11040 28648 11048 28712
rect 11112 28648 11120 28712
rect 11040 28552 11120 28648
rect 11040 28488 11048 28552
rect 11112 28488 11120 28552
rect 11040 28392 11120 28488
rect 11040 28328 11048 28392
rect 11112 28328 11120 28392
rect 11040 28232 11120 28328
rect 11040 28168 11048 28232
rect 11112 28168 11120 28232
rect 11040 28072 11120 28168
rect 11040 28008 11048 28072
rect 11112 28008 11120 28072
rect 11040 27912 11120 28008
rect 11040 27848 11048 27912
rect 11112 27848 11120 27912
rect 11040 27752 11120 27848
rect 11040 27688 11048 27752
rect 11112 27688 11120 27752
rect 11040 27592 11120 27688
rect 11040 27528 11048 27592
rect 11112 27528 11120 27592
rect 11040 27432 11120 27528
rect 11040 27368 11048 27432
rect 11112 27368 11120 27432
rect 11040 27272 11120 27368
rect 11040 27208 11048 27272
rect 11112 27208 11120 27272
rect 11040 27112 11120 27208
rect 11040 27048 11048 27112
rect 11112 27048 11120 27112
rect 11040 26952 11120 27048
rect 11040 26888 11048 26952
rect 11112 26888 11120 26952
rect 11040 26792 11120 26888
rect 11040 26728 11048 26792
rect 11112 26728 11120 26792
rect 11040 26632 11120 26728
rect 11040 26568 11048 26632
rect 11112 26568 11120 26632
rect 11040 26472 11120 26568
rect 11040 26408 11048 26472
rect 11112 26408 11120 26472
rect 11040 26312 11120 26408
rect 11040 26248 11048 26312
rect 11112 26248 11120 26312
rect 11040 26152 11120 26248
rect 11040 26088 11048 26152
rect 11112 26088 11120 26152
rect 11040 25992 11120 26088
rect 11040 25928 11048 25992
rect 11112 25928 11120 25992
rect 11040 25832 11120 25928
rect 11040 25768 11048 25832
rect 11112 25768 11120 25832
rect 11040 25672 11120 25768
rect 11040 25608 11048 25672
rect 11112 25608 11120 25672
rect 11040 25512 11120 25608
rect 11040 25448 11048 25512
rect 11112 25448 11120 25512
rect 11040 25352 11120 25448
rect 11040 25288 11048 25352
rect 11112 25288 11120 25352
rect 11040 25192 11120 25288
rect 11040 25128 11048 25192
rect 11112 25128 11120 25192
rect 11040 25032 11120 25128
rect 11040 24968 11048 25032
rect 11112 24968 11120 25032
rect 11040 24872 11120 24968
rect 11040 24808 11048 24872
rect 11112 24808 11120 24872
rect 11040 24712 11120 24808
rect 11040 24648 11048 24712
rect 11112 24648 11120 24712
rect 11040 24552 11120 24648
rect 11040 24488 11048 24552
rect 11112 24488 11120 24552
rect 11040 24392 11120 24488
rect 11040 24328 11048 24392
rect 11112 24328 11120 24392
rect 11040 24232 11120 24328
rect 11040 24168 11048 24232
rect 11112 24168 11120 24232
rect 11040 24072 11120 24168
rect 11040 24008 11048 24072
rect 11112 24008 11120 24072
rect 11040 23912 11120 24008
rect 11040 23848 11048 23912
rect 11112 23848 11120 23912
rect 11040 23752 11120 23848
rect 11040 23688 11048 23752
rect 11112 23688 11120 23752
rect 11040 23592 11120 23688
rect 11040 23528 11048 23592
rect 11112 23528 11120 23592
rect 11040 23432 11120 23528
rect 11040 23368 11048 23432
rect 11112 23368 11120 23432
rect 11040 23272 11120 23368
rect 11040 23208 11048 23272
rect 11112 23208 11120 23272
rect 11040 23112 11120 23208
rect 11040 23048 11048 23112
rect 11112 23048 11120 23112
rect 11040 22952 11120 23048
rect 11040 22888 11048 22952
rect 11112 22888 11120 22952
rect 11040 22792 11120 22888
rect 11040 22728 11048 22792
rect 11112 22728 11120 22792
rect 11040 22632 11120 22728
rect 11040 22568 11048 22632
rect 11112 22568 11120 22632
rect 11040 22472 11120 22568
rect 11040 22408 11048 22472
rect 11112 22408 11120 22472
rect 11040 22312 11120 22408
rect 11040 22248 11048 22312
rect 11112 22248 11120 22312
rect 11040 22152 11120 22248
rect 11040 22088 11048 22152
rect 11112 22088 11120 22152
rect 11040 21992 11120 22088
rect 11040 21928 11048 21992
rect 11112 21928 11120 21992
rect 11040 21832 11120 21928
rect 11040 21768 11048 21832
rect 11112 21768 11120 21832
rect 11040 21672 11120 21768
rect 11040 21608 11048 21672
rect 11112 21608 11120 21672
rect 11040 21512 11120 21608
rect 11040 21448 11048 21512
rect 11112 21448 11120 21512
rect 11040 21352 11120 21448
rect 11040 21288 11048 21352
rect 11112 21288 11120 21352
rect 11040 21192 11120 21288
rect 11040 21128 11048 21192
rect 11112 21128 11120 21192
rect 11040 21032 11120 21128
rect 11040 20968 11048 21032
rect 11112 20968 11120 21032
rect 11040 20872 11120 20968
rect 11040 20808 11048 20872
rect 11112 20808 11120 20872
rect 11040 20712 11120 20808
rect 11040 20648 11048 20712
rect 11112 20648 11120 20712
rect 11040 20552 11120 20648
rect 11040 20488 11048 20552
rect 11112 20488 11120 20552
rect 11040 20392 11120 20488
rect 11040 20328 11048 20392
rect 11112 20328 11120 20392
rect 11040 20232 11120 20328
rect 11040 20168 11048 20232
rect 11112 20168 11120 20232
rect 11040 20072 11120 20168
rect 11040 20008 11048 20072
rect 11112 20008 11120 20072
rect 11040 19912 11120 20008
rect 11040 19848 11048 19912
rect 11112 19848 11120 19912
rect 11040 19752 11120 19848
rect 11040 19688 11048 19752
rect 11112 19688 11120 19752
rect 11040 19592 11120 19688
rect 11040 19528 11048 19592
rect 11112 19528 11120 19592
rect 11040 19432 11120 19528
rect 11040 19368 11048 19432
rect 11112 19368 11120 19432
rect 11040 19272 11120 19368
rect 11040 19208 11048 19272
rect 11112 19208 11120 19272
rect 11040 19112 11120 19208
rect 11040 19048 11048 19112
rect 11112 19048 11120 19112
rect 11040 18952 11120 19048
rect 11040 18888 11048 18952
rect 11112 18888 11120 18952
rect 11040 18792 11120 18888
rect 11040 18728 11048 18792
rect 11112 18728 11120 18792
rect 11040 18632 11120 18728
rect 11040 18568 11048 18632
rect 11112 18568 11120 18632
rect 11040 18472 11120 18568
rect 11040 18408 11048 18472
rect 11112 18408 11120 18472
rect 11040 18312 11120 18408
rect 11040 18248 11048 18312
rect 11112 18248 11120 18312
rect 11040 18152 11120 18248
rect 11040 18088 11048 18152
rect 11112 18088 11120 18152
rect 11040 17992 11120 18088
rect 11040 17928 11048 17992
rect 11112 17928 11120 17992
rect 11040 17832 11120 17928
rect 11040 17768 11048 17832
rect 11112 17768 11120 17832
rect 11040 17672 11120 17768
rect 11040 17608 11048 17672
rect 11112 17608 11120 17672
rect 11040 17512 11120 17608
rect 11040 17448 11048 17512
rect 11112 17448 11120 17512
rect 11040 17352 11120 17448
rect 11040 17288 11048 17352
rect 11112 17288 11120 17352
rect 11040 17192 11120 17288
rect 11040 17128 11048 17192
rect 11112 17128 11120 17192
rect 11040 17032 11120 17128
rect 11040 16968 11048 17032
rect 11112 16968 11120 17032
rect 11040 16872 11120 16968
rect 11040 16808 11048 16872
rect 11112 16808 11120 16872
rect 11040 16712 11120 16808
rect 11040 16648 11048 16712
rect 11112 16648 11120 16712
rect 11040 16552 11120 16648
rect 11040 16488 11048 16552
rect 11112 16488 11120 16552
rect 11040 16392 11120 16488
rect 11040 16328 11048 16392
rect 11112 16328 11120 16392
rect 11040 16232 11120 16328
rect 11040 16168 11048 16232
rect 11112 16168 11120 16232
rect 11040 16072 11120 16168
rect 11040 16008 11048 16072
rect 11112 16008 11120 16072
rect 11040 15912 11120 16008
rect 11040 15848 11048 15912
rect 11112 15848 11120 15912
rect 11040 15752 11120 15848
rect 11040 15688 11048 15752
rect 11112 15688 11120 15752
rect 11040 15592 11120 15688
rect 11040 15528 11048 15592
rect 11112 15528 11120 15592
rect 11040 15432 11120 15528
rect 11040 15368 11048 15432
rect 11112 15368 11120 15432
rect 11040 15272 11120 15368
rect 11040 15208 11048 15272
rect 11112 15208 11120 15272
rect 11040 15112 11120 15208
rect 11040 15048 11048 15112
rect 11112 15048 11120 15112
rect 11040 14952 11120 15048
rect 11040 14888 11048 14952
rect 11112 14888 11120 14952
rect 11040 14792 11120 14888
rect 11040 14728 11048 14792
rect 11112 14728 11120 14792
rect 11040 14632 11120 14728
rect 11040 14568 11048 14632
rect 11112 14568 11120 14632
rect 11040 14472 11120 14568
rect 11040 14408 11048 14472
rect 11112 14408 11120 14472
rect 11040 14312 11120 14408
rect 11040 14248 11048 14312
rect 11112 14248 11120 14312
rect 11040 14152 11120 14248
rect 11040 14088 11048 14152
rect 11112 14088 11120 14152
rect 11040 13992 11120 14088
rect 11040 13928 11048 13992
rect 11112 13928 11120 13992
rect 11040 13832 11120 13928
rect 11040 13768 11048 13832
rect 11112 13768 11120 13832
rect 11040 13672 11120 13768
rect 11040 13608 11048 13672
rect 11112 13608 11120 13672
rect 11040 13512 11120 13608
rect 11040 13448 11048 13512
rect 11112 13448 11120 13512
rect 11040 13352 11120 13448
rect 11040 13288 11048 13352
rect 11112 13288 11120 13352
rect 11040 13192 11120 13288
rect 11040 13128 11048 13192
rect 11112 13128 11120 13192
rect 11040 13032 11120 13128
rect 11040 12968 11048 13032
rect 11112 12968 11120 13032
rect 11040 12872 11120 12968
rect 11040 12808 11048 12872
rect 11112 12808 11120 12872
rect 11040 12712 11120 12808
rect 11040 12648 11048 12712
rect 11112 12648 11120 12712
rect 11040 12552 11120 12648
rect 11040 12488 11048 12552
rect 11112 12488 11120 12552
rect 11040 12392 11120 12488
rect 11040 12328 11048 12392
rect 11112 12328 11120 12392
rect 11040 12232 11120 12328
rect 11040 12168 11048 12232
rect 11112 12168 11120 12232
rect 11040 12072 11120 12168
rect 11040 12008 11048 12072
rect 11112 12008 11120 12072
rect 11040 11912 11120 12008
rect 11040 11848 11048 11912
rect 11112 11848 11120 11912
rect 11040 11752 11120 11848
rect 11040 11688 11048 11752
rect 11112 11688 11120 11752
rect 11040 11592 11120 11688
rect 11040 11528 11048 11592
rect 11112 11528 11120 11592
rect 11040 11432 11120 11528
rect 11040 11368 11048 11432
rect 11112 11368 11120 11432
rect 11040 11272 11120 11368
rect 11040 11208 11048 11272
rect 11112 11208 11120 11272
rect 11040 11112 11120 11208
rect 11040 11048 11048 11112
rect 11112 11048 11120 11112
rect 11040 10952 11120 11048
rect 11040 10888 11048 10952
rect 11112 10888 11120 10952
rect 11040 10792 11120 10888
rect 11040 10728 11048 10792
rect 11112 10728 11120 10792
rect 11040 10632 11120 10728
rect 11040 10568 11048 10632
rect 11112 10568 11120 10632
rect 11040 10472 11120 10568
rect 11040 10408 11048 10472
rect 11112 10408 11120 10472
rect 11040 10312 11120 10408
rect 11040 10248 11048 10312
rect 11112 10248 11120 10312
rect 11040 10152 11120 10248
rect 11040 10088 11048 10152
rect 11112 10088 11120 10152
rect 11040 9992 11120 10088
rect 11040 9928 11048 9992
rect 11112 9928 11120 9992
rect 11040 9832 11120 9928
rect 11040 9768 11048 9832
rect 11112 9768 11120 9832
rect 11040 9672 11120 9768
rect 11040 9608 11048 9672
rect 11112 9608 11120 9672
rect 11040 9512 11120 9608
rect 11040 9448 11048 9512
rect 11112 9448 11120 9512
rect 11040 9352 11120 9448
rect 11040 9288 11048 9352
rect 11112 9288 11120 9352
rect 11040 9192 11120 9288
rect 11040 9128 11048 9192
rect 11112 9128 11120 9192
rect 11040 9032 11120 9128
rect 11040 8968 11048 9032
rect 11112 8968 11120 9032
rect 11040 8872 11120 8968
rect 11040 8808 11048 8872
rect 11112 8808 11120 8872
rect 11040 8712 11120 8808
rect 11040 8648 11048 8712
rect 11112 8648 11120 8712
rect 11040 8552 11120 8648
rect 11040 8488 11048 8552
rect 11112 8488 11120 8552
rect 11040 8392 11120 8488
rect 11040 8328 11048 8392
rect 11112 8328 11120 8392
rect 11040 8232 11120 8328
rect 11040 8168 11048 8232
rect 11112 8168 11120 8232
rect 11040 8072 11120 8168
rect 11040 8008 11048 8072
rect 11112 8008 11120 8072
rect 11040 7912 11120 8008
rect 11040 7848 11048 7912
rect 11112 7848 11120 7912
rect 11040 7752 11120 7848
rect 11040 7688 11048 7752
rect 11112 7688 11120 7752
rect 11040 7592 11120 7688
rect 11040 7528 11048 7592
rect 11112 7528 11120 7592
rect 11040 7432 11120 7528
rect 11040 7368 11048 7432
rect 11112 7368 11120 7432
rect 11040 7272 11120 7368
rect 11040 7208 11048 7272
rect 11112 7208 11120 7272
rect 11040 7112 11120 7208
rect 11040 7048 11048 7112
rect 11112 7048 11120 7112
rect 11040 6952 11120 7048
rect 11040 6888 11048 6952
rect 11112 6888 11120 6952
rect 11040 6792 11120 6888
rect 11040 6728 11048 6792
rect 11112 6728 11120 6792
rect 11040 6632 11120 6728
rect 11040 6568 11048 6632
rect 11112 6568 11120 6632
rect 11040 6472 11120 6568
rect 11040 6408 11048 6472
rect 11112 6408 11120 6472
rect 11040 6312 11120 6408
rect 11040 6248 11048 6312
rect 11112 6248 11120 6312
rect 11040 6152 11120 6248
rect 11040 6088 11048 6152
rect 11112 6088 11120 6152
rect 11040 5992 11120 6088
rect 11040 5928 11048 5992
rect 11112 5928 11120 5992
rect 11040 5832 11120 5928
rect 11040 5768 11048 5832
rect 11112 5768 11120 5832
rect 11040 5672 11120 5768
rect 11040 5608 11048 5672
rect 11112 5608 11120 5672
rect 11040 5512 11120 5608
rect 11040 5448 11048 5512
rect 11112 5448 11120 5512
rect 11040 5352 11120 5448
rect 11040 5288 11048 5352
rect 11112 5288 11120 5352
rect 11040 5192 11120 5288
rect 11040 5128 11048 5192
rect 11112 5128 11120 5192
rect 11040 5032 11120 5128
rect 11040 4968 11048 5032
rect 11112 4968 11120 5032
rect 11040 4872 11120 4968
rect 11040 4808 11048 4872
rect 11112 4808 11120 4872
rect 11040 4712 11120 4808
rect 11040 4648 11048 4712
rect 11112 4648 11120 4712
rect 11040 4552 11120 4648
rect 11040 4488 11048 4552
rect 11112 4488 11120 4552
rect 11040 4392 11120 4488
rect 11040 4328 11048 4392
rect 11112 4328 11120 4392
rect 11040 4232 11120 4328
rect 11040 4168 11048 4232
rect 11112 4168 11120 4232
rect 11040 4072 11120 4168
rect 11040 4008 11048 4072
rect 11112 4008 11120 4072
rect 11040 3912 11120 4008
rect 11040 3848 11048 3912
rect 11112 3848 11120 3912
rect 11040 3752 11120 3848
rect 11040 3688 11048 3752
rect 11112 3688 11120 3752
rect 11040 3592 11120 3688
rect 11040 3528 11048 3592
rect 11112 3528 11120 3592
rect 11040 3432 11120 3528
rect 11040 3368 11048 3432
rect 11112 3368 11120 3432
rect 11040 3272 11120 3368
rect 11040 3208 11048 3272
rect 11112 3208 11120 3272
rect 11040 3112 11120 3208
rect 11040 3048 11048 3112
rect 11112 3048 11120 3112
rect 11040 2952 11120 3048
rect 11040 2888 11048 2952
rect 11112 2888 11120 2952
rect 11040 2792 11120 2888
rect 11040 2728 11048 2792
rect 11112 2728 11120 2792
rect 11040 2632 11120 2728
rect 11040 2568 11048 2632
rect 11112 2568 11120 2632
rect 11040 2472 11120 2568
rect 11040 2408 11048 2472
rect 11112 2408 11120 2472
rect 11040 2312 11120 2408
rect 11040 2248 11048 2312
rect 11112 2248 11120 2312
rect 11040 2152 11120 2248
rect 11040 2088 11048 2152
rect 11112 2088 11120 2152
rect 11040 1992 11120 2088
rect 11040 1928 11048 1992
rect 11112 1928 11120 1992
rect 11040 1832 11120 1928
rect 11040 1768 11048 1832
rect 11112 1768 11120 1832
rect 11040 1672 11120 1768
rect 11040 1608 11048 1672
rect 11112 1608 11120 1672
rect 11040 1512 11120 1608
rect 11040 1448 11048 1512
rect 11112 1448 11120 1512
rect 11040 1352 11120 1448
rect 11040 1288 11048 1352
rect 11112 1288 11120 1352
rect 11040 1192 11120 1288
rect 11040 1128 11048 1192
rect 11112 1128 11120 1192
rect 11040 1032 11120 1128
rect 11040 968 11048 1032
rect 11112 968 11120 1032
rect 11040 872 11120 968
rect 11040 808 11048 872
rect 11112 808 11120 872
rect 11040 712 11120 808
rect 11040 648 11048 712
rect 11112 648 11120 712
rect 11040 552 11120 648
rect 11040 488 11048 552
rect 11112 488 11120 552
rect 11040 392 11120 488
rect 11040 328 11048 392
rect 11112 328 11120 392
rect 11040 232 11120 328
rect 11040 168 11048 232
rect 11112 168 11120 232
rect 11040 72 11120 168
rect 11040 8 11048 72
rect 11112 8 11120 72
rect 10720 -1112 10728 -1048
rect 10792 -1112 10800 -1048
rect 10720 -1128 10800 -1112
rect 10720 -1192 10728 -1128
rect 10792 -1192 10800 -1128
rect 10720 -1208 10800 -1192
rect 10720 -1272 10728 -1208
rect 10792 -1272 10800 -1208
rect 10720 -1288 10800 -1272
rect 10720 -1352 10728 -1288
rect 10792 -1352 10800 -1288
rect 10720 -1368 10800 -1352
rect 10720 -1432 10728 -1368
rect 10792 -1432 10800 -1368
rect 10720 -1920 10800 -1432
rect 11040 -1048 11120 8
rect 11200 12308 11280 31520
rect 11200 12252 11212 12308
rect 11268 12252 11280 12308
rect 11200 0 11280 12252
rect 11360 31432 11440 31520
rect 11360 31368 11368 31432
rect 11432 31368 11440 31432
rect 11360 31272 11440 31368
rect 11360 31208 11368 31272
rect 11432 31208 11440 31272
rect 11360 31112 11440 31208
rect 11360 31048 11368 31112
rect 11432 31048 11440 31112
rect 11360 30952 11440 31048
rect 11360 30888 11368 30952
rect 11432 30888 11440 30952
rect 11360 30792 11440 30888
rect 11360 30728 11368 30792
rect 11432 30728 11440 30792
rect 11360 30632 11440 30728
rect 11360 30568 11368 30632
rect 11432 30568 11440 30632
rect 11360 30472 11440 30568
rect 11360 30408 11368 30472
rect 11432 30408 11440 30472
rect 11360 30312 11440 30408
rect 11360 30248 11368 30312
rect 11432 30248 11440 30312
rect 11360 30152 11440 30248
rect 11360 30088 11368 30152
rect 11432 30088 11440 30152
rect 11360 29992 11440 30088
rect 11360 29928 11368 29992
rect 11432 29928 11440 29992
rect 11360 29832 11440 29928
rect 11360 29768 11368 29832
rect 11432 29768 11440 29832
rect 11360 29672 11440 29768
rect 11360 29608 11368 29672
rect 11432 29608 11440 29672
rect 11360 29512 11440 29608
rect 11360 29448 11368 29512
rect 11432 29448 11440 29512
rect 11360 29352 11440 29448
rect 11360 29288 11368 29352
rect 11432 29288 11440 29352
rect 11360 29192 11440 29288
rect 11360 29128 11368 29192
rect 11432 29128 11440 29192
rect 11360 29032 11440 29128
rect 11360 28968 11368 29032
rect 11432 28968 11440 29032
rect 11360 28872 11440 28968
rect 11360 28808 11368 28872
rect 11432 28808 11440 28872
rect 11360 28712 11440 28808
rect 11360 28648 11368 28712
rect 11432 28648 11440 28712
rect 11360 28552 11440 28648
rect 11360 28488 11368 28552
rect 11432 28488 11440 28552
rect 11360 28392 11440 28488
rect 11360 28328 11368 28392
rect 11432 28328 11440 28392
rect 11360 28232 11440 28328
rect 11360 28168 11368 28232
rect 11432 28168 11440 28232
rect 11360 28072 11440 28168
rect 11360 28008 11368 28072
rect 11432 28008 11440 28072
rect 11360 27912 11440 28008
rect 11360 27848 11368 27912
rect 11432 27848 11440 27912
rect 11360 27752 11440 27848
rect 11360 27688 11368 27752
rect 11432 27688 11440 27752
rect 11360 27592 11440 27688
rect 11360 27528 11368 27592
rect 11432 27528 11440 27592
rect 11360 27432 11440 27528
rect 11360 27368 11368 27432
rect 11432 27368 11440 27432
rect 11360 27272 11440 27368
rect 11360 27208 11368 27272
rect 11432 27208 11440 27272
rect 11360 27112 11440 27208
rect 11360 27048 11368 27112
rect 11432 27048 11440 27112
rect 11360 26952 11440 27048
rect 11360 26888 11368 26952
rect 11432 26888 11440 26952
rect 11360 26792 11440 26888
rect 11360 26728 11368 26792
rect 11432 26728 11440 26792
rect 11360 26632 11440 26728
rect 11360 26568 11368 26632
rect 11432 26568 11440 26632
rect 11360 26472 11440 26568
rect 11360 26408 11368 26472
rect 11432 26408 11440 26472
rect 11360 26312 11440 26408
rect 11360 26248 11368 26312
rect 11432 26248 11440 26312
rect 11360 26152 11440 26248
rect 11360 26088 11368 26152
rect 11432 26088 11440 26152
rect 11360 25992 11440 26088
rect 11360 25928 11368 25992
rect 11432 25928 11440 25992
rect 11360 25832 11440 25928
rect 11360 25768 11368 25832
rect 11432 25768 11440 25832
rect 11360 25672 11440 25768
rect 11360 25608 11368 25672
rect 11432 25608 11440 25672
rect 11360 25512 11440 25608
rect 11360 25448 11368 25512
rect 11432 25448 11440 25512
rect 11360 25352 11440 25448
rect 11360 25288 11368 25352
rect 11432 25288 11440 25352
rect 11360 25192 11440 25288
rect 11360 25128 11368 25192
rect 11432 25128 11440 25192
rect 11360 25032 11440 25128
rect 11360 24968 11368 25032
rect 11432 24968 11440 25032
rect 11360 24872 11440 24968
rect 11360 24808 11368 24872
rect 11432 24808 11440 24872
rect 11360 24712 11440 24808
rect 11360 24648 11368 24712
rect 11432 24648 11440 24712
rect 11360 24552 11440 24648
rect 11360 24488 11368 24552
rect 11432 24488 11440 24552
rect 11360 24392 11440 24488
rect 11360 24328 11368 24392
rect 11432 24328 11440 24392
rect 11360 24232 11440 24328
rect 11360 24168 11368 24232
rect 11432 24168 11440 24232
rect 11360 24072 11440 24168
rect 11360 24008 11368 24072
rect 11432 24008 11440 24072
rect 11360 23912 11440 24008
rect 11360 23848 11368 23912
rect 11432 23848 11440 23912
rect 11360 23752 11440 23848
rect 11360 23688 11368 23752
rect 11432 23688 11440 23752
rect 11360 23592 11440 23688
rect 11360 23528 11368 23592
rect 11432 23528 11440 23592
rect 11360 23432 11440 23528
rect 11360 23368 11368 23432
rect 11432 23368 11440 23432
rect 11360 23272 11440 23368
rect 11360 23208 11368 23272
rect 11432 23208 11440 23272
rect 11360 23112 11440 23208
rect 11360 23048 11368 23112
rect 11432 23048 11440 23112
rect 11360 22952 11440 23048
rect 11360 22888 11368 22952
rect 11432 22888 11440 22952
rect 11360 22792 11440 22888
rect 11360 22728 11368 22792
rect 11432 22728 11440 22792
rect 11360 22632 11440 22728
rect 11360 22568 11368 22632
rect 11432 22568 11440 22632
rect 11360 22472 11440 22568
rect 11360 22408 11368 22472
rect 11432 22408 11440 22472
rect 11360 22312 11440 22408
rect 11360 22248 11368 22312
rect 11432 22248 11440 22312
rect 11360 22152 11440 22248
rect 11360 22088 11368 22152
rect 11432 22088 11440 22152
rect 11360 21992 11440 22088
rect 11360 21928 11368 21992
rect 11432 21928 11440 21992
rect 11360 21832 11440 21928
rect 11360 21768 11368 21832
rect 11432 21768 11440 21832
rect 11360 21672 11440 21768
rect 11360 21608 11368 21672
rect 11432 21608 11440 21672
rect 11360 21512 11440 21608
rect 11360 21448 11368 21512
rect 11432 21448 11440 21512
rect 11360 21352 11440 21448
rect 11360 21288 11368 21352
rect 11432 21288 11440 21352
rect 11360 21192 11440 21288
rect 11360 21128 11368 21192
rect 11432 21128 11440 21192
rect 11360 21032 11440 21128
rect 11360 20968 11368 21032
rect 11432 20968 11440 21032
rect 11360 20872 11440 20968
rect 11360 20808 11368 20872
rect 11432 20808 11440 20872
rect 11360 20712 11440 20808
rect 11360 20648 11368 20712
rect 11432 20648 11440 20712
rect 11360 20552 11440 20648
rect 11360 20488 11368 20552
rect 11432 20488 11440 20552
rect 11360 20392 11440 20488
rect 11360 20328 11368 20392
rect 11432 20328 11440 20392
rect 11360 20232 11440 20328
rect 11360 20168 11368 20232
rect 11432 20168 11440 20232
rect 11360 20072 11440 20168
rect 11360 20008 11368 20072
rect 11432 20008 11440 20072
rect 11360 19912 11440 20008
rect 11360 19848 11368 19912
rect 11432 19848 11440 19912
rect 11360 19752 11440 19848
rect 11360 19688 11368 19752
rect 11432 19688 11440 19752
rect 11360 19592 11440 19688
rect 11360 19528 11368 19592
rect 11432 19528 11440 19592
rect 11360 19432 11440 19528
rect 11360 19368 11368 19432
rect 11432 19368 11440 19432
rect 11360 19272 11440 19368
rect 11360 19208 11368 19272
rect 11432 19208 11440 19272
rect 11360 19112 11440 19208
rect 11360 19048 11368 19112
rect 11432 19048 11440 19112
rect 11360 18952 11440 19048
rect 11360 18888 11368 18952
rect 11432 18888 11440 18952
rect 11360 18792 11440 18888
rect 11360 18728 11368 18792
rect 11432 18728 11440 18792
rect 11360 18632 11440 18728
rect 11360 18568 11368 18632
rect 11432 18568 11440 18632
rect 11360 18472 11440 18568
rect 11360 18408 11368 18472
rect 11432 18408 11440 18472
rect 11360 18312 11440 18408
rect 11360 18248 11368 18312
rect 11432 18248 11440 18312
rect 11360 18152 11440 18248
rect 11360 18088 11368 18152
rect 11432 18088 11440 18152
rect 11360 17992 11440 18088
rect 11360 17928 11368 17992
rect 11432 17928 11440 17992
rect 11360 17832 11440 17928
rect 11360 17768 11368 17832
rect 11432 17768 11440 17832
rect 11360 17672 11440 17768
rect 11360 17608 11368 17672
rect 11432 17608 11440 17672
rect 11360 17512 11440 17608
rect 11360 17448 11368 17512
rect 11432 17448 11440 17512
rect 11360 17352 11440 17448
rect 11360 17288 11368 17352
rect 11432 17288 11440 17352
rect 11360 17192 11440 17288
rect 11360 17128 11368 17192
rect 11432 17128 11440 17192
rect 11360 17032 11440 17128
rect 11360 16968 11368 17032
rect 11432 16968 11440 17032
rect 11360 16872 11440 16968
rect 11360 16808 11368 16872
rect 11432 16808 11440 16872
rect 11360 16712 11440 16808
rect 11360 16648 11368 16712
rect 11432 16648 11440 16712
rect 11360 16552 11440 16648
rect 11360 16488 11368 16552
rect 11432 16488 11440 16552
rect 11360 16392 11440 16488
rect 11360 16328 11368 16392
rect 11432 16328 11440 16392
rect 11360 16232 11440 16328
rect 11360 16168 11368 16232
rect 11432 16168 11440 16232
rect 11360 16072 11440 16168
rect 11360 16008 11368 16072
rect 11432 16008 11440 16072
rect 11360 15912 11440 16008
rect 11360 15848 11368 15912
rect 11432 15848 11440 15912
rect 11360 15752 11440 15848
rect 11360 15688 11368 15752
rect 11432 15688 11440 15752
rect 11360 15592 11440 15688
rect 11360 15528 11368 15592
rect 11432 15528 11440 15592
rect 11360 15432 11440 15528
rect 11360 15368 11368 15432
rect 11432 15368 11440 15432
rect 11360 15272 11440 15368
rect 11360 15208 11368 15272
rect 11432 15208 11440 15272
rect 11360 15112 11440 15208
rect 11360 15048 11368 15112
rect 11432 15048 11440 15112
rect 11360 14952 11440 15048
rect 11360 14888 11368 14952
rect 11432 14888 11440 14952
rect 11360 14792 11440 14888
rect 11360 14728 11368 14792
rect 11432 14728 11440 14792
rect 11360 14632 11440 14728
rect 11360 14568 11368 14632
rect 11432 14568 11440 14632
rect 11360 14472 11440 14568
rect 11360 14408 11368 14472
rect 11432 14408 11440 14472
rect 11360 14312 11440 14408
rect 11360 14248 11368 14312
rect 11432 14248 11440 14312
rect 11360 14152 11440 14248
rect 11360 14088 11368 14152
rect 11432 14088 11440 14152
rect 11360 13992 11440 14088
rect 11360 13928 11368 13992
rect 11432 13928 11440 13992
rect 11360 13832 11440 13928
rect 11360 13768 11368 13832
rect 11432 13768 11440 13832
rect 11360 13672 11440 13768
rect 11360 13608 11368 13672
rect 11432 13608 11440 13672
rect 11360 13512 11440 13608
rect 11360 13448 11368 13512
rect 11432 13448 11440 13512
rect 11360 13352 11440 13448
rect 11360 13288 11368 13352
rect 11432 13288 11440 13352
rect 11360 13192 11440 13288
rect 11360 13128 11368 13192
rect 11432 13128 11440 13192
rect 11360 13032 11440 13128
rect 11360 12968 11368 13032
rect 11432 12968 11440 13032
rect 11360 12872 11440 12968
rect 11360 12808 11368 12872
rect 11432 12808 11440 12872
rect 11360 12712 11440 12808
rect 11360 12648 11368 12712
rect 11432 12648 11440 12712
rect 11360 12552 11440 12648
rect 11360 12488 11368 12552
rect 11432 12488 11440 12552
rect 11360 12392 11440 12488
rect 11360 12328 11368 12392
rect 11432 12328 11440 12392
rect 11360 12232 11440 12328
rect 11360 12168 11368 12232
rect 11432 12168 11440 12232
rect 11360 12072 11440 12168
rect 11360 12008 11368 12072
rect 11432 12008 11440 12072
rect 11360 11912 11440 12008
rect 11360 11848 11368 11912
rect 11432 11848 11440 11912
rect 11360 11752 11440 11848
rect 11360 11688 11368 11752
rect 11432 11688 11440 11752
rect 11360 11592 11440 11688
rect 11360 11528 11368 11592
rect 11432 11528 11440 11592
rect 11360 11432 11440 11528
rect 11360 11368 11368 11432
rect 11432 11368 11440 11432
rect 11360 11272 11440 11368
rect 11360 11208 11368 11272
rect 11432 11208 11440 11272
rect 11360 11112 11440 11208
rect 11360 11048 11368 11112
rect 11432 11048 11440 11112
rect 11360 10952 11440 11048
rect 11360 10888 11368 10952
rect 11432 10888 11440 10952
rect 11360 10792 11440 10888
rect 11360 10728 11368 10792
rect 11432 10728 11440 10792
rect 11360 10632 11440 10728
rect 11360 10568 11368 10632
rect 11432 10568 11440 10632
rect 11360 10472 11440 10568
rect 11360 10408 11368 10472
rect 11432 10408 11440 10472
rect 11360 10312 11440 10408
rect 11360 10248 11368 10312
rect 11432 10248 11440 10312
rect 11360 10152 11440 10248
rect 11360 10088 11368 10152
rect 11432 10088 11440 10152
rect 11360 9992 11440 10088
rect 11360 9928 11368 9992
rect 11432 9928 11440 9992
rect 11360 9832 11440 9928
rect 11360 9768 11368 9832
rect 11432 9768 11440 9832
rect 11360 9672 11440 9768
rect 11360 9608 11368 9672
rect 11432 9608 11440 9672
rect 11360 9512 11440 9608
rect 11360 9448 11368 9512
rect 11432 9448 11440 9512
rect 11360 9352 11440 9448
rect 11360 9288 11368 9352
rect 11432 9288 11440 9352
rect 11360 9192 11440 9288
rect 11360 9128 11368 9192
rect 11432 9128 11440 9192
rect 11360 9032 11440 9128
rect 11360 8968 11368 9032
rect 11432 8968 11440 9032
rect 11360 8872 11440 8968
rect 11360 8808 11368 8872
rect 11432 8808 11440 8872
rect 11360 8712 11440 8808
rect 11360 8648 11368 8712
rect 11432 8648 11440 8712
rect 11360 8552 11440 8648
rect 11360 8488 11368 8552
rect 11432 8488 11440 8552
rect 11360 8392 11440 8488
rect 11360 8328 11368 8392
rect 11432 8328 11440 8392
rect 11360 8232 11440 8328
rect 11360 8168 11368 8232
rect 11432 8168 11440 8232
rect 11360 8072 11440 8168
rect 11360 8008 11368 8072
rect 11432 8008 11440 8072
rect 11360 7912 11440 8008
rect 11360 7848 11368 7912
rect 11432 7848 11440 7912
rect 11360 7752 11440 7848
rect 11360 7688 11368 7752
rect 11432 7688 11440 7752
rect 11360 7592 11440 7688
rect 11360 7528 11368 7592
rect 11432 7528 11440 7592
rect 11360 7432 11440 7528
rect 11360 7368 11368 7432
rect 11432 7368 11440 7432
rect 11360 7272 11440 7368
rect 11360 7208 11368 7272
rect 11432 7208 11440 7272
rect 11360 7112 11440 7208
rect 11360 7048 11368 7112
rect 11432 7048 11440 7112
rect 11360 6952 11440 7048
rect 11360 6888 11368 6952
rect 11432 6888 11440 6952
rect 11360 6792 11440 6888
rect 11360 6728 11368 6792
rect 11432 6728 11440 6792
rect 11360 6632 11440 6728
rect 11360 6568 11368 6632
rect 11432 6568 11440 6632
rect 11360 6472 11440 6568
rect 11360 6408 11368 6472
rect 11432 6408 11440 6472
rect 11360 6312 11440 6408
rect 11360 6248 11368 6312
rect 11432 6248 11440 6312
rect 11360 6152 11440 6248
rect 11360 6088 11368 6152
rect 11432 6088 11440 6152
rect 11360 5992 11440 6088
rect 11360 5928 11368 5992
rect 11432 5928 11440 5992
rect 11360 5832 11440 5928
rect 11360 5768 11368 5832
rect 11432 5768 11440 5832
rect 11360 5672 11440 5768
rect 11360 5608 11368 5672
rect 11432 5608 11440 5672
rect 11360 5512 11440 5608
rect 11360 5448 11368 5512
rect 11432 5448 11440 5512
rect 11360 5352 11440 5448
rect 11360 5288 11368 5352
rect 11432 5288 11440 5352
rect 11360 5192 11440 5288
rect 11360 5128 11368 5192
rect 11432 5128 11440 5192
rect 11360 5032 11440 5128
rect 11360 4968 11368 5032
rect 11432 4968 11440 5032
rect 11360 4872 11440 4968
rect 11360 4808 11368 4872
rect 11432 4808 11440 4872
rect 11360 4712 11440 4808
rect 11360 4648 11368 4712
rect 11432 4648 11440 4712
rect 11360 4552 11440 4648
rect 11360 4488 11368 4552
rect 11432 4488 11440 4552
rect 11360 4392 11440 4488
rect 11360 4328 11368 4392
rect 11432 4328 11440 4392
rect 11360 4232 11440 4328
rect 11360 4168 11368 4232
rect 11432 4168 11440 4232
rect 11360 4072 11440 4168
rect 11360 4008 11368 4072
rect 11432 4008 11440 4072
rect 11360 3912 11440 4008
rect 11360 3848 11368 3912
rect 11432 3848 11440 3912
rect 11360 3752 11440 3848
rect 11360 3688 11368 3752
rect 11432 3688 11440 3752
rect 11360 3592 11440 3688
rect 11360 3528 11368 3592
rect 11432 3528 11440 3592
rect 11360 3432 11440 3528
rect 11360 3368 11368 3432
rect 11432 3368 11440 3432
rect 11360 3272 11440 3368
rect 11360 3208 11368 3272
rect 11432 3208 11440 3272
rect 11360 3112 11440 3208
rect 11360 3048 11368 3112
rect 11432 3048 11440 3112
rect 11360 2952 11440 3048
rect 11360 2888 11368 2952
rect 11432 2888 11440 2952
rect 11360 2792 11440 2888
rect 11360 2728 11368 2792
rect 11432 2728 11440 2792
rect 11360 2632 11440 2728
rect 11360 2568 11368 2632
rect 11432 2568 11440 2632
rect 11360 2472 11440 2568
rect 11360 2408 11368 2472
rect 11432 2408 11440 2472
rect 11360 2312 11440 2408
rect 11360 2248 11368 2312
rect 11432 2248 11440 2312
rect 11360 2152 11440 2248
rect 11360 2088 11368 2152
rect 11432 2088 11440 2152
rect 11360 1992 11440 2088
rect 11360 1928 11368 1992
rect 11432 1928 11440 1992
rect 11360 1832 11440 1928
rect 11360 1768 11368 1832
rect 11432 1768 11440 1832
rect 11360 1672 11440 1768
rect 11360 1608 11368 1672
rect 11432 1608 11440 1672
rect 11360 1512 11440 1608
rect 11360 1448 11368 1512
rect 11432 1448 11440 1512
rect 11360 1352 11440 1448
rect 11360 1288 11368 1352
rect 11432 1288 11440 1352
rect 11360 1192 11440 1288
rect 11360 1128 11368 1192
rect 11432 1128 11440 1192
rect 11360 1032 11440 1128
rect 11360 968 11368 1032
rect 11432 968 11440 1032
rect 11360 872 11440 968
rect 11360 808 11368 872
rect 11432 808 11440 872
rect 11360 712 11440 808
rect 11360 648 11368 712
rect 11432 648 11440 712
rect 11360 552 11440 648
rect 11360 488 11368 552
rect 11432 488 11440 552
rect 11360 392 11440 488
rect 11360 328 11368 392
rect 11432 328 11440 392
rect 11360 232 11440 328
rect 11360 168 11368 232
rect 11432 168 11440 232
rect 11360 72 11440 168
rect 11360 8 11368 72
rect 11432 8 11440 72
rect 11040 -1112 11048 -1048
rect 11112 -1112 11120 -1048
rect 11040 -1128 11120 -1112
rect 11040 -1192 11048 -1128
rect 11112 -1192 11120 -1128
rect 11040 -1208 11120 -1192
rect 11040 -1272 11048 -1208
rect 11112 -1272 11120 -1208
rect 11040 -1288 11120 -1272
rect 11040 -1352 11048 -1288
rect 11112 -1352 11120 -1288
rect 11040 -1368 11120 -1352
rect 11040 -1432 11048 -1368
rect 11112 -1432 11120 -1368
rect 11040 -1920 11120 -1432
rect 11360 -1048 11440 8
rect 11360 -1112 11368 -1048
rect 11432 -1112 11440 -1048
rect 11360 -1128 11440 -1112
rect 11360 -1192 11368 -1128
rect 11432 -1192 11440 -1128
rect 11360 -1208 11440 -1192
rect 11360 -1272 11368 -1208
rect 11432 -1272 11440 -1208
rect 11360 -1288 11440 -1272
rect 11360 -1352 11368 -1288
rect 11432 -1352 11440 -1288
rect 11360 -1368 11440 -1352
rect 11360 -1432 11368 -1368
rect 11432 -1432 11440 -1368
rect 11360 -1920 11440 -1432
rect 11520 31432 11600 31520
rect 11520 31368 11528 31432
rect 11592 31368 11600 31432
rect 11520 31272 11600 31368
rect 11520 31208 11528 31272
rect 11592 31208 11600 31272
rect 11520 31112 11600 31208
rect 11520 31048 11528 31112
rect 11592 31048 11600 31112
rect 11520 30952 11600 31048
rect 11520 30888 11528 30952
rect 11592 30888 11600 30952
rect 11520 30792 11600 30888
rect 11520 30728 11528 30792
rect 11592 30728 11600 30792
rect 11520 30632 11600 30728
rect 11520 30568 11528 30632
rect 11592 30568 11600 30632
rect 11520 30472 11600 30568
rect 11520 30408 11528 30472
rect 11592 30408 11600 30472
rect 11520 30312 11600 30408
rect 11520 30248 11528 30312
rect 11592 30248 11600 30312
rect 11520 30152 11600 30248
rect 11520 30088 11528 30152
rect 11592 30088 11600 30152
rect 11520 29992 11600 30088
rect 11520 29928 11528 29992
rect 11592 29928 11600 29992
rect 11520 29832 11600 29928
rect 11520 29768 11528 29832
rect 11592 29768 11600 29832
rect 11520 29672 11600 29768
rect 11520 29608 11528 29672
rect 11592 29608 11600 29672
rect 11520 29512 11600 29608
rect 11520 29448 11528 29512
rect 11592 29448 11600 29512
rect 11520 29352 11600 29448
rect 11520 29288 11528 29352
rect 11592 29288 11600 29352
rect 11520 29192 11600 29288
rect 11520 29128 11528 29192
rect 11592 29128 11600 29192
rect 11520 29032 11600 29128
rect 11520 28968 11528 29032
rect 11592 28968 11600 29032
rect 11520 28872 11600 28968
rect 11520 28808 11528 28872
rect 11592 28808 11600 28872
rect 11520 28712 11600 28808
rect 11520 28648 11528 28712
rect 11592 28648 11600 28712
rect 11520 28552 11600 28648
rect 11520 28488 11528 28552
rect 11592 28488 11600 28552
rect 11520 28392 11600 28488
rect 11520 28328 11528 28392
rect 11592 28328 11600 28392
rect 11520 28232 11600 28328
rect 11520 28168 11528 28232
rect 11592 28168 11600 28232
rect 11520 28072 11600 28168
rect 11520 28008 11528 28072
rect 11592 28008 11600 28072
rect 11520 27912 11600 28008
rect 11520 27848 11528 27912
rect 11592 27848 11600 27912
rect 11520 27752 11600 27848
rect 11520 27688 11528 27752
rect 11592 27688 11600 27752
rect 11520 27592 11600 27688
rect 11520 27528 11528 27592
rect 11592 27528 11600 27592
rect 11520 27432 11600 27528
rect 11520 27368 11528 27432
rect 11592 27368 11600 27432
rect 11520 27272 11600 27368
rect 11520 27208 11528 27272
rect 11592 27208 11600 27272
rect 11520 27112 11600 27208
rect 11520 27048 11528 27112
rect 11592 27048 11600 27112
rect 11520 26952 11600 27048
rect 11520 26888 11528 26952
rect 11592 26888 11600 26952
rect 11520 26792 11600 26888
rect 11520 26728 11528 26792
rect 11592 26728 11600 26792
rect 11520 26632 11600 26728
rect 11520 26568 11528 26632
rect 11592 26568 11600 26632
rect 11520 26472 11600 26568
rect 11520 26408 11528 26472
rect 11592 26408 11600 26472
rect 11520 26312 11600 26408
rect 11520 26248 11528 26312
rect 11592 26248 11600 26312
rect 11520 26152 11600 26248
rect 11520 26088 11528 26152
rect 11592 26088 11600 26152
rect 11520 25992 11600 26088
rect 11520 25928 11528 25992
rect 11592 25928 11600 25992
rect 11520 25832 11600 25928
rect 11520 25768 11528 25832
rect 11592 25768 11600 25832
rect 11520 25672 11600 25768
rect 11520 25608 11528 25672
rect 11592 25608 11600 25672
rect 11520 25512 11600 25608
rect 11520 25448 11528 25512
rect 11592 25448 11600 25512
rect 11520 25352 11600 25448
rect 11520 25288 11528 25352
rect 11592 25288 11600 25352
rect 11520 25192 11600 25288
rect 11520 25128 11528 25192
rect 11592 25128 11600 25192
rect 11520 25032 11600 25128
rect 11520 24968 11528 25032
rect 11592 24968 11600 25032
rect 11520 24872 11600 24968
rect 11520 24808 11528 24872
rect 11592 24808 11600 24872
rect 11520 24712 11600 24808
rect 11520 24648 11528 24712
rect 11592 24648 11600 24712
rect 11520 24552 11600 24648
rect 11520 24488 11528 24552
rect 11592 24488 11600 24552
rect 11520 24392 11600 24488
rect 11520 24328 11528 24392
rect 11592 24328 11600 24392
rect 11520 24232 11600 24328
rect 11520 24168 11528 24232
rect 11592 24168 11600 24232
rect 11520 24072 11600 24168
rect 11520 24008 11528 24072
rect 11592 24008 11600 24072
rect 11520 23912 11600 24008
rect 11520 23848 11528 23912
rect 11592 23848 11600 23912
rect 11520 23752 11600 23848
rect 11520 23688 11528 23752
rect 11592 23688 11600 23752
rect 11520 23592 11600 23688
rect 11520 23528 11528 23592
rect 11592 23528 11600 23592
rect 11520 23432 11600 23528
rect 11520 23368 11528 23432
rect 11592 23368 11600 23432
rect 11520 23272 11600 23368
rect 11520 23208 11528 23272
rect 11592 23208 11600 23272
rect 11520 23112 11600 23208
rect 11520 23048 11528 23112
rect 11592 23048 11600 23112
rect 11520 22952 11600 23048
rect 11520 22888 11528 22952
rect 11592 22888 11600 22952
rect 11520 22792 11600 22888
rect 11520 22728 11528 22792
rect 11592 22728 11600 22792
rect 11520 22632 11600 22728
rect 11520 22568 11528 22632
rect 11592 22568 11600 22632
rect 11520 22472 11600 22568
rect 11520 22408 11528 22472
rect 11592 22408 11600 22472
rect 11520 22312 11600 22408
rect 11520 22248 11528 22312
rect 11592 22248 11600 22312
rect 11520 22152 11600 22248
rect 11520 22088 11528 22152
rect 11592 22088 11600 22152
rect 11520 21992 11600 22088
rect 11520 21928 11528 21992
rect 11592 21928 11600 21992
rect 11520 21832 11600 21928
rect 11520 21768 11528 21832
rect 11592 21768 11600 21832
rect 11520 21672 11600 21768
rect 11520 21608 11528 21672
rect 11592 21608 11600 21672
rect 11520 21512 11600 21608
rect 11520 21448 11528 21512
rect 11592 21448 11600 21512
rect 11520 21352 11600 21448
rect 11520 21288 11528 21352
rect 11592 21288 11600 21352
rect 11520 21192 11600 21288
rect 11520 21128 11528 21192
rect 11592 21128 11600 21192
rect 11520 21032 11600 21128
rect 11520 20968 11528 21032
rect 11592 20968 11600 21032
rect 11520 20872 11600 20968
rect 11520 20808 11528 20872
rect 11592 20808 11600 20872
rect 11520 20712 11600 20808
rect 11520 20648 11528 20712
rect 11592 20648 11600 20712
rect 11520 20552 11600 20648
rect 11520 20488 11528 20552
rect 11592 20488 11600 20552
rect 11520 20392 11600 20488
rect 11520 20328 11528 20392
rect 11592 20328 11600 20392
rect 11520 20232 11600 20328
rect 11520 20168 11528 20232
rect 11592 20168 11600 20232
rect 11520 20072 11600 20168
rect 11520 20008 11528 20072
rect 11592 20008 11600 20072
rect 11520 19912 11600 20008
rect 11520 19848 11528 19912
rect 11592 19848 11600 19912
rect 11520 19752 11600 19848
rect 11520 19688 11528 19752
rect 11592 19688 11600 19752
rect 11520 19592 11600 19688
rect 11520 19528 11528 19592
rect 11592 19528 11600 19592
rect 11520 19432 11600 19528
rect 11520 19368 11528 19432
rect 11592 19368 11600 19432
rect 11520 19272 11600 19368
rect 11520 19208 11528 19272
rect 11592 19208 11600 19272
rect 11520 19112 11600 19208
rect 11520 19048 11528 19112
rect 11592 19048 11600 19112
rect 11520 18952 11600 19048
rect 11520 18888 11528 18952
rect 11592 18888 11600 18952
rect 11520 18792 11600 18888
rect 11520 18728 11528 18792
rect 11592 18728 11600 18792
rect 11520 18632 11600 18728
rect 11520 18568 11528 18632
rect 11592 18568 11600 18632
rect 11520 18472 11600 18568
rect 11520 18408 11528 18472
rect 11592 18408 11600 18472
rect 11520 18312 11600 18408
rect 11520 18248 11528 18312
rect 11592 18248 11600 18312
rect 11520 18152 11600 18248
rect 11520 18088 11528 18152
rect 11592 18088 11600 18152
rect 11520 17992 11600 18088
rect 11520 17928 11528 17992
rect 11592 17928 11600 17992
rect 11520 17832 11600 17928
rect 11520 17768 11528 17832
rect 11592 17768 11600 17832
rect 11520 17672 11600 17768
rect 11520 17608 11528 17672
rect 11592 17608 11600 17672
rect 11520 17512 11600 17608
rect 11520 17448 11528 17512
rect 11592 17448 11600 17512
rect 11520 17352 11600 17448
rect 11520 17288 11528 17352
rect 11592 17288 11600 17352
rect 11520 17192 11600 17288
rect 11520 17128 11528 17192
rect 11592 17128 11600 17192
rect 11520 17032 11600 17128
rect 11520 16968 11528 17032
rect 11592 16968 11600 17032
rect 11520 16872 11600 16968
rect 11520 16808 11528 16872
rect 11592 16808 11600 16872
rect 11520 16712 11600 16808
rect 11520 16648 11528 16712
rect 11592 16648 11600 16712
rect 11520 16552 11600 16648
rect 11520 16488 11528 16552
rect 11592 16488 11600 16552
rect 11520 16392 11600 16488
rect 11520 16328 11528 16392
rect 11592 16328 11600 16392
rect 11520 16232 11600 16328
rect 11520 16168 11528 16232
rect 11592 16168 11600 16232
rect 11520 16072 11600 16168
rect 11520 16008 11528 16072
rect 11592 16008 11600 16072
rect 11520 15912 11600 16008
rect 11520 15848 11528 15912
rect 11592 15848 11600 15912
rect 11520 15752 11600 15848
rect 11520 15688 11528 15752
rect 11592 15688 11600 15752
rect 11520 15592 11600 15688
rect 11520 15528 11528 15592
rect 11592 15528 11600 15592
rect 11520 15432 11600 15528
rect 11520 15368 11528 15432
rect 11592 15368 11600 15432
rect 11520 15272 11600 15368
rect 11520 15208 11528 15272
rect 11592 15208 11600 15272
rect 11520 15112 11600 15208
rect 11520 15048 11528 15112
rect 11592 15048 11600 15112
rect 11520 14952 11600 15048
rect 11520 14888 11528 14952
rect 11592 14888 11600 14952
rect 11520 14792 11600 14888
rect 11520 14728 11528 14792
rect 11592 14728 11600 14792
rect 11520 14632 11600 14728
rect 11520 14568 11528 14632
rect 11592 14568 11600 14632
rect 11520 14472 11600 14568
rect 11520 14408 11528 14472
rect 11592 14408 11600 14472
rect 11520 14312 11600 14408
rect 11520 14248 11528 14312
rect 11592 14248 11600 14312
rect 11520 14152 11600 14248
rect 11520 14088 11528 14152
rect 11592 14088 11600 14152
rect 11520 13992 11600 14088
rect 11520 13928 11528 13992
rect 11592 13928 11600 13992
rect 11520 13832 11600 13928
rect 11520 13768 11528 13832
rect 11592 13768 11600 13832
rect 11520 13672 11600 13768
rect 11520 13608 11528 13672
rect 11592 13608 11600 13672
rect 11520 13512 11600 13608
rect 11520 13448 11528 13512
rect 11592 13448 11600 13512
rect 11520 13352 11600 13448
rect 11520 13288 11528 13352
rect 11592 13288 11600 13352
rect 11520 13192 11600 13288
rect 11520 13128 11528 13192
rect 11592 13128 11600 13192
rect 11520 13032 11600 13128
rect 11520 12968 11528 13032
rect 11592 12968 11600 13032
rect 11520 12872 11600 12968
rect 11520 12808 11528 12872
rect 11592 12808 11600 12872
rect 11520 12712 11600 12808
rect 11520 12648 11528 12712
rect 11592 12648 11600 12712
rect 11520 12552 11600 12648
rect 11520 12488 11528 12552
rect 11592 12488 11600 12552
rect 11520 12392 11600 12488
rect 11520 12328 11528 12392
rect 11592 12328 11600 12392
rect 11520 12232 11600 12328
rect 11520 12168 11528 12232
rect 11592 12168 11600 12232
rect 11520 12072 11600 12168
rect 11520 12008 11528 12072
rect 11592 12008 11600 12072
rect 11520 11912 11600 12008
rect 11520 11848 11528 11912
rect 11592 11848 11600 11912
rect 11520 11752 11600 11848
rect 11520 11688 11528 11752
rect 11592 11688 11600 11752
rect 11520 11592 11600 11688
rect 11520 11528 11528 11592
rect 11592 11528 11600 11592
rect 11520 11432 11600 11528
rect 11520 11368 11528 11432
rect 11592 11368 11600 11432
rect 11520 11272 11600 11368
rect 11520 11208 11528 11272
rect 11592 11208 11600 11272
rect 11520 11112 11600 11208
rect 11520 11048 11528 11112
rect 11592 11048 11600 11112
rect 11520 10952 11600 11048
rect 11520 10888 11528 10952
rect 11592 10888 11600 10952
rect 11520 10792 11600 10888
rect 11520 10728 11528 10792
rect 11592 10728 11600 10792
rect 11520 10632 11600 10728
rect 11520 10568 11528 10632
rect 11592 10568 11600 10632
rect 11520 10472 11600 10568
rect 11520 10408 11528 10472
rect 11592 10408 11600 10472
rect 11520 10312 11600 10408
rect 11520 10248 11528 10312
rect 11592 10248 11600 10312
rect 11520 10152 11600 10248
rect 11520 10088 11528 10152
rect 11592 10088 11600 10152
rect 11520 9992 11600 10088
rect 11520 9928 11528 9992
rect 11592 9928 11600 9992
rect 11520 9832 11600 9928
rect 11520 9768 11528 9832
rect 11592 9768 11600 9832
rect 11520 9672 11600 9768
rect 11520 9608 11528 9672
rect 11592 9608 11600 9672
rect 11520 9512 11600 9608
rect 11520 9448 11528 9512
rect 11592 9448 11600 9512
rect 11520 9352 11600 9448
rect 11520 9288 11528 9352
rect 11592 9288 11600 9352
rect 11520 9192 11600 9288
rect 11520 9128 11528 9192
rect 11592 9128 11600 9192
rect 11520 9032 11600 9128
rect 11520 8968 11528 9032
rect 11592 8968 11600 9032
rect 11520 8872 11600 8968
rect 11520 8808 11528 8872
rect 11592 8808 11600 8872
rect 11520 8712 11600 8808
rect 11520 8648 11528 8712
rect 11592 8648 11600 8712
rect 11520 8552 11600 8648
rect 11520 8488 11528 8552
rect 11592 8488 11600 8552
rect 11520 8392 11600 8488
rect 11520 8328 11528 8392
rect 11592 8328 11600 8392
rect 11520 8232 11600 8328
rect 11520 8168 11528 8232
rect 11592 8168 11600 8232
rect 11520 8072 11600 8168
rect 11520 8008 11528 8072
rect 11592 8008 11600 8072
rect 11520 7912 11600 8008
rect 11520 7848 11528 7912
rect 11592 7848 11600 7912
rect 11520 7752 11600 7848
rect 11520 7688 11528 7752
rect 11592 7688 11600 7752
rect 11520 7592 11600 7688
rect 11520 7528 11528 7592
rect 11592 7528 11600 7592
rect 11520 7432 11600 7528
rect 11520 7368 11528 7432
rect 11592 7368 11600 7432
rect 11520 7272 11600 7368
rect 11520 7208 11528 7272
rect 11592 7208 11600 7272
rect 11520 7112 11600 7208
rect 11520 7048 11528 7112
rect 11592 7048 11600 7112
rect 11520 6952 11600 7048
rect 11520 6888 11528 6952
rect 11592 6888 11600 6952
rect 11520 6792 11600 6888
rect 11520 6728 11528 6792
rect 11592 6728 11600 6792
rect 11520 6632 11600 6728
rect 11520 6568 11528 6632
rect 11592 6568 11600 6632
rect 11520 6472 11600 6568
rect 11520 6408 11528 6472
rect 11592 6408 11600 6472
rect 11520 6312 11600 6408
rect 11520 6248 11528 6312
rect 11592 6248 11600 6312
rect 11520 6152 11600 6248
rect 11520 6088 11528 6152
rect 11592 6088 11600 6152
rect 11520 5992 11600 6088
rect 11520 5928 11528 5992
rect 11592 5928 11600 5992
rect 11520 5832 11600 5928
rect 11520 5768 11528 5832
rect 11592 5768 11600 5832
rect 11520 5672 11600 5768
rect 11520 5608 11528 5672
rect 11592 5608 11600 5672
rect 11520 5512 11600 5608
rect 11520 5448 11528 5512
rect 11592 5448 11600 5512
rect 11520 5352 11600 5448
rect 11520 5288 11528 5352
rect 11592 5288 11600 5352
rect 11520 5192 11600 5288
rect 11520 5128 11528 5192
rect 11592 5128 11600 5192
rect 11520 5032 11600 5128
rect 11520 4968 11528 5032
rect 11592 4968 11600 5032
rect 11520 4872 11600 4968
rect 11520 4808 11528 4872
rect 11592 4808 11600 4872
rect 11520 4712 11600 4808
rect 11520 4648 11528 4712
rect 11592 4648 11600 4712
rect 11520 4552 11600 4648
rect 11520 4488 11528 4552
rect 11592 4488 11600 4552
rect 11520 4392 11600 4488
rect 11520 4328 11528 4392
rect 11592 4328 11600 4392
rect 11520 4232 11600 4328
rect 11520 4168 11528 4232
rect 11592 4168 11600 4232
rect 11520 4072 11600 4168
rect 11520 4008 11528 4072
rect 11592 4008 11600 4072
rect 11520 3912 11600 4008
rect 11520 3848 11528 3912
rect 11592 3848 11600 3912
rect 11520 3752 11600 3848
rect 11520 3688 11528 3752
rect 11592 3688 11600 3752
rect 11520 3592 11600 3688
rect 11520 3528 11528 3592
rect 11592 3528 11600 3592
rect 11520 3432 11600 3528
rect 11520 3368 11528 3432
rect 11592 3368 11600 3432
rect 11520 3272 11600 3368
rect 11520 3208 11528 3272
rect 11592 3208 11600 3272
rect 11520 3112 11600 3208
rect 11520 3048 11528 3112
rect 11592 3048 11600 3112
rect 11520 2952 11600 3048
rect 11520 2888 11528 2952
rect 11592 2888 11600 2952
rect 11520 2792 11600 2888
rect 11520 2728 11528 2792
rect 11592 2728 11600 2792
rect 11520 2632 11600 2728
rect 11520 2568 11528 2632
rect 11592 2568 11600 2632
rect 11520 2472 11600 2568
rect 11520 2408 11528 2472
rect 11592 2408 11600 2472
rect 11520 2312 11600 2408
rect 11520 2248 11528 2312
rect 11592 2248 11600 2312
rect 11520 2152 11600 2248
rect 11520 2088 11528 2152
rect 11592 2088 11600 2152
rect 11520 1992 11600 2088
rect 11520 1928 11528 1992
rect 11592 1928 11600 1992
rect 11520 1832 11600 1928
rect 11520 1768 11528 1832
rect 11592 1768 11600 1832
rect 11520 1672 11600 1768
rect 11520 1608 11528 1672
rect 11592 1608 11600 1672
rect 11520 1512 11600 1608
rect 11520 1448 11528 1512
rect 11592 1448 11600 1512
rect 11520 1352 11600 1448
rect 11520 1288 11528 1352
rect 11592 1288 11600 1352
rect 11520 1192 11600 1288
rect 11520 1128 11528 1192
rect 11592 1128 11600 1192
rect 11520 1032 11600 1128
rect 11520 968 11528 1032
rect 11592 968 11600 1032
rect 11520 872 11600 968
rect 11520 808 11528 872
rect 11592 808 11600 872
rect 11520 712 11600 808
rect 11520 648 11528 712
rect 11592 648 11600 712
rect 11520 552 11600 648
rect 11520 488 11528 552
rect 11592 488 11600 552
rect 11520 392 11600 488
rect 11520 328 11528 392
rect 11592 328 11600 392
rect 11520 232 11600 328
rect 11520 168 11528 232
rect 11592 168 11600 232
rect 11520 72 11600 168
rect 11520 8 11528 72
rect 11592 8 11600 72
rect 11520 -88 11600 8
rect 11680 9668 11760 31520
rect 11680 9612 11692 9668
rect 11748 9612 11760 9668
rect 11680 6628 11760 9612
rect 11680 6572 11692 6628
rect 11748 6572 11760 6628
rect 11680 0 11760 6572
rect 11840 31432 11920 31520
rect 11840 31368 11848 31432
rect 11912 31368 11920 31432
rect 11840 31272 11920 31368
rect 11840 31208 11848 31272
rect 11912 31208 11920 31272
rect 11840 31112 11920 31208
rect 11840 31048 11848 31112
rect 11912 31048 11920 31112
rect 11840 30952 11920 31048
rect 11840 30888 11848 30952
rect 11912 30888 11920 30952
rect 11840 30792 11920 30888
rect 11840 30728 11848 30792
rect 11912 30728 11920 30792
rect 11840 30632 11920 30728
rect 11840 30568 11848 30632
rect 11912 30568 11920 30632
rect 11840 30472 11920 30568
rect 11840 30408 11848 30472
rect 11912 30408 11920 30472
rect 11840 30312 11920 30408
rect 11840 30248 11848 30312
rect 11912 30248 11920 30312
rect 11840 30152 11920 30248
rect 11840 30088 11848 30152
rect 11912 30088 11920 30152
rect 11840 29992 11920 30088
rect 11840 29928 11848 29992
rect 11912 29928 11920 29992
rect 11840 29832 11920 29928
rect 11840 29768 11848 29832
rect 11912 29768 11920 29832
rect 11840 29672 11920 29768
rect 11840 29608 11848 29672
rect 11912 29608 11920 29672
rect 11840 29512 11920 29608
rect 11840 29448 11848 29512
rect 11912 29448 11920 29512
rect 11840 29352 11920 29448
rect 11840 29288 11848 29352
rect 11912 29288 11920 29352
rect 11840 29192 11920 29288
rect 11840 29128 11848 29192
rect 11912 29128 11920 29192
rect 11840 29032 11920 29128
rect 11840 28968 11848 29032
rect 11912 28968 11920 29032
rect 11840 28872 11920 28968
rect 11840 28808 11848 28872
rect 11912 28808 11920 28872
rect 11840 28712 11920 28808
rect 11840 28648 11848 28712
rect 11912 28648 11920 28712
rect 11840 28552 11920 28648
rect 11840 28488 11848 28552
rect 11912 28488 11920 28552
rect 11840 28392 11920 28488
rect 11840 28328 11848 28392
rect 11912 28328 11920 28392
rect 11840 28232 11920 28328
rect 11840 28168 11848 28232
rect 11912 28168 11920 28232
rect 11840 28072 11920 28168
rect 11840 28008 11848 28072
rect 11912 28008 11920 28072
rect 11840 27912 11920 28008
rect 11840 27848 11848 27912
rect 11912 27848 11920 27912
rect 11840 27752 11920 27848
rect 11840 27688 11848 27752
rect 11912 27688 11920 27752
rect 11840 27592 11920 27688
rect 11840 27528 11848 27592
rect 11912 27528 11920 27592
rect 11840 27432 11920 27528
rect 11840 27368 11848 27432
rect 11912 27368 11920 27432
rect 11840 27272 11920 27368
rect 11840 27208 11848 27272
rect 11912 27208 11920 27272
rect 11840 27112 11920 27208
rect 11840 27048 11848 27112
rect 11912 27048 11920 27112
rect 11840 26952 11920 27048
rect 11840 26888 11848 26952
rect 11912 26888 11920 26952
rect 11840 26792 11920 26888
rect 11840 26728 11848 26792
rect 11912 26728 11920 26792
rect 11840 26632 11920 26728
rect 11840 26568 11848 26632
rect 11912 26568 11920 26632
rect 11840 26472 11920 26568
rect 11840 26408 11848 26472
rect 11912 26408 11920 26472
rect 11840 26312 11920 26408
rect 11840 26248 11848 26312
rect 11912 26248 11920 26312
rect 11840 26152 11920 26248
rect 11840 26088 11848 26152
rect 11912 26088 11920 26152
rect 11840 25992 11920 26088
rect 11840 25928 11848 25992
rect 11912 25928 11920 25992
rect 11840 25832 11920 25928
rect 11840 25768 11848 25832
rect 11912 25768 11920 25832
rect 11840 25672 11920 25768
rect 11840 25608 11848 25672
rect 11912 25608 11920 25672
rect 11840 25512 11920 25608
rect 11840 25448 11848 25512
rect 11912 25448 11920 25512
rect 11840 25352 11920 25448
rect 11840 25288 11848 25352
rect 11912 25288 11920 25352
rect 11840 25192 11920 25288
rect 11840 25128 11848 25192
rect 11912 25128 11920 25192
rect 11840 25032 11920 25128
rect 11840 24968 11848 25032
rect 11912 24968 11920 25032
rect 11840 24872 11920 24968
rect 11840 24808 11848 24872
rect 11912 24808 11920 24872
rect 11840 24712 11920 24808
rect 11840 24648 11848 24712
rect 11912 24648 11920 24712
rect 11840 24552 11920 24648
rect 11840 24488 11848 24552
rect 11912 24488 11920 24552
rect 11840 24392 11920 24488
rect 11840 24328 11848 24392
rect 11912 24328 11920 24392
rect 11840 24232 11920 24328
rect 11840 24168 11848 24232
rect 11912 24168 11920 24232
rect 11840 24072 11920 24168
rect 11840 24008 11848 24072
rect 11912 24008 11920 24072
rect 11840 23912 11920 24008
rect 11840 23848 11848 23912
rect 11912 23848 11920 23912
rect 11840 23752 11920 23848
rect 11840 23688 11848 23752
rect 11912 23688 11920 23752
rect 11840 23592 11920 23688
rect 11840 23528 11848 23592
rect 11912 23528 11920 23592
rect 11840 23432 11920 23528
rect 11840 23368 11848 23432
rect 11912 23368 11920 23432
rect 11840 23272 11920 23368
rect 11840 23208 11848 23272
rect 11912 23208 11920 23272
rect 11840 23112 11920 23208
rect 11840 23048 11848 23112
rect 11912 23048 11920 23112
rect 11840 22952 11920 23048
rect 11840 22888 11848 22952
rect 11912 22888 11920 22952
rect 11840 22792 11920 22888
rect 11840 22728 11848 22792
rect 11912 22728 11920 22792
rect 11840 22632 11920 22728
rect 11840 22568 11848 22632
rect 11912 22568 11920 22632
rect 11840 22472 11920 22568
rect 11840 22408 11848 22472
rect 11912 22408 11920 22472
rect 11840 22312 11920 22408
rect 11840 22248 11848 22312
rect 11912 22248 11920 22312
rect 11840 22152 11920 22248
rect 11840 22088 11848 22152
rect 11912 22088 11920 22152
rect 11840 21992 11920 22088
rect 11840 21928 11848 21992
rect 11912 21928 11920 21992
rect 11840 21832 11920 21928
rect 11840 21768 11848 21832
rect 11912 21768 11920 21832
rect 11840 21672 11920 21768
rect 11840 21608 11848 21672
rect 11912 21608 11920 21672
rect 11840 21512 11920 21608
rect 11840 21448 11848 21512
rect 11912 21448 11920 21512
rect 11840 21352 11920 21448
rect 11840 21288 11848 21352
rect 11912 21288 11920 21352
rect 11840 21192 11920 21288
rect 11840 21128 11848 21192
rect 11912 21128 11920 21192
rect 11840 21032 11920 21128
rect 11840 20968 11848 21032
rect 11912 20968 11920 21032
rect 11840 20872 11920 20968
rect 11840 20808 11848 20872
rect 11912 20808 11920 20872
rect 11840 20712 11920 20808
rect 11840 20648 11848 20712
rect 11912 20648 11920 20712
rect 11840 20552 11920 20648
rect 11840 20488 11848 20552
rect 11912 20488 11920 20552
rect 11840 20392 11920 20488
rect 11840 20328 11848 20392
rect 11912 20328 11920 20392
rect 11840 20232 11920 20328
rect 11840 20168 11848 20232
rect 11912 20168 11920 20232
rect 11840 20072 11920 20168
rect 11840 20008 11848 20072
rect 11912 20008 11920 20072
rect 11840 19912 11920 20008
rect 11840 19848 11848 19912
rect 11912 19848 11920 19912
rect 11840 19752 11920 19848
rect 11840 19688 11848 19752
rect 11912 19688 11920 19752
rect 11840 19592 11920 19688
rect 11840 19528 11848 19592
rect 11912 19528 11920 19592
rect 11840 19432 11920 19528
rect 11840 19368 11848 19432
rect 11912 19368 11920 19432
rect 11840 19272 11920 19368
rect 11840 19208 11848 19272
rect 11912 19208 11920 19272
rect 11840 19112 11920 19208
rect 11840 19048 11848 19112
rect 11912 19048 11920 19112
rect 11840 18952 11920 19048
rect 11840 18888 11848 18952
rect 11912 18888 11920 18952
rect 11840 18792 11920 18888
rect 11840 18728 11848 18792
rect 11912 18728 11920 18792
rect 11840 18632 11920 18728
rect 11840 18568 11848 18632
rect 11912 18568 11920 18632
rect 11840 18472 11920 18568
rect 11840 18408 11848 18472
rect 11912 18408 11920 18472
rect 11840 18312 11920 18408
rect 11840 18248 11848 18312
rect 11912 18248 11920 18312
rect 11840 18152 11920 18248
rect 11840 18088 11848 18152
rect 11912 18088 11920 18152
rect 11840 17992 11920 18088
rect 11840 17928 11848 17992
rect 11912 17928 11920 17992
rect 11840 17832 11920 17928
rect 11840 17768 11848 17832
rect 11912 17768 11920 17832
rect 11840 17672 11920 17768
rect 11840 17608 11848 17672
rect 11912 17608 11920 17672
rect 11840 17512 11920 17608
rect 11840 17448 11848 17512
rect 11912 17448 11920 17512
rect 11840 17352 11920 17448
rect 11840 17288 11848 17352
rect 11912 17288 11920 17352
rect 11840 17192 11920 17288
rect 11840 17128 11848 17192
rect 11912 17128 11920 17192
rect 11840 17032 11920 17128
rect 11840 16968 11848 17032
rect 11912 16968 11920 17032
rect 11840 16872 11920 16968
rect 11840 16808 11848 16872
rect 11912 16808 11920 16872
rect 11840 16712 11920 16808
rect 11840 16648 11848 16712
rect 11912 16648 11920 16712
rect 11840 16552 11920 16648
rect 11840 16488 11848 16552
rect 11912 16488 11920 16552
rect 11840 16392 11920 16488
rect 11840 16328 11848 16392
rect 11912 16328 11920 16392
rect 11840 16232 11920 16328
rect 11840 16168 11848 16232
rect 11912 16168 11920 16232
rect 11840 16072 11920 16168
rect 11840 16008 11848 16072
rect 11912 16008 11920 16072
rect 11840 15912 11920 16008
rect 11840 15848 11848 15912
rect 11912 15848 11920 15912
rect 11840 15752 11920 15848
rect 11840 15688 11848 15752
rect 11912 15688 11920 15752
rect 11840 15592 11920 15688
rect 11840 15528 11848 15592
rect 11912 15528 11920 15592
rect 11840 15432 11920 15528
rect 11840 15368 11848 15432
rect 11912 15368 11920 15432
rect 11840 15272 11920 15368
rect 11840 15208 11848 15272
rect 11912 15208 11920 15272
rect 11840 15112 11920 15208
rect 11840 15048 11848 15112
rect 11912 15048 11920 15112
rect 11840 14952 11920 15048
rect 11840 14888 11848 14952
rect 11912 14888 11920 14952
rect 11840 14792 11920 14888
rect 11840 14728 11848 14792
rect 11912 14728 11920 14792
rect 11840 14632 11920 14728
rect 11840 14568 11848 14632
rect 11912 14568 11920 14632
rect 11840 14472 11920 14568
rect 11840 14408 11848 14472
rect 11912 14408 11920 14472
rect 11840 14312 11920 14408
rect 11840 14248 11848 14312
rect 11912 14248 11920 14312
rect 11840 14152 11920 14248
rect 11840 14088 11848 14152
rect 11912 14088 11920 14152
rect 11840 13992 11920 14088
rect 11840 13928 11848 13992
rect 11912 13928 11920 13992
rect 11840 13832 11920 13928
rect 11840 13768 11848 13832
rect 11912 13768 11920 13832
rect 11840 13672 11920 13768
rect 11840 13608 11848 13672
rect 11912 13608 11920 13672
rect 11840 13512 11920 13608
rect 11840 13448 11848 13512
rect 11912 13448 11920 13512
rect 11840 13352 11920 13448
rect 11840 13288 11848 13352
rect 11912 13288 11920 13352
rect 11840 13192 11920 13288
rect 11840 13128 11848 13192
rect 11912 13128 11920 13192
rect 11840 13032 11920 13128
rect 11840 12968 11848 13032
rect 11912 12968 11920 13032
rect 11840 12872 11920 12968
rect 11840 12808 11848 12872
rect 11912 12808 11920 12872
rect 11840 12712 11920 12808
rect 11840 12648 11848 12712
rect 11912 12648 11920 12712
rect 11840 12552 11920 12648
rect 11840 12488 11848 12552
rect 11912 12488 11920 12552
rect 11840 12392 11920 12488
rect 11840 12328 11848 12392
rect 11912 12328 11920 12392
rect 11840 12232 11920 12328
rect 11840 12168 11848 12232
rect 11912 12168 11920 12232
rect 11840 12072 11920 12168
rect 11840 12008 11848 12072
rect 11912 12008 11920 12072
rect 11840 11912 11920 12008
rect 11840 11848 11848 11912
rect 11912 11848 11920 11912
rect 11840 11752 11920 11848
rect 11840 11688 11848 11752
rect 11912 11688 11920 11752
rect 11840 11592 11920 11688
rect 11840 11528 11848 11592
rect 11912 11528 11920 11592
rect 11840 11432 11920 11528
rect 11840 11368 11848 11432
rect 11912 11368 11920 11432
rect 11840 11272 11920 11368
rect 11840 11208 11848 11272
rect 11912 11208 11920 11272
rect 11840 11112 11920 11208
rect 11840 11048 11848 11112
rect 11912 11048 11920 11112
rect 11840 10952 11920 11048
rect 11840 10888 11848 10952
rect 11912 10888 11920 10952
rect 11840 10792 11920 10888
rect 11840 10728 11848 10792
rect 11912 10728 11920 10792
rect 11840 10632 11920 10728
rect 11840 10568 11848 10632
rect 11912 10568 11920 10632
rect 11840 10472 11920 10568
rect 11840 10408 11848 10472
rect 11912 10408 11920 10472
rect 11840 10312 11920 10408
rect 11840 10248 11848 10312
rect 11912 10248 11920 10312
rect 11840 10152 11920 10248
rect 11840 10088 11848 10152
rect 11912 10088 11920 10152
rect 11840 9992 11920 10088
rect 11840 9928 11848 9992
rect 11912 9928 11920 9992
rect 11840 9832 11920 9928
rect 11840 9768 11848 9832
rect 11912 9768 11920 9832
rect 11840 9672 11920 9768
rect 11840 9608 11848 9672
rect 11912 9608 11920 9672
rect 11840 9512 11920 9608
rect 11840 9448 11848 9512
rect 11912 9448 11920 9512
rect 11840 9352 11920 9448
rect 11840 9288 11848 9352
rect 11912 9288 11920 9352
rect 11840 9192 11920 9288
rect 11840 9128 11848 9192
rect 11912 9128 11920 9192
rect 11840 9032 11920 9128
rect 11840 8968 11848 9032
rect 11912 8968 11920 9032
rect 11840 8872 11920 8968
rect 11840 8808 11848 8872
rect 11912 8808 11920 8872
rect 11840 8712 11920 8808
rect 11840 8648 11848 8712
rect 11912 8648 11920 8712
rect 11840 8552 11920 8648
rect 11840 8488 11848 8552
rect 11912 8488 11920 8552
rect 11840 8392 11920 8488
rect 11840 8328 11848 8392
rect 11912 8328 11920 8392
rect 11840 8232 11920 8328
rect 11840 8168 11848 8232
rect 11912 8168 11920 8232
rect 11840 8072 11920 8168
rect 11840 8008 11848 8072
rect 11912 8008 11920 8072
rect 11840 7912 11920 8008
rect 11840 7848 11848 7912
rect 11912 7848 11920 7912
rect 11840 7752 11920 7848
rect 11840 7688 11848 7752
rect 11912 7688 11920 7752
rect 11840 7592 11920 7688
rect 11840 7528 11848 7592
rect 11912 7528 11920 7592
rect 11840 7432 11920 7528
rect 11840 7368 11848 7432
rect 11912 7368 11920 7432
rect 11840 7272 11920 7368
rect 11840 7208 11848 7272
rect 11912 7208 11920 7272
rect 11840 7112 11920 7208
rect 11840 7048 11848 7112
rect 11912 7048 11920 7112
rect 11840 6952 11920 7048
rect 11840 6888 11848 6952
rect 11912 6888 11920 6952
rect 11840 6792 11920 6888
rect 11840 6728 11848 6792
rect 11912 6728 11920 6792
rect 11840 6632 11920 6728
rect 11840 6568 11848 6632
rect 11912 6568 11920 6632
rect 11840 6472 11920 6568
rect 11840 6408 11848 6472
rect 11912 6408 11920 6472
rect 11840 6312 11920 6408
rect 11840 6248 11848 6312
rect 11912 6248 11920 6312
rect 11840 6152 11920 6248
rect 11840 6088 11848 6152
rect 11912 6088 11920 6152
rect 11840 5992 11920 6088
rect 11840 5928 11848 5992
rect 11912 5928 11920 5992
rect 11840 5832 11920 5928
rect 11840 5768 11848 5832
rect 11912 5768 11920 5832
rect 11840 5672 11920 5768
rect 11840 5608 11848 5672
rect 11912 5608 11920 5672
rect 11840 5512 11920 5608
rect 11840 5448 11848 5512
rect 11912 5448 11920 5512
rect 11840 5352 11920 5448
rect 11840 5288 11848 5352
rect 11912 5288 11920 5352
rect 11840 5192 11920 5288
rect 11840 5128 11848 5192
rect 11912 5128 11920 5192
rect 11840 5032 11920 5128
rect 11840 4968 11848 5032
rect 11912 4968 11920 5032
rect 11840 4872 11920 4968
rect 11840 4808 11848 4872
rect 11912 4808 11920 4872
rect 11840 4712 11920 4808
rect 11840 4648 11848 4712
rect 11912 4648 11920 4712
rect 11840 4552 11920 4648
rect 11840 4488 11848 4552
rect 11912 4488 11920 4552
rect 11840 4392 11920 4488
rect 11840 4328 11848 4392
rect 11912 4328 11920 4392
rect 11840 4232 11920 4328
rect 11840 4168 11848 4232
rect 11912 4168 11920 4232
rect 11840 4072 11920 4168
rect 11840 4008 11848 4072
rect 11912 4008 11920 4072
rect 11840 3912 11920 4008
rect 11840 3848 11848 3912
rect 11912 3848 11920 3912
rect 11840 3752 11920 3848
rect 11840 3688 11848 3752
rect 11912 3688 11920 3752
rect 11840 3592 11920 3688
rect 11840 3528 11848 3592
rect 11912 3528 11920 3592
rect 11840 3432 11920 3528
rect 11840 3368 11848 3432
rect 11912 3368 11920 3432
rect 11840 3272 11920 3368
rect 11840 3208 11848 3272
rect 11912 3208 11920 3272
rect 11840 3112 11920 3208
rect 11840 3048 11848 3112
rect 11912 3048 11920 3112
rect 11840 2952 11920 3048
rect 11840 2888 11848 2952
rect 11912 2888 11920 2952
rect 11840 2792 11920 2888
rect 11840 2728 11848 2792
rect 11912 2728 11920 2792
rect 11840 2632 11920 2728
rect 11840 2568 11848 2632
rect 11912 2568 11920 2632
rect 11840 2472 11920 2568
rect 11840 2408 11848 2472
rect 11912 2408 11920 2472
rect 11840 2312 11920 2408
rect 11840 2248 11848 2312
rect 11912 2248 11920 2312
rect 11840 2152 11920 2248
rect 11840 2088 11848 2152
rect 11912 2088 11920 2152
rect 11840 1992 11920 2088
rect 11840 1928 11848 1992
rect 11912 1928 11920 1992
rect 11840 1832 11920 1928
rect 11840 1768 11848 1832
rect 11912 1768 11920 1832
rect 11840 1672 11920 1768
rect 11840 1608 11848 1672
rect 11912 1608 11920 1672
rect 11840 1512 11920 1608
rect 11840 1448 11848 1512
rect 11912 1448 11920 1512
rect 11840 1352 11920 1448
rect 11840 1288 11848 1352
rect 11912 1288 11920 1352
rect 11840 1192 11920 1288
rect 11840 1128 11848 1192
rect 11912 1128 11920 1192
rect 11840 1032 11920 1128
rect 11840 968 11848 1032
rect 11912 968 11920 1032
rect 11840 872 11920 968
rect 11840 808 11848 872
rect 11912 808 11920 872
rect 11840 712 11920 808
rect 11840 648 11848 712
rect 11912 648 11920 712
rect 11840 552 11920 648
rect 11840 488 11848 552
rect 11912 488 11920 552
rect 11840 392 11920 488
rect 11840 328 11848 392
rect 11912 328 11920 392
rect 11840 232 11920 328
rect 11840 168 11848 232
rect 11912 168 11920 232
rect 11840 72 11920 168
rect 11840 8 11848 72
rect 11912 8 11920 72
rect 11520 -152 11528 -88
rect 11592 -152 11600 -88
rect 11520 -168 11600 -152
rect 11520 -232 11528 -168
rect 11592 -232 11600 -168
rect 11520 -248 11600 -232
rect 11520 -312 11528 -248
rect 11592 -312 11600 -248
rect 11520 -328 11600 -312
rect 11520 -392 11528 -328
rect 11592 -392 11600 -328
rect 11520 -408 11600 -392
rect 11520 -472 11528 -408
rect 11592 -472 11600 -408
rect 11520 -1920 11600 -472
rect 11840 -88 11920 8
rect 11840 -152 11848 -88
rect 11912 -152 11920 -88
rect 11840 -168 11920 -152
rect 11840 -232 11848 -168
rect 11912 -232 11920 -168
rect 11840 -248 11920 -232
rect 11840 -312 11848 -248
rect 11912 -312 11920 -248
rect 11840 -328 11920 -312
rect 11840 -392 11848 -328
rect 11912 -392 11920 -328
rect 11840 -408 11920 -392
rect 11840 -472 11848 -408
rect 11912 -472 11920 -408
rect 11840 -1920 11920 -472
rect 12000 31432 12080 31520
rect 12000 31368 12008 31432
rect 12072 31368 12080 31432
rect 12000 31272 12080 31368
rect 12000 31208 12008 31272
rect 12072 31208 12080 31272
rect 12000 31112 12080 31208
rect 12000 31048 12008 31112
rect 12072 31048 12080 31112
rect 12000 30952 12080 31048
rect 12000 30888 12008 30952
rect 12072 30888 12080 30952
rect 12000 30792 12080 30888
rect 12000 30728 12008 30792
rect 12072 30728 12080 30792
rect 12000 30632 12080 30728
rect 12000 30568 12008 30632
rect 12072 30568 12080 30632
rect 12000 30472 12080 30568
rect 12000 30408 12008 30472
rect 12072 30408 12080 30472
rect 12000 30312 12080 30408
rect 12000 30248 12008 30312
rect 12072 30248 12080 30312
rect 12000 30152 12080 30248
rect 12000 30088 12008 30152
rect 12072 30088 12080 30152
rect 12000 29992 12080 30088
rect 12000 29928 12008 29992
rect 12072 29928 12080 29992
rect 12000 29832 12080 29928
rect 12000 29768 12008 29832
rect 12072 29768 12080 29832
rect 12000 29672 12080 29768
rect 12000 29608 12008 29672
rect 12072 29608 12080 29672
rect 12000 29512 12080 29608
rect 12000 29448 12008 29512
rect 12072 29448 12080 29512
rect 12000 29352 12080 29448
rect 12000 29288 12008 29352
rect 12072 29288 12080 29352
rect 12000 29192 12080 29288
rect 12000 29128 12008 29192
rect 12072 29128 12080 29192
rect 12000 29032 12080 29128
rect 12000 28968 12008 29032
rect 12072 28968 12080 29032
rect 12000 28872 12080 28968
rect 12000 28808 12008 28872
rect 12072 28808 12080 28872
rect 12000 28712 12080 28808
rect 12000 28648 12008 28712
rect 12072 28648 12080 28712
rect 12000 28552 12080 28648
rect 12000 28488 12008 28552
rect 12072 28488 12080 28552
rect 12000 28392 12080 28488
rect 12000 28328 12008 28392
rect 12072 28328 12080 28392
rect 12000 28232 12080 28328
rect 12000 28168 12008 28232
rect 12072 28168 12080 28232
rect 12000 28072 12080 28168
rect 12000 28008 12008 28072
rect 12072 28008 12080 28072
rect 12000 27912 12080 28008
rect 12000 27848 12008 27912
rect 12072 27848 12080 27912
rect 12000 27752 12080 27848
rect 12000 27688 12008 27752
rect 12072 27688 12080 27752
rect 12000 27592 12080 27688
rect 12000 27528 12008 27592
rect 12072 27528 12080 27592
rect 12000 27432 12080 27528
rect 12000 27368 12008 27432
rect 12072 27368 12080 27432
rect 12000 27272 12080 27368
rect 12000 27208 12008 27272
rect 12072 27208 12080 27272
rect 12000 27112 12080 27208
rect 12000 27048 12008 27112
rect 12072 27048 12080 27112
rect 12000 26952 12080 27048
rect 12000 26888 12008 26952
rect 12072 26888 12080 26952
rect 12000 26792 12080 26888
rect 12000 26728 12008 26792
rect 12072 26728 12080 26792
rect 12000 26632 12080 26728
rect 12000 26568 12008 26632
rect 12072 26568 12080 26632
rect 12000 26472 12080 26568
rect 12000 26408 12008 26472
rect 12072 26408 12080 26472
rect 12000 26312 12080 26408
rect 12000 26248 12008 26312
rect 12072 26248 12080 26312
rect 12000 26152 12080 26248
rect 12000 26088 12008 26152
rect 12072 26088 12080 26152
rect 12000 25992 12080 26088
rect 12000 25928 12008 25992
rect 12072 25928 12080 25992
rect 12000 25832 12080 25928
rect 12000 25768 12008 25832
rect 12072 25768 12080 25832
rect 12000 25672 12080 25768
rect 12000 25608 12008 25672
rect 12072 25608 12080 25672
rect 12000 25512 12080 25608
rect 12000 25448 12008 25512
rect 12072 25448 12080 25512
rect 12000 25352 12080 25448
rect 12000 25288 12008 25352
rect 12072 25288 12080 25352
rect 12000 25192 12080 25288
rect 12000 25128 12008 25192
rect 12072 25128 12080 25192
rect 12000 25032 12080 25128
rect 12000 24968 12008 25032
rect 12072 24968 12080 25032
rect 12000 24872 12080 24968
rect 12000 24808 12008 24872
rect 12072 24808 12080 24872
rect 12000 24712 12080 24808
rect 12000 24648 12008 24712
rect 12072 24648 12080 24712
rect 12000 24552 12080 24648
rect 12000 24488 12008 24552
rect 12072 24488 12080 24552
rect 12000 24392 12080 24488
rect 12000 24328 12008 24392
rect 12072 24328 12080 24392
rect 12000 24232 12080 24328
rect 12000 24168 12008 24232
rect 12072 24168 12080 24232
rect 12000 24072 12080 24168
rect 12000 24008 12008 24072
rect 12072 24008 12080 24072
rect 12000 23912 12080 24008
rect 12000 23848 12008 23912
rect 12072 23848 12080 23912
rect 12000 23752 12080 23848
rect 12000 23688 12008 23752
rect 12072 23688 12080 23752
rect 12000 23592 12080 23688
rect 12000 23528 12008 23592
rect 12072 23528 12080 23592
rect 12000 23432 12080 23528
rect 12000 23368 12008 23432
rect 12072 23368 12080 23432
rect 12000 23272 12080 23368
rect 12000 23208 12008 23272
rect 12072 23208 12080 23272
rect 12000 23112 12080 23208
rect 12000 23048 12008 23112
rect 12072 23048 12080 23112
rect 12000 22952 12080 23048
rect 12000 22888 12008 22952
rect 12072 22888 12080 22952
rect 12000 22792 12080 22888
rect 12000 22728 12008 22792
rect 12072 22728 12080 22792
rect 12000 22632 12080 22728
rect 12000 22568 12008 22632
rect 12072 22568 12080 22632
rect 12000 22472 12080 22568
rect 12000 22408 12008 22472
rect 12072 22408 12080 22472
rect 12000 22312 12080 22408
rect 12000 22248 12008 22312
rect 12072 22248 12080 22312
rect 12000 22152 12080 22248
rect 12000 22088 12008 22152
rect 12072 22088 12080 22152
rect 12000 21992 12080 22088
rect 12000 21928 12008 21992
rect 12072 21928 12080 21992
rect 12000 21832 12080 21928
rect 12000 21768 12008 21832
rect 12072 21768 12080 21832
rect 12000 21672 12080 21768
rect 12000 21608 12008 21672
rect 12072 21608 12080 21672
rect 12000 21512 12080 21608
rect 12000 21448 12008 21512
rect 12072 21448 12080 21512
rect 12000 21352 12080 21448
rect 12000 21288 12008 21352
rect 12072 21288 12080 21352
rect 12000 21192 12080 21288
rect 12000 21128 12008 21192
rect 12072 21128 12080 21192
rect 12000 21032 12080 21128
rect 12000 20968 12008 21032
rect 12072 20968 12080 21032
rect 12000 20872 12080 20968
rect 12000 20808 12008 20872
rect 12072 20808 12080 20872
rect 12000 20712 12080 20808
rect 12000 20648 12008 20712
rect 12072 20648 12080 20712
rect 12000 20552 12080 20648
rect 12000 20488 12008 20552
rect 12072 20488 12080 20552
rect 12000 20392 12080 20488
rect 12000 20328 12008 20392
rect 12072 20328 12080 20392
rect 12000 20232 12080 20328
rect 12000 20168 12008 20232
rect 12072 20168 12080 20232
rect 12000 20072 12080 20168
rect 12000 20008 12008 20072
rect 12072 20008 12080 20072
rect 12000 19912 12080 20008
rect 12000 19848 12008 19912
rect 12072 19848 12080 19912
rect 12000 19752 12080 19848
rect 12000 19688 12008 19752
rect 12072 19688 12080 19752
rect 12000 19592 12080 19688
rect 12000 19528 12008 19592
rect 12072 19528 12080 19592
rect 12000 19432 12080 19528
rect 12000 19368 12008 19432
rect 12072 19368 12080 19432
rect 12000 19272 12080 19368
rect 12000 19208 12008 19272
rect 12072 19208 12080 19272
rect 12000 19112 12080 19208
rect 12000 19048 12008 19112
rect 12072 19048 12080 19112
rect 12000 18952 12080 19048
rect 12000 18888 12008 18952
rect 12072 18888 12080 18952
rect 12000 18792 12080 18888
rect 12000 18728 12008 18792
rect 12072 18728 12080 18792
rect 12000 18632 12080 18728
rect 12000 18568 12008 18632
rect 12072 18568 12080 18632
rect 12000 18472 12080 18568
rect 12000 18408 12008 18472
rect 12072 18408 12080 18472
rect 12000 18312 12080 18408
rect 12000 18248 12008 18312
rect 12072 18248 12080 18312
rect 12000 18152 12080 18248
rect 12000 18088 12008 18152
rect 12072 18088 12080 18152
rect 12000 17992 12080 18088
rect 12000 17928 12008 17992
rect 12072 17928 12080 17992
rect 12000 17832 12080 17928
rect 12000 17768 12008 17832
rect 12072 17768 12080 17832
rect 12000 17672 12080 17768
rect 12000 17608 12008 17672
rect 12072 17608 12080 17672
rect 12000 17512 12080 17608
rect 12000 17448 12008 17512
rect 12072 17448 12080 17512
rect 12000 17352 12080 17448
rect 12000 17288 12008 17352
rect 12072 17288 12080 17352
rect 12000 17192 12080 17288
rect 12000 17128 12008 17192
rect 12072 17128 12080 17192
rect 12000 17032 12080 17128
rect 12000 16968 12008 17032
rect 12072 16968 12080 17032
rect 12000 16872 12080 16968
rect 12000 16808 12008 16872
rect 12072 16808 12080 16872
rect 12000 16712 12080 16808
rect 12000 16648 12008 16712
rect 12072 16648 12080 16712
rect 12000 16552 12080 16648
rect 12000 16488 12008 16552
rect 12072 16488 12080 16552
rect 12000 16392 12080 16488
rect 12000 16328 12008 16392
rect 12072 16328 12080 16392
rect 12000 16232 12080 16328
rect 12000 16168 12008 16232
rect 12072 16168 12080 16232
rect 12000 16072 12080 16168
rect 12000 16008 12008 16072
rect 12072 16008 12080 16072
rect 12000 15912 12080 16008
rect 12000 15848 12008 15912
rect 12072 15848 12080 15912
rect 12000 15752 12080 15848
rect 12000 15688 12008 15752
rect 12072 15688 12080 15752
rect 12000 15592 12080 15688
rect 12000 15528 12008 15592
rect 12072 15528 12080 15592
rect 12000 15432 12080 15528
rect 12000 15368 12008 15432
rect 12072 15368 12080 15432
rect 12000 15272 12080 15368
rect 12000 15208 12008 15272
rect 12072 15208 12080 15272
rect 12000 15112 12080 15208
rect 12000 15048 12008 15112
rect 12072 15048 12080 15112
rect 12000 14952 12080 15048
rect 12000 14888 12008 14952
rect 12072 14888 12080 14952
rect 12000 14792 12080 14888
rect 12000 14728 12008 14792
rect 12072 14728 12080 14792
rect 12000 14632 12080 14728
rect 12000 14568 12008 14632
rect 12072 14568 12080 14632
rect 12000 14472 12080 14568
rect 12000 14408 12008 14472
rect 12072 14408 12080 14472
rect 12000 14312 12080 14408
rect 12000 14248 12008 14312
rect 12072 14248 12080 14312
rect 12000 14152 12080 14248
rect 12000 14088 12008 14152
rect 12072 14088 12080 14152
rect 12000 13992 12080 14088
rect 12000 13928 12008 13992
rect 12072 13928 12080 13992
rect 12000 13832 12080 13928
rect 12000 13768 12008 13832
rect 12072 13768 12080 13832
rect 12000 13672 12080 13768
rect 12000 13608 12008 13672
rect 12072 13608 12080 13672
rect 12000 13512 12080 13608
rect 12000 13448 12008 13512
rect 12072 13448 12080 13512
rect 12000 13352 12080 13448
rect 12000 13288 12008 13352
rect 12072 13288 12080 13352
rect 12000 13192 12080 13288
rect 12000 13128 12008 13192
rect 12072 13128 12080 13192
rect 12000 13032 12080 13128
rect 12000 12968 12008 13032
rect 12072 12968 12080 13032
rect 12000 12872 12080 12968
rect 12000 12808 12008 12872
rect 12072 12808 12080 12872
rect 12000 12712 12080 12808
rect 12000 12648 12008 12712
rect 12072 12648 12080 12712
rect 12000 12552 12080 12648
rect 12000 12488 12008 12552
rect 12072 12488 12080 12552
rect 12000 12392 12080 12488
rect 12000 12328 12008 12392
rect 12072 12328 12080 12392
rect 12000 12232 12080 12328
rect 12000 12168 12008 12232
rect 12072 12168 12080 12232
rect 12000 12072 12080 12168
rect 12000 12008 12008 12072
rect 12072 12008 12080 12072
rect 12000 11912 12080 12008
rect 12000 11848 12008 11912
rect 12072 11848 12080 11912
rect 12000 11752 12080 11848
rect 12000 11688 12008 11752
rect 12072 11688 12080 11752
rect 12000 11592 12080 11688
rect 12000 11528 12008 11592
rect 12072 11528 12080 11592
rect 12000 11432 12080 11528
rect 12000 11368 12008 11432
rect 12072 11368 12080 11432
rect 12000 11272 12080 11368
rect 12000 11208 12008 11272
rect 12072 11208 12080 11272
rect 12000 11112 12080 11208
rect 12000 11048 12008 11112
rect 12072 11048 12080 11112
rect 12000 10952 12080 11048
rect 12000 10888 12008 10952
rect 12072 10888 12080 10952
rect 12000 10792 12080 10888
rect 12000 10728 12008 10792
rect 12072 10728 12080 10792
rect 12000 10632 12080 10728
rect 12000 10568 12008 10632
rect 12072 10568 12080 10632
rect 12000 10472 12080 10568
rect 12000 10408 12008 10472
rect 12072 10408 12080 10472
rect 12000 10312 12080 10408
rect 12000 10248 12008 10312
rect 12072 10248 12080 10312
rect 12000 10152 12080 10248
rect 12000 10088 12008 10152
rect 12072 10088 12080 10152
rect 12000 9992 12080 10088
rect 12000 9928 12008 9992
rect 12072 9928 12080 9992
rect 12000 9832 12080 9928
rect 12000 9768 12008 9832
rect 12072 9768 12080 9832
rect 12000 9672 12080 9768
rect 12000 9608 12008 9672
rect 12072 9608 12080 9672
rect 12000 9512 12080 9608
rect 12000 9448 12008 9512
rect 12072 9448 12080 9512
rect 12000 9352 12080 9448
rect 12000 9288 12008 9352
rect 12072 9288 12080 9352
rect 12000 9192 12080 9288
rect 12000 9128 12008 9192
rect 12072 9128 12080 9192
rect 12000 9032 12080 9128
rect 12000 8968 12008 9032
rect 12072 8968 12080 9032
rect 12000 8872 12080 8968
rect 12000 8808 12008 8872
rect 12072 8808 12080 8872
rect 12000 8712 12080 8808
rect 12000 8648 12008 8712
rect 12072 8648 12080 8712
rect 12000 8552 12080 8648
rect 12000 8488 12008 8552
rect 12072 8488 12080 8552
rect 12000 8392 12080 8488
rect 12000 8328 12008 8392
rect 12072 8328 12080 8392
rect 12000 8232 12080 8328
rect 12000 8168 12008 8232
rect 12072 8168 12080 8232
rect 12000 8072 12080 8168
rect 12000 8008 12008 8072
rect 12072 8008 12080 8072
rect 12000 7912 12080 8008
rect 12000 7848 12008 7912
rect 12072 7848 12080 7912
rect 12000 7752 12080 7848
rect 12000 7688 12008 7752
rect 12072 7688 12080 7752
rect 12000 7592 12080 7688
rect 12000 7528 12008 7592
rect 12072 7528 12080 7592
rect 12000 7432 12080 7528
rect 12000 7368 12008 7432
rect 12072 7368 12080 7432
rect 12000 7272 12080 7368
rect 12000 7208 12008 7272
rect 12072 7208 12080 7272
rect 12000 7112 12080 7208
rect 12000 7048 12008 7112
rect 12072 7048 12080 7112
rect 12000 6952 12080 7048
rect 12000 6888 12008 6952
rect 12072 6888 12080 6952
rect 12000 6792 12080 6888
rect 12000 6728 12008 6792
rect 12072 6728 12080 6792
rect 12000 6632 12080 6728
rect 12000 6568 12008 6632
rect 12072 6568 12080 6632
rect 12000 6472 12080 6568
rect 12000 6408 12008 6472
rect 12072 6408 12080 6472
rect 12000 6312 12080 6408
rect 12000 6248 12008 6312
rect 12072 6248 12080 6312
rect 12000 6152 12080 6248
rect 12000 6088 12008 6152
rect 12072 6088 12080 6152
rect 12000 5992 12080 6088
rect 12000 5928 12008 5992
rect 12072 5928 12080 5992
rect 12000 5832 12080 5928
rect 12000 5768 12008 5832
rect 12072 5768 12080 5832
rect 12000 5672 12080 5768
rect 12000 5608 12008 5672
rect 12072 5608 12080 5672
rect 12000 5512 12080 5608
rect 12000 5448 12008 5512
rect 12072 5448 12080 5512
rect 12000 5352 12080 5448
rect 12000 5288 12008 5352
rect 12072 5288 12080 5352
rect 12000 5192 12080 5288
rect 12000 5128 12008 5192
rect 12072 5128 12080 5192
rect 12000 5032 12080 5128
rect 12000 4968 12008 5032
rect 12072 4968 12080 5032
rect 12000 4872 12080 4968
rect 12000 4808 12008 4872
rect 12072 4808 12080 4872
rect 12000 4712 12080 4808
rect 12000 4648 12008 4712
rect 12072 4648 12080 4712
rect 12000 4552 12080 4648
rect 12000 4488 12008 4552
rect 12072 4488 12080 4552
rect 12000 4392 12080 4488
rect 12000 4328 12008 4392
rect 12072 4328 12080 4392
rect 12000 4232 12080 4328
rect 12000 4168 12008 4232
rect 12072 4168 12080 4232
rect 12000 4072 12080 4168
rect 12000 4008 12008 4072
rect 12072 4008 12080 4072
rect 12000 3912 12080 4008
rect 12000 3848 12008 3912
rect 12072 3848 12080 3912
rect 12000 3752 12080 3848
rect 12000 3688 12008 3752
rect 12072 3688 12080 3752
rect 12000 3592 12080 3688
rect 12000 3528 12008 3592
rect 12072 3528 12080 3592
rect 12000 3432 12080 3528
rect 12000 3368 12008 3432
rect 12072 3368 12080 3432
rect 12000 3272 12080 3368
rect 12000 3208 12008 3272
rect 12072 3208 12080 3272
rect 12000 3112 12080 3208
rect 12000 3048 12008 3112
rect 12072 3048 12080 3112
rect 12000 2952 12080 3048
rect 12000 2888 12008 2952
rect 12072 2888 12080 2952
rect 12000 2792 12080 2888
rect 12000 2728 12008 2792
rect 12072 2728 12080 2792
rect 12000 2632 12080 2728
rect 12000 2568 12008 2632
rect 12072 2568 12080 2632
rect 12000 2472 12080 2568
rect 12000 2408 12008 2472
rect 12072 2408 12080 2472
rect 12000 2312 12080 2408
rect 12000 2248 12008 2312
rect 12072 2248 12080 2312
rect 12000 2152 12080 2248
rect 12000 2088 12008 2152
rect 12072 2088 12080 2152
rect 12000 1992 12080 2088
rect 12000 1928 12008 1992
rect 12072 1928 12080 1992
rect 12000 1832 12080 1928
rect 12000 1768 12008 1832
rect 12072 1768 12080 1832
rect 12000 1672 12080 1768
rect 12000 1608 12008 1672
rect 12072 1608 12080 1672
rect 12000 1512 12080 1608
rect 12000 1448 12008 1512
rect 12072 1448 12080 1512
rect 12000 1352 12080 1448
rect 12000 1288 12008 1352
rect 12072 1288 12080 1352
rect 12000 1192 12080 1288
rect 12000 1128 12008 1192
rect 12072 1128 12080 1192
rect 12000 1032 12080 1128
rect 12000 968 12008 1032
rect 12072 968 12080 1032
rect 12000 872 12080 968
rect 12000 808 12008 872
rect 12072 808 12080 872
rect 12000 712 12080 808
rect 12000 648 12008 712
rect 12072 648 12080 712
rect 12000 552 12080 648
rect 12000 488 12008 552
rect 12072 488 12080 552
rect 12000 392 12080 488
rect 12000 328 12008 392
rect 12072 328 12080 392
rect 12000 232 12080 328
rect 12000 168 12008 232
rect 12072 168 12080 232
rect 12000 72 12080 168
rect 12000 8 12008 72
rect 12072 8 12080 72
rect 12000 -1048 12080 8
rect 12160 9188 12240 31520
rect 12160 9132 12172 9188
rect 12228 9132 12240 9188
rect 12160 1828 12240 9132
rect 12160 1772 12172 1828
rect 12228 1772 12240 1828
rect 12160 0 12240 1772
rect 12320 31432 12400 31520
rect 12320 31368 12328 31432
rect 12392 31368 12400 31432
rect 12320 31272 12400 31368
rect 12320 31208 12328 31272
rect 12392 31208 12400 31272
rect 12320 31112 12400 31208
rect 12320 31048 12328 31112
rect 12392 31048 12400 31112
rect 12320 30952 12400 31048
rect 12320 30888 12328 30952
rect 12392 30888 12400 30952
rect 12320 30792 12400 30888
rect 12320 30728 12328 30792
rect 12392 30728 12400 30792
rect 12320 30632 12400 30728
rect 12320 30568 12328 30632
rect 12392 30568 12400 30632
rect 12320 30472 12400 30568
rect 12320 30408 12328 30472
rect 12392 30408 12400 30472
rect 12320 30312 12400 30408
rect 12320 30248 12328 30312
rect 12392 30248 12400 30312
rect 12320 30152 12400 30248
rect 12320 30088 12328 30152
rect 12392 30088 12400 30152
rect 12320 29992 12400 30088
rect 12320 29928 12328 29992
rect 12392 29928 12400 29992
rect 12320 29832 12400 29928
rect 12320 29768 12328 29832
rect 12392 29768 12400 29832
rect 12320 29672 12400 29768
rect 12320 29608 12328 29672
rect 12392 29608 12400 29672
rect 12320 29512 12400 29608
rect 12320 29448 12328 29512
rect 12392 29448 12400 29512
rect 12320 29352 12400 29448
rect 12320 29288 12328 29352
rect 12392 29288 12400 29352
rect 12320 29192 12400 29288
rect 12320 29128 12328 29192
rect 12392 29128 12400 29192
rect 12320 29032 12400 29128
rect 12320 28968 12328 29032
rect 12392 28968 12400 29032
rect 12320 28872 12400 28968
rect 12320 28808 12328 28872
rect 12392 28808 12400 28872
rect 12320 28712 12400 28808
rect 12320 28648 12328 28712
rect 12392 28648 12400 28712
rect 12320 28552 12400 28648
rect 12320 28488 12328 28552
rect 12392 28488 12400 28552
rect 12320 28392 12400 28488
rect 12320 28328 12328 28392
rect 12392 28328 12400 28392
rect 12320 28232 12400 28328
rect 12320 28168 12328 28232
rect 12392 28168 12400 28232
rect 12320 28072 12400 28168
rect 12320 28008 12328 28072
rect 12392 28008 12400 28072
rect 12320 27912 12400 28008
rect 12320 27848 12328 27912
rect 12392 27848 12400 27912
rect 12320 27752 12400 27848
rect 12320 27688 12328 27752
rect 12392 27688 12400 27752
rect 12320 27592 12400 27688
rect 12320 27528 12328 27592
rect 12392 27528 12400 27592
rect 12320 27432 12400 27528
rect 12320 27368 12328 27432
rect 12392 27368 12400 27432
rect 12320 27272 12400 27368
rect 12320 27208 12328 27272
rect 12392 27208 12400 27272
rect 12320 27112 12400 27208
rect 12320 27048 12328 27112
rect 12392 27048 12400 27112
rect 12320 26952 12400 27048
rect 12320 26888 12328 26952
rect 12392 26888 12400 26952
rect 12320 26792 12400 26888
rect 12320 26728 12328 26792
rect 12392 26728 12400 26792
rect 12320 26632 12400 26728
rect 12320 26568 12328 26632
rect 12392 26568 12400 26632
rect 12320 26472 12400 26568
rect 12320 26408 12328 26472
rect 12392 26408 12400 26472
rect 12320 26312 12400 26408
rect 12320 26248 12328 26312
rect 12392 26248 12400 26312
rect 12320 26152 12400 26248
rect 12320 26088 12328 26152
rect 12392 26088 12400 26152
rect 12320 25992 12400 26088
rect 12320 25928 12328 25992
rect 12392 25928 12400 25992
rect 12320 25832 12400 25928
rect 12320 25768 12328 25832
rect 12392 25768 12400 25832
rect 12320 25672 12400 25768
rect 12320 25608 12328 25672
rect 12392 25608 12400 25672
rect 12320 25512 12400 25608
rect 12320 25448 12328 25512
rect 12392 25448 12400 25512
rect 12320 25352 12400 25448
rect 12320 25288 12328 25352
rect 12392 25288 12400 25352
rect 12320 25192 12400 25288
rect 12320 25128 12328 25192
rect 12392 25128 12400 25192
rect 12320 25032 12400 25128
rect 12320 24968 12328 25032
rect 12392 24968 12400 25032
rect 12320 24872 12400 24968
rect 12320 24808 12328 24872
rect 12392 24808 12400 24872
rect 12320 24712 12400 24808
rect 12320 24648 12328 24712
rect 12392 24648 12400 24712
rect 12320 24552 12400 24648
rect 12320 24488 12328 24552
rect 12392 24488 12400 24552
rect 12320 24392 12400 24488
rect 12320 24328 12328 24392
rect 12392 24328 12400 24392
rect 12320 24232 12400 24328
rect 12320 24168 12328 24232
rect 12392 24168 12400 24232
rect 12320 24072 12400 24168
rect 12320 24008 12328 24072
rect 12392 24008 12400 24072
rect 12320 23912 12400 24008
rect 12320 23848 12328 23912
rect 12392 23848 12400 23912
rect 12320 23752 12400 23848
rect 12320 23688 12328 23752
rect 12392 23688 12400 23752
rect 12320 23592 12400 23688
rect 12320 23528 12328 23592
rect 12392 23528 12400 23592
rect 12320 23432 12400 23528
rect 12320 23368 12328 23432
rect 12392 23368 12400 23432
rect 12320 23272 12400 23368
rect 12320 23208 12328 23272
rect 12392 23208 12400 23272
rect 12320 23112 12400 23208
rect 12320 23048 12328 23112
rect 12392 23048 12400 23112
rect 12320 22952 12400 23048
rect 12320 22888 12328 22952
rect 12392 22888 12400 22952
rect 12320 22792 12400 22888
rect 12320 22728 12328 22792
rect 12392 22728 12400 22792
rect 12320 22632 12400 22728
rect 12320 22568 12328 22632
rect 12392 22568 12400 22632
rect 12320 22472 12400 22568
rect 12320 22408 12328 22472
rect 12392 22408 12400 22472
rect 12320 22312 12400 22408
rect 12320 22248 12328 22312
rect 12392 22248 12400 22312
rect 12320 22152 12400 22248
rect 12320 22088 12328 22152
rect 12392 22088 12400 22152
rect 12320 21992 12400 22088
rect 12320 21928 12328 21992
rect 12392 21928 12400 21992
rect 12320 21832 12400 21928
rect 12320 21768 12328 21832
rect 12392 21768 12400 21832
rect 12320 21672 12400 21768
rect 12320 21608 12328 21672
rect 12392 21608 12400 21672
rect 12320 21512 12400 21608
rect 12320 21448 12328 21512
rect 12392 21448 12400 21512
rect 12320 21352 12400 21448
rect 12320 21288 12328 21352
rect 12392 21288 12400 21352
rect 12320 21192 12400 21288
rect 12320 21128 12328 21192
rect 12392 21128 12400 21192
rect 12320 21032 12400 21128
rect 12320 20968 12328 21032
rect 12392 20968 12400 21032
rect 12320 20872 12400 20968
rect 12320 20808 12328 20872
rect 12392 20808 12400 20872
rect 12320 20712 12400 20808
rect 12320 20648 12328 20712
rect 12392 20648 12400 20712
rect 12320 20552 12400 20648
rect 12320 20488 12328 20552
rect 12392 20488 12400 20552
rect 12320 20392 12400 20488
rect 12320 20328 12328 20392
rect 12392 20328 12400 20392
rect 12320 20232 12400 20328
rect 12320 20168 12328 20232
rect 12392 20168 12400 20232
rect 12320 20072 12400 20168
rect 12320 20008 12328 20072
rect 12392 20008 12400 20072
rect 12320 19912 12400 20008
rect 12320 19848 12328 19912
rect 12392 19848 12400 19912
rect 12320 19752 12400 19848
rect 12320 19688 12328 19752
rect 12392 19688 12400 19752
rect 12320 19592 12400 19688
rect 12320 19528 12328 19592
rect 12392 19528 12400 19592
rect 12320 19432 12400 19528
rect 12320 19368 12328 19432
rect 12392 19368 12400 19432
rect 12320 19272 12400 19368
rect 12320 19208 12328 19272
rect 12392 19208 12400 19272
rect 12320 19112 12400 19208
rect 12320 19048 12328 19112
rect 12392 19048 12400 19112
rect 12320 18952 12400 19048
rect 12320 18888 12328 18952
rect 12392 18888 12400 18952
rect 12320 18792 12400 18888
rect 12320 18728 12328 18792
rect 12392 18728 12400 18792
rect 12320 18632 12400 18728
rect 12320 18568 12328 18632
rect 12392 18568 12400 18632
rect 12320 18472 12400 18568
rect 12320 18408 12328 18472
rect 12392 18408 12400 18472
rect 12320 18312 12400 18408
rect 12320 18248 12328 18312
rect 12392 18248 12400 18312
rect 12320 18152 12400 18248
rect 12320 18088 12328 18152
rect 12392 18088 12400 18152
rect 12320 17992 12400 18088
rect 12320 17928 12328 17992
rect 12392 17928 12400 17992
rect 12320 17832 12400 17928
rect 12320 17768 12328 17832
rect 12392 17768 12400 17832
rect 12320 17672 12400 17768
rect 12320 17608 12328 17672
rect 12392 17608 12400 17672
rect 12320 17512 12400 17608
rect 12320 17448 12328 17512
rect 12392 17448 12400 17512
rect 12320 17352 12400 17448
rect 12320 17288 12328 17352
rect 12392 17288 12400 17352
rect 12320 17192 12400 17288
rect 12320 17128 12328 17192
rect 12392 17128 12400 17192
rect 12320 17032 12400 17128
rect 12320 16968 12328 17032
rect 12392 16968 12400 17032
rect 12320 16872 12400 16968
rect 12320 16808 12328 16872
rect 12392 16808 12400 16872
rect 12320 16712 12400 16808
rect 12320 16648 12328 16712
rect 12392 16648 12400 16712
rect 12320 16552 12400 16648
rect 12320 16488 12328 16552
rect 12392 16488 12400 16552
rect 12320 16392 12400 16488
rect 12320 16328 12328 16392
rect 12392 16328 12400 16392
rect 12320 16232 12400 16328
rect 12320 16168 12328 16232
rect 12392 16168 12400 16232
rect 12320 16072 12400 16168
rect 12320 16008 12328 16072
rect 12392 16008 12400 16072
rect 12320 15912 12400 16008
rect 12320 15848 12328 15912
rect 12392 15848 12400 15912
rect 12320 15752 12400 15848
rect 12320 15688 12328 15752
rect 12392 15688 12400 15752
rect 12320 15592 12400 15688
rect 12320 15528 12328 15592
rect 12392 15528 12400 15592
rect 12320 15432 12400 15528
rect 12320 15368 12328 15432
rect 12392 15368 12400 15432
rect 12320 15272 12400 15368
rect 12320 15208 12328 15272
rect 12392 15208 12400 15272
rect 12320 15112 12400 15208
rect 12320 15048 12328 15112
rect 12392 15048 12400 15112
rect 12320 14952 12400 15048
rect 12320 14888 12328 14952
rect 12392 14888 12400 14952
rect 12320 14792 12400 14888
rect 12320 14728 12328 14792
rect 12392 14728 12400 14792
rect 12320 14632 12400 14728
rect 12320 14568 12328 14632
rect 12392 14568 12400 14632
rect 12320 14472 12400 14568
rect 12320 14408 12328 14472
rect 12392 14408 12400 14472
rect 12320 14312 12400 14408
rect 12320 14248 12328 14312
rect 12392 14248 12400 14312
rect 12320 14152 12400 14248
rect 12320 14088 12328 14152
rect 12392 14088 12400 14152
rect 12320 13992 12400 14088
rect 12320 13928 12328 13992
rect 12392 13928 12400 13992
rect 12320 13832 12400 13928
rect 12320 13768 12328 13832
rect 12392 13768 12400 13832
rect 12320 13672 12400 13768
rect 12320 13608 12328 13672
rect 12392 13608 12400 13672
rect 12320 13512 12400 13608
rect 12320 13448 12328 13512
rect 12392 13448 12400 13512
rect 12320 13352 12400 13448
rect 12320 13288 12328 13352
rect 12392 13288 12400 13352
rect 12320 13192 12400 13288
rect 12320 13128 12328 13192
rect 12392 13128 12400 13192
rect 12320 13032 12400 13128
rect 12320 12968 12328 13032
rect 12392 12968 12400 13032
rect 12320 12872 12400 12968
rect 12320 12808 12328 12872
rect 12392 12808 12400 12872
rect 12320 12712 12400 12808
rect 12320 12648 12328 12712
rect 12392 12648 12400 12712
rect 12320 12552 12400 12648
rect 12320 12488 12328 12552
rect 12392 12488 12400 12552
rect 12320 12392 12400 12488
rect 12320 12328 12328 12392
rect 12392 12328 12400 12392
rect 12320 12232 12400 12328
rect 12320 12168 12328 12232
rect 12392 12168 12400 12232
rect 12320 12072 12400 12168
rect 12320 12008 12328 12072
rect 12392 12008 12400 12072
rect 12320 11912 12400 12008
rect 12320 11848 12328 11912
rect 12392 11848 12400 11912
rect 12320 11752 12400 11848
rect 12320 11688 12328 11752
rect 12392 11688 12400 11752
rect 12320 11592 12400 11688
rect 12320 11528 12328 11592
rect 12392 11528 12400 11592
rect 12320 11432 12400 11528
rect 12320 11368 12328 11432
rect 12392 11368 12400 11432
rect 12320 11272 12400 11368
rect 12320 11208 12328 11272
rect 12392 11208 12400 11272
rect 12320 11112 12400 11208
rect 12320 11048 12328 11112
rect 12392 11048 12400 11112
rect 12320 10952 12400 11048
rect 12320 10888 12328 10952
rect 12392 10888 12400 10952
rect 12320 10792 12400 10888
rect 12320 10728 12328 10792
rect 12392 10728 12400 10792
rect 12320 10632 12400 10728
rect 12320 10568 12328 10632
rect 12392 10568 12400 10632
rect 12320 10472 12400 10568
rect 12320 10408 12328 10472
rect 12392 10408 12400 10472
rect 12320 10312 12400 10408
rect 12320 10248 12328 10312
rect 12392 10248 12400 10312
rect 12320 10152 12400 10248
rect 12320 10088 12328 10152
rect 12392 10088 12400 10152
rect 12320 9992 12400 10088
rect 12320 9928 12328 9992
rect 12392 9928 12400 9992
rect 12320 9832 12400 9928
rect 12320 9768 12328 9832
rect 12392 9768 12400 9832
rect 12320 9672 12400 9768
rect 12320 9608 12328 9672
rect 12392 9608 12400 9672
rect 12320 9512 12400 9608
rect 12320 9448 12328 9512
rect 12392 9448 12400 9512
rect 12320 9352 12400 9448
rect 12320 9288 12328 9352
rect 12392 9288 12400 9352
rect 12320 9192 12400 9288
rect 12320 9128 12328 9192
rect 12392 9128 12400 9192
rect 12320 9032 12400 9128
rect 12320 8968 12328 9032
rect 12392 8968 12400 9032
rect 12320 8872 12400 8968
rect 12320 8808 12328 8872
rect 12392 8808 12400 8872
rect 12320 8712 12400 8808
rect 12320 8648 12328 8712
rect 12392 8648 12400 8712
rect 12320 8552 12400 8648
rect 12320 8488 12328 8552
rect 12392 8488 12400 8552
rect 12320 8392 12400 8488
rect 12320 8328 12328 8392
rect 12392 8328 12400 8392
rect 12320 8232 12400 8328
rect 12320 8168 12328 8232
rect 12392 8168 12400 8232
rect 12320 8072 12400 8168
rect 12320 8008 12328 8072
rect 12392 8008 12400 8072
rect 12320 7912 12400 8008
rect 12320 7848 12328 7912
rect 12392 7848 12400 7912
rect 12320 7752 12400 7848
rect 12320 7688 12328 7752
rect 12392 7688 12400 7752
rect 12320 7592 12400 7688
rect 12320 7528 12328 7592
rect 12392 7528 12400 7592
rect 12320 7432 12400 7528
rect 12320 7368 12328 7432
rect 12392 7368 12400 7432
rect 12320 7272 12400 7368
rect 12320 7208 12328 7272
rect 12392 7208 12400 7272
rect 12320 7112 12400 7208
rect 12320 7048 12328 7112
rect 12392 7048 12400 7112
rect 12320 6952 12400 7048
rect 12320 6888 12328 6952
rect 12392 6888 12400 6952
rect 12320 6792 12400 6888
rect 12320 6728 12328 6792
rect 12392 6728 12400 6792
rect 12320 6632 12400 6728
rect 12320 6568 12328 6632
rect 12392 6568 12400 6632
rect 12320 6472 12400 6568
rect 12320 6408 12328 6472
rect 12392 6408 12400 6472
rect 12320 6312 12400 6408
rect 12320 6248 12328 6312
rect 12392 6248 12400 6312
rect 12320 6152 12400 6248
rect 12320 6088 12328 6152
rect 12392 6088 12400 6152
rect 12320 5992 12400 6088
rect 12320 5928 12328 5992
rect 12392 5928 12400 5992
rect 12320 5832 12400 5928
rect 12320 5768 12328 5832
rect 12392 5768 12400 5832
rect 12320 5672 12400 5768
rect 12320 5608 12328 5672
rect 12392 5608 12400 5672
rect 12320 5512 12400 5608
rect 12320 5448 12328 5512
rect 12392 5448 12400 5512
rect 12320 5352 12400 5448
rect 12320 5288 12328 5352
rect 12392 5288 12400 5352
rect 12320 5192 12400 5288
rect 12320 5128 12328 5192
rect 12392 5128 12400 5192
rect 12320 5032 12400 5128
rect 12320 4968 12328 5032
rect 12392 4968 12400 5032
rect 12320 4872 12400 4968
rect 12320 4808 12328 4872
rect 12392 4808 12400 4872
rect 12320 4712 12400 4808
rect 12320 4648 12328 4712
rect 12392 4648 12400 4712
rect 12320 4552 12400 4648
rect 12320 4488 12328 4552
rect 12392 4488 12400 4552
rect 12320 4392 12400 4488
rect 12320 4328 12328 4392
rect 12392 4328 12400 4392
rect 12320 4232 12400 4328
rect 12320 4168 12328 4232
rect 12392 4168 12400 4232
rect 12320 4072 12400 4168
rect 12320 4008 12328 4072
rect 12392 4008 12400 4072
rect 12320 3912 12400 4008
rect 12320 3848 12328 3912
rect 12392 3848 12400 3912
rect 12320 3752 12400 3848
rect 12320 3688 12328 3752
rect 12392 3688 12400 3752
rect 12320 3592 12400 3688
rect 12320 3528 12328 3592
rect 12392 3528 12400 3592
rect 12320 3432 12400 3528
rect 12320 3368 12328 3432
rect 12392 3368 12400 3432
rect 12320 3272 12400 3368
rect 12320 3208 12328 3272
rect 12392 3208 12400 3272
rect 12320 3112 12400 3208
rect 12320 3048 12328 3112
rect 12392 3048 12400 3112
rect 12320 2952 12400 3048
rect 12320 2888 12328 2952
rect 12392 2888 12400 2952
rect 12320 2792 12400 2888
rect 12320 2728 12328 2792
rect 12392 2728 12400 2792
rect 12320 2632 12400 2728
rect 12320 2568 12328 2632
rect 12392 2568 12400 2632
rect 12320 2472 12400 2568
rect 12320 2408 12328 2472
rect 12392 2408 12400 2472
rect 12320 2312 12400 2408
rect 12320 2248 12328 2312
rect 12392 2248 12400 2312
rect 12320 2152 12400 2248
rect 12320 2088 12328 2152
rect 12392 2088 12400 2152
rect 12320 1992 12400 2088
rect 12320 1928 12328 1992
rect 12392 1928 12400 1992
rect 12320 1832 12400 1928
rect 12320 1768 12328 1832
rect 12392 1768 12400 1832
rect 12320 1672 12400 1768
rect 12320 1608 12328 1672
rect 12392 1608 12400 1672
rect 12320 1512 12400 1608
rect 12320 1448 12328 1512
rect 12392 1448 12400 1512
rect 12320 1352 12400 1448
rect 12320 1288 12328 1352
rect 12392 1288 12400 1352
rect 12320 1192 12400 1288
rect 12320 1128 12328 1192
rect 12392 1128 12400 1192
rect 12320 1032 12400 1128
rect 12320 968 12328 1032
rect 12392 968 12400 1032
rect 12320 872 12400 968
rect 12320 808 12328 872
rect 12392 808 12400 872
rect 12320 712 12400 808
rect 12320 648 12328 712
rect 12392 648 12400 712
rect 12320 552 12400 648
rect 12320 488 12328 552
rect 12392 488 12400 552
rect 12320 392 12400 488
rect 12320 328 12328 392
rect 12392 328 12400 392
rect 12320 232 12400 328
rect 12320 168 12328 232
rect 12392 168 12400 232
rect 12320 72 12400 168
rect 12320 8 12328 72
rect 12392 8 12400 72
rect 12000 -1112 12008 -1048
rect 12072 -1112 12080 -1048
rect 12000 -1128 12080 -1112
rect 12000 -1192 12008 -1128
rect 12072 -1192 12080 -1128
rect 12000 -1208 12080 -1192
rect 12000 -1272 12008 -1208
rect 12072 -1272 12080 -1208
rect 12000 -1288 12080 -1272
rect 12000 -1352 12008 -1288
rect 12072 -1352 12080 -1288
rect 12000 -1368 12080 -1352
rect 12000 -1432 12008 -1368
rect 12072 -1432 12080 -1368
rect 12000 -1920 12080 -1432
rect 12320 -1048 12400 8
rect 12320 -1112 12328 -1048
rect 12392 -1112 12400 -1048
rect 12320 -1128 12400 -1112
rect 12320 -1192 12328 -1128
rect 12392 -1192 12400 -1128
rect 12320 -1208 12400 -1192
rect 12320 -1272 12328 -1208
rect 12392 -1272 12400 -1208
rect 12320 -1288 12400 -1272
rect 12320 -1352 12328 -1288
rect 12392 -1352 12400 -1288
rect 12320 -1368 12400 -1352
rect 12320 -1432 12328 -1368
rect 12392 -1432 12400 -1368
rect 12320 -1920 12400 -1432
rect 9280 -2072 9288 -2008
rect 9352 -2072 9360 -2008
rect 9280 -2080 9360 -2072
rect 20560 -2008 20640 -2000
rect 20560 -2072 20568 -2008
rect 20632 -2072 20640 -2008
rect 400 -2168 480 -2160
rect 400 -2232 408 -2168
rect 472 -2232 480 -2168
rect 400 -2320 480 -2232
rect 2480 -2168 2560 -2160
rect 2480 -2232 2488 -2168
rect 2552 -2232 2560 -2168
rect 2480 -2320 2560 -2232
rect 400 -4480 2560 -2320
rect 2640 -2168 2720 -2160
rect 2640 -2232 2648 -2168
rect 2712 -2232 2720 -2168
rect 2640 -2320 2720 -2232
rect 4720 -2168 4800 -2160
rect 4720 -2232 4728 -2168
rect 4792 -2232 4800 -2168
rect 4720 -2320 4800 -2232
rect 2640 -4480 4800 -2320
rect 4880 -2168 4960 -2160
rect 4880 -2232 4888 -2168
rect 4952 -2232 4960 -2168
rect 4880 -2320 4960 -2232
rect 6960 -2168 7040 -2160
rect 6960 -2232 6968 -2168
rect 7032 -2232 7040 -2168
rect 6960 -2320 7040 -2232
rect 4880 -4480 7040 -2320
rect 7120 -2168 7200 -2160
rect 7120 -2232 7128 -2168
rect 7192 -2232 7200 -2168
rect 7120 -2320 7200 -2232
rect 9120 -2168 9280 -2160
rect 9120 -2232 9208 -2168
rect 9272 -2232 9280 -2168
rect 9120 -2240 9280 -2232
rect 9200 -2320 9280 -2240
rect 7120 -4480 9280 -2320
rect 9360 -2168 9440 -2160
rect 9360 -2232 9368 -2168
rect 9432 -2232 9440 -2168
rect 9360 -2320 9440 -2232
rect 11440 -2168 11520 -2160
rect 11440 -2232 11448 -2168
rect 11512 -2232 11520 -2168
rect 11440 -2320 11520 -2232
rect 9360 -4480 11520 -2320
rect 11600 -2168 11680 -2160
rect 11600 -2232 11608 -2168
rect 11672 -2232 11680 -2168
rect 11600 -2320 11680 -2232
rect 13680 -2168 13760 -2160
rect 13680 -2232 13688 -2168
rect 13752 -2232 13760 -2168
rect 13680 -2320 13760 -2232
rect 11600 -4480 13760 -2320
rect 13840 -2168 13920 -2160
rect 13840 -2232 13848 -2168
rect 13912 -2232 13920 -2168
rect 13840 -2320 13920 -2232
rect 15920 -2168 16000 -2160
rect 15920 -2232 15928 -2168
rect 15992 -2232 16000 -2168
rect 15920 -2320 16000 -2232
rect 13840 -4480 16000 -2320
rect 16080 -2168 16160 -2160
rect 16080 -2232 16088 -2168
rect 16152 -2232 16160 -2168
rect 16080 -2320 16160 -2232
rect 18160 -2168 18240 -2160
rect 18160 -2232 18168 -2168
rect 18232 -2232 18240 -2168
rect 18160 -2320 18240 -2232
rect 16080 -4480 18240 -2320
rect 18320 -2168 18400 -2160
rect 18320 -2232 18328 -2168
rect 18392 -2232 18400 -2168
rect 18320 -2320 18400 -2232
rect 20400 -2168 20480 -2160
rect 20400 -2232 20408 -2168
rect 20472 -2232 20480 -2168
rect 20400 -2320 20480 -2232
rect 18320 -4480 20480 -2320
rect 240 -4632 248 -4568
rect 312 -4632 320 -4568
rect 240 -4640 320 -4632
rect 20560 -4568 20640 -2072
rect 20560 -4632 20568 -4568
rect 20632 -4632 20640 -4568
rect 20560 -4640 20640 -4632
<< via3 >>
rect 8488 31428 8552 31432
rect 8488 31372 8492 31428
rect 8492 31372 8548 31428
rect 8548 31372 8552 31428
rect 8488 31368 8552 31372
rect 8488 31268 8552 31272
rect 8488 31212 8492 31268
rect 8492 31212 8548 31268
rect 8548 31212 8552 31268
rect 8488 31208 8552 31212
rect 8488 31108 8552 31112
rect 8488 31052 8492 31108
rect 8492 31052 8548 31108
rect 8548 31052 8552 31108
rect 8488 31048 8552 31052
rect 8488 30948 8552 30952
rect 8488 30892 8492 30948
rect 8492 30892 8548 30948
rect 8548 30892 8552 30948
rect 8488 30888 8552 30892
rect 8488 30788 8552 30792
rect 8488 30732 8492 30788
rect 8492 30732 8548 30788
rect 8548 30732 8552 30788
rect 8488 30728 8552 30732
rect 8488 30628 8552 30632
rect 8488 30572 8492 30628
rect 8492 30572 8548 30628
rect 8548 30572 8552 30628
rect 8488 30568 8552 30572
rect 8488 30468 8552 30472
rect 8488 30412 8492 30468
rect 8492 30412 8548 30468
rect 8548 30412 8552 30468
rect 8488 30408 8552 30412
rect 8488 30308 8552 30312
rect 8488 30252 8492 30308
rect 8492 30252 8548 30308
rect 8548 30252 8552 30308
rect 8488 30248 8552 30252
rect 8488 30088 8552 30152
rect 8488 29988 8552 29992
rect 8488 29932 8492 29988
rect 8492 29932 8548 29988
rect 8548 29932 8552 29988
rect 8488 29928 8552 29932
rect 8488 29828 8552 29832
rect 8488 29772 8492 29828
rect 8492 29772 8548 29828
rect 8548 29772 8552 29828
rect 8488 29768 8552 29772
rect 8488 29668 8552 29672
rect 8488 29612 8492 29668
rect 8492 29612 8548 29668
rect 8548 29612 8552 29668
rect 8488 29608 8552 29612
rect 8488 29508 8552 29512
rect 8488 29452 8492 29508
rect 8492 29452 8548 29508
rect 8548 29452 8552 29508
rect 8488 29448 8552 29452
rect 8488 29348 8552 29352
rect 8488 29292 8492 29348
rect 8492 29292 8548 29348
rect 8548 29292 8552 29348
rect 8488 29288 8552 29292
rect 8488 29188 8552 29192
rect 8488 29132 8492 29188
rect 8492 29132 8548 29188
rect 8548 29132 8552 29188
rect 8488 29128 8552 29132
rect 8488 29028 8552 29032
rect 8488 28972 8492 29028
rect 8492 28972 8548 29028
rect 8548 28972 8552 29028
rect 8488 28968 8552 28972
rect 8488 28868 8552 28872
rect 8488 28812 8492 28868
rect 8492 28812 8548 28868
rect 8548 28812 8552 28868
rect 8488 28808 8552 28812
rect 8488 28648 8552 28712
rect 8488 28488 8552 28552
rect 8488 28328 8552 28392
rect 8488 28168 8552 28232
rect 8488 28068 8552 28072
rect 8488 28012 8492 28068
rect 8492 28012 8548 28068
rect 8548 28012 8552 28068
rect 8488 28008 8552 28012
rect 8488 27908 8552 27912
rect 8488 27852 8492 27908
rect 8492 27852 8548 27908
rect 8548 27852 8552 27908
rect 8488 27848 8552 27852
rect 8488 27748 8552 27752
rect 8488 27692 8492 27748
rect 8492 27692 8548 27748
rect 8548 27692 8552 27748
rect 8488 27688 8552 27692
rect 8488 27588 8552 27592
rect 8488 27532 8492 27588
rect 8492 27532 8548 27588
rect 8548 27532 8552 27588
rect 8488 27528 8552 27532
rect 8488 27428 8552 27432
rect 8488 27372 8492 27428
rect 8492 27372 8548 27428
rect 8548 27372 8552 27428
rect 8488 27368 8552 27372
rect 8488 27268 8552 27272
rect 8488 27212 8492 27268
rect 8492 27212 8548 27268
rect 8548 27212 8552 27268
rect 8488 27208 8552 27212
rect 8488 27108 8552 27112
rect 8488 27052 8492 27108
rect 8492 27052 8548 27108
rect 8548 27052 8552 27108
rect 8488 27048 8552 27052
rect 8488 26948 8552 26952
rect 8488 26892 8492 26948
rect 8492 26892 8548 26948
rect 8548 26892 8552 26948
rect 8488 26888 8552 26892
rect 8488 26728 8552 26792
rect 8488 26568 8552 26632
rect 8488 26408 8552 26472
rect 8488 26248 8552 26312
rect 8488 26148 8552 26152
rect 8488 26092 8492 26148
rect 8492 26092 8548 26148
rect 8548 26092 8552 26148
rect 8488 26088 8552 26092
rect 8488 25988 8552 25992
rect 8488 25932 8492 25988
rect 8492 25932 8548 25988
rect 8548 25932 8552 25988
rect 8488 25928 8552 25932
rect 8488 25828 8552 25832
rect 8488 25772 8492 25828
rect 8492 25772 8548 25828
rect 8548 25772 8552 25828
rect 8488 25768 8552 25772
rect 8488 25668 8552 25672
rect 8488 25612 8492 25668
rect 8492 25612 8548 25668
rect 8548 25612 8552 25668
rect 8488 25608 8552 25612
rect 8488 25508 8552 25512
rect 8488 25452 8492 25508
rect 8492 25452 8548 25508
rect 8548 25452 8552 25508
rect 8488 25448 8552 25452
rect 8488 25348 8552 25352
rect 8488 25292 8492 25348
rect 8492 25292 8548 25348
rect 8548 25292 8552 25348
rect 8488 25288 8552 25292
rect 8488 25188 8552 25192
rect 8488 25132 8492 25188
rect 8492 25132 8548 25188
rect 8548 25132 8552 25188
rect 8488 25128 8552 25132
rect 8488 25028 8552 25032
rect 8488 24972 8492 25028
rect 8492 24972 8548 25028
rect 8548 24972 8552 25028
rect 8488 24968 8552 24972
rect 8488 24808 8552 24872
rect 8488 24708 8552 24712
rect 8488 24652 8492 24708
rect 8492 24652 8548 24708
rect 8548 24652 8552 24708
rect 8488 24648 8552 24652
rect 8488 24548 8552 24552
rect 8488 24492 8492 24548
rect 8492 24492 8548 24548
rect 8548 24492 8552 24548
rect 8488 24488 8552 24492
rect 8488 24388 8552 24392
rect 8488 24332 8492 24388
rect 8492 24332 8548 24388
rect 8548 24332 8552 24388
rect 8488 24328 8552 24332
rect 8488 24228 8552 24232
rect 8488 24172 8492 24228
rect 8492 24172 8548 24228
rect 8548 24172 8552 24228
rect 8488 24168 8552 24172
rect 8488 24068 8552 24072
rect 8488 24012 8492 24068
rect 8492 24012 8548 24068
rect 8548 24012 8552 24068
rect 8488 24008 8552 24012
rect 8488 23908 8552 23912
rect 8488 23852 8492 23908
rect 8492 23852 8548 23908
rect 8548 23852 8552 23908
rect 8488 23848 8552 23852
rect 8488 23748 8552 23752
rect 8488 23692 8492 23748
rect 8492 23692 8548 23748
rect 8548 23692 8552 23748
rect 8488 23688 8552 23692
rect 8488 23588 8552 23592
rect 8488 23532 8492 23588
rect 8492 23532 8548 23588
rect 8548 23532 8552 23588
rect 8488 23528 8552 23532
rect 8488 23428 8552 23432
rect 8488 23372 8492 23428
rect 8492 23372 8548 23428
rect 8548 23372 8552 23428
rect 8488 23368 8552 23372
rect 8488 23268 8552 23272
rect 8488 23212 8492 23268
rect 8492 23212 8548 23268
rect 8548 23212 8552 23268
rect 8488 23208 8552 23212
rect 8488 23108 8552 23112
rect 8488 23052 8492 23108
rect 8492 23052 8548 23108
rect 8548 23052 8552 23108
rect 8488 23048 8552 23052
rect 8488 22948 8552 22952
rect 8488 22892 8492 22948
rect 8492 22892 8548 22948
rect 8548 22892 8552 22948
rect 8488 22888 8552 22892
rect 8488 22788 8552 22792
rect 8488 22732 8492 22788
rect 8492 22732 8548 22788
rect 8548 22732 8552 22788
rect 8488 22728 8552 22732
rect 8488 22628 8552 22632
rect 8488 22572 8492 22628
rect 8492 22572 8548 22628
rect 8548 22572 8552 22628
rect 8488 22568 8552 22572
rect 8488 22468 8552 22472
rect 8488 22412 8492 22468
rect 8492 22412 8548 22468
rect 8548 22412 8552 22468
rect 8488 22408 8552 22412
rect 8488 22308 8552 22312
rect 8488 22252 8492 22308
rect 8492 22252 8548 22308
rect 8548 22252 8552 22308
rect 8488 22248 8552 22252
rect 8488 22148 8552 22152
rect 8488 22092 8492 22148
rect 8492 22092 8548 22148
rect 8548 22092 8552 22148
rect 8488 22088 8552 22092
rect 8488 21928 8552 21992
rect 8488 21828 8552 21832
rect 8488 21772 8492 21828
rect 8492 21772 8548 21828
rect 8548 21772 8552 21828
rect 8488 21768 8552 21772
rect 8488 21668 8552 21672
rect 8488 21612 8492 21668
rect 8492 21612 8548 21668
rect 8548 21612 8552 21668
rect 8488 21608 8552 21612
rect 8488 21508 8552 21512
rect 8488 21452 8492 21508
rect 8492 21452 8548 21508
rect 8548 21452 8552 21508
rect 8488 21448 8552 21452
rect 8488 21348 8552 21352
rect 8488 21292 8492 21348
rect 8492 21292 8548 21348
rect 8548 21292 8552 21348
rect 8488 21288 8552 21292
rect 8488 21188 8552 21192
rect 8488 21132 8492 21188
rect 8492 21132 8548 21188
rect 8548 21132 8552 21188
rect 8488 21128 8552 21132
rect 8488 21028 8552 21032
rect 8488 20972 8492 21028
rect 8492 20972 8548 21028
rect 8548 20972 8552 21028
rect 8488 20968 8552 20972
rect 8488 20868 8552 20872
rect 8488 20812 8492 20868
rect 8492 20812 8548 20868
rect 8548 20812 8552 20868
rect 8488 20808 8552 20812
rect 8488 20708 8552 20712
rect 8488 20652 8492 20708
rect 8492 20652 8548 20708
rect 8548 20652 8552 20708
rect 8488 20648 8552 20652
rect 8488 20488 8552 20552
rect 8488 20328 8552 20392
rect 8488 20168 8552 20232
rect 8488 20008 8552 20072
rect 8488 19908 8552 19912
rect 8488 19852 8492 19908
rect 8492 19852 8548 19908
rect 8548 19852 8552 19908
rect 8488 19848 8552 19852
rect 8488 19748 8552 19752
rect 8488 19692 8492 19748
rect 8492 19692 8548 19748
rect 8548 19692 8552 19748
rect 8488 19688 8552 19692
rect 8488 19588 8552 19592
rect 8488 19532 8492 19588
rect 8492 19532 8548 19588
rect 8548 19532 8552 19588
rect 8488 19528 8552 19532
rect 8488 19428 8552 19432
rect 8488 19372 8492 19428
rect 8492 19372 8548 19428
rect 8548 19372 8552 19428
rect 8488 19368 8552 19372
rect 8488 19268 8552 19272
rect 8488 19212 8492 19268
rect 8492 19212 8548 19268
rect 8548 19212 8552 19268
rect 8488 19208 8552 19212
rect 8488 19108 8552 19112
rect 8488 19052 8492 19108
rect 8492 19052 8548 19108
rect 8548 19052 8552 19108
rect 8488 19048 8552 19052
rect 8488 18948 8552 18952
rect 8488 18892 8492 18948
rect 8492 18892 8548 18948
rect 8548 18892 8552 18948
rect 8488 18888 8552 18892
rect 8488 18788 8552 18792
rect 8488 18732 8492 18788
rect 8492 18732 8548 18788
rect 8548 18732 8552 18788
rect 8488 18728 8552 18732
rect 8488 18568 8552 18632
rect 8488 18408 8552 18472
rect 8488 18248 8552 18312
rect 8488 18088 8552 18152
rect 8488 17988 8552 17992
rect 8488 17932 8492 17988
rect 8492 17932 8548 17988
rect 8548 17932 8552 17988
rect 8488 17928 8552 17932
rect 8488 17828 8552 17832
rect 8488 17772 8492 17828
rect 8492 17772 8548 17828
rect 8548 17772 8552 17828
rect 8488 17768 8552 17772
rect 8488 17668 8552 17672
rect 8488 17612 8492 17668
rect 8492 17612 8548 17668
rect 8548 17612 8552 17668
rect 8488 17608 8552 17612
rect 8488 17508 8552 17512
rect 8488 17452 8492 17508
rect 8492 17452 8548 17508
rect 8548 17452 8552 17508
rect 8488 17448 8552 17452
rect 8488 17348 8552 17352
rect 8488 17292 8492 17348
rect 8492 17292 8548 17348
rect 8548 17292 8552 17348
rect 8488 17288 8552 17292
rect 8488 17188 8552 17192
rect 8488 17132 8492 17188
rect 8492 17132 8548 17188
rect 8548 17132 8552 17188
rect 8488 17128 8552 17132
rect 8488 17028 8552 17032
rect 8488 16972 8492 17028
rect 8492 16972 8548 17028
rect 8548 16972 8552 17028
rect 8488 16968 8552 16972
rect 8488 16868 8552 16872
rect 8488 16812 8492 16868
rect 8492 16812 8548 16868
rect 8548 16812 8552 16868
rect 8488 16808 8552 16812
rect 8488 16648 8552 16712
rect 8488 16548 8552 16552
rect 8488 16492 8492 16548
rect 8492 16492 8548 16548
rect 8548 16492 8552 16548
rect 8488 16488 8552 16492
rect 8488 16388 8552 16392
rect 8488 16332 8492 16388
rect 8492 16332 8548 16388
rect 8548 16332 8552 16388
rect 8488 16328 8552 16332
rect 8488 16228 8552 16232
rect 8488 16172 8492 16228
rect 8492 16172 8548 16228
rect 8548 16172 8552 16228
rect 8488 16168 8552 16172
rect 8488 16068 8552 16072
rect 8488 16012 8492 16068
rect 8492 16012 8548 16068
rect 8548 16012 8552 16068
rect 8488 16008 8552 16012
rect 8488 15908 8552 15912
rect 8488 15852 8492 15908
rect 8492 15852 8548 15908
rect 8548 15852 8552 15908
rect 8488 15848 8552 15852
rect 8488 15748 8552 15752
rect 8488 15692 8492 15748
rect 8492 15692 8548 15748
rect 8548 15692 8552 15748
rect 8488 15688 8552 15692
rect 8488 15588 8552 15592
rect 8488 15532 8492 15588
rect 8492 15532 8548 15588
rect 8548 15532 8552 15588
rect 8488 15528 8552 15532
rect 8488 15428 8552 15432
rect 8488 15372 8492 15428
rect 8492 15372 8548 15428
rect 8548 15372 8552 15428
rect 8488 15368 8552 15372
rect 8488 15268 8552 15272
rect 8488 15212 8492 15268
rect 8492 15212 8548 15268
rect 8548 15212 8552 15268
rect 8488 15208 8552 15212
rect 8488 15108 8552 15112
rect 8488 15052 8492 15108
rect 8492 15052 8548 15108
rect 8548 15052 8552 15108
rect 8488 15048 8552 15052
rect 8488 14948 8552 14952
rect 8488 14892 8492 14948
rect 8492 14892 8548 14948
rect 8548 14892 8552 14948
rect 8488 14888 8552 14892
rect 8488 14788 8552 14792
rect 8488 14732 8492 14788
rect 8492 14732 8548 14788
rect 8548 14732 8552 14788
rect 8488 14728 8552 14732
rect 8488 14628 8552 14632
rect 8488 14572 8492 14628
rect 8492 14572 8548 14628
rect 8548 14572 8552 14628
rect 8488 14568 8552 14572
rect 8488 14468 8552 14472
rect 8488 14412 8492 14468
rect 8492 14412 8548 14468
rect 8548 14412 8552 14468
rect 8488 14408 8552 14412
rect 8488 14308 8552 14312
rect 8488 14252 8492 14308
rect 8492 14252 8548 14308
rect 8548 14252 8552 14308
rect 8488 14248 8552 14252
rect 8488 14148 8552 14152
rect 8488 14092 8492 14148
rect 8492 14092 8548 14148
rect 8548 14092 8552 14148
rect 8488 14088 8552 14092
rect 8488 13988 8552 13992
rect 8488 13932 8492 13988
rect 8492 13932 8548 13988
rect 8548 13932 8552 13988
rect 8488 13928 8552 13932
rect 8488 13768 8552 13832
rect 8488 13668 8552 13672
rect 8488 13612 8492 13668
rect 8492 13612 8548 13668
rect 8548 13612 8552 13668
rect 8488 13608 8552 13612
rect 8488 13508 8552 13512
rect 8488 13452 8492 13508
rect 8492 13452 8548 13508
rect 8548 13452 8552 13508
rect 8488 13448 8552 13452
rect 8488 13348 8552 13352
rect 8488 13292 8492 13348
rect 8492 13292 8548 13348
rect 8548 13292 8552 13348
rect 8488 13288 8552 13292
rect 8488 13188 8552 13192
rect 8488 13132 8492 13188
rect 8492 13132 8548 13188
rect 8548 13132 8552 13188
rect 8488 13128 8552 13132
rect 8488 13028 8552 13032
rect 8488 12972 8492 13028
rect 8492 12972 8548 13028
rect 8548 12972 8552 13028
rect 8488 12968 8552 12972
rect 8488 12868 8552 12872
rect 8488 12812 8492 12868
rect 8492 12812 8548 12868
rect 8548 12812 8552 12868
rect 8488 12808 8552 12812
rect 8488 12708 8552 12712
rect 8488 12652 8492 12708
rect 8492 12652 8548 12708
rect 8548 12652 8552 12708
rect 8488 12648 8552 12652
rect 8488 12548 8552 12552
rect 8488 12492 8492 12548
rect 8492 12492 8548 12548
rect 8548 12492 8552 12548
rect 8488 12488 8552 12492
rect 8488 12328 8552 12392
rect 8488 12168 8552 12232
rect 8488 12008 8552 12072
rect 8488 11848 8552 11912
rect 8488 11748 8552 11752
rect 8488 11692 8492 11748
rect 8492 11692 8548 11748
rect 8548 11692 8552 11748
rect 8488 11688 8552 11692
rect 8488 11588 8552 11592
rect 8488 11532 8492 11588
rect 8492 11532 8548 11588
rect 8548 11532 8552 11588
rect 8488 11528 8552 11532
rect 8488 11428 8552 11432
rect 8488 11372 8492 11428
rect 8492 11372 8548 11428
rect 8548 11372 8552 11428
rect 8488 11368 8552 11372
rect 8488 11268 8552 11272
rect 8488 11212 8492 11268
rect 8492 11212 8548 11268
rect 8548 11212 8552 11268
rect 8488 11208 8552 11212
rect 8488 11108 8552 11112
rect 8488 11052 8492 11108
rect 8492 11052 8548 11108
rect 8548 11052 8552 11108
rect 8488 11048 8552 11052
rect 8488 10948 8552 10952
rect 8488 10892 8492 10948
rect 8492 10892 8548 10948
rect 8548 10892 8552 10948
rect 8488 10888 8552 10892
rect 8488 10788 8552 10792
rect 8488 10732 8492 10788
rect 8492 10732 8548 10788
rect 8548 10732 8552 10788
rect 8488 10728 8552 10732
rect 8488 10628 8552 10632
rect 8488 10572 8492 10628
rect 8492 10572 8548 10628
rect 8548 10572 8552 10628
rect 8488 10568 8552 10572
rect 8488 10468 8552 10472
rect 8488 10412 8492 10468
rect 8492 10412 8548 10468
rect 8548 10412 8552 10468
rect 8488 10408 8552 10412
rect 8488 10308 8552 10312
rect 8488 10252 8492 10308
rect 8492 10252 8548 10308
rect 8548 10252 8552 10308
rect 8488 10248 8552 10252
rect 8488 10148 8552 10152
rect 8488 10092 8492 10148
rect 8492 10092 8548 10148
rect 8548 10092 8552 10148
rect 8488 10088 8552 10092
rect 8488 9988 8552 9992
rect 8488 9932 8492 9988
rect 8492 9932 8548 9988
rect 8548 9932 8552 9988
rect 8488 9928 8552 9932
rect 8488 9828 8552 9832
rect 8488 9772 8492 9828
rect 8492 9772 8548 9828
rect 8548 9772 8552 9828
rect 8488 9768 8552 9772
rect 8488 9608 8552 9672
rect 8488 9508 8552 9512
rect 8488 9452 8492 9508
rect 8492 9452 8548 9508
rect 8548 9452 8552 9508
rect 8488 9448 8552 9452
rect 8488 9348 8552 9352
rect 8488 9292 8492 9348
rect 8492 9292 8548 9348
rect 8548 9292 8552 9348
rect 8488 9288 8552 9292
rect 8488 9128 8552 9192
rect 8488 9028 8552 9032
rect 8488 8972 8492 9028
rect 8492 8972 8548 9028
rect 8548 8972 8552 9028
rect 8488 8968 8552 8972
rect 8488 8868 8552 8872
rect 8488 8812 8492 8868
rect 8492 8812 8548 8868
rect 8548 8812 8552 8868
rect 8488 8808 8552 8812
rect 8488 8708 8552 8712
rect 8488 8652 8492 8708
rect 8492 8652 8548 8708
rect 8548 8652 8552 8708
rect 8488 8648 8552 8652
rect 8488 8548 8552 8552
rect 8488 8492 8492 8548
rect 8492 8492 8548 8548
rect 8548 8492 8552 8548
rect 8488 8488 8552 8492
rect 8488 8388 8552 8392
rect 8488 8332 8492 8388
rect 8492 8332 8548 8388
rect 8548 8332 8552 8388
rect 8488 8328 8552 8332
rect 8488 8228 8552 8232
rect 8488 8172 8492 8228
rect 8492 8172 8548 8228
rect 8548 8172 8552 8228
rect 8488 8168 8552 8172
rect 8488 8068 8552 8072
rect 8488 8012 8492 8068
rect 8492 8012 8548 8068
rect 8548 8012 8552 8068
rect 8488 8008 8552 8012
rect 8488 7908 8552 7912
rect 8488 7852 8492 7908
rect 8492 7852 8548 7908
rect 8548 7852 8552 7908
rect 8488 7848 8552 7852
rect 8488 7748 8552 7752
rect 8488 7692 8492 7748
rect 8492 7692 8548 7748
rect 8548 7692 8552 7748
rect 8488 7688 8552 7692
rect 8488 7528 8552 7592
rect 8488 7428 8552 7432
rect 8488 7372 8492 7428
rect 8492 7372 8548 7428
rect 8548 7372 8552 7428
rect 8488 7368 8552 7372
rect 8488 7268 8552 7272
rect 8488 7212 8492 7268
rect 8492 7212 8548 7268
rect 8548 7212 8552 7268
rect 8488 7208 8552 7212
rect 8488 7048 8552 7112
rect 8488 6948 8552 6952
rect 8488 6892 8492 6948
rect 8492 6892 8548 6948
rect 8548 6892 8552 6948
rect 8488 6888 8552 6892
rect 8488 6788 8552 6792
rect 8488 6732 8492 6788
rect 8492 6732 8548 6788
rect 8548 6732 8552 6788
rect 8488 6728 8552 6732
rect 8488 6568 8552 6632
rect 8488 6468 8552 6472
rect 8488 6412 8492 6468
rect 8492 6412 8548 6468
rect 8548 6412 8552 6468
rect 8488 6408 8552 6412
rect 8488 6308 8552 6312
rect 8488 6252 8492 6308
rect 8492 6252 8548 6308
rect 8548 6252 8552 6308
rect 8488 6248 8552 6252
rect 8488 6148 8552 6152
rect 8488 6092 8492 6148
rect 8492 6092 8548 6148
rect 8548 6092 8552 6148
rect 8488 6088 8552 6092
rect 8488 5988 8552 5992
rect 8488 5932 8492 5988
rect 8492 5932 8548 5988
rect 8548 5932 8552 5988
rect 8488 5928 8552 5932
rect 8488 5828 8552 5832
rect 8488 5772 8492 5828
rect 8492 5772 8548 5828
rect 8548 5772 8552 5828
rect 8488 5768 8552 5772
rect 8488 5668 8552 5672
rect 8488 5612 8492 5668
rect 8492 5612 8548 5668
rect 8548 5612 8552 5668
rect 8488 5608 8552 5612
rect 8488 5508 8552 5512
rect 8488 5452 8492 5508
rect 8492 5452 8548 5508
rect 8548 5452 8552 5508
rect 8488 5448 8552 5452
rect 8488 5348 8552 5352
rect 8488 5292 8492 5348
rect 8492 5292 8548 5348
rect 8548 5292 8552 5348
rect 8488 5288 8552 5292
rect 8488 5188 8552 5192
rect 8488 5132 8492 5188
rect 8492 5132 8548 5188
rect 8548 5132 8552 5188
rect 8488 5128 8552 5132
rect 8488 5028 8552 5032
rect 8488 4972 8492 5028
rect 8492 4972 8548 5028
rect 8548 4972 8552 5028
rect 8488 4968 8552 4972
rect 8488 4868 8552 4872
rect 8488 4812 8492 4868
rect 8492 4812 8548 4868
rect 8548 4812 8552 4868
rect 8488 4808 8552 4812
rect 8488 4708 8552 4712
rect 8488 4652 8492 4708
rect 8492 4652 8548 4708
rect 8548 4652 8552 4708
rect 8488 4648 8552 4652
rect 8488 4548 8552 4552
rect 8488 4492 8492 4548
rect 8492 4492 8548 4548
rect 8548 4492 8552 4548
rect 8488 4488 8552 4492
rect 8488 4388 8552 4392
rect 8488 4332 8492 4388
rect 8492 4332 8548 4388
rect 8548 4332 8552 4388
rect 8488 4328 8552 4332
rect 8488 4228 8552 4232
rect 8488 4172 8492 4228
rect 8492 4172 8548 4228
rect 8548 4172 8552 4228
rect 8488 4168 8552 4172
rect 8488 4068 8552 4072
rect 8488 4012 8492 4068
rect 8492 4012 8548 4068
rect 8548 4012 8552 4068
rect 8488 4008 8552 4012
rect 8488 3908 8552 3912
rect 8488 3852 8492 3908
rect 8492 3852 8548 3908
rect 8548 3852 8552 3908
rect 8488 3848 8552 3852
rect 8488 3688 8552 3752
rect 8488 3528 8552 3592
rect 8488 3428 8552 3432
rect 8488 3372 8492 3428
rect 8492 3372 8548 3428
rect 8548 3372 8552 3428
rect 8488 3368 8552 3372
rect 8488 3268 8552 3272
rect 8488 3212 8492 3268
rect 8492 3212 8548 3268
rect 8548 3212 8552 3268
rect 8488 3208 8552 3212
rect 8488 3108 8552 3112
rect 8488 3052 8492 3108
rect 8492 3052 8548 3108
rect 8548 3052 8552 3108
rect 8488 3048 8552 3052
rect 8488 2948 8552 2952
rect 8488 2892 8492 2948
rect 8492 2892 8548 2948
rect 8548 2892 8552 2948
rect 8488 2888 8552 2892
rect 8488 2788 8552 2792
rect 8488 2732 8492 2788
rect 8492 2732 8548 2788
rect 8548 2732 8552 2788
rect 8488 2728 8552 2732
rect 8488 2628 8552 2632
rect 8488 2572 8492 2628
rect 8492 2572 8548 2628
rect 8548 2572 8552 2628
rect 8488 2568 8552 2572
rect 8488 2468 8552 2472
rect 8488 2412 8492 2468
rect 8492 2412 8548 2468
rect 8548 2412 8552 2468
rect 8488 2408 8552 2412
rect 8488 2308 8552 2312
rect 8488 2252 8492 2308
rect 8492 2252 8548 2308
rect 8548 2252 8552 2308
rect 8488 2248 8552 2252
rect 8488 2148 8552 2152
rect 8488 2092 8492 2148
rect 8492 2092 8548 2148
rect 8548 2092 8552 2148
rect 8488 2088 8552 2092
rect 8488 1988 8552 1992
rect 8488 1932 8492 1988
rect 8492 1932 8548 1988
rect 8548 1932 8552 1988
rect 8488 1928 8552 1932
rect 8488 1768 8552 1832
rect 8488 1668 8552 1672
rect 8488 1612 8492 1668
rect 8492 1612 8548 1668
rect 8548 1612 8552 1668
rect 8488 1608 8552 1612
rect 8488 1508 8552 1512
rect 8488 1452 8492 1508
rect 8492 1452 8548 1508
rect 8548 1452 8552 1508
rect 8488 1448 8552 1452
rect 8488 1348 8552 1352
rect 8488 1292 8492 1348
rect 8492 1292 8548 1348
rect 8548 1292 8552 1348
rect 8488 1288 8552 1292
rect 8488 1188 8552 1192
rect 8488 1132 8492 1188
rect 8492 1132 8548 1188
rect 8548 1132 8552 1188
rect 8488 1128 8552 1132
rect 8488 1028 8552 1032
rect 8488 972 8492 1028
rect 8492 972 8548 1028
rect 8548 972 8552 1028
rect 8488 968 8552 972
rect 8488 808 8552 872
rect 8488 648 8552 712
rect 8488 548 8552 552
rect 8488 492 8492 548
rect 8492 492 8548 548
rect 8548 492 8552 548
rect 8488 488 8552 492
rect 8488 388 8552 392
rect 8488 332 8492 388
rect 8492 332 8548 388
rect 8548 332 8552 388
rect 8488 328 8552 332
rect 8488 228 8552 232
rect 8488 172 8492 228
rect 8492 172 8548 228
rect 8548 172 8552 228
rect 8488 168 8552 172
rect 8488 68 8552 72
rect 8488 12 8492 68
rect 8492 12 8548 68
rect 8548 12 8552 68
rect 8488 8 8552 12
rect 8808 31428 8872 31432
rect 8808 31372 8812 31428
rect 8812 31372 8868 31428
rect 8868 31372 8872 31428
rect 8808 31368 8872 31372
rect 8808 31268 8872 31272
rect 8808 31212 8812 31268
rect 8812 31212 8868 31268
rect 8868 31212 8872 31268
rect 8808 31208 8872 31212
rect 8808 31108 8872 31112
rect 8808 31052 8812 31108
rect 8812 31052 8868 31108
rect 8868 31052 8872 31108
rect 8808 31048 8872 31052
rect 8808 30948 8872 30952
rect 8808 30892 8812 30948
rect 8812 30892 8868 30948
rect 8868 30892 8872 30948
rect 8808 30888 8872 30892
rect 8808 30788 8872 30792
rect 8808 30732 8812 30788
rect 8812 30732 8868 30788
rect 8868 30732 8872 30788
rect 8808 30728 8872 30732
rect 8808 30628 8872 30632
rect 8808 30572 8812 30628
rect 8812 30572 8868 30628
rect 8868 30572 8872 30628
rect 8808 30568 8872 30572
rect 8808 30468 8872 30472
rect 8808 30412 8812 30468
rect 8812 30412 8868 30468
rect 8868 30412 8872 30468
rect 8808 30408 8872 30412
rect 8808 30308 8872 30312
rect 8808 30252 8812 30308
rect 8812 30252 8868 30308
rect 8868 30252 8872 30308
rect 8808 30248 8872 30252
rect 8808 30088 8872 30152
rect 8808 29988 8872 29992
rect 8808 29932 8812 29988
rect 8812 29932 8868 29988
rect 8868 29932 8872 29988
rect 8808 29928 8872 29932
rect 8808 29828 8872 29832
rect 8808 29772 8812 29828
rect 8812 29772 8868 29828
rect 8868 29772 8872 29828
rect 8808 29768 8872 29772
rect 8808 29668 8872 29672
rect 8808 29612 8812 29668
rect 8812 29612 8868 29668
rect 8868 29612 8872 29668
rect 8808 29608 8872 29612
rect 8808 29508 8872 29512
rect 8808 29452 8812 29508
rect 8812 29452 8868 29508
rect 8868 29452 8872 29508
rect 8808 29448 8872 29452
rect 8808 29348 8872 29352
rect 8808 29292 8812 29348
rect 8812 29292 8868 29348
rect 8868 29292 8872 29348
rect 8808 29288 8872 29292
rect 8808 29188 8872 29192
rect 8808 29132 8812 29188
rect 8812 29132 8868 29188
rect 8868 29132 8872 29188
rect 8808 29128 8872 29132
rect 8808 29028 8872 29032
rect 8808 28972 8812 29028
rect 8812 28972 8868 29028
rect 8868 28972 8872 29028
rect 8808 28968 8872 28972
rect 8808 28868 8872 28872
rect 8808 28812 8812 28868
rect 8812 28812 8868 28868
rect 8868 28812 8872 28868
rect 8808 28808 8872 28812
rect 8808 28648 8872 28712
rect 8808 28488 8872 28552
rect 8808 28328 8872 28392
rect 8808 28168 8872 28232
rect 8808 28068 8872 28072
rect 8808 28012 8812 28068
rect 8812 28012 8868 28068
rect 8868 28012 8872 28068
rect 8808 28008 8872 28012
rect 8808 27908 8872 27912
rect 8808 27852 8812 27908
rect 8812 27852 8868 27908
rect 8868 27852 8872 27908
rect 8808 27848 8872 27852
rect 8808 27748 8872 27752
rect 8808 27692 8812 27748
rect 8812 27692 8868 27748
rect 8868 27692 8872 27748
rect 8808 27688 8872 27692
rect 8808 27588 8872 27592
rect 8808 27532 8812 27588
rect 8812 27532 8868 27588
rect 8868 27532 8872 27588
rect 8808 27528 8872 27532
rect 8808 27428 8872 27432
rect 8808 27372 8812 27428
rect 8812 27372 8868 27428
rect 8868 27372 8872 27428
rect 8808 27368 8872 27372
rect 8808 27268 8872 27272
rect 8808 27212 8812 27268
rect 8812 27212 8868 27268
rect 8868 27212 8872 27268
rect 8808 27208 8872 27212
rect 8808 27108 8872 27112
rect 8808 27052 8812 27108
rect 8812 27052 8868 27108
rect 8868 27052 8872 27108
rect 8808 27048 8872 27052
rect 8808 26948 8872 26952
rect 8808 26892 8812 26948
rect 8812 26892 8868 26948
rect 8868 26892 8872 26948
rect 8808 26888 8872 26892
rect 8808 26728 8872 26792
rect 8808 26568 8872 26632
rect 8808 26408 8872 26472
rect 8808 26248 8872 26312
rect 8808 26148 8872 26152
rect 8808 26092 8812 26148
rect 8812 26092 8868 26148
rect 8868 26092 8872 26148
rect 8808 26088 8872 26092
rect 8808 25988 8872 25992
rect 8808 25932 8812 25988
rect 8812 25932 8868 25988
rect 8868 25932 8872 25988
rect 8808 25928 8872 25932
rect 8808 25828 8872 25832
rect 8808 25772 8812 25828
rect 8812 25772 8868 25828
rect 8868 25772 8872 25828
rect 8808 25768 8872 25772
rect 8808 25668 8872 25672
rect 8808 25612 8812 25668
rect 8812 25612 8868 25668
rect 8868 25612 8872 25668
rect 8808 25608 8872 25612
rect 8808 25508 8872 25512
rect 8808 25452 8812 25508
rect 8812 25452 8868 25508
rect 8868 25452 8872 25508
rect 8808 25448 8872 25452
rect 8808 25348 8872 25352
rect 8808 25292 8812 25348
rect 8812 25292 8868 25348
rect 8868 25292 8872 25348
rect 8808 25288 8872 25292
rect 8808 25188 8872 25192
rect 8808 25132 8812 25188
rect 8812 25132 8868 25188
rect 8868 25132 8872 25188
rect 8808 25128 8872 25132
rect 8808 25028 8872 25032
rect 8808 24972 8812 25028
rect 8812 24972 8868 25028
rect 8868 24972 8872 25028
rect 8808 24968 8872 24972
rect 8808 24808 8872 24872
rect 8808 24708 8872 24712
rect 8808 24652 8812 24708
rect 8812 24652 8868 24708
rect 8868 24652 8872 24708
rect 8808 24648 8872 24652
rect 8808 24548 8872 24552
rect 8808 24492 8812 24548
rect 8812 24492 8868 24548
rect 8868 24492 8872 24548
rect 8808 24488 8872 24492
rect 8808 24388 8872 24392
rect 8808 24332 8812 24388
rect 8812 24332 8868 24388
rect 8868 24332 8872 24388
rect 8808 24328 8872 24332
rect 8808 24228 8872 24232
rect 8808 24172 8812 24228
rect 8812 24172 8868 24228
rect 8868 24172 8872 24228
rect 8808 24168 8872 24172
rect 8808 24068 8872 24072
rect 8808 24012 8812 24068
rect 8812 24012 8868 24068
rect 8868 24012 8872 24068
rect 8808 24008 8872 24012
rect 8808 23908 8872 23912
rect 8808 23852 8812 23908
rect 8812 23852 8868 23908
rect 8868 23852 8872 23908
rect 8808 23848 8872 23852
rect 8808 23748 8872 23752
rect 8808 23692 8812 23748
rect 8812 23692 8868 23748
rect 8868 23692 8872 23748
rect 8808 23688 8872 23692
rect 8808 23588 8872 23592
rect 8808 23532 8812 23588
rect 8812 23532 8868 23588
rect 8868 23532 8872 23588
rect 8808 23528 8872 23532
rect 8808 23428 8872 23432
rect 8808 23372 8812 23428
rect 8812 23372 8868 23428
rect 8868 23372 8872 23428
rect 8808 23368 8872 23372
rect 8808 23268 8872 23272
rect 8808 23212 8812 23268
rect 8812 23212 8868 23268
rect 8868 23212 8872 23268
rect 8808 23208 8872 23212
rect 8808 23108 8872 23112
rect 8808 23052 8812 23108
rect 8812 23052 8868 23108
rect 8868 23052 8872 23108
rect 8808 23048 8872 23052
rect 8808 22948 8872 22952
rect 8808 22892 8812 22948
rect 8812 22892 8868 22948
rect 8868 22892 8872 22948
rect 8808 22888 8872 22892
rect 8808 22788 8872 22792
rect 8808 22732 8812 22788
rect 8812 22732 8868 22788
rect 8868 22732 8872 22788
rect 8808 22728 8872 22732
rect 8808 22628 8872 22632
rect 8808 22572 8812 22628
rect 8812 22572 8868 22628
rect 8868 22572 8872 22628
rect 8808 22568 8872 22572
rect 8808 22468 8872 22472
rect 8808 22412 8812 22468
rect 8812 22412 8868 22468
rect 8868 22412 8872 22468
rect 8808 22408 8872 22412
rect 8808 22308 8872 22312
rect 8808 22252 8812 22308
rect 8812 22252 8868 22308
rect 8868 22252 8872 22308
rect 8808 22248 8872 22252
rect 8808 22148 8872 22152
rect 8808 22092 8812 22148
rect 8812 22092 8868 22148
rect 8868 22092 8872 22148
rect 8808 22088 8872 22092
rect 8808 21928 8872 21992
rect 8808 21828 8872 21832
rect 8808 21772 8812 21828
rect 8812 21772 8868 21828
rect 8868 21772 8872 21828
rect 8808 21768 8872 21772
rect 8808 21668 8872 21672
rect 8808 21612 8812 21668
rect 8812 21612 8868 21668
rect 8868 21612 8872 21668
rect 8808 21608 8872 21612
rect 8808 21508 8872 21512
rect 8808 21452 8812 21508
rect 8812 21452 8868 21508
rect 8868 21452 8872 21508
rect 8808 21448 8872 21452
rect 8808 21348 8872 21352
rect 8808 21292 8812 21348
rect 8812 21292 8868 21348
rect 8868 21292 8872 21348
rect 8808 21288 8872 21292
rect 8808 21188 8872 21192
rect 8808 21132 8812 21188
rect 8812 21132 8868 21188
rect 8868 21132 8872 21188
rect 8808 21128 8872 21132
rect 8808 21028 8872 21032
rect 8808 20972 8812 21028
rect 8812 20972 8868 21028
rect 8868 20972 8872 21028
rect 8808 20968 8872 20972
rect 8808 20868 8872 20872
rect 8808 20812 8812 20868
rect 8812 20812 8868 20868
rect 8868 20812 8872 20868
rect 8808 20808 8872 20812
rect 8808 20708 8872 20712
rect 8808 20652 8812 20708
rect 8812 20652 8868 20708
rect 8868 20652 8872 20708
rect 8808 20648 8872 20652
rect 8808 20488 8872 20552
rect 8808 20328 8872 20392
rect 8808 20168 8872 20232
rect 8808 20008 8872 20072
rect 8808 19908 8872 19912
rect 8808 19852 8812 19908
rect 8812 19852 8868 19908
rect 8868 19852 8872 19908
rect 8808 19848 8872 19852
rect 8808 19748 8872 19752
rect 8808 19692 8812 19748
rect 8812 19692 8868 19748
rect 8868 19692 8872 19748
rect 8808 19688 8872 19692
rect 8808 19588 8872 19592
rect 8808 19532 8812 19588
rect 8812 19532 8868 19588
rect 8868 19532 8872 19588
rect 8808 19528 8872 19532
rect 8808 19428 8872 19432
rect 8808 19372 8812 19428
rect 8812 19372 8868 19428
rect 8868 19372 8872 19428
rect 8808 19368 8872 19372
rect 8808 19268 8872 19272
rect 8808 19212 8812 19268
rect 8812 19212 8868 19268
rect 8868 19212 8872 19268
rect 8808 19208 8872 19212
rect 8808 19108 8872 19112
rect 8808 19052 8812 19108
rect 8812 19052 8868 19108
rect 8868 19052 8872 19108
rect 8808 19048 8872 19052
rect 8808 18948 8872 18952
rect 8808 18892 8812 18948
rect 8812 18892 8868 18948
rect 8868 18892 8872 18948
rect 8808 18888 8872 18892
rect 8808 18788 8872 18792
rect 8808 18732 8812 18788
rect 8812 18732 8868 18788
rect 8868 18732 8872 18788
rect 8808 18728 8872 18732
rect 8808 18568 8872 18632
rect 8808 18408 8872 18472
rect 8808 18248 8872 18312
rect 8808 18088 8872 18152
rect 8808 17988 8872 17992
rect 8808 17932 8812 17988
rect 8812 17932 8868 17988
rect 8868 17932 8872 17988
rect 8808 17928 8872 17932
rect 8808 17828 8872 17832
rect 8808 17772 8812 17828
rect 8812 17772 8868 17828
rect 8868 17772 8872 17828
rect 8808 17768 8872 17772
rect 8808 17668 8872 17672
rect 8808 17612 8812 17668
rect 8812 17612 8868 17668
rect 8868 17612 8872 17668
rect 8808 17608 8872 17612
rect 8808 17508 8872 17512
rect 8808 17452 8812 17508
rect 8812 17452 8868 17508
rect 8868 17452 8872 17508
rect 8808 17448 8872 17452
rect 8808 17348 8872 17352
rect 8808 17292 8812 17348
rect 8812 17292 8868 17348
rect 8868 17292 8872 17348
rect 8808 17288 8872 17292
rect 8808 17188 8872 17192
rect 8808 17132 8812 17188
rect 8812 17132 8868 17188
rect 8868 17132 8872 17188
rect 8808 17128 8872 17132
rect 8808 17028 8872 17032
rect 8808 16972 8812 17028
rect 8812 16972 8868 17028
rect 8868 16972 8872 17028
rect 8808 16968 8872 16972
rect 8808 16868 8872 16872
rect 8808 16812 8812 16868
rect 8812 16812 8868 16868
rect 8868 16812 8872 16868
rect 8808 16808 8872 16812
rect 8808 16648 8872 16712
rect 8808 16548 8872 16552
rect 8808 16492 8812 16548
rect 8812 16492 8868 16548
rect 8868 16492 8872 16548
rect 8808 16488 8872 16492
rect 8808 16388 8872 16392
rect 8808 16332 8812 16388
rect 8812 16332 8868 16388
rect 8868 16332 8872 16388
rect 8808 16328 8872 16332
rect 8808 16228 8872 16232
rect 8808 16172 8812 16228
rect 8812 16172 8868 16228
rect 8868 16172 8872 16228
rect 8808 16168 8872 16172
rect 8808 16068 8872 16072
rect 8808 16012 8812 16068
rect 8812 16012 8868 16068
rect 8868 16012 8872 16068
rect 8808 16008 8872 16012
rect 8808 15908 8872 15912
rect 8808 15852 8812 15908
rect 8812 15852 8868 15908
rect 8868 15852 8872 15908
rect 8808 15848 8872 15852
rect 8808 15748 8872 15752
rect 8808 15692 8812 15748
rect 8812 15692 8868 15748
rect 8868 15692 8872 15748
rect 8808 15688 8872 15692
rect 8808 15588 8872 15592
rect 8808 15532 8812 15588
rect 8812 15532 8868 15588
rect 8868 15532 8872 15588
rect 8808 15528 8872 15532
rect 8808 15428 8872 15432
rect 8808 15372 8812 15428
rect 8812 15372 8868 15428
rect 8868 15372 8872 15428
rect 8808 15368 8872 15372
rect 8808 15268 8872 15272
rect 8808 15212 8812 15268
rect 8812 15212 8868 15268
rect 8868 15212 8872 15268
rect 8808 15208 8872 15212
rect 8808 15108 8872 15112
rect 8808 15052 8812 15108
rect 8812 15052 8868 15108
rect 8868 15052 8872 15108
rect 8808 15048 8872 15052
rect 8808 14948 8872 14952
rect 8808 14892 8812 14948
rect 8812 14892 8868 14948
rect 8868 14892 8872 14948
rect 8808 14888 8872 14892
rect 8808 14788 8872 14792
rect 8808 14732 8812 14788
rect 8812 14732 8868 14788
rect 8868 14732 8872 14788
rect 8808 14728 8872 14732
rect 8808 14628 8872 14632
rect 8808 14572 8812 14628
rect 8812 14572 8868 14628
rect 8868 14572 8872 14628
rect 8808 14568 8872 14572
rect 8808 14468 8872 14472
rect 8808 14412 8812 14468
rect 8812 14412 8868 14468
rect 8868 14412 8872 14468
rect 8808 14408 8872 14412
rect 8808 14308 8872 14312
rect 8808 14252 8812 14308
rect 8812 14252 8868 14308
rect 8868 14252 8872 14308
rect 8808 14248 8872 14252
rect 8808 14148 8872 14152
rect 8808 14092 8812 14148
rect 8812 14092 8868 14148
rect 8868 14092 8872 14148
rect 8808 14088 8872 14092
rect 8808 13988 8872 13992
rect 8808 13932 8812 13988
rect 8812 13932 8868 13988
rect 8868 13932 8872 13988
rect 8808 13928 8872 13932
rect 8808 13768 8872 13832
rect 8808 13668 8872 13672
rect 8808 13612 8812 13668
rect 8812 13612 8868 13668
rect 8868 13612 8872 13668
rect 8808 13608 8872 13612
rect 8808 13508 8872 13512
rect 8808 13452 8812 13508
rect 8812 13452 8868 13508
rect 8868 13452 8872 13508
rect 8808 13448 8872 13452
rect 8808 13348 8872 13352
rect 8808 13292 8812 13348
rect 8812 13292 8868 13348
rect 8868 13292 8872 13348
rect 8808 13288 8872 13292
rect 8808 13188 8872 13192
rect 8808 13132 8812 13188
rect 8812 13132 8868 13188
rect 8868 13132 8872 13188
rect 8808 13128 8872 13132
rect 8808 13028 8872 13032
rect 8808 12972 8812 13028
rect 8812 12972 8868 13028
rect 8868 12972 8872 13028
rect 8808 12968 8872 12972
rect 8808 12868 8872 12872
rect 8808 12812 8812 12868
rect 8812 12812 8868 12868
rect 8868 12812 8872 12868
rect 8808 12808 8872 12812
rect 8808 12708 8872 12712
rect 8808 12652 8812 12708
rect 8812 12652 8868 12708
rect 8868 12652 8872 12708
rect 8808 12648 8872 12652
rect 8808 12548 8872 12552
rect 8808 12492 8812 12548
rect 8812 12492 8868 12548
rect 8868 12492 8872 12548
rect 8808 12488 8872 12492
rect 8808 12328 8872 12392
rect 8808 12168 8872 12232
rect 8808 12008 8872 12072
rect 8808 11848 8872 11912
rect 8808 11748 8872 11752
rect 8808 11692 8812 11748
rect 8812 11692 8868 11748
rect 8868 11692 8872 11748
rect 8808 11688 8872 11692
rect 8808 11588 8872 11592
rect 8808 11532 8812 11588
rect 8812 11532 8868 11588
rect 8868 11532 8872 11588
rect 8808 11528 8872 11532
rect 8808 11428 8872 11432
rect 8808 11372 8812 11428
rect 8812 11372 8868 11428
rect 8868 11372 8872 11428
rect 8808 11368 8872 11372
rect 8808 11268 8872 11272
rect 8808 11212 8812 11268
rect 8812 11212 8868 11268
rect 8868 11212 8872 11268
rect 8808 11208 8872 11212
rect 8808 11108 8872 11112
rect 8808 11052 8812 11108
rect 8812 11052 8868 11108
rect 8868 11052 8872 11108
rect 8808 11048 8872 11052
rect 8808 10948 8872 10952
rect 8808 10892 8812 10948
rect 8812 10892 8868 10948
rect 8868 10892 8872 10948
rect 8808 10888 8872 10892
rect 8808 10788 8872 10792
rect 8808 10732 8812 10788
rect 8812 10732 8868 10788
rect 8868 10732 8872 10788
rect 8808 10728 8872 10732
rect 8808 10628 8872 10632
rect 8808 10572 8812 10628
rect 8812 10572 8868 10628
rect 8868 10572 8872 10628
rect 8808 10568 8872 10572
rect 8808 10468 8872 10472
rect 8808 10412 8812 10468
rect 8812 10412 8868 10468
rect 8868 10412 8872 10468
rect 8808 10408 8872 10412
rect 8808 10308 8872 10312
rect 8808 10252 8812 10308
rect 8812 10252 8868 10308
rect 8868 10252 8872 10308
rect 8808 10248 8872 10252
rect 8808 10148 8872 10152
rect 8808 10092 8812 10148
rect 8812 10092 8868 10148
rect 8868 10092 8872 10148
rect 8808 10088 8872 10092
rect 8808 9988 8872 9992
rect 8808 9932 8812 9988
rect 8812 9932 8868 9988
rect 8868 9932 8872 9988
rect 8808 9928 8872 9932
rect 8808 9828 8872 9832
rect 8808 9772 8812 9828
rect 8812 9772 8868 9828
rect 8868 9772 8872 9828
rect 8808 9768 8872 9772
rect 8808 9608 8872 9672
rect 8808 9508 8872 9512
rect 8808 9452 8812 9508
rect 8812 9452 8868 9508
rect 8868 9452 8872 9508
rect 8808 9448 8872 9452
rect 8808 9348 8872 9352
rect 8808 9292 8812 9348
rect 8812 9292 8868 9348
rect 8868 9292 8872 9348
rect 8808 9288 8872 9292
rect 8808 9128 8872 9192
rect 8808 9028 8872 9032
rect 8808 8972 8812 9028
rect 8812 8972 8868 9028
rect 8868 8972 8872 9028
rect 8808 8968 8872 8972
rect 8808 8868 8872 8872
rect 8808 8812 8812 8868
rect 8812 8812 8868 8868
rect 8868 8812 8872 8868
rect 8808 8808 8872 8812
rect 8808 8708 8872 8712
rect 8808 8652 8812 8708
rect 8812 8652 8868 8708
rect 8868 8652 8872 8708
rect 8808 8648 8872 8652
rect 8808 8548 8872 8552
rect 8808 8492 8812 8548
rect 8812 8492 8868 8548
rect 8868 8492 8872 8548
rect 8808 8488 8872 8492
rect 8808 8388 8872 8392
rect 8808 8332 8812 8388
rect 8812 8332 8868 8388
rect 8868 8332 8872 8388
rect 8808 8328 8872 8332
rect 8808 8228 8872 8232
rect 8808 8172 8812 8228
rect 8812 8172 8868 8228
rect 8868 8172 8872 8228
rect 8808 8168 8872 8172
rect 8808 8068 8872 8072
rect 8808 8012 8812 8068
rect 8812 8012 8868 8068
rect 8868 8012 8872 8068
rect 8808 8008 8872 8012
rect 8808 7908 8872 7912
rect 8808 7852 8812 7908
rect 8812 7852 8868 7908
rect 8868 7852 8872 7908
rect 8808 7848 8872 7852
rect 8808 7748 8872 7752
rect 8808 7692 8812 7748
rect 8812 7692 8868 7748
rect 8868 7692 8872 7748
rect 8808 7688 8872 7692
rect 8808 7528 8872 7592
rect 8808 7428 8872 7432
rect 8808 7372 8812 7428
rect 8812 7372 8868 7428
rect 8868 7372 8872 7428
rect 8808 7368 8872 7372
rect 8808 7268 8872 7272
rect 8808 7212 8812 7268
rect 8812 7212 8868 7268
rect 8868 7212 8872 7268
rect 8808 7208 8872 7212
rect 8808 7048 8872 7112
rect 8808 6948 8872 6952
rect 8808 6892 8812 6948
rect 8812 6892 8868 6948
rect 8868 6892 8872 6948
rect 8808 6888 8872 6892
rect 8808 6788 8872 6792
rect 8808 6732 8812 6788
rect 8812 6732 8868 6788
rect 8868 6732 8872 6788
rect 8808 6728 8872 6732
rect 8808 6568 8872 6632
rect 8808 6468 8872 6472
rect 8808 6412 8812 6468
rect 8812 6412 8868 6468
rect 8868 6412 8872 6468
rect 8808 6408 8872 6412
rect 8808 6308 8872 6312
rect 8808 6252 8812 6308
rect 8812 6252 8868 6308
rect 8868 6252 8872 6308
rect 8808 6248 8872 6252
rect 8808 6148 8872 6152
rect 8808 6092 8812 6148
rect 8812 6092 8868 6148
rect 8868 6092 8872 6148
rect 8808 6088 8872 6092
rect 8808 5988 8872 5992
rect 8808 5932 8812 5988
rect 8812 5932 8868 5988
rect 8868 5932 8872 5988
rect 8808 5928 8872 5932
rect 8808 5828 8872 5832
rect 8808 5772 8812 5828
rect 8812 5772 8868 5828
rect 8868 5772 8872 5828
rect 8808 5768 8872 5772
rect 8808 5668 8872 5672
rect 8808 5612 8812 5668
rect 8812 5612 8868 5668
rect 8868 5612 8872 5668
rect 8808 5608 8872 5612
rect 8808 5508 8872 5512
rect 8808 5452 8812 5508
rect 8812 5452 8868 5508
rect 8868 5452 8872 5508
rect 8808 5448 8872 5452
rect 8808 5348 8872 5352
rect 8808 5292 8812 5348
rect 8812 5292 8868 5348
rect 8868 5292 8872 5348
rect 8808 5288 8872 5292
rect 8808 5188 8872 5192
rect 8808 5132 8812 5188
rect 8812 5132 8868 5188
rect 8868 5132 8872 5188
rect 8808 5128 8872 5132
rect 8808 5028 8872 5032
rect 8808 4972 8812 5028
rect 8812 4972 8868 5028
rect 8868 4972 8872 5028
rect 8808 4968 8872 4972
rect 8808 4868 8872 4872
rect 8808 4812 8812 4868
rect 8812 4812 8868 4868
rect 8868 4812 8872 4868
rect 8808 4808 8872 4812
rect 8808 4708 8872 4712
rect 8808 4652 8812 4708
rect 8812 4652 8868 4708
rect 8868 4652 8872 4708
rect 8808 4648 8872 4652
rect 8808 4548 8872 4552
rect 8808 4492 8812 4548
rect 8812 4492 8868 4548
rect 8868 4492 8872 4548
rect 8808 4488 8872 4492
rect 8808 4388 8872 4392
rect 8808 4332 8812 4388
rect 8812 4332 8868 4388
rect 8868 4332 8872 4388
rect 8808 4328 8872 4332
rect 8808 4228 8872 4232
rect 8808 4172 8812 4228
rect 8812 4172 8868 4228
rect 8868 4172 8872 4228
rect 8808 4168 8872 4172
rect 8808 4068 8872 4072
rect 8808 4012 8812 4068
rect 8812 4012 8868 4068
rect 8868 4012 8872 4068
rect 8808 4008 8872 4012
rect 8808 3908 8872 3912
rect 8808 3852 8812 3908
rect 8812 3852 8868 3908
rect 8868 3852 8872 3908
rect 8808 3848 8872 3852
rect 8808 3688 8872 3752
rect 8808 3528 8872 3592
rect 8808 3428 8872 3432
rect 8808 3372 8812 3428
rect 8812 3372 8868 3428
rect 8868 3372 8872 3428
rect 8808 3368 8872 3372
rect 8808 3268 8872 3272
rect 8808 3212 8812 3268
rect 8812 3212 8868 3268
rect 8868 3212 8872 3268
rect 8808 3208 8872 3212
rect 8808 3108 8872 3112
rect 8808 3052 8812 3108
rect 8812 3052 8868 3108
rect 8868 3052 8872 3108
rect 8808 3048 8872 3052
rect 8808 2948 8872 2952
rect 8808 2892 8812 2948
rect 8812 2892 8868 2948
rect 8868 2892 8872 2948
rect 8808 2888 8872 2892
rect 8808 2788 8872 2792
rect 8808 2732 8812 2788
rect 8812 2732 8868 2788
rect 8868 2732 8872 2788
rect 8808 2728 8872 2732
rect 8808 2628 8872 2632
rect 8808 2572 8812 2628
rect 8812 2572 8868 2628
rect 8868 2572 8872 2628
rect 8808 2568 8872 2572
rect 8808 2468 8872 2472
rect 8808 2412 8812 2468
rect 8812 2412 8868 2468
rect 8868 2412 8872 2468
rect 8808 2408 8872 2412
rect 8808 2308 8872 2312
rect 8808 2252 8812 2308
rect 8812 2252 8868 2308
rect 8868 2252 8872 2308
rect 8808 2248 8872 2252
rect 8808 2148 8872 2152
rect 8808 2092 8812 2148
rect 8812 2092 8868 2148
rect 8868 2092 8872 2148
rect 8808 2088 8872 2092
rect 8808 1988 8872 1992
rect 8808 1932 8812 1988
rect 8812 1932 8868 1988
rect 8868 1932 8872 1988
rect 8808 1928 8872 1932
rect 8808 1768 8872 1832
rect 8808 1668 8872 1672
rect 8808 1612 8812 1668
rect 8812 1612 8868 1668
rect 8868 1612 8872 1668
rect 8808 1608 8872 1612
rect 8808 1508 8872 1512
rect 8808 1452 8812 1508
rect 8812 1452 8868 1508
rect 8868 1452 8872 1508
rect 8808 1448 8872 1452
rect 8808 1348 8872 1352
rect 8808 1292 8812 1348
rect 8812 1292 8868 1348
rect 8868 1292 8872 1348
rect 8808 1288 8872 1292
rect 8808 1188 8872 1192
rect 8808 1132 8812 1188
rect 8812 1132 8868 1188
rect 8868 1132 8872 1188
rect 8808 1128 8872 1132
rect 8808 1028 8872 1032
rect 8808 972 8812 1028
rect 8812 972 8868 1028
rect 8868 972 8872 1028
rect 8808 968 8872 972
rect 8808 808 8872 872
rect 8808 648 8872 712
rect 8808 548 8872 552
rect 8808 492 8812 548
rect 8812 492 8868 548
rect 8868 492 8872 548
rect 8808 488 8872 492
rect 8808 388 8872 392
rect 8808 332 8812 388
rect 8812 332 8868 388
rect 8868 332 8872 388
rect 8808 328 8872 332
rect 8808 228 8872 232
rect 8808 172 8812 228
rect 8812 172 8868 228
rect 8868 172 8872 228
rect 8808 168 8872 172
rect 8808 68 8872 72
rect 8808 12 8812 68
rect 8812 12 8868 68
rect 8868 12 8872 68
rect 8808 8 8872 12
rect 8488 -1592 8552 -1528
rect 8488 -1672 8552 -1608
rect 8488 -1752 8552 -1688
rect 8488 -1832 8552 -1768
rect 8488 -1912 8552 -1848
rect 8808 -1592 8872 -1528
rect 8808 -1672 8872 -1608
rect 8808 -1752 8872 -1688
rect 8808 -1832 8872 -1768
rect 8808 -1912 8872 -1848
rect 8968 31428 9032 31432
rect 8968 31372 8972 31428
rect 8972 31372 9028 31428
rect 9028 31372 9032 31428
rect 8968 31368 9032 31372
rect 8968 31268 9032 31272
rect 8968 31212 8972 31268
rect 8972 31212 9028 31268
rect 9028 31212 9032 31268
rect 8968 31208 9032 31212
rect 8968 31108 9032 31112
rect 8968 31052 8972 31108
rect 8972 31052 9028 31108
rect 9028 31052 9032 31108
rect 8968 31048 9032 31052
rect 8968 30948 9032 30952
rect 8968 30892 8972 30948
rect 8972 30892 9028 30948
rect 9028 30892 9032 30948
rect 8968 30888 9032 30892
rect 8968 30788 9032 30792
rect 8968 30732 8972 30788
rect 8972 30732 9028 30788
rect 9028 30732 9032 30788
rect 8968 30728 9032 30732
rect 8968 30628 9032 30632
rect 8968 30572 8972 30628
rect 8972 30572 9028 30628
rect 9028 30572 9032 30628
rect 8968 30568 9032 30572
rect 8968 30468 9032 30472
rect 8968 30412 8972 30468
rect 8972 30412 9028 30468
rect 9028 30412 9032 30468
rect 8968 30408 9032 30412
rect 8968 30308 9032 30312
rect 8968 30252 8972 30308
rect 8972 30252 9028 30308
rect 9028 30252 9032 30308
rect 8968 30248 9032 30252
rect 8968 30088 9032 30152
rect 8968 29988 9032 29992
rect 8968 29932 8972 29988
rect 8972 29932 9028 29988
rect 9028 29932 9032 29988
rect 8968 29928 9032 29932
rect 8968 29828 9032 29832
rect 8968 29772 8972 29828
rect 8972 29772 9028 29828
rect 9028 29772 9032 29828
rect 8968 29768 9032 29772
rect 8968 29668 9032 29672
rect 8968 29612 8972 29668
rect 8972 29612 9028 29668
rect 9028 29612 9032 29668
rect 8968 29608 9032 29612
rect 8968 29508 9032 29512
rect 8968 29452 8972 29508
rect 8972 29452 9028 29508
rect 9028 29452 9032 29508
rect 8968 29448 9032 29452
rect 8968 29348 9032 29352
rect 8968 29292 8972 29348
rect 8972 29292 9028 29348
rect 9028 29292 9032 29348
rect 8968 29288 9032 29292
rect 8968 29188 9032 29192
rect 8968 29132 8972 29188
rect 8972 29132 9028 29188
rect 9028 29132 9032 29188
rect 8968 29128 9032 29132
rect 8968 29028 9032 29032
rect 8968 28972 8972 29028
rect 8972 28972 9028 29028
rect 9028 28972 9032 29028
rect 8968 28968 9032 28972
rect 8968 28868 9032 28872
rect 8968 28812 8972 28868
rect 8972 28812 9028 28868
rect 9028 28812 9032 28868
rect 8968 28808 9032 28812
rect 8968 28648 9032 28712
rect 8968 28488 9032 28552
rect 8968 28328 9032 28392
rect 8968 28168 9032 28232
rect 8968 28068 9032 28072
rect 8968 28012 8972 28068
rect 8972 28012 9028 28068
rect 9028 28012 9032 28068
rect 8968 28008 9032 28012
rect 8968 27908 9032 27912
rect 8968 27852 8972 27908
rect 8972 27852 9028 27908
rect 9028 27852 9032 27908
rect 8968 27848 9032 27852
rect 8968 27748 9032 27752
rect 8968 27692 8972 27748
rect 8972 27692 9028 27748
rect 9028 27692 9032 27748
rect 8968 27688 9032 27692
rect 8968 27588 9032 27592
rect 8968 27532 8972 27588
rect 8972 27532 9028 27588
rect 9028 27532 9032 27588
rect 8968 27528 9032 27532
rect 8968 27428 9032 27432
rect 8968 27372 8972 27428
rect 8972 27372 9028 27428
rect 9028 27372 9032 27428
rect 8968 27368 9032 27372
rect 8968 27268 9032 27272
rect 8968 27212 8972 27268
rect 8972 27212 9028 27268
rect 9028 27212 9032 27268
rect 8968 27208 9032 27212
rect 8968 27108 9032 27112
rect 8968 27052 8972 27108
rect 8972 27052 9028 27108
rect 9028 27052 9032 27108
rect 8968 27048 9032 27052
rect 8968 26948 9032 26952
rect 8968 26892 8972 26948
rect 8972 26892 9028 26948
rect 9028 26892 9032 26948
rect 8968 26888 9032 26892
rect 8968 26728 9032 26792
rect 8968 26568 9032 26632
rect 8968 26408 9032 26472
rect 8968 26248 9032 26312
rect 8968 26148 9032 26152
rect 8968 26092 8972 26148
rect 8972 26092 9028 26148
rect 9028 26092 9032 26148
rect 8968 26088 9032 26092
rect 8968 25988 9032 25992
rect 8968 25932 8972 25988
rect 8972 25932 9028 25988
rect 9028 25932 9032 25988
rect 8968 25928 9032 25932
rect 8968 25828 9032 25832
rect 8968 25772 8972 25828
rect 8972 25772 9028 25828
rect 9028 25772 9032 25828
rect 8968 25768 9032 25772
rect 8968 25668 9032 25672
rect 8968 25612 8972 25668
rect 8972 25612 9028 25668
rect 9028 25612 9032 25668
rect 8968 25608 9032 25612
rect 8968 25508 9032 25512
rect 8968 25452 8972 25508
rect 8972 25452 9028 25508
rect 9028 25452 9032 25508
rect 8968 25448 9032 25452
rect 8968 25348 9032 25352
rect 8968 25292 8972 25348
rect 8972 25292 9028 25348
rect 9028 25292 9032 25348
rect 8968 25288 9032 25292
rect 8968 25188 9032 25192
rect 8968 25132 8972 25188
rect 8972 25132 9028 25188
rect 9028 25132 9032 25188
rect 8968 25128 9032 25132
rect 8968 25028 9032 25032
rect 8968 24972 8972 25028
rect 8972 24972 9028 25028
rect 9028 24972 9032 25028
rect 8968 24968 9032 24972
rect 8968 24808 9032 24872
rect 8968 24708 9032 24712
rect 8968 24652 8972 24708
rect 8972 24652 9028 24708
rect 9028 24652 9032 24708
rect 8968 24648 9032 24652
rect 8968 24548 9032 24552
rect 8968 24492 8972 24548
rect 8972 24492 9028 24548
rect 9028 24492 9032 24548
rect 8968 24488 9032 24492
rect 8968 24388 9032 24392
rect 8968 24332 8972 24388
rect 8972 24332 9028 24388
rect 9028 24332 9032 24388
rect 8968 24328 9032 24332
rect 8968 24228 9032 24232
rect 8968 24172 8972 24228
rect 8972 24172 9028 24228
rect 9028 24172 9032 24228
rect 8968 24168 9032 24172
rect 8968 24068 9032 24072
rect 8968 24012 8972 24068
rect 8972 24012 9028 24068
rect 9028 24012 9032 24068
rect 8968 24008 9032 24012
rect 8968 23908 9032 23912
rect 8968 23852 8972 23908
rect 8972 23852 9028 23908
rect 9028 23852 9032 23908
rect 8968 23848 9032 23852
rect 8968 23748 9032 23752
rect 8968 23692 8972 23748
rect 8972 23692 9028 23748
rect 9028 23692 9032 23748
rect 8968 23688 9032 23692
rect 8968 23588 9032 23592
rect 8968 23532 8972 23588
rect 8972 23532 9028 23588
rect 9028 23532 9032 23588
rect 8968 23528 9032 23532
rect 8968 23428 9032 23432
rect 8968 23372 8972 23428
rect 8972 23372 9028 23428
rect 9028 23372 9032 23428
rect 8968 23368 9032 23372
rect 8968 23268 9032 23272
rect 8968 23212 8972 23268
rect 8972 23212 9028 23268
rect 9028 23212 9032 23268
rect 8968 23208 9032 23212
rect 8968 23108 9032 23112
rect 8968 23052 8972 23108
rect 8972 23052 9028 23108
rect 9028 23052 9032 23108
rect 8968 23048 9032 23052
rect 8968 22948 9032 22952
rect 8968 22892 8972 22948
rect 8972 22892 9028 22948
rect 9028 22892 9032 22948
rect 8968 22888 9032 22892
rect 8968 22788 9032 22792
rect 8968 22732 8972 22788
rect 8972 22732 9028 22788
rect 9028 22732 9032 22788
rect 8968 22728 9032 22732
rect 8968 22628 9032 22632
rect 8968 22572 8972 22628
rect 8972 22572 9028 22628
rect 9028 22572 9032 22628
rect 8968 22568 9032 22572
rect 8968 22468 9032 22472
rect 8968 22412 8972 22468
rect 8972 22412 9028 22468
rect 9028 22412 9032 22468
rect 8968 22408 9032 22412
rect 8968 22308 9032 22312
rect 8968 22252 8972 22308
rect 8972 22252 9028 22308
rect 9028 22252 9032 22308
rect 8968 22248 9032 22252
rect 8968 22148 9032 22152
rect 8968 22092 8972 22148
rect 8972 22092 9028 22148
rect 9028 22092 9032 22148
rect 8968 22088 9032 22092
rect 8968 21928 9032 21992
rect 8968 21828 9032 21832
rect 8968 21772 8972 21828
rect 8972 21772 9028 21828
rect 9028 21772 9032 21828
rect 8968 21768 9032 21772
rect 8968 21668 9032 21672
rect 8968 21612 8972 21668
rect 8972 21612 9028 21668
rect 9028 21612 9032 21668
rect 8968 21608 9032 21612
rect 8968 21508 9032 21512
rect 8968 21452 8972 21508
rect 8972 21452 9028 21508
rect 9028 21452 9032 21508
rect 8968 21448 9032 21452
rect 8968 21348 9032 21352
rect 8968 21292 8972 21348
rect 8972 21292 9028 21348
rect 9028 21292 9032 21348
rect 8968 21288 9032 21292
rect 8968 21188 9032 21192
rect 8968 21132 8972 21188
rect 8972 21132 9028 21188
rect 9028 21132 9032 21188
rect 8968 21128 9032 21132
rect 8968 21028 9032 21032
rect 8968 20972 8972 21028
rect 8972 20972 9028 21028
rect 9028 20972 9032 21028
rect 8968 20968 9032 20972
rect 8968 20868 9032 20872
rect 8968 20812 8972 20868
rect 8972 20812 9028 20868
rect 9028 20812 9032 20868
rect 8968 20808 9032 20812
rect 8968 20708 9032 20712
rect 8968 20652 8972 20708
rect 8972 20652 9028 20708
rect 9028 20652 9032 20708
rect 8968 20648 9032 20652
rect 8968 20488 9032 20552
rect 8968 20328 9032 20392
rect 8968 20168 9032 20232
rect 8968 20008 9032 20072
rect 8968 19908 9032 19912
rect 8968 19852 8972 19908
rect 8972 19852 9028 19908
rect 9028 19852 9032 19908
rect 8968 19848 9032 19852
rect 8968 19748 9032 19752
rect 8968 19692 8972 19748
rect 8972 19692 9028 19748
rect 9028 19692 9032 19748
rect 8968 19688 9032 19692
rect 8968 19588 9032 19592
rect 8968 19532 8972 19588
rect 8972 19532 9028 19588
rect 9028 19532 9032 19588
rect 8968 19528 9032 19532
rect 8968 19428 9032 19432
rect 8968 19372 8972 19428
rect 8972 19372 9028 19428
rect 9028 19372 9032 19428
rect 8968 19368 9032 19372
rect 8968 19268 9032 19272
rect 8968 19212 8972 19268
rect 8972 19212 9028 19268
rect 9028 19212 9032 19268
rect 8968 19208 9032 19212
rect 8968 19108 9032 19112
rect 8968 19052 8972 19108
rect 8972 19052 9028 19108
rect 9028 19052 9032 19108
rect 8968 19048 9032 19052
rect 8968 18948 9032 18952
rect 8968 18892 8972 18948
rect 8972 18892 9028 18948
rect 9028 18892 9032 18948
rect 8968 18888 9032 18892
rect 8968 18788 9032 18792
rect 8968 18732 8972 18788
rect 8972 18732 9028 18788
rect 9028 18732 9032 18788
rect 8968 18728 9032 18732
rect 8968 18568 9032 18632
rect 8968 18408 9032 18472
rect 8968 18248 9032 18312
rect 8968 18088 9032 18152
rect 8968 17988 9032 17992
rect 8968 17932 8972 17988
rect 8972 17932 9028 17988
rect 9028 17932 9032 17988
rect 8968 17928 9032 17932
rect 8968 17828 9032 17832
rect 8968 17772 8972 17828
rect 8972 17772 9028 17828
rect 9028 17772 9032 17828
rect 8968 17768 9032 17772
rect 8968 17668 9032 17672
rect 8968 17612 8972 17668
rect 8972 17612 9028 17668
rect 9028 17612 9032 17668
rect 8968 17608 9032 17612
rect 8968 17508 9032 17512
rect 8968 17452 8972 17508
rect 8972 17452 9028 17508
rect 9028 17452 9032 17508
rect 8968 17448 9032 17452
rect 8968 17348 9032 17352
rect 8968 17292 8972 17348
rect 8972 17292 9028 17348
rect 9028 17292 9032 17348
rect 8968 17288 9032 17292
rect 8968 17188 9032 17192
rect 8968 17132 8972 17188
rect 8972 17132 9028 17188
rect 9028 17132 9032 17188
rect 8968 17128 9032 17132
rect 8968 17028 9032 17032
rect 8968 16972 8972 17028
rect 8972 16972 9028 17028
rect 9028 16972 9032 17028
rect 8968 16968 9032 16972
rect 8968 16868 9032 16872
rect 8968 16812 8972 16868
rect 8972 16812 9028 16868
rect 9028 16812 9032 16868
rect 8968 16808 9032 16812
rect 8968 16648 9032 16712
rect 8968 16548 9032 16552
rect 8968 16492 8972 16548
rect 8972 16492 9028 16548
rect 9028 16492 9032 16548
rect 8968 16488 9032 16492
rect 8968 16388 9032 16392
rect 8968 16332 8972 16388
rect 8972 16332 9028 16388
rect 9028 16332 9032 16388
rect 8968 16328 9032 16332
rect 8968 16228 9032 16232
rect 8968 16172 8972 16228
rect 8972 16172 9028 16228
rect 9028 16172 9032 16228
rect 8968 16168 9032 16172
rect 8968 16068 9032 16072
rect 8968 16012 8972 16068
rect 8972 16012 9028 16068
rect 9028 16012 9032 16068
rect 8968 16008 9032 16012
rect 8968 15908 9032 15912
rect 8968 15852 8972 15908
rect 8972 15852 9028 15908
rect 9028 15852 9032 15908
rect 8968 15848 9032 15852
rect 8968 15748 9032 15752
rect 8968 15692 8972 15748
rect 8972 15692 9028 15748
rect 9028 15692 9032 15748
rect 8968 15688 9032 15692
rect 8968 15588 9032 15592
rect 8968 15532 8972 15588
rect 8972 15532 9028 15588
rect 9028 15532 9032 15588
rect 8968 15528 9032 15532
rect 8968 15428 9032 15432
rect 8968 15372 8972 15428
rect 8972 15372 9028 15428
rect 9028 15372 9032 15428
rect 8968 15368 9032 15372
rect 8968 15268 9032 15272
rect 8968 15212 8972 15268
rect 8972 15212 9028 15268
rect 9028 15212 9032 15268
rect 8968 15208 9032 15212
rect 8968 15108 9032 15112
rect 8968 15052 8972 15108
rect 8972 15052 9028 15108
rect 9028 15052 9032 15108
rect 8968 15048 9032 15052
rect 8968 14948 9032 14952
rect 8968 14892 8972 14948
rect 8972 14892 9028 14948
rect 9028 14892 9032 14948
rect 8968 14888 9032 14892
rect 8968 14788 9032 14792
rect 8968 14732 8972 14788
rect 8972 14732 9028 14788
rect 9028 14732 9032 14788
rect 8968 14728 9032 14732
rect 8968 14628 9032 14632
rect 8968 14572 8972 14628
rect 8972 14572 9028 14628
rect 9028 14572 9032 14628
rect 8968 14568 9032 14572
rect 8968 14468 9032 14472
rect 8968 14412 8972 14468
rect 8972 14412 9028 14468
rect 9028 14412 9032 14468
rect 8968 14408 9032 14412
rect 8968 14308 9032 14312
rect 8968 14252 8972 14308
rect 8972 14252 9028 14308
rect 9028 14252 9032 14308
rect 8968 14248 9032 14252
rect 8968 14148 9032 14152
rect 8968 14092 8972 14148
rect 8972 14092 9028 14148
rect 9028 14092 9032 14148
rect 8968 14088 9032 14092
rect 8968 13988 9032 13992
rect 8968 13932 8972 13988
rect 8972 13932 9028 13988
rect 9028 13932 9032 13988
rect 8968 13928 9032 13932
rect 8968 13768 9032 13832
rect 8968 13668 9032 13672
rect 8968 13612 8972 13668
rect 8972 13612 9028 13668
rect 9028 13612 9032 13668
rect 8968 13608 9032 13612
rect 8968 13508 9032 13512
rect 8968 13452 8972 13508
rect 8972 13452 9028 13508
rect 9028 13452 9032 13508
rect 8968 13448 9032 13452
rect 8968 13348 9032 13352
rect 8968 13292 8972 13348
rect 8972 13292 9028 13348
rect 9028 13292 9032 13348
rect 8968 13288 9032 13292
rect 8968 13188 9032 13192
rect 8968 13132 8972 13188
rect 8972 13132 9028 13188
rect 9028 13132 9032 13188
rect 8968 13128 9032 13132
rect 8968 13028 9032 13032
rect 8968 12972 8972 13028
rect 8972 12972 9028 13028
rect 9028 12972 9032 13028
rect 8968 12968 9032 12972
rect 8968 12868 9032 12872
rect 8968 12812 8972 12868
rect 8972 12812 9028 12868
rect 9028 12812 9032 12868
rect 8968 12808 9032 12812
rect 8968 12708 9032 12712
rect 8968 12652 8972 12708
rect 8972 12652 9028 12708
rect 9028 12652 9032 12708
rect 8968 12648 9032 12652
rect 8968 12548 9032 12552
rect 8968 12492 8972 12548
rect 8972 12492 9028 12548
rect 9028 12492 9032 12548
rect 8968 12488 9032 12492
rect 8968 12328 9032 12392
rect 8968 12168 9032 12232
rect 8968 12008 9032 12072
rect 8968 11848 9032 11912
rect 8968 11748 9032 11752
rect 8968 11692 8972 11748
rect 8972 11692 9028 11748
rect 9028 11692 9032 11748
rect 8968 11688 9032 11692
rect 8968 11588 9032 11592
rect 8968 11532 8972 11588
rect 8972 11532 9028 11588
rect 9028 11532 9032 11588
rect 8968 11528 9032 11532
rect 8968 11428 9032 11432
rect 8968 11372 8972 11428
rect 8972 11372 9028 11428
rect 9028 11372 9032 11428
rect 8968 11368 9032 11372
rect 8968 11268 9032 11272
rect 8968 11212 8972 11268
rect 8972 11212 9028 11268
rect 9028 11212 9032 11268
rect 8968 11208 9032 11212
rect 8968 11108 9032 11112
rect 8968 11052 8972 11108
rect 8972 11052 9028 11108
rect 9028 11052 9032 11108
rect 8968 11048 9032 11052
rect 8968 10948 9032 10952
rect 8968 10892 8972 10948
rect 8972 10892 9028 10948
rect 9028 10892 9032 10948
rect 8968 10888 9032 10892
rect 8968 10788 9032 10792
rect 8968 10732 8972 10788
rect 8972 10732 9028 10788
rect 9028 10732 9032 10788
rect 8968 10728 9032 10732
rect 8968 10628 9032 10632
rect 8968 10572 8972 10628
rect 8972 10572 9028 10628
rect 9028 10572 9032 10628
rect 8968 10568 9032 10572
rect 8968 10468 9032 10472
rect 8968 10412 8972 10468
rect 8972 10412 9028 10468
rect 9028 10412 9032 10468
rect 8968 10408 9032 10412
rect 8968 10308 9032 10312
rect 8968 10252 8972 10308
rect 8972 10252 9028 10308
rect 9028 10252 9032 10308
rect 8968 10248 9032 10252
rect 8968 10148 9032 10152
rect 8968 10092 8972 10148
rect 8972 10092 9028 10148
rect 9028 10092 9032 10148
rect 8968 10088 9032 10092
rect 8968 9988 9032 9992
rect 8968 9932 8972 9988
rect 8972 9932 9028 9988
rect 9028 9932 9032 9988
rect 8968 9928 9032 9932
rect 8968 9828 9032 9832
rect 8968 9772 8972 9828
rect 8972 9772 9028 9828
rect 9028 9772 9032 9828
rect 8968 9768 9032 9772
rect 8968 9608 9032 9672
rect 8968 9508 9032 9512
rect 8968 9452 8972 9508
rect 8972 9452 9028 9508
rect 9028 9452 9032 9508
rect 8968 9448 9032 9452
rect 8968 9348 9032 9352
rect 8968 9292 8972 9348
rect 8972 9292 9028 9348
rect 9028 9292 9032 9348
rect 8968 9288 9032 9292
rect 8968 9128 9032 9192
rect 8968 9028 9032 9032
rect 8968 8972 8972 9028
rect 8972 8972 9028 9028
rect 9028 8972 9032 9028
rect 8968 8968 9032 8972
rect 8968 8868 9032 8872
rect 8968 8812 8972 8868
rect 8972 8812 9028 8868
rect 9028 8812 9032 8868
rect 8968 8808 9032 8812
rect 8968 8708 9032 8712
rect 8968 8652 8972 8708
rect 8972 8652 9028 8708
rect 9028 8652 9032 8708
rect 8968 8648 9032 8652
rect 8968 8548 9032 8552
rect 8968 8492 8972 8548
rect 8972 8492 9028 8548
rect 9028 8492 9032 8548
rect 8968 8488 9032 8492
rect 8968 8388 9032 8392
rect 8968 8332 8972 8388
rect 8972 8332 9028 8388
rect 9028 8332 9032 8388
rect 8968 8328 9032 8332
rect 8968 8228 9032 8232
rect 8968 8172 8972 8228
rect 8972 8172 9028 8228
rect 9028 8172 9032 8228
rect 8968 8168 9032 8172
rect 8968 8068 9032 8072
rect 8968 8012 8972 8068
rect 8972 8012 9028 8068
rect 9028 8012 9032 8068
rect 8968 8008 9032 8012
rect 8968 7908 9032 7912
rect 8968 7852 8972 7908
rect 8972 7852 9028 7908
rect 9028 7852 9032 7908
rect 8968 7848 9032 7852
rect 8968 7748 9032 7752
rect 8968 7692 8972 7748
rect 8972 7692 9028 7748
rect 9028 7692 9032 7748
rect 8968 7688 9032 7692
rect 8968 7528 9032 7592
rect 8968 7428 9032 7432
rect 8968 7372 8972 7428
rect 8972 7372 9028 7428
rect 9028 7372 9032 7428
rect 8968 7368 9032 7372
rect 8968 7268 9032 7272
rect 8968 7212 8972 7268
rect 8972 7212 9028 7268
rect 9028 7212 9032 7268
rect 8968 7208 9032 7212
rect 8968 7048 9032 7112
rect 8968 6948 9032 6952
rect 8968 6892 8972 6948
rect 8972 6892 9028 6948
rect 9028 6892 9032 6948
rect 8968 6888 9032 6892
rect 8968 6788 9032 6792
rect 8968 6732 8972 6788
rect 8972 6732 9028 6788
rect 9028 6732 9032 6788
rect 8968 6728 9032 6732
rect 8968 6568 9032 6632
rect 8968 6468 9032 6472
rect 8968 6412 8972 6468
rect 8972 6412 9028 6468
rect 9028 6412 9032 6468
rect 8968 6408 9032 6412
rect 8968 6308 9032 6312
rect 8968 6252 8972 6308
rect 8972 6252 9028 6308
rect 9028 6252 9032 6308
rect 8968 6248 9032 6252
rect 8968 6148 9032 6152
rect 8968 6092 8972 6148
rect 8972 6092 9028 6148
rect 9028 6092 9032 6148
rect 8968 6088 9032 6092
rect 8968 5988 9032 5992
rect 8968 5932 8972 5988
rect 8972 5932 9028 5988
rect 9028 5932 9032 5988
rect 8968 5928 9032 5932
rect 8968 5828 9032 5832
rect 8968 5772 8972 5828
rect 8972 5772 9028 5828
rect 9028 5772 9032 5828
rect 8968 5768 9032 5772
rect 8968 5668 9032 5672
rect 8968 5612 8972 5668
rect 8972 5612 9028 5668
rect 9028 5612 9032 5668
rect 8968 5608 9032 5612
rect 8968 5508 9032 5512
rect 8968 5452 8972 5508
rect 8972 5452 9028 5508
rect 9028 5452 9032 5508
rect 8968 5448 9032 5452
rect 8968 5348 9032 5352
rect 8968 5292 8972 5348
rect 8972 5292 9028 5348
rect 9028 5292 9032 5348
rect 8968 5288 9032 5292
rect 8968 5188 9032 5192
rect 8968 5132 8972 5188
rect 8972 5132 9028 5188
rect 9028 5132 9032 5188
rect 8968 5128 9032 5132
rect 8968 5028 9032 5032
rect 8968 4972 8972 5028
rect 8972 4972 9028 5028
rect 9028 4972 9032 5028
rect 8968 4968 9032 4972
rect 8968 4868 9032 4872
rect 8968 4812 8972 4868
rect 8972 4812 9028 4868
rect 9028 4812 9032 4868
rect 8968 4808 9032 4812
rect 8968 4708 9032 4712
rect 8968 4652 8972 4708
rect 8972 4652 9028 4708
rect 9028 4652 9032 4708
rect 8968 4648 9032 4652
rect 8968 4548 9032 4552
rect 8968 4492 8972 4548
rect 8972 4492 9028 4548
rect 9028 4492 9032 4548
rect 8968 4488 9032 4492
rect 8968 4388 9032 4392
rect 8968 4332 8972 4388
rect 8972 4332 9028 4388
rect 9028 4332 9032 4388
rect 8968 4328 9032 4332
rect 8968 4228 9032 4232
rect 8968 4172 8972 4228
rect 8972 4172 9028 4228
rect 9028 4172 9032 4228
rect 8968 4168 9032 4172
rect 8968 4068 9032 4072
rect 8968 4012 8972 4068
rect 8972 4012 9028 4068
rect 9028 4012 9032 4068
rect 8968 4008 9032 4012
rect 8968 3908 9032 3912
rect 8968 3852 8972 3908
rect 8972 3852 9028 3908
rect 9028 3852 9032 3908
rect 8968 3848 9032 3852
rect 8968 3688 9032 3752
rect 8968 3528 9032 3592
rect 8968 3428 9032 3432
rect 8968 3372 8972 3428
rect 8972 3372 9028 3428
rect 9028 3372 9032 3428
rect 8968 3368 9032 3372
rect 8968 3268 9032 3272
rect 8968 3212 8972 3268
rect 8972 3212 9028 3268
rect 9028 3212 9032 3268
rect 8968 3208 9032 3212
rect 8968 3108 9032 3112
rect 8968 3052 8972 3108
rect 8972 3052 9028 3108
rect 9028 3052 9032 3108
rect 8968 3048 9032 3052
rect 8968 2948 9032 2952
rect 8968 2892 8972 2948
rect 8972 2892 9028 2948
rect 9028 2892 9032 2948
rect 8968 2888 9032 2892
rect 8968 2788 9032 2792
rect 8968 2732 8972 2788
rect 8972 2732 9028 2788
rect 9028 2732 9032 2788
rect 8968 2728 9032 2732
rect 8968 2628 9032 2632
rect 8968 2572 8972 2628
rect 8972 2572 9028 2628
rect 9028 2572 9032 2628
rect 8968 2568 9032 2572
rect 8968 2468 9032 2472
rect 8968 2412 8972 2468
rect 8972 2412 9028 2468
rect 9028 2412 9032 2468
rect 8968 2408 9032 2412
rect 8968 2308 9032 2312
rect 8968 2252 8972 2308
rect 8972 2252 9028 2308
rect 9028 2252 9032 2308
rect 8968 2248 9032 2252
rect 8968 2148 9032 2152
rect 8968 2092 8972 2148
rect 8972 2092 9028 2148
rect 9028 2092 9032 2148
rect 8968 2088 9032 2092
rect 8968 1988 9032 1992
rect 8968 1932 8972 1988
rect 8972 1932 9028 1988
rect 9028 1932 9032 1988
rect 8968 1928 9032 1932
rect 8968 1768 9032 1832
rect 8968 1668 9032 1672
rect 8968 1612 8972 1668
rect 8972 1612 9028 1668
rect 9028 1612 9032 1668
rect 8968 1608 9032 1612
rect 8968 1508 9032 1512
rect 8968 1452 8972 1508
rect 8972 1452 9028 1508
rect 9028 1452 9032 1508
rect 8968 1448 9032 1452
rect 8968 1348 9032 1352
rect 8968 1292 8972 1348
rect 8972 1292 9028 1348
rect 9028 1292 9032 1348
rect 8968 1288 9032 1292
rect 8968 1188 9032 1192
rect 8968 1132 8972 1188
rect 8972 1132 9028 1188
rect 9028 1132 9032 1188
rect 8968 1128 9032 1132
rect 8968 1028 9032 1032
rect 8968 972 8972 1028
rect 8972 972 9028 1028
rect 9028 972 9032 1028
rect 8968 968 9032 972
rect 8968 808 9032 872
rect 8968 648 9032 712
rect 8968 548 9032 552
rect 8968 492 8972 548
rect 8972 492 9028 548
rect 9028 492 9032 548
rect 8968 488 9032 492
rect 8968 388 9032 392
rect 8968 332 8972 388
rect 8972 332 9028 388
rect 9028 332 9032 388
rect 8968 328 9032 332
rect 8968 228 9032 232
rect 8968 172 8972 228
rect 8972 172 9028 228
rect 9028 172 9032 228
rect 8968 168 9032 172
rect 8968 68 9032 72
rect 8968 12 8972 68
rect 8972 12 9028 68
rect 9028 12 9032 68
rect 8968 8 9032 12
rect 8968 -632 9032 -568
rect 8968 -712 9032 -648
rect 8968 -792 9032 -728
rect 8968 -872 9032 -808
rect 8968 -952 9032 -888
rect 248 -2072 312 -2008
rect 8968 -2072 9032 -2008
rect 9288 31428 9352 31432
rect 9288 31372 9292 31428
rect 9292 31372 9348 31428
rect 9348 31372 9352 31428
rect 9288 31368 9352 31372
rect 9288 31268 9352 31272
rect 9288 31212 9292 31268
rect 9292 31212 9348 31268
rect 9348 31212 9352 31268
rect 9288 31208 9352 31212
rect 9288 31108 9352 31112
rect 9288 31052 9292 31108
rect 9292 31052 9348 31108
rect 9348 31052 9352 31108
rect 9288 31048 9352 31052
rect 9288 30948 9352 30952
rect 9288 30892 9292 30948
rect 9292 30892 9348 30948
rect 9348 30892 9352 30948
rect 9288 30888 9352 30892
rect 9288 30788 9352 30792
rect 9288 30732 9292 30788
rect 9292 30732 9348 30788
rect 9348 30732 9352 30788
rect 9288 30728 9352 30732
rect 9288 30628 9352 30632
rect 9288 30572 9292 30628
rect 9292 30572 9348 30628
rect 9348 30572 9352 30628
rect 9288 30568 9352 30572
rect 9288 30468 9352 30472
rect 9288 30412 9292 30468
rect 9292 30412 9348 30468
rect 9348 30412 9352 30468
rect 9288 30408 9352 30412
rect 9288 30308 9352 30312
rect 9288 30252 9292 30308
rect 9292 30252 9348 30308
rect 9348 30252 9352 30308
rect 9288 30248 9352 30252
rect 9288 30088 9352 30152
rect 9288 29988 9352 29992
rect 9288 29932 9292 29988
rect 9292 29932 9348 29988
rect 9348 29932 9352 29988
rect 9288 29928 9352 29932
rect 9288 29828 9352 29832
rect 9288 29772 9292 29828
rect 9292 29772 9348 29828
rect 9348 29772 9352 29828
rect 9288 29768 9352 29772
rect 9288 29668 9352 29672
rect 9288 29612 9292 29668
rect 9292 29612 9348 29668
rect 9348 29612 9352 29668
rect 9288 29608 9352 29612
rect 9288 29508 9352 29512
rect 9288 29452 9292 29508
rect 9292 29452 9348 29508
rect 9348 29452 9352 29508
rect 9288 29448 9352 29452
rect 9288 29348 9352 29352
rect 9288 29292 9292 29348
rect 9292 29292 9348 29348
rect 9348 29292 9352 29348
rect 9288 29288 9352 29292
rect 9288 29188 9352 29192
rect 9288 29132 9292 29188
rect 9292 29132 9348 29188
rect 9348 29132 9352 29188
rect 9288 29128 9352 29132
rect 9288 29028 9352 29032
rect 9288 28972 9292 29028
rect 9292 28972 9348 29028
rect 9348 28972 9352 29028
rect 9288 28968 9352 28972
rect 9288 28868 9352 28872
rect 9288 28812 9292 28868
rect 9292 28812 9348 28868
rect 9348 28812 9352 28868
rect 9288 28808 9352 28812
rect 9288 28648 9352 28712
rect 9288 28488 9352 28552
rect 9288 28328 9352 28392
rect 9288 28168 9352 28232
rect 9288 28068 9352 28072
rect 9288 28012 9292 28068
rect 9292 28012 9348 28068
rect 9348 28012 9352 28068
rect 9288 28008 9352 28012
rect 9288 27908 9352 27912
rect 9288 27852 9292 27908
rect 9292 27852 9348 27908
rect 9348 27852 9352 27908
rect 9288 27848 9352 27852
rect 9288 27748 9352 27752
rect 9288 27692 9292 27748
rect 9292 27692 9348 27748
rect 9348 27692 9352 27748
rect 9288 27688 9352 27692
rect 9288 27588 9352 27592
rect 9288 27532 9292 27588
rect 9292 27532 9348 27588
rect 9348 27532 9352 27588
rect 9288 27528 9352 27532
rect 9288 27428 9352 27432
rect 9288 27372 9292 27428
rect 9292 27372 9348 27428
rect 9348 27372 9352 27428
rect 9288 27368 9352 27372
rect 9288 27268 9352 27272
rect 9288 27212 9292 27268
rect 9292 27212 9348 27268
rect 9348 27212 9352 27268
rect 9288 27208 9352 27212
rect 9288 27108 9352 27112
rect 9288 27052 9292 27108
rect 9292 27052 9348 27108
rect 9348 27052 9352 27108
rect 9288 27048 9352 27052
rect 9288 26948 9352 26952
rect 9288 26892 9292 26948
rect 9292 26892 9348 26948
rect 9348 26892 9352 26948
rect 9288 26888 9352 26892
rect 9288 26728 9352 26792
rect 9288 26568 9352 26632
rect 9288 26408 9352 26472
rect 9288 26248 9352 26312
rect 9288 26148 9352 26152
rect 9288 26092 9292 26148
rect 9292 26092 9348 26148
rect 9348 26092 9352 26148
rect 9288 26088 9352 26092
rect 9288 25988 9352 25992
rect 9288 25932 9292 25988
rect 9292 25932 9348 25988
rect 9348 25932 9352 25988
rect 9288 25928 9352 25932
rect 9288 25828 9352 25832
rect 9288 25772 9292 25828
rect 9292 25772 9348 25828
rect 9348 25772 9352 25828
rect 9288 25768 9352 25772
rect 9288 25668 9352 25672
rect 9288 25612 9292 25668
rect 9292 25612 9348 25668
rect 9348 25612 9352 25668
rect 9288 25608 9352 25612
rect 9288 25508 9352 25512
rect 9288 25452 9292 25508
rect 9292 25452 9348 25508
rect 9348 25452 9352 25508
rect 9288 25448 9352 25452
rect 9288 25348 9352 25352
rect 9288 25292 9292 25348
rect 9292 25292 9348 25348
rect 9348 25292 9352 25348
rect 9288 25288 9352 25292
rect 9288 25188 9352 25192
rect 9288 25132 9292 25188
rect 9292 25132 9348 25188
rect 9348 25132 9352 25188
rect 9288 25128 9352 25132
rect 9288 25028 9352 25032
rect 9288 24972 9292 25028
rect 9292 24972 9348 25028
rect 9348 24972 9352 25028
rect 9288 24968 9352 24972
rect 9288 24808 9352 24872
rect 9288 24708 9352 24712
rect 9288 24652 9292 24708
rect 9292 24652 9348 24708
rect 9348 24652 9352 24708
rect 9288 24648 9352 24652
rect 9288 24548 9352 24552
rect 9288 24492 9292 24548
rect 9292 24492 9348 24548
rect 9348 24492 9352 24548
rect 9288 24488 9352 24492
rect 9288 24388 9352 24392
rect 9288 24332 9292 24388
rect 9292 24332 9348 24388
rect 9348 24332 9352 24388
rect 9288 24328 9352 24332
rect 9288 24228 9352 24232
rect 9288 24172 9292 24228
rect 9292 24172 9348 24228
rect 9348 24172 9352 24228
rect 9288 24168 9352 24172
rect 9288 24068 9352 24072
rect 9288 24012 9292 24068
rect 9292 24012 9348 24068
rect 9348 24012 9352 24068
rect 9288 24008 9352 24012
rect 9288 23908 9352 23912
rect 9288 23852 9292 23908
rect 9292 23852 9348 23908
rect 9348 23852 9352 23908
rect 9288 23848 9352 23852
rect 9288 23748 9352 23752
rect 9288 23692 9292 23748
rect 9292 23692 9348 23748
rect 9348 23692 9352 23748
rect 9288 23688 9352 23692
rect 9288 23588 9352 23592
rect 9288 23532 9292 23588
rect 9292 23532 9348 23588
rect 9348 23532 9352 23588
rect 9288 23528 9352 23532
rect 9288 23428 9352 23432
rect 9288 23372 9292 23428
rect 9292 23372 9348 23428
rect 9348 23372 9352 23428
rect 9288 23368 9352 23372
rect 9288 23268 9352 23272
rect 9288 23212 9292 23268
rect 9292 23212 9348 23268
rect 9348 23212 9352 23268
rect 9288 23208 9352 23212
rect 9288 23108 9352 23112
rect 9288 23052 9292 23108
rect 9292 23052 9348 23108
rect 9348 23052 9352 23108
rect 9288 23048 9352 23052
rect 9288 22948 9352 22952
rect 9288 22892 9292 22948
rect 9292 22892 9348 22948
rect 9348 22892 9352 22948
rect 9288 22888 9352 22892
rect 9288 22788 9352 22792
rect 9288 22732 9292 22788
rect 9292 22732 9348 22788
rect 9348 22732 9352 22788
rect 9288 22728 9352 22732
rect 9288 22628 9352 22632
rect 9288 22572 9292 22628
rect 9292 22572 9348 22628
rect 9348 22572 9352 22628
rect 9288 22568 9352 22572
rect 9288 22468 9352 22472
rect 9288 22412 9292 22468
rect 9292 22412 9348 22468
rect 9348 22412 9352 22468
rect 9288 22408 9352 22412
rect 9288 22308 9352 22312
rect 9288 22252 9292 22308
rect 9292 22252 9348 22308
rect 9348 22252 9352 22308
rect 9288 22248 9352 22252
rect 9288 22148 9352 22152
rect 9288 22092 9292 22148
rect 9292 22092 9348 22148
rect 9348 22092 9352 22148
rect 9288 22088 9352 22092
rect 9288 21928 9352 21992
rect 9288 21828 9352 21832
rect 9288 21772 9292 21828
rect 9292 21772 9348 21828
rect 9348 21772 9352 21828
rect 9288 21768 9352 21772
rect 9288 21668 9352 21672
rect 9288 21612 9292 21668
rect 9292 21612 9348 21668
rect 9348 21612 9352 21668
rect 9288 21608 9352 21612
rect 9288 21508 9352 21512
rect 9288 21452 9292 21508
rect 9292 21452 9348 21508
rect 9348 21452 9352 21508
rect 9288 21448 9352 21452
rect 9288 21348 9352 21352
rect 9288 21292 9292 21348
rect 9292 21292 9348 21348
rect 9348 21292 9352 21348
rect 9288 21288 9352 21292
rect 9288 21188 9352 21192
rect 9288 21132 9292 21188
rect 9292 21132 9348 21188
rect 9348 21132 9352 21188
rect 9288 21128 9352 21132
rect 9288 21028 9352 21032
rect 9288 20972 9292 21028
rect 9292 20972 9348 21028
rect 9348 20972 9352 21028
rect 9288 20968 9352 20972
rect 9288 20868 9352 20872
rect 9288 20812 9292 20868
rect 9292 20812 9348 20868
rect 9348 20812 9352 20868
rect 9288 20808 9352 20812
rect 9288 20708 9352 20712
rect 9288 20652 9292 20708
rect 9292 20652 9348 20708
rect 9348 20652 9352 20708
rect 9288 20648 9352 20652
rect 9288 20488 9352 20552
rect 9288 20328 9352 20392
rect 9288 20168 9352 20232
rect 9288 20008 9352 20072
rect 9288 19908 9352 19912
rect 9288 19852 9292 19908
rect 9292 19852 9348 19908
rect 9348 19852 9352 19908
rect 9288 19848 9352 19852
rect 9288 19748 9352 19752
rect 9288 19692 9292 19748
rect 9292 19692 9348 19748
rect 9348 19692 9352 19748
rect 9288 19688 9352 19692
rect 9288 19588 9352 19592
rect 9288 19532 9292 19588
rect 9292 19532 9348 19588
rect 9348 19532 9352 19588
rect 9288 19528 9352 19532
rect 9288 19428 9352 19432
rect 9288 19372 9292 19428
rect 9292 19372 9348 19428
rect 9348 19372 9352 19428
rect 9288 19368 9352 19372
rect 9288 19268 9352 19272
rect 9288 19212 9292 19268
rect 9292 19212 9348 19268
rect 9348 19212 9352 19268
rect 9288 19208 9352 19212
rect 9288 19108 9352 19112
rect 9288 19052 9292 19108
rect 9292 19052 9348 19108
rect 9348 19052 9352 19108
rect 9288 19048 9352 19052
rect 9288 18948 9352 18952
rect 9288 18892 9292 18948
rect 9292 18892 9348 18948
rect 9348 18892 9352 18948
rect 9288 18888 9352 18892
rect 9288 18788 9352 18792
rect 9288 18732 9292 18788
rect 9292 18732 9348 18788
rect 9348 18732 9352 18788
rect 9288 18728 9352 18732
rect 9288 18568 9352 18632
rect 9288 18408 9352 18472
rect 9288 18248 9352 18312
rect 9288 18088 9352 18152
rect 9288 17988 9352 17992
rect 9288 17932 9292 17988
rect 9292 17932 9348 17988
rect 9348 17932 9352 17988
rect 9288 17928 9352 17932
rect 9288 17828 9352 17832
rect 9288 17772 9292 17828
rect 9292 17772 9348 17828
rect 9348 17772 9352 17828
rect 9288 17768 9352 17772
rect 9288 17668 9352 17672
rect 9288 17612 9292 17668
rect 9292 17612 9348 17668
rect 9348 17612 9352 17668
rect 9288 17608 9352 17612
rect 9288 17508 9352 17512
rect 9288 17452 9292 17508
rect 9292 17452 9348 17508
rect 9348 17452 9352 17508
rect 9288 17448 9352 17452
rect 9288 17348 9352 17352
rect 9288 17292 9292 17348
rect 9292 17292 9348 17348
rect 9348 17292 9352 17348
rect 9288 17288 9352 17292
rect 9288 17188 9352 17192
rect 9288 17132 9292 17188
rect 9292 17132 9348 17188
rect 9348 17132 9352 17188
rect 9288 17128 9352 17132
rect 9288 17028 9352 17032
rect 9288 16972 9292 17028
rect 9292 16972 9348 17028
rect 9348 16972 9352 17028
rect 9288 16968 9352 16972
rect 9288 16868 9352 16872
rect 9288 16812 9292 16868
rect 9292 16812 9348 16868
rect 9348 16812 9352 16868
rect 9288 16808 9352 16812
rect 9288 16648 9352 16712
rect 9288 16548 9352 16552
rect 9288 16492 9292 16548
rect 9292 16492 9348 16548
rect 9348 16492 9352 16548
rect 9288 16488 9352 16492
rect 9288 16388 9352 16392
rect 9288 16332 9292 16388
rect 9292 16332 9348 16388
rect 9348 16332 9352 16388
rect 9288 16328 9352 16332
rect 9288 16228 9352 16232
rect 9288 16172 9292 16228
rect 9292 16172 9348 16228
rect 9348 16172 9352 16228
rect 9288 16168 9352 16172
rect 9288 16068 9352 16072
rect 9288 16012 9292 16068
rect 9292 16012 9348 16068
rect 9348 16012 9352 16068
rect 9288 16008 9352 16012
rect 9288 15908 9352 15912
rect 9288 15852 9292 15908
rect 9292 15852 9348 15908
rect 9348 15852 9352 15908
rect 9288 15848 9352 15852
rect 9288 15748 9352 15752
rect 9288 15692 9292 15748
rect 9292 15692 9348 15748
rect 9348 15692 9352 15748
rect 9288 15688 9352 15692
rect 9288 15588 9352 15592
rect 9288 15532 9292 15588
rect 9292 15532 9348 15588
rect 9348 15532 9352 15588
rect 9288 15528 9352 15532
rect 9288 15428 9352 15432
rect 9288 15372 9292 15428
rect 9292 15372 9348 15428
rect 9348 15372 9352 15428
rect 9288 15368 9352 15372
rect 9288 15268 9352 15272
rect 9288 15212 9292 15268
rect 9292 15212 9348 15268
rect 9348 15212 9352 15268
rect 9288 15208 9352 15212
rect 9288 15108 9352 15112
rect 9288 15052 9292 15108
rect 9292 15052 9348 15108
rect 9348 15052 9352 15108
rect 9288 15048 9352 15052
rect 9288 14948 9352 14952
rect 9288 14892 9292 14948
rect 9292 14892 9348 14948
rect 9348 14892 9352 14948
rect 9288 14888 9352 14892
rect 9288 14788 9352 14792
rect 9288 14732 9292 14788
rect 9292 14732 9348 14788
rect 9348 14732 9352 14788
rect 9288 14728 9352 14732
rect 9288 14628 9352 14632
rect 9288 14572 9292 14628
rect 9292 14572 9348 14628
rect 9348 14572 9352 14628
rect 9288 14568 9352 14572
rect 9288 14468 9352 14472
rect 9288 14412 9292 14468
rect 9292 14412 9348 14468
rect 9348 14412 9352 14468
rect 9288 14408 9352 14412
rect 9288 14308 9352 14312
rect 9288 14252 9292 14308
rect 9292 14252 9348 14308
rect 9348 14252 9352 14308
rect 9288 14248 9352 14252
rect 9288 14148 9352 14152
rect 9288 14092 9292 14148
rect 9292 14092 9348 14148
rect 9348 14092 9352 14148
rect 9288 14088 9352 14092
rect 9288 13988 9352 13992
rect 9288 13932 9292 13988
rect 9292 13932 9348 13988
rect 9348 13932 9352 13988
rect 9288 13928 9352 13932
rect 9288 13768 9352 13832
rect 9288 13668 9352 13672
rect 9288 13612 9292 13668
rect 9292 13612 9348 13668
rect 9348 13612 9352 13668
rect 9288 13608 9352 13612
rect 9288 13508 9352 13512
rect 9288 13452 9292 13508
rect 9292 13452 9348 13508
rect 9348 13452 9352 13508
rect 9288 13448 9352 13452
rect 9288 13348 9352 13352
rect 9288 13292 9292 13348
rect 9292 13292 9348 13348
rect 9348 13292 9352 13348
rect 9288 13288 9352 13292
rect 9288 13188 9352 13192
rect 9288 13132 9292 13188
rect 9292 13132 9348 13188
rect 9348 13132 9352 13188
rect 9288 13128 9352 13132
rect 9288 13028 9352 13032
rect 9288 12972 9292 13028
rect 9292 12972 9348 13028
rect 9348 12972 9352 13028
rect 9288 12968 9352 12972
rect 9288 12868 9352 12872
rect 9288 12812 9292 12868
rect 9292 12812 9348 12868
rect 9348 12812 9352 12868
rect 9288 12808 9352 12812
rect 9288 12708 9352 12712
rect 9288 12652 9292 12708
rect 9292 12652 9348 12708
rect 9348 12652 9352 12708
rect 9288 12648 9352 12652
rect 9288 12548 9352 12552
rect 9288 12492 9292 12548
rect 9292 12492 9348 12548
rect 9348 12492 9352 12548
rect 9288 12488 9352 12492
rect 9288 12328 9352 12392
rect 9288 12168 9352 12232
rect 9288 12008 9352 12072
rect 9288 11848 9352 11912
rect 9288 11748 9352 11752
rect 9288 11692 9292 11748
rect 9292 11692 9348 11748
rect 9348 11692 9352 11748
rect 9288 11688 9352 11692
rect 9288 11588 9352 11592
rect 9288 11532 9292 11588
rect 9292 11532 9348 11588
rect 9348 11532 9352 11588
rect 9288 11528 9352 11532
rect 9288 11428 9352 11432
rect 9288 11372 9292 11428
rect 9292 11372 9348 11428
rect 9348 11372 9352 11428
rect 9288 11368 9352 11372
rect 9288 11268 9352 11272
rect 9288 11212 9292 11268
rect 9292 11212 9348 11268
rect 9348 11212 9352 11268
rect 9288 11208 9352 11212
rect 9288 11108 9352 11112
rect 9288 11052 9292 11108
rect 9292 11052 9348 11108
rect 9348 11052 9352 11108
rect 9288 11048 9352 11052
rect 9288 10948 9352 10952
rect 9288 10892 9292 10948
rect 9292 10892 9348 10948
rect 9348 10892 9352 10948
rect 9288 10888 9352 10892
rect 9288 10788 9352 10792
rect 9288 10732 9292 10788
rect 9292 10732 9348 10788
rect 9348 10732 9352 10788
rect 9288 10728 9352 10732
rect 9288 10628 9352 10632
rect 9288 10572 9292 10628
rect 9292 10572 9348 10628
rect 9348 10572 9352 10628
rect 9288 10568 9352 10572
rect 9288 10468 9352 10472
rect 9288 10412 9292 10468
rect 9292 10412 9348 10468
rect 9348 10412 9352 10468
rect 9288 10408 9352 10412
rect 9288 10308 9352 10312
rect 9288 10252 9292 10308
rect 9292 10252 9348 10308
rect 9348 10252 9352 10308
rect 9288 10248 9352 10252
rect 9288 10148 9352 10152
rect 9288 10092 9292 10148
rect 9292 10092 9348 10148
rect 9348 10092 9352 10148
rect 9288 10088 9352 10092
rect 9288 9988 9352 9992
rect 9288 9932 9292 9988
rect 9292 9932 9348 9988
rect 9348 9932 9352 9988
rect 9288 9928 9352 9932
rect 9288 9828 9352 9832
rect 9288 9772 9292 9828
rect 9292 9772 9348 9828
rect 9348 9772 9352 9828
rect 9288 9768 9352 9772
rect 9288 9608 9352 9672
rect 9288 9508 9352 9512
rect 9288 9452 9292 9508
rect 9292 9452 9348 9508
rect 9348 9452 9352 9508
rect 9288 9448 9352 9452
rect 9288 9348 9352 9352
rect 9288 9292 9292 9348
rect 9292 9292 9348 9348
rect 9348 9292 9352 9348
rect 9288 9288 9352 9292
rect 9288 9128 9352 9192
rect 9288 9028 9352 9032
rect 9288 8972 9292 9028
rect 9292 8972 9348 9028
rect 9348 8972 9352 9028
rect 9288 8968 9352 8972
rect 9288 8868 9352 8872
rect 9288 8812 9292 8868
rect 9292 8812 9348 8868
rect 9348 8812 9352 8868
rect 9288 8808 9352 8812
rect 9288 8708 9352 8712
rect 9288 8652 9292 8708
rect 9292 8652 9348 8708
rect 9348 8652 9352 8708
rect 9288 8648 9352 8652
rect 9288 8548 9352 8552
rect 9288 8492 9292 8548
rect 9292 8492 9348 8548
rect 9348 8492 9352 8548
rect 9288 8488 9352 8492
rect 9288 8388 9352 8392
rect 9288 8332 9292 8388
rect 9292 8332 9348 8388
rect 9348 8332 9352 8388
rect 9288 8328 9352 8332
rect 9288 8228 9352 8232
rect 9288 8172 9292 8228
rect 9292 8172 9348 8228
rect 9348 8172 9352 8228
rect 9288 8168 9352 8172
rect 9288 8068 9352 8072
rect 9288 8012 9292 8068
rect 9292 8012 9348 8068
rect 9348 8012 9352 8068
rect 9288 8008 9352 8012
rect 9288 7908 9352 7912
rect 9288 7852 9292 7908
rect 9292 7852 9348 7908
rect 9348 7852 9352 7908
rect 9288 7848 9352 7852
rect 9288 7748 9352 7752
rect 9288 7692 9292 7748
rect 9292 7692 9348 7748
rect 9348 7692 9352 7748
rect 9288 7688 9352 7692
rect 9288 7528 9352 7592
rect 9288 7428 9352 7432
rect 9288 7372 9292 7428
rect 9292 7372 9348 7428
rect 9348 7372 9352 7428
rect 9288 7368 9352 7372
rect 9288 7268 9352 7272
rect 9288 7212 9292 7268
rect 9292 7212 9348 7268
rect 9348 7212 9352 7268
rect 9288 7208 9352 7212
rect 9288 7048 9352 7112
rect 9288 6948 9352 6952
rect 9288 6892 9292 6948
rect 9292 6892 9348 6948
rect 9348 6892 9352 6948
rect 9288 6888 9352 6892
rect 9288 6788 9352 6792
rect 9288 6732 9292 6788
rect 9292 6732 9348 6788
rect 9348 6732 9352 6788
rect 9288 6728 9352 6732
rect 9288 6568 9352 6632
rect 9288 6468 9352 6472
rect 9288 6412 9292 6468
rect 9292 6412 9348 6468
rect 9348 6412 9352 6468
rect 9288 6408 9352 6412
rect 9288 6308 9352 6312
rect 9288 6252 9292 6308
rect 9292 6252 9348 6308
rect 9348 6252 9352 6308
rect 9288 6248 9352 6252
rect 9288 6148 9352 6152
rect 9288 6092 9292 6148
rect 9292 6092 9348 6148
rect 9348 6092 9352 6148
rect 9288 6088 9352 6092
rect 9288 5988 9352 5992
rect 9288 5932 9292 5988
rect 9292 5932 9348 5988
rect 9348 5932 9352 5988
rect 9288 5928 9352 5932
rect 9288 5828 9352 5832
rect 9288 5772 9292 5828
rect 9292 5772 9348 5828
rect 9348 5772 9352 5828
rect 9288 5768 9352 5772
rect 9288 5668 9352 5672
rect 9288 5612 9292 5668
rect 9292 5612 9348 5668
rect 9348 5612 9352 5668
rect 9288 5608 9352 5612
rect 9288 5508 9352 5512
rect 9288 5452 9292 5508
rect 9292 5452 9348 5508
rect 9348 5452 9352 5508
rect 9288 5448 9352 5452
rect 9288 5348 9352 5352
rect 9288 5292 9292 5348
rect 9292 5292 9348 5348
rect 9348 5292 9352 5348
rect 9288 5288 9352 5292
rect 9288 5188 9352 5192
rect 9288 5132 9292 5188
rect 9292 5132 9348 5188
rect 9348 5132 9352 5188
rect 9288 5128 9352 5132
rect 9288 5028 9352 5032
rect 9288 4972 9292 5028
rect 9292 4972 9348 5028
rect 9348 4972 9352 5028
rect 9288 4968 9352 4972
rect 9288 4868 9352 4872
rect 9288 4812 9292 4868
rect 9292 4812 9348 4868
rect 9348 4812 9352 4868
rect 9288 4808 9352 4812
rect 9288 4708 9352 4712
rect 9288 4652 9292 4708
rect 9292 4652 9348 4708
rect 9348 4652 9352 4708
rect 9288 4648 9352 4652
rect 9288 4548 9352 4552
rect 9288 4492 9292 4548
rect 9292 4492 9348 4548
rect 9348 4492 9352 4548
rect 9288 4488 9352 4492
rect 9288 4388 9352 4392
rect 9288 4332 9292 4388
rect 9292 4332 9348 4388
rect 9348 4332 9352 4388
rect 9288 4328 9352 4332
rect 9288 4228 9352 4232
rect 9288 4172 9292 4228
rect 9292 4172 9348 4228
rect 9348 4172 9352 4228
rect 9288 4168 9352 4172
rect 9288 4068 9352 4072
rect 9288 4012 9292 4068
rect 9292 4012 9348 4068
rect 9348 4012 9352 4068
rect 9288 4008 9352 4012
rect 9288 3908 9352 3912
rect 9288 3852 9292 3908
rect 9292 3852 9348 3908
rect 9348 3852 9352 3908
rect 9288 3848 9352 3852
rect 9288 3688 9352 3752
rect 9288 3528 9352 3592
rect 9288 3428 9352 3432
rect 9288 3372 9292 3428
rect 9292 3372 9348 3428
rect 9348 3372 9352 3428
rect 9288 3368 9352 3372
rect 9288 3268 9352 3272
rect 9288 3212 9292 3268
rect 9292 3212 9348 3268
rect 9348 3212 9352 3268
rect 9288 3208 9352 3212
rect 9288 3108 9352 3112
rect 9288 3052 9292 3108
rect 9292 3052 9348 3108
rect 9348 3052 9352 3108
rect 9288 3048 9352 3052
rect 9288 2948 9352 2952
rect 9288 2892 9292 2948
rect 9292 2892 9348 2948
rect 9348 2892 9352 2948
rect 9288 2888 9352 2892
rect 9288 2788 9352 2792
rect 9288 2732 9292 2788
rect 9292 2732 9348 2788
rect 9348 2732 9352 2788
rect 9288 2728 9352 2732
rect 9288 2628 9352 2632
rect 9288 2572 9292 2628
rect 9292 2572 9348 2628
rect 9348 2572 9352 2628
rect 9288 2568 9352 2572
rect 9288 2468 9352 2472
rect 9288 2412 9292 2468
rect 9292 2412 9348 2468
rect 9348 2412 9352 2468
rect 9288 2408 9352 2412
rect 9288 2308 9352 2312
rect 9288 2252 9292 2308
rect 9292 2252 9348 2308
rect 9348 2252 9352 2308
rect 9288 2248 9352 2252
rect 9288 2148 9352 2152
rect 9288 2092 9292 2148
rect 9292 2092 9348 2148
rect 9348 2092 9352 2148
rect 9288 2088 9352 2092
rect 9288 1988 9352 1992
rect 9288 1932 9292 1988
rect 9292 1932 9348 1988
rect 9348 1932 9352 1988
rect 9288 1928 9352 1932
rect 9288 1768 9352 1832
rect 9288 1668 9352 1672
rect 9288 1612 9292 1668
rect 9292 1612 9348 1668
rect 9348 1612 9352 1668
rect 9288 1608 9352 1612
rect 9288 1508 9352 1512
rect 9288 1452 9292 1508
rect 9292 1452 9348 1508
rect 9348 1452 9352 1508
rect 9288 1448 9352 1452
rect 9288 1348 9352 1352
rect 9288 1292 9292 1348
rect 9292 1292 9348 1348
rect 9348 1292 9352 1348
rect 9288 1288 9352 1292
rect 9288 1188 9352 1192
rect 9288 1132 9292 1188
rect 9292 1132 9348 1188
rect 9348 1132 9352 1188
rect 9288 1128 9352 1132
rect 9288 1028 9352 1032
rect 9288 972 9292 1028
rect 9292 972 9348 1028
rect 9348 972 9352 1028
rect 9288 968 9352 972
rect 9288 808 9352 872
rect 9288 648 9352 712
rect 9288 548 9352 552
rect 9288 492 9292 548
rect 9292 492 9348 548
rect 9348 492 9352 548
rect 9288 488 9352 492
rect 9288 388 9352 392
rect 9288 332 9292 388
rect 9292 332 9348 388
rect 9348 332 9352 388
rect 9288 328 9352 332
rect 9288 228 9352 232
rect 9288 172 9292 228
rect 9292 172 9348 228
rect 9348 172 9352 228
rect 9288 168 9352 172
rect 9288 68 9352 72
rect 9288 12 9292 68
rect 9292 12 9348 68
rect 9348 12 9352 68
rect 9288 8 9352 12
rect 9288 -632 9352 -568
rect 9288 -712 9352 -648
rect 9288 -792 9352 -728
rect 9288 -872 9352 -808
rect 9288 -952 9352 -888
rect 9448 31428 9512 31432
rect 9448 31372 9452 31428
rect 9452 31372 9508 31428
rect 9508 31372 9512 31428
rect 9448 31368 9512 31372
rect 9448 31268 9512 31272
rect 9448 31212 9452 31268
rect 9452 31212 9508 31268
rect 9508 31212 9512 31268
rect 9448 31208 9512 31212
rect 9448 31108 9512 31112
rect 9448 31052 9452 31108
rect 9452 31052 9508 31108
rect 9508 31052 9512 31108
rect 9448 31048 9512 31052
rect 9448 30948 9512 30952
rect 9448 30892 9452 30948
rect 9452 30892 9508 30948
rect 9508 30892 9512 30948
rect 9448 30888 9512 30892
rect 9448 30788 9512 30792
rect 9448 30732 9452 30788
rect 9452 30732 9508 30788
rect 9508 30732 9512 30788
rect 9448 30728 9512 30732
rect 9448 30628 9512 30632
rect 9448 30572 9452 30628
rect 9452 30572 9508 30628
rect 9508 30572 9512 30628
rect 9448 30568 9512 30572
rect 9448 30468 9512 30472
rect 9448 30412 9452 30468
rect 9452 30412 9508 30468
rect 9508 30412 9512 30468
rect 9448 30408 9512 30412
rect 9448 30308 9512 30312
rect 9448 30252 9452 30308
rect 9452 30252 9508 30308
rect 9508 30252 9512 30308
rect 9448 30248 9512 30252
rect 9448 30088 9512 30152
rect 9448 29988 9512 29992
rect 9448 29932 9452 29988
rect 9452 29932 9508 29988
rect 9508 29932 9512 29988
rect 9448 29928 9512 29932
rect 9448 29828 9512 29832
rect 9448 29772 9452 29828
rect 9452 29772 9508 29828
rect 9508 29772 9512 29828
rect 9448 29768 9512 29772
rect 9448 29668 9512 29672
rect 9448 29612 9452 29668
rect 9452 29612 9508 29668
rect 9508 29612 9512 29668
rect 9448 29608 9512 29612
rect 9448 29508 9512 29512
rect 9448 29452 9452 29508
rect 9452 29452 9508 29508
rect 9508 29452 9512 29508
rect 9448 29448 9512 29452
rect 9448 29348 9512 29352
rect 9448 29292 9452 29348
rect 9452 29292 9508 29348
rect 9508 29292 9512 29348
rect 9448 29288 9512 29292
rect 9448 29188 9512 29192
rect 9448 29132 9452 29188
rect 9452 29132 9508 29188
rect 9508 29132 9512 29188
rect 9448 29128 9512 29132
rect 9448 29028 9512 29032
rect 9448 28972 9452 29028
rect 9452 28972 9508 29028
rect 9508 28972 9512 29028
rect 9448 28968 9512 28972
rect 9448 28868 9512 28872
rect 9448 28812 9452 28868
rect 9452 28812 9508 28868
rect 9508 28812 9512 28868
rect 9448 28808 9512 28812
rect 9448 28648 9512 28712
rect 9448 28488 9512 28552
rect 9448 28328 9512 28392
rect 9448 28168 9512 28232
rect 9448 28068 9512 28072
rect 9448 28012 9452 28068
rect 9452 28012 9508 28068
rect 9508 28012 9512 28068
rect 9448 28008 9512 28012
rect 9448 27908 9512 27912
rect 9448 27852 9452 27908
rect 9452 27852 9508 27908
rect 9508 27852 9512 27908
rect 9448 27848 9512 27852
rect 9448 27748 9512 27752
rect 9448 27692 9452 27748
rect 9452 27692 9508 27748
rect 9508 27692 9512 27748
rect 9448 27688 9512 27692
rect 9448 27588 9512 27592
rect 9448 27532 9452 27588
rect 9452 27532 9508 27588
rect 9508 27532 9512 27588
rect 9448 27528 9512 27532
rect 9448 27428 9512 27432
rect 9448 27372 9452 27428
rect 9452 27372 9508 27428
rect 9508 27372 9512 27428
rect 9448 27368 9512 27372
rect 9448 27268 9512 27272
rect 9448 27212 9452 27268
rect 9452 27212 9508 27268
rect 9508 27212 9512 27268
rect 9448 27208 9512 27212
rect 9448 27108 9512 27112
rect 9448 27052 9452 27108
rect 9452 27052 9508 27108
rect 9508 27052 9512 27108
rect 9448 27048 9512 27052
rect 9448 26948 9512 26952
rect 9448 26892 9452 26948
rect 9452 26892 9508 26948
rect 9508 26892 9512 26948
rect 9448 26888 9512 26892
rect 9448 26728 9512 26792
rect 9448 26568 9512 26632
rect 9448 26408 9512 26472
rect 9448 26248 9512 26312
rect 9448 26148 9512 26152
rect 9448 26092 9452 26148
rect 9452 26092 9508 26148
rect 9508 26092 9512 26148
rect 9448 26088 9512 26092
rect 9448 25988 9512 25992
rect 9448 25932 9452 25988
rect 9452 25932 9508 25988
rect 9508 25932 9512 25988
rect 9448 25928 9512 25932
rect 9448 25828 9512 25832
rect 9448 25772 9452 25828
rect 9452 25772 9508 25828
rect 9508 25772 9512 25828
rect 9448 25768 9512 25772
rect 9448 25668 9512 25672
rect 9448 25612 9452 25668
rect 9452 25612 9508 25668
rect 9508 25612 9512 25668
rect 9448 25608 9512 25612
rect 9448 25508 9512 25512
rect 9448 25452 9452 25508
rect 9452 25452 9508 25508
rect 9508 25452 9512 25508
rect 9448 25448 9512 25452
rect 9448 25348 9512 25352
rect 9448 25292 9452 25348
rect 9452 25292 9508 25348
rect 9508 25292 9512 25348
rect 9448 25288 9512 25292
rect 9448 25188 9512 25192
rect 9448 25132 9452 25188
rect 9452 25132 9508 25188
rect 9508 25132 9512 25188
rect 9448 25128 9512 25132
rect 9448 25028 9512 25032
rect 9448 24972 9452 25028
rect 9452 24972 9508 25028
rect 9508 24972 9512 25028
rect 9448 24968 9512 24972
rect 9448 24808 9512 24872
rect 9448 24708 9512 24712
rect 9448 24652 9452 24708
rect 9452 24652 9508 24708
rect 9508 24652 9512 24708
rect 9448 24648 9512 24652
rect 9448 24548 9512 24552
rect 9448 24492 9452 24548
rect 9452 24492 9508 24548
rect 9508 24492 9512 24548
rect 9448 24488 9512 24492
rect 9448 24388 9512 24392
rect 9448 24332 9452 24388
rect 9452 24332 9508 24388
rect 9508 24332 9512 24388
rect 9448 24328 9512 24332
rect 9448 24228 9512 24232
rect 9448 24172 9452 24228
rect 9452 24172 9508 24228
rect 9508 24172 9512 24228
rect 9448 24168 9512 24172
rect 9448 24068 9512 24072
rect 9448 24012 9452 24068
rect 9452 24012 9508 24068
rect 9508 24012 9512 24068
rect 9448 24008 9512 24012
rect 9448 23908 9512 23912
rect 9448 23852 9452 23908
rect 9452 23852 9508 23908
rect 9508 23852 9512 23908
rect 9448 23848 9512 23852
rect 9448 23748 9512 23752
rect 9448 23692 9452 23748
rect 9452 23692 9508 23748
rect 9508 23692 9512 23748
rect 9448 23688 9512 23692
rect 9448 23588 9512 23592
rect 9448 23532 9452 23588
rect 9452 23532 9508 23588
rect 9508 23532 9512 23588
rect 9448 23528 9512 23532
rect 9448 23428 9512 23432
rect 9448 23372 9452 23428
rect 9452 23372 9508 23428
rect 9508 23372 9512 23428
rect 9448 23368 9512 23372
rect 9448 23268 9512 23272
rect 9448 23212 9452 23268
rect 9452 23212 9508 23268
rect 9508 23212 9512 23268
rect 9448 23208 9512 23212
rect 9448 23108 9512 23112
rect 9448 23052 9452 23108
rect 9452 23052 9508 23108
rect 9508 23052 9512 23108
rect 9448 23048 9512 23052
rect 9448 22948 9512 22952
rect 9448 22892 9452 22948
rect 9452 22892 9508 22948
rect 9508 22892 9512 22948
rect 9448 22888 9512 22892
rect 9448 22788 9512 22792
rect 9448 22732 9452 22788
rect 9452 22732 9508 22788
rect 9508 22732 9512 22788
rect 9448 22728 9512 22732
rect 9448 22628 9512 22632
rect 9448 22572 9452 22628
rect 9452 22572 9508 22628
rect 9508 22572 9512 22628
rect 9448 22568 9512 22572
rect 9448 22468 9512 22472
rect 9448 22412 9452 22468
rect 9452 22412 9508 22468
rect 9508 22412 9512 22468
rect 9448 22408 9512 22412
rect 9448 22308 9512 22312
rect 9448 22252 9452 22308
rect 9452 22252 9508 22308
rect 9508 22252 9512 22308
rect 9448 22248 9512 22252
rect 9448 22148 9512 22152
rect 9448 22092 9452 22148
rect 9452 22092 9508 22148
rect 9508 22092 9512 22148
rect 9448 22088 9512 22092
rect 9448 21928 9512 21992
rect 9448 21828 9512 21832
rect 9448 21772 9452 21828
rect 9452 21772 9508 21828
rect 9508 21772 9512 21828
rect 9448 21768 9512 21772
rect 9448 21668 9512 21672
rect 9448 21612 9452 21668
rect 9452 21612 9508 21668
rect 9508 21612 9512 21668
rect 9448 21608 9512 21612
rect 9448 21508 9512 21512
rect 9448 21452 9452 21508
rect 9452 21452 9508 21508
rect 9508 21452 9512 21508
rect 9448 21448 9512 21452
rect 9448 21348 9512 21352
rect 9448 21292 9452 21348
rect 9452 21292 9508 21348
rect 9508 21292 9512 21348
rect 9448 21288 9512 21292
rect 9448 21188 9512 21192
rect 9448 21132 9452 21188
rect 9452 21132 9508 21188
rect 9508 21132 9512 21188
rect 9448 21128 9512 21132
rect 9448 21028 9512 21032
rect 9448 20972 9452 21028
rect 9452 20972 9508 21028
rect 9508 20972 9512 21028
rect 9448 20968 9512 20972
rect 9448 20868 9512 20872
rect 9448 20812 9452 20868
rect 9452 20812 9508 20868
rect 9508 20812 9512 20868
rect 9448 20808 9512 20812
rect 9448 20708 9512 20712
rect 9448 20652 9452 20708
rect 9452 20652 9508 20708
rect 9508 20652 9512 20708
rect 9448 20648 9512 20652
rect 9448 20488 9512 20552
rect 9448 20328 9512 20392
rect 9448 20168 9512 20232
rect 9448 20008 9512 20072
rect 9448 19908 9512 19912
rect 9448 19852 9452 19908
rect 9452 19852 9508 19908
rect 9508 19852 9512 19908
rect 9448 19848 9512 19852
rect 9448 19748 9512 19752
rect 9448 19692 9452 19748
rect 9452 19692 9508 19748
rect 9508 19692 9512 19748
rect 9448 19688 9512 19692
rect 9448 19588 9512 19592
rect 9448 19532 9452 19588
rect 9452 19532 9508 19588
rect 9508 19532 9512 19588
rect 9448 19528 9512 19532
rect 9448 19428 9512 19432
rect 9448 19372 9452 19428
rect 9452 19372 9508 19428
rect 9508 19372 9512 19428
rect 9448 19368 9512 19372
rect 9448 19268 9512 19272
rect 9448 19212 9452 19268
rect 9452 19212 9508 19268
rect 9508 19212 9512 19268
rect 9448 19208 9512 19212
rect 9448 19108 9512 19112
rect 9448 19052 9452 19108
rect 9452 19052 9508 19108
rect 9508 19052 9512 19108
rect 9448 19048 9512 19052
rect 9448 18948 9512 18952
rect 9448 18892 9452 18948
rect 9452 18892 9508 18948
rect 9508 18892 9512 18948
rect 9448 18888 9512 18892
rect 9448 18788 9512 18792
rect 9448 18732 9452 18788
rect 9452 18732 9508 18788
rect 9508 18732 9512 18788
rect 9448 18728 9512 18732
rect 9448 18568 9512 18632
rect 9448 18408 9512 18472
rect 9448 18248 9512 18312
rect 9448 18088 9512 18152
rect 9448 17988 9512 17992
rect 9448 17932 9452 17988
rect 9452 17932 9508 17988
rect 9508 17932 9512 17988
rect 9448 17928 9512 17932
rect 9448 17828 9512 17832
rect 9448 17772 9452 17828
rect 9452 17772 9508 17828
rect 9508 17772 9512 17828
rect 9448 17768 9512 17772
rect 9448 17668 9512 17672
rect 9448 17612 9452 17668
rect 9452 17612 9508 17668
rect 9508 17612 9512 17668
rect 9448 17608 9512 17612
rect 9448 17508 9512 17512
rect 9448 17452 9452 17508
rect 9452 17452 9508 17508
rect 9508 17452 9512 17508
rect 9448 17448 9512 17452
rect 9448 17348 9512 17352
rect 9448 17292 9452 17348
rect 9452 17292 9508 17348
rect 9508 17292 9512 17348
rect 9448 17288 9512 17292
rect 9448 17188 9512 17192
rect 9448 17132 9452 17188
rect 9452 17132 9508 17188
rect 9508 17132 9512 17188
rect 9448 17128 9512 17132
rect 9448 17028 9512 17032
rect 9448 16972 9452 17028
rect 9452 16972 9508 17028
rect 9508 16972 9512 17028
rect 9448 16968 9512 16972
rect 9448 16868 9512 16872
rect 9448 16812 9452 16868
rect 9452 16812 9508 16868
rect 9508 16812 9512 16868
rect 9448 16808 9512 16812
rect 9448 16648 9512 16712
rect 9448 16548 9512 16552
rect 9448 16492 9452 16548
rect 9452 16492 9508 16548
rect 9508 16492 9512 16548
rect 9448 16488 9512 16492
rect 9448 16388 9512 16392
rect 9448 16332 9452 16388
rect 9452 16332 9508 16388
rect 9508 16332 9512 16388
rect 9448 16328 9512 16332
rect 9448 16228 9512 16232
rect 9448 16172 9452 16228
rect 9452 16172 9508 16228
rect 9508 16172 9512 16228
rect 9448 16168 9512 16172
rect 9448 16068 9512 16072
rect 9448 16012 9452 16068
rect 9452 16012 9508 16068
rect 9508 16012 9512 16068
rect 9448 16008 9512 16012
rect 9448 15908 9512 15912
rect 9448 15852 9452 15908
rect 9452 15852 9508 15908
rect 9508 15852 9512 15908
rect 9448 15848 9512 15852
rect 9448 15748 9512 15752
rect 9448 15692 9452 15748
rect 9452 15692 9508 15748
rect 9508 15692 9512 15748
rect 9448 15688 9512 15692
rect 9448 15588 9512 15592
rect 9448 15532 9452 15588
rect 9452 15532 9508 15588
rect 9508 15532 9512 15588
rect 9448 15528 9512 15532
rect 9448 15428 9512 15432
rect 9448 15372 9452 15428
rect 9452 15372 9508 15428
rect 9508 15372 9512 15428
rect 9448 15368 9512 15372
rect 9448 15268 9512 15272
rect 9448 15212 9452 15268
rect 9452 15212 9508 15268
rect 9508 15212 9512 15268
rect 9448 15208 9512 15212
rect 9448 15108 9512 15112
rect 9448 15052 9452 15108
rect 9452 15052 9508 15108
rect 9508 15052 9512 15108
rect 9448 15048 9512 15052
rect 9448 14948 9512 14952
rect 9448 14892 9452 14948
rect 9452 14892 9508 14948
rect 9508 14892 9512 14948
rect 9448 14888 9512 14892
rect 9448 14788 9512 14792
rect 9448 14732 9452 14788
rect 9452 14732 9508 14788
rect 9508 14732 9512 14788
rect 9448 14728 9512 14732
rect 9448 14628 9512 14632
rect 9448 14572 9452 14628
rect 9452 14572 9508 14628
rect 9508 14572 9512 14628
rect 9448 14568 9512 14572
rect 9448 14468 9512 14472
rect 9448 14412 9452 14468
rect 9452 14412 9508 14468
rect 9508 14412 9512 14468
rect 9448 14408 9512 14412
rect 9448 14308 9512 14312
rect 9448 14252 9452 14308
rect 9452 14252 9508 14308
rect 9508 14252 9512 14308
rect 9448 14248 9512 14252
rect 9448 14148 9512 14152
rect 9448 14092 9452 14148
rect 9452 14092 9508 14148
rect 9508 14092 9512 14148
rect 9448 14088 9512 14092
rect 9448 13988 9512 13992
rect 9448 13932 9452 13988
rect 9452 13932 9508 13988
rect 9508 13932 9512 13988
rect 9448 13928 9512 13932
rect 9448 13768 9512 13832
rect 9448 13668 9512 13672
rect 9448 13612 9452 13668
rect 9452 13612 9508 13668
rect 9508 13612 9512 13668
rect 9448 13608 9512 13612
rect 9448 13508 9512 13512
rect 9448 13452 9452 13508
rect 9452 13452 9508 13508
rect 9508 13452 9512 13508
rect 9448 13448 9512 13452
rect 9448 13348 9512 13352
rect 9448 13292 9452 13348
rect 9452 13292 9508 13348
rect 9508 13292 9512 13348
rect 9448 13288 9512 13292
rect 9448 13188 9512 13192
rect 9448 13132 9452 13188
rect 9452 13132 9508 13188
rect 9508 13132 9512 13188
rect 9448 13128 9512 13132
rect 9448 13028 9512 13032
rect 9448 12972 9452 13028
rect 9452 12972 9508 13028
rect 9508 12972 9512 13028
rect 9448 12968 9512 12972
rect 9448 12868 9512 12872
rect 9448 12812 9452 12868
rect 9452 12812 9508 12868
rect 9508 12812 9512 12868
rect 9448 12808 9512 12812
rect 9448 12708 9512 12712
rect 9448 12652 9452 12708
rect 9452 12652 9508 12708
rect 9508 12652 9512 12708
rect 9448 12648 9512 12652
rect 9448 12548 9512 12552
rect 9448 12492 9452 12548
rect 9452 12492 9508 12548
rect 9508 12492 9512 12548
rect 9448 12488 9512 12492
rect 9448 12328 9512 12392
rect 9448 12168 9512 12232
rect 9448 12008 9512 12072
rect 9448 11848 9512 11912
rect 9448 11748 9512 11752
rect 9448 11692 9452 11748
rect 9452 11692 9508 11748
rect 9508 11692 9512 11748
rect 9448 11688 9512 11692
rect 9448 11588 9512 11592
rect 9448 11532 9452 11588
rect 9452 11532 9508 11588
rect 9508 11532 9512 11588
rect 9448 11528 9512 11532
rect 9448 11428 9512 11432
rect 9448 11372 9452 11428
rect 9452 11372 9508 11428
rect 9508 11372 9512 11428
rect 9448 11368 9512 11372
rect 9448 11268 9512 11272
rect 9448 11212 9452 11268
rect 9452 11212 9508 11268
rect 9508 11212 9512 11268
rect 9448 11208 9512 11212
rect 9448 11108 9512 11112
rect 9448 11052 9452 11108
rect 9452 11052 9508 11108
rect 9508 11052 9512 11108
rect 9448 11048 9512 11052
rect 9448 10948 9512 10952
rect 9448 10892 9452 10948
rect 9452 10892 9508 10948
rect 9508 10892 9512 10948
rect 9448 10888 9512 10892
rect 9448 10788 9512 10792
rect 9448 10732 9452 10788
rect 9452 10732 9508 10788
rect 9508 10732 9512 10788
rect 9448 10728 9512 10732
rect 9448 10628 9512 10632
rect 9448 10572 9452 10628
rect 9452 10572 9508 10628
rect 9508 10572 9512 10628
rect 9448 10568 9512 10572
rect 9448 10468 9512 10472
rect 9448 10412 9452 10468
rect 9452 10412 9508 10468
rect 9508 10412 9512 10468
rect 9448 10408 9512 10412
rect 9448 10308 9512 10312
rect 9448 10252 9452 10308
rect 9452 10252 9508 10308
rect 9508 10252 9512 10308
rect 9448 10248 9512 10252
rect 9448 10148 9512 10152
rect 9448 10092 9452 10148
rect 9452 10092 9508 10148
rect 9508 10092 9512 10148
rect 9448 10088 9512 10092
rect 9448 9988 9512 9992
rect 9448 9932 9452 9988
rect 9452 9932 9508 9988
rect 9508 9932 9512 9988
rect 9448 9928 9512 9932
rect 9448 9828 9512 9832
rect 9448 9772 9452 9828
rect 9452 9772 9508 9828
rect 9508 9772 9512 9828
rect 9448 9768 9512 9772
rect 9448 9608 9512 9672
rect 9448 9508 9512 9512
rect 9448 9452 9452 9508
rect 9452 9452 9508 9508
rect 9508 9452 9512 9508
rect 9448 9448 9512 9452
rect 9448 9348 9512 9352
rect 9448 9292 9452 9348
rect 9452 9292 9508 9348
rect 9508 9292 9512 9348
rect 9448 9288 9512 9292
rect 9448 9128 9512 9192
rect 9448 9028 9512 9032
rect 9448 8972 9452 9028
rect 9452 8972 9508 9028
rect 9508 8972 9512 9028
rect 9448 8968 9512 8972
rect 9448 8868 9512 8872
rect 9448 8812 9452 8868
rect 9452 8812 9508 8868
rect 9508 8812 9512 8868
rect 9448 8808 9512 8812
rect 9448 8708 9512 8712
rect 9448 8652 9452 8708
rect 9452 8652 9508 8708
rect 9508 8652 9512 8708
rect 9448 8648 9512 8652
rect 9448 8548 9512 8552
rect 9448 8492 9452 8548
rect 9452 8492 9508 8548
rect 9508 8492 9512 8548
rect 9448 8488 9512 8492
rect 9448 8388 9512 8392
rect 9448 8332 9452 8388
rect 9452 8332 9508 8388
rect 9508 8332 9512 8388
rect 9448 8328 9512 8332
rect 9448 8228 9512 8232
rect 9448 8172 9452 8228
rect 9452 8172 9508 8228
rect 9508 8172 9512 8228
rect 9448 8168 9512 8172
rect 9448 8068 9512 8072
rect 9448 8012 9452 8068
rect 9452 8012 9508 8068
rect 9508 8012 9512 8068
rect 9448 8008 9512 8012
rect 9448 7908 9512 7912
rect 9448 7852 9452 7908
rect 9452 7852 9508 7908
rect 9508 7852 9512 7908
rect 9448 7848 9512 7852
rect 9448 7748 9512 7752
rect 9448 7692 9452 7748
rect 9452 7692 9508 7748
rect 9508 7692 9512 7748
rect 9448 7688 9512 7692
rect 9448 7528 9512 7592
rect 9448 7428 9512 7432
rect 9448 7372 9452 7428
rect 9452 7372 9508 7428
rect 9508 7372 9512 7428
rect 9448 7368 9512 7372
rect 9448 7268 9512 7272
rect 9448 7212 9452 7268
rect 9452 7212 9508 7268
rect 9508 7212 9512 7268
rect 9448 7208 9512 7212
rect 9448 7048 9512 7112
rect 9448 6948 9512 6952
rect 9448 6892 9452 6948
rect 9452 6892 9508 6948
rect 9508 6892 9512 6948
rect 9448 6888 9512 6892
rect 9448 6788 9512 6792
rect 9448 6732 9452 6788
rect 9452 6732 9508 6788
rect 9508 6732 9512 6788
rect 9448 6728 9512 6732
rect 9448 6568 9512 6632
rect 9448 6468 9512 6472
rect 9448 6412 9452 6468
rect 9452 6412 9508 6468
rect 9508 6412 9512 6468
rect 9448 6408 9512 6412
rect 9448 6308 9512 6312
rect 9448 6252 9452 6308
rect 9452 6252 9508 6308
rect 9508 6252 9512 6308
rect 9448 6248 9512 6252
rect 9448 6148 9512 6152
rect 9448 6092 9452 6148
rect 9452 6092 9508 6148
rect 9508 6092 9512 6148
rect 9448 6088 9512 6092
rect 9448 5988 9512 5992
rect 9448 5932 9452 5988
rect 9452 5932 9508 5988
rect 9508 5932 9512 5988
rect 9448 5928 9512 5932
rect 9448 5828 9512 5832
rect 9448 5772 9452 5828
rect 9452 5772 9508 5828
rect 9508 5772 9512 5828
rect 9448 5768 9512 5772
rect 9448 5668 9512 5672
rect 9448 5612 9452 5668
rect 9452 5612 9508 5668
rect 9508 5612 9512 5668
rect 9448 5608 9512 5612
rect 9448 5508 9512 5512
rect 9448 5452 9452 5508
rect 9452 5452 9508 5508
rect 9508 5452 9512 5508
rect 9448 5448 9512 5452
rect 9448 5348 9512 5352
rect 9448 5292 9452 5348
rect 9452 5292 9508 5348
rect 9508 5292 9512 5348
rect 9448 5288 9512 5292
rect 9448 5188 9512 5192
rect 9448 5132 9452 5188
rect 9452 5132 9508 5188
rect 9508 5132 9512 5188
rect 9448 5128 9512 5132
rect 9448 5028 9512 5032
rect 9448 4972 9452 5028
rect 9452 4972 9508 5028
rect 9508 4972 9512 5028
rect 9448 4968 9512 4972
rect 9448 4868 9512 4872
rect 9448 4812 9452 4868
rect 9452 4812 9508 4868
rect 9508 4812 9512 4868
rect 9448 4808 9512 4812
rect 9448 4708 9512 4712
rect 9448 4652 9452 4708
rect 9452 4652 9508 4708
rect 9508 4652 9512 4708
rect 9448 4648 9512 4652
rect 9448 4548 9512 4552
rect 9448 4492 9452 4548
rect 9452 4492 9508 4548
rect 9508 4492 9512 4548
rect 9448 4488 9512 4492
rect 9448 4388 9512 4392
rect 9448 4332 9452 4388
rect 9452 4332 9508 4388
rect 9508 4332 9512 4388
rect 9448 4328 9512 4332
rect 9448 4228 9512 4232
rect 9448 4172 9452 4228
rect 9452 4172 9508 4228
rect 9508 4172 9512 4228
rect 9448 4168 9512 4172
rect 9448 4068 9512 4072
rect 9448 4012 9452 4068
rect 9452 4012 9508 4068
rect 9508 4012 9512 4068
rect 9448 4008 9512 4012
rect 9448 3908 9512 3912
rect 9448 3852 9452 3908
rect 9452 3852 9508 3908
rect 9508 3852 9512 3908
rect 9448 3848 9512 3852
rect 9448 3688 9512 3752
rect 9448 3528 9512 3592
rect 9448 3428 9512 3432
rect 9448 3372 9452 3428
rect 9452 3372 9508 3428
rect 9508 3372 9512 3428
rect 9448 3368 9512 3372
rect 9448 3268 9512 3272
rect 9448 3212 9452 3268
rect 9452 3212 9508 3268
rect 9508 3212 9512 3268
rect 9448 3208 9512 3212
rect 9448 3108 9512 3112
rect 9448 3052 9452 3108
rect 9452 3052 9508 3108
rect 9508 3052 9512 3108
rect 9448 3048 9512 3052
rect 9448 2948 9512 2952
rect 9448 2892 9452 2948
rect 9452 2892 9508 2948
rect 9508 2892 9512 2948
rect 9448 2888 9512 2892
rect 9448 2788 9512 2792
rect 9448 2732 9452 2788
rect 9452 2732 9508 2788
rect 9508 2732 9512 2788
rect 9448 2728 9512 2732
rect 9448 2628 9512 2632
rect 9448 2572 9452 2628
rect 9452 2572 9508 2628
rect 9508 2572 9512 2628
rect 9448 2568 9512 2572
rect 9448 2468 9512 2472
rect 9448 2412 9452 2468
rect 9452 2412 9508 2468
rect 9508 2412 9512 2468
rect 9448 2408 9512 2412
rect 9448 2308 9512 2312
rect 9448 2252 9452 2308
rect 9452 2252 9508 2308
rect 9508 2252 9512 2308
rect 9448 2248 9512 2252
rect 9448 2148 9512 2152
rect 9448 2092 9452 2148
rect 9452 2092 9508 2148
rect 9508 2092 9512 2148
rect 9448 2088 9512 2092
rect 9448 1988 9512 1992
rect 9448 1932 9452 1988
rect 9452 1932 9508 1988
rect 9508 1932 9512 1988
rect 9448 1928 9512 1932
rect 9448 1768 9512 1832
rect 9448 1668 9512 1672
rect 9448 1612 9452 1668
rect 9452 1612 9508 1668
rect 9508 1612 9512 1668
rect 9448 1608 9512 1612
rect 9448 1508 9512 1512
rect 9448 1452 9452 1508
rect 9452 1452 9508 1508
rect 9508 1452 9512 1508
rect 9448 1448 9512 1452
rect 9448 1348 9512 1352
rect 9448 1292 9452 1348
rect 9452 1292 9508 1348
rect 9508 1292 9512 1348
rect 9448 1288 9512 1292
rect 9448 1188 9512 1192
rect 9448 1132 9452 1188
rect 9452 1132 9508 1188
rect 9508 1132 9512 1188
rect 9448 1128 9512 1132
rect 9448 1028 9512 1032
rect 9448 972 9452 1028
rect 9452 972 9508 1028
rect 9508 972 9512 1028
rect 9448 968 9512 972
rect 9448 808 9512 872
rect 9448 648 9512 712
rect 9448 548 9512 552
rect 9448 492 9452 548
rect 9452 492 9508 548
rect 9508 492 9512 548
rect 9448 488 9512 492
rect 9448 388 9512 392
rect 9448 332 9452 388
rect 9452 332 9508 388
rect 9508 332 9512 388
rect 9448 328 9512 332
rect 9448 228 9512 232
rect 9448 172 9452 228
rect 9452 172 9508 228
rect 9508 172 9512 228
rect 9448 168 9512 172
rect 9448 68 9512 72
rect 9448 12 9452 68
rect 9452 12 9508 68
rect 9508 12 9512 68
rect 9448 8 9512 12
rect 9768 31428 9832 31432
rect 9768 31372 9772 31428
rect 9772 31372 9828 31428
rect 9828 31372 9832 31428
rect 9768 31368 9832 31372
rect 9768 31268 9832 31272
rect 9768 31212 9772 31268
rect 9772 31212 9828 31268
rect 9828 31212 9832 31268
rect 9768 31208 9832 31212
rect 9768 31108 9832 31112
rect 9768 31052 9772 31108
rect 9772 31052 9828 31108
rect 9828 31052 9832 31108
rect 9768 31048 9832 31052
rect 9768 30948 9832 30952
rect 9768 30892 9772 30948
rect 9772 30892 9828 30948
rect 9828 30892 9832 30948
rect 9768 30888 9832 30892
rect 9768 30788 9832 30792
rect 9768 30732 9772 30788
rect 9772 30732 9828 30788
rect 9828 30732 9832 30788
rect 9768 30728 9832 30732
rect 9768 30628 9832 30632
rect 9768 30572 9772 30628
rect 9772 30572 9828 30628
rect 9828 30572 9832 30628
rect 9768 30568 9832 30572
rect 9768 30468 9832 30472
rect 9768 30412 9772 30468
rect 9772 30412 9828 30468
rect 9828 30412 9832 30468
rect 9768 30408 9832 30412
rect 9768 30308 9832 30312
rect 9768 30252 9772 30308
rect 9772 30252 9828 30308
rect 9828 30252 9832 30308
rect 9768 30248 9832 30252
rect 9768 30088 9832 30152
rect 9768 29988 9832 29992
rect 9768 29932 9772 29988
rect 9772 29932 9828 29988
rect 9828 29932 9832 29988
rect 9768 29928 9832 29932
rect 9768 29828 9832 29832
rect 9768 29772 9772 29828
rect 9772 29772 9828 29828
rect 9828 29772 9832 29828
rect 9768 29768 9832 29772
rect 9768 29668 9832 29672
rect 9768 29612 9772 29668
rect 9772 29612 9828 29668
rect 9828 29612 9832 29668
rect 9768 29608 9832 29612
rect 9768 29508 9832 29512
rect 9768 29452 9772 29508
rect 9772 29452 9828 29508
rect 9828 29452 9832 29508
rect 9768 29448 9832 29452
rect 9768 29348 9832 29352
rect 9768 29292 9772 29348
rect 9772 29292 9828 29348
rect 9828 29292 9832 29348
rect 9768 29288 9832 29292
rect 9768 29188 9832 29192
rect 9768 29132 9772 29188
rect 9772 29132 9828 29188
rect 9828 29132 9832 29188
rect 9768 29128 9832 29132
rect 9768 29028 9832 29032
rect 9768 28972 9772 29028
rect 9772 28972 9828 29028
rect 9828 28972 9832 29028
rect 9768 28968 9832 28972
rect 9768 28868 9832 28872
rect 9768 28812 9772 28868
rect 9772 28812 9828 28868
rect 9828 28812 9832 28868
rect 9768 28808 9832 28812
rect 9768 28648 9832 28712
rect 9768 28488 9832 28552
rect 9768 28328 9832 28392
rect 9768 28168 9832 28232
rect 9768 28068 9832 28072
rect 9768 28012 9772 28068
rect 9772 28012 9828 28068
rect 9828 28012 9832 28068
rect 9768 28008 9832 28012
rect 9768 27908 9832 27912
rect 9768 27852 9772 27908
rect 9772 27852 9828 27908
rect 9828 27852 9832 27908
rect 9768 27848 9832 27852
rect 9768 27748 9832 27752
rect 9768 27692 9772 27748
rect 9772 27692 9828 27748
rect 9828 27692 9832 27748
rect 9768 27688 9832 27692
rect 9768 27588 9832 27592
rect 9768 27532 9772 27588
rect 9772 27532 9828 27588
rect 9828 27532 9832 27588
rect 9768 27528 9832 27532
rect 9768 27428 9832 27432
rect 9768 27372 9772 27428
rect 9772 27372 9828 27428
rect 9828 27372 9832 27428
rect 9768 27368 9832 27372
rect 9768 27268 9832 27272
rect 9768 27212 9772 27268
rect 9772 27212 9828 27268
rect 9828 27212 9832 27268
rect 9768 27208 9832 27212
rect 9768 27108 9832 27112
rect 9768 27052 9772 27108
rect 9772 27052 9828 27108
rect 9828 27052 9832 27108
rect 9768 27048 9832 27052
rect 9768 26948 9832 26952
rect 9768 26892 9772 26948
rect 9772 26892 9828 26948
rect 9828 26892 9832 26948
rect 9768 26888 9832 26892
rect 9768 26728 9832 26792
rect 9768 26568 9832 26632
rect 9768 26408 9832 26472
rect 9768 26248 9832 26312
rect 9768 26148 9832 26152
rect 9768 26092 9772 26148
rect 9772 26092 9828 26148
rect 9828 26092 9832 26148
rect 9768 26088 9832 26092
rect 9768 25988 9832 25992
rect 9768 25932 9772 25988
rect 9772 25932 9828 25988
rect 9828 25932 9832 25988
rect 9768 25928 9832 25932
rect 9768 25828 9832 25832
rect 9768 25772 9772 25828
rect 9772 25772 9828 25828
rect 9828 25772 9832 25828
rect 9768 25768 9832 25772
rect 9768 25668 9832 25672
rect 9768 25612 9772 25668
rect 9772 25612 9828 25668
rect 9828 25612 9832 25668
rect 9768 25608 9832 25612
rect 9768 25508 9832 25512
rect 9768 25452 9772 25508
rect 9772 25452 9828 25508
rect 9828 25452 9832 25508
rect 9768 25448 9832 25452
rect 9768 25348 9832 25352
rect 9768 25292 9772 25348
rect 9772 25292 9828 25348
rect 9828 25292 9832 25348
rect 9768 25288 9832 25292
rect 9768 25188 9832 25192
rect 9768 25132 9772 25188
rect 9772 25132 9828 25188
rect 9828 25132 9832 25188
rect 9768 25128 9832 25132
rect 9768 25028 9832 25032
rect 9768 24972 9772 25028
rect 9772 24972 9828 25028
rect 9828 24972 9832 25028
rect 9768 24968 9832 24972
rect 9768 24808 9832 24872
rect 9768 24708 9832 24712
rect 9768 24652 9772 24708
rect 9772 24652 9828 24708
rect 9828 24652 9832 24708
rect 9768 24648 9832 24652
rect 9768 24548 9832 24552
rect 9768 24492 9772 24548
rect 9772 24492 9828 24548
rect 9828 24492 9832 24548
rect 9768 24488 9832 24492
rect 9768 24388 9832 24392
rect 9768 24332 9772 24388
rect 9772 24332 9828 24388
rect 9828 24332 9832 24388
rect 9768 24328 9832 24332
rect 9768 24228 9832 24232
rect 9768 24172 9772 24228
rect 9772 24172 9828 24228
rect 9828 24172 9832 24228
rect 9768 24168 9832 24172
rect 9768 24068 9832 24072
rect 9768 24012 9772 24068
rect 9772 24012 9828 24068
rect 9828 24012 9832 24068
rect 9768 24008 9832 24012
rect 9768 23908 9832 23912
rect 9768 23852 9772 23908
rect 9772 23852 9828 23908
rect 9828 23852 9832 23908
rect 9768 23848 9832 23852
rect 9768 23748 9832 23752
rect 9768 23692 9772 23748
rect 9772 23692 9828 23748
rect 9828 23692 9832 23748
rect 9768 23688 9832 23692
rect 9768 23588 9832 23592
rect 9768 23532 9772 23588
rect 9772 23532 9828 23588
rect 9828 23532 9832 23588
rect 9768 23528 9832 23532
rect 9768 23428 9832 23432
rect 9768 23372 9772 23428
rect 9772 23372 9828 23428
rect 9828 23372 9832 23428
rect 9768 23368 9832 23372
rect 9768 23268 9832 23272
rect 9768 23212 9772 23268
rect 9772 23212 9828 23268
rect 9828 23212 9832 23268
rect 9768 23208 9832 23212
rect 9768 23108 9832 23112
rect 9768 23052 9772 23108
rect 9772 23052 9828 23108
rect 9828 23052 9832 23108
rect 9768 23048 9832 23052
rect 9768 22948 9832 22952
rect 9768 22892 9772 22948
rect 9772 22892 9828 22948
rect 9828 22892 9832 22948
rect 9768 22888 9832 22892
rect 9768 22788 9832 22792
rect 9768 22732 9772 22788
rect 9772 22732 9828 22788
rect 9828 22732 9832 22788
rect 9768 22728 9832 22732
rect 9768 22628 9832 22632
rect 9768 22572 9772 22628
rect 9772 22572 9828 22628
rect 9828 22572 9832 22628
rect 9768 22568 9832 22572
rect 9768 22468 9832 22472
rect 9768 22412 9772 22468
rect 9772 22412 9828 22468
rect 9828 22412 9832 22468
rect 9768 22408 9832 22412
rect 9768 22308 9832 22312
rect 9768 22252 9772 22308
rect 9772 22252 9828 22308
rect 9828 22252 9832 22308
rect 9768 22248 9832 22252
rect 9768 22148 9832 22152
rect 9768 22092 9772 22148
rect 9772 22092 9828 22148
rect 9828 22092 9832 22148
rect 9768 22088 9832 22092
rect 9768 21928 9832 21992
rect 9768 21828 9832 21832
rect 9768 21772 9772 21828
rect 9772 21772 9828 21828
rect 9828 21772 9832 21828
rect 9768 21768 9832 21772
rect 9768 21668 9832 21672
rect 9768 21612 9772 21668
rect 9772 21612 9828 21668
rect 9828 21612 9832 21668
rect 9768 21608 9832 21612
rect 9768 21508 9832 21512
rect 9768 21452 9772 21508
rect 9772 21452 9828 21508
rect 9828 21452 9832 21508
rect 9768 21448 9832 21452
rect 9768 21348 9832 21352
rect 9768 21292 9772 21348
rect 9772 21292 9828 21348
rect 9828 21292 9832 21348
rect 9768 21288 9832 21292
rect 9768 21188 9832 21192
rect 9768 21132 9772 21188
rect 9772 21132 9828 21188
rect 9828 21132 9832 21188
rect 9768 21128 9832 21132
rect 9768 21028 9832 21032
rect 9768 20972 9772 21028
rect 9772 20972 9828 21028
rect 9828 20972 9832 21028
rect 9768 20968 9832 20972
rect 9768 20868 9832 20872
rect 9768 20812 9772 20868
rect 9772 20812 9828 20868
rect 9828 20812 9832 20868
rect 9768 20808 9832 20812
rect 9768 20708 9832 20712
rect 9768 20652 9772 20708
rect 9772 20652 9828 20708
rect 9828 20652 9832 20708
rect 9768 20648 9832 20652
rect 9768 20488 9832 20552
rect 9768 20328 9832 20392
rect 9768 20168 9832 20232
rect 9768 20008 9832 20072
rect 9768 19908 9832 19912
rect 9768 19852 9772 19908
rect 9772 19852 9828 19908
rect 9828 19852 9832 19908
rect 9768 19848 9832 19852
rect 9768 19748 9832 19752
rect 9768 19692 9772 19748
rect 9772 19692 9828 19748
rect 9828 19692 9832 19748
rect 9768 19688 9832 19692
rect 9768 19588 9832 19592
rect 9768 19532 9772 19588
rect 9772 19532 9828 19588
rect 9828 19532 9832 19588
rect 9768 19528 9832 19532
rect 9768 19428 9832 19432
rect 9768 19372 9772 19428
rect 9772 19372 9828 19428
rect 9828 19372 9832 19428
rect 9768 19368 9832 19372
rect 9768 19268 9832 19272
rect 9768 19212 9772 19268
rect 9772 19212 9828 19268
rect 9828 19212 9832 19268
rect 9768 19208 9832 19212
rect 9768 19108 9832 19112
rect 9768 19052 9772 19108
rect 9772 19052 9828 19108
rect 9828 19052 9832 19108
rect 9768 19048 9832 19052
rect 9768 18948 9832 18952
rect 9768 18892 9772 18948
rect 9772 18892 9828 18948
rect 9828 18892 9832 18948
rect 9768 18888 9832 18892
rect 9768 18788 9832 18792
rect 9768 18732 9772 18788
rect 9772 18732 9828 18788
rect 9828 18732 9832 18788
rect 9768 18728 9832 18732
rect 9768 18568 9832 18632
rect 9768 18408 9832 18472
rect 9768 18248 9832 18312
rect 9768 18088 9832 18152
rect 9768 17988 9832 17992
rect 9768 17932 9772 17988
rect 9772 17932 9828 17988
rect 9828 17932 9832 17988
rect 9768 17928 9832 17932
rect 9768 17828 9832 17832
rect 9768 17772 9772 17828
rect 9772 17772 9828 17828
rect 9828 17772 9832 17828
rect 9768 17768 9832 17772
rect 9768 17668 9832 17672
rect 9768 17612 9772 17668
rect 9772 17612 9828 17668
rect 9828 17612 9832 17668
rect 9768 17608 9832 17612
rect 9768 17508 9832 17512
rect 9768 17452 9772 17508
rect 9772 17452 9828 17508
rect 9828 17452 9832 17508
rect 9768 17448 9832 17452
rect 9768 17348 9832 17352
rect 9768 17292 9772 17348
rect 9772 17292 9828 17348
rect 9828 17292 9832 17348
rect 9768 17288 9832 17292
rect 9768 17188 9832 17192
rect 9768 17132 9772 17188
rect 9772 17132 9828 17188
rect 9828 17132 9832 17188
rect 9768 17128 9832 17132
rect 9768 17028 9832 17032
rect 9768 16972 9772 17028
rect 9772 16972 9828 17028
rect 9828 16972 9832 17028
rect 9768 16968 9832 16972
rect 9768 16868 9832 16872
rect 9768 16812 9772 16868
rect 9772 16812 9828 16868
rect 9828 16812 9832 16868
rect 9768 16808 9832 16812
rect 9768 16648 9832 16712
rect 9768 16548 9832 16552
rect 9768 16492 9772 16548
rect 9772 16492 9828 16548
rect 9828 16492 9832 16548
rect 9768 16488 9832 16492
rect 9768 16388 9832 16392
rect 9768 16332 9772 16388
rect 9772 16332 9828 16388
rect 9828 16332 9832 16388
rect 9768 16328 9832 16332
rect 9768 16228 9832 16232
rect 9768 16172 9772 16228
rect 9772 16172 9828 16228
rect 9828 16172 9832 16228
rect 9768 16168 9832 16172
rect 9768 16068 9832 16072
rect 9768 16012 9772 16068
rect 9772 16012 9828 16068
rect 9828 16012 9832 16068
rect 9768 16008 9832 16012
rect 9768 15908 9832 15912
rect 9768 15852 9772 15908
rect 9772 15852 9828 15908
rect 9828 15852 9832 15908
rect 9768 15848 9832 15852
rect 9768 15748 9832 15752
rect 9768 15692 9772 15748
rect 9772 15692 9828 15748
rect 9828 15692 9832 15748
rect 9768 15688 9832 15692
rect 9768 15588 9832 15592
rect 9768 15532 9772 15588
rect 9772 15532 9828 15588
rect 9828 15532 9832 15588
rect 9768 15528 9832 15532
rect 9768 15428 9832 15432
rect 9768 15372 9772 15428
rect 9772 15372 9828 15428
rect 9828 15372 9832 15428
rect 9768 15368 9832 15372
rect 9768 15268 9832 15272
rect 9768 15212 9772 15268
rect 9772 15212 9828 15268
rect 9828 15212 9832 15268
rect 9768 15208 9832 15212
rect 9768 15108 9832 15112
rect 9768 15052 9772 15108
rect 9772 15052 9828 15108
rect 9828 15052 9832 15108
rect 9768 15048 9832 15052
rect 9768 14948 9832 14952
rect 9768 14892 9772 14948
rect 9772 14892 9828 14948
rect 9828 14892 9832 14948
rect 9768 14888 9832 14892
rect 9768 14788 9832 14792
rect 9768 14732 9772 14788
rect 9772 14732 9828 14788
rect 9828 14732 9832 14788
rect 9768 14728 9832 14732
rect 9768 14628 9832 14632
rect 9768 14572 9772 14628
rect 9772 14572 9828 14628
rect 9828 14572 9832 14628
rect 9768 14568 9832 14572
rect 9768 14468 9832 14472
rect 9768 14412 9772 14468
rect 9772 14412 9828 14468
rect 9828 14412 9832 14468
rect 9768 14408 9832 14412
rect 9768 14308 9832 14312
rect 9768 14252 9772 14308
rect 9772 14252 9828 14308
rect 9828 14252 9832 14308
rect 9768 14248 9832 14252
rect 9768 14148 9832 14152
rect 9768 14092 9772 14148
rect 9772 14092 9828 14148
rect 9828 14092 9832 14148
rect 9768 14088 9832 14092
rect 9768 13988 9832 13992
rect 9768 13932 9772 13988
rect 9772 13932 9828 13988
rect 9828 13932 9832 13988
rect 9768 13928 9832 13932
rect 9768 13768 9832 13832
rect 9768 13668 9832 13672
rect 9768 13612 9772 13668
rect 9772 13612 9828 13668
rect 9828 13612 9832 13668
rect 9768 13608 9832 13612
rect 9768 13508 9832 13512
rect 9768 13452 9772 13508
rect 9772 13452 9828 13508
rect 9828 13452 9832 13508
rect 9768 13448 9832 13452
rect 9768 13348 9832 13352
rect 9768 13292 9772 13348
rect 9772 13292 9828 13348
rect 9828 13292 9832 13348
rect 9768 13288 9832 13292
rect 9768 13188 9832 13192
rect 9768 13132 9772 13188
rect 9772 13132 9828 13188
rect 9828 13132 9832 13188
rect 9768 13128 9832 13132
rect 9768 13028 9832 13032
rect 9768 12972 9772 13028
rect 9772 12972 9828 13028
rect 9828 12972 9832 13028
rect 9768 12968 9832 12972
rect 9768 12868 9832 12872
rect 9768 12812 9772 12868
rect 9772 12812 9828 12868
rect 9828 12812 9832 12868
rect 9768 12808 9832 12812
rect 9768 12708 9832 12712
rect 9768 12652 9772 12708
rect 9772 12652 9828 12708
rect 9828 12652 9832 12708
rect 9768 12648 9832 12652
rect 9768 12548 9832 12552
rect 9768 12492 9772 12548
rect 9772 12492 9828 12548
rect 9828 12492 9832 12548
rect 9768 12488 9832 12492
rect 9768 12328 9832 12392
rect 9768 12168 9832 12232
rect 9768 12008 9832 12072
rect 9768 11848 9832 11912
rect 9768 11748 9832 11752
rect 9768 11692 9772 11748
rect 9772 11692 9828 11748
rect 9828 11692 9832 11748
rect 9768 11688 9832 11692
rect 9768 11588 9832 11592
rect 9768 11532 9772 11588
rect 9772 11532 9828 11588
rect 9828 11532 9832 11588
rect 9768 11528 9832 11532
rect 9768 11428 9832 11432
rect 9768 11372 9772 11428
rect 9772 11372 9828 11428
rect 9828 11372 9832 11428
rect 9768 11368 9832 11372
rect 9768 11268 9832 11272
rect 9768 11212 9772 11268
rect 9772 11212 9828 11268
rect 9828 11212 9832 11268
rect 9768 11208 9832 11212
rect 9768 11108 9832 11112
rect 9768 11052 9772 11108
rect 9772 11052 9828 11108
rect 9828 11052 9832 11108
rect 9768 11048 9832 11052
rect 9768 10948 9832 10952
rect 9768 10892 9772 10948
rect 9772 10892 9828 10948
rect 9828 10892 9832 10948
rect 9768 10888 9832 10892
rect 9768 10788 9832 10792
rect 9768 10732 9772 10788
rect 9772 10732 9828 10788
rect 9828 10732 9832 10788
rect 9768 10728 9832 10732
rect 9768 10628 9832 10632
rect 9768 10572 9772 10628
rect 9772 10572 9828 10628
rect 9828 10572 9832 10628
rect 9768 10568 9832 10572
rect 9768 10468 9832 10472
rect 9768 10412 9772 10468
rect 9772 10412 9828 10468
rect 9828 10412 9832 10468
rect 9768 10408 9832 10412
rect 9768 10308 9832 10312
rect 9768 10252 9772 10308
rect 9772 10252 9828 10308
rect 9828 10252 9832 10308
rect 9768 10248 9832 10252
rect 9768 10148 9832 10152
rect 9768 10092 9772 10148
rect 9772 10092 9828 10148
rect 9828 10092 9832 10148
rect 9768 10088 9832 10092
rect 9768 9988 9832 9992
rect 9768 9932 9772 9988
rect 9772 9932 9828 9988
rect 9828 9932 9832 9988
rect 9768 9928 9832 9932
rect 9768 9828 9832 9832
rect 9768 9772 9772 9828
rect 9772 9772 9828 9828
rect 9828 9772 9832 9828
rect 9768 9768 9832 9772
rect 9768 9608 9832 9672
rect 9768 9508 9832 9512
rect 9768 9452 9772 9508
rect 9772 9452 9828 9508
rect 9828 9452 9832 9508
rect 9768 9448 9832 9452
rect 9768 9348 9832 9352
rect 9768 9292 9772 9348
rect 9772 9292 9828 9348
rect 9828 9292 9832 9348
rect 9768 9288 9832 9292
rect 9768 9128 9832 9192
rect 9768 9028 9832 9032
rect 9768 8972 9772 9028
rect 9772 8972 9828 9028
rect 9828 8972 9832 9028
rect 9768 8968 9832 8972
rect 9768 8868 9832 8872
rect 9768 8812 9772 8868
rect 9772 8812 9828 8868
rect 9828 8812 9832 8868
rect 9768 8808 9832 8812
rect 9768 8708 9832 8712
rect 9768 8652 9772 8708
rect 9772 8652 9828 8708
rect 9828 8652 9832 8708
rect 9768 8648 9832 8652
rect 9768 8548 9832 8552
rect 9768 8492 9772 8548
rect 9772 8492 9828 8548
rect 9828 8492 9832 8548
rect 9768 8488 9832 8492
rect 9768 8388 9832 8392
rect 9768 8332 9772 8388
rect 9772 8332 9828 8388
rect 9828 8332 9832 8388
rect 9768 8328 9832 8332
rect 9768 8228 9832 8232
rect 9768 8172 9772 8228
rect 9772 8172 9828 8228
rect 9828 8172 9832 8228
rect 9768 8168 9832 8172
rect 9768 8068 9832 8072
rect 9768 8012 9772 8068
rect 9772 8012 9828 8068
rect 9828 8012 9832 8068
rect 9768 8008 9832 8012
rect 9768 7908 9832 7912
rect 9768 7852 9772 7908
rect 9772 7852 9828 7908
rect 9828 7852 9832 7908
rect 9768 7848 9832 7852
rect 9768 7748 9832 7752
rect 9768 7692 9772 7748
rect 9772 7692 9828 7748
rect 9828 7692 9832 7748
rect 9768 7688 9832 7692
rect 9768 7528 9832 7592
rect 9768 7428 9832 7432
rect 9768 7372 9772 7428
rect 9772 7372 9828 7428
rect 9828 7372 9832 7428
rect 9768 7368 9832 7372
rect 9768 7268 9832 7272
rect 9768 7212 9772 7268
rect 9772 7212 9828 7268
rect 9828 7212 9832 7268
rect 9768 7208 9832 7212
rect 9768 7048 9832 7112
rect 9768 6948 9832 6952
rect 9768 6892 9772 6948
rect 9772 6892 9828 6948
rect 9828 6892 9832 6948
rect 9768 6888 9832 6892
rect 9768 6788 9832 6792
rect 9768 6732 9772 6788
rect 9772 6732 9828 6788
rect 9828 6732 9832 6788
rect 9768 6728 9832 6732
rect 9768 6568 9832 6632
rect 9768 6468 9832 6472
rect 9768 6412 9772 6468
rect 9772 6412 9828 6468
rect 9828 6412 9832 6468
rect 9768 6408 9832 6412
rect 9768 6308 9832 6312
rect 9768 6252 9772 6308
rect 9772 6252 9828 6308
rect 9828 6252 9832 6308
rect 9768 6248 9832 6252
rect 9768 6148 9832 6152
rect 9768 6092 9772 6148
rect 9772 6092 9828 6148
rect 9828 6092 9832 6148
rect 9768 6088 9832 6092
rect 9768 5988 9832 5992
rect 9768 5932 9772 5988
rect 9772 5932 9828 5988
rect 9828 5932 9832 5988
rect 9768 5928 9832 5932
rect 9768 5828 9832 5832
rect 9768 5772 9772 5828
rect 9772 5772 9828 5828
rect 9828 5772 9832 5828
rect 9768 5768 9832 5772
rect 9768 5668 9832 5672
rect 9768 5612 9772 5668
rect 9772 5612 9828 5668
rect 9828 5612 9832 5668
rect 9768 5608 9832 5612
rect 9768 5508 9832 5512
rect 9768 5452 9772 5508
rect 9772 5452 9828 5508
rect 9828 5452 9832 5508
rect 9768 5448 9832 5452
rect 9768 5348 9832 5352
rect 9768 5292 9772 5348
rect 9772 5292 9828 5348
rect 9828 5292 9832 5348
rect 9768 5288 9832 5292
rect 9768 5188 9832 5192
rect 9768 5132 9772 5188
rect 9772 5132 9828 5188
rect 9828 5132 9832 5188
rect 9768 5128 9832 5132
rect 9768 5028 9832 5032
rect 9768 4972 9772 5028
rect 9772 4972 9828 5028
rect 9828 4972 9832 5028
rect 9768 4968 9832 4972
rect 9768 4868 9832 4872
rect 9768 4812 9772 4868
rect 9772 4812 9828 4868
rect 9828 4812 9832 4868
rect 9768 4808 9832 4812
rect 9768 4708 9832 4712
rect 9768 4652 9772 4708
rect 9772 4652 9828 4708
rect 9828 4652 9832 4708
rect 9768 4648 9832 4652
rect 9768 4548 9832 4552
rect 9768 4492 9772 4548
rect 9772 4492 9828 4548
rect 9828 4492 9832 4548
rect 9768 4488 9832 4492
rect 9768 4388 9832 4392
rect 9768 4332 9772 4388
rect 9772 4332 9828 4388
rect 9828 4332 9832 4388
rect 9768 4328 9832 4332
rect 9768 4228 9832 4232
rect 9768 4172 9772 4228
rect 9772 4172 9828 4228
rect 9828 4172 9832 4228
rect 9768 4168 9832 4172
rect 9768 4068 9832 4072
rect 9768 4012 9772 4068
rect 9772 4012 9828 4068
rect 9828 4012 9832 4068
rect 9768 4008 9832 4012
rect 9768 3908 9832 3912
rect 9768 3852 9772 3908
rect 9772 3852 9828 3908
rect 9828 3852 9832 3908
rect 9768 3848 9832 3852
rect 9768 3688 9832 3752
rect 9768 3528 9832 3592
rect 9768 3428 9832 3432
rect 9768 3372 9772 3428
rect 9772 3372 9828 3428
rect 9828 3372 9832 3428
rect 9768 3368 9832 3372
rect 9768 3268 9832 3272
rect 9768 3212 9772 3268
rect 9772 3212 9828 3268
rect 9828 3212 9832 3268
rect 9768 3208 9832 3212
rect 9768 3108 9832 3112
rect 9768 3052 9772 3108
rect 9772 3052 9828 3108
rect 9828 3052 9832 3108
rect 9768 3048 9832 3052
rect 9768 2948 9832 2952
rect 9768 2892 9772 2948
rect 9772 2892 9828 2948
rect 9828 2892 9832 2948
rect 9768 2888 9832 2892
rect 9768 2788 9832 2792
rect 9768 2732 9772 2788
rect 9772 2732 9828 2788
rect 9828 2732 9832 2788
rect 9768 2728 9832 2732
rect 9768 2628 9832 2632
rect 9768 2572 9772 2628
rect 9772 2572 9828 2628
rect 9828 2572 9832 2628
rect 9768 2568 9832 2572
rect 9768 2468 9832 2472
rect 9768 2412 9772 2468
rect 9772 2412 9828 2468
rect 9828 2412 9832 2468
rect 9768 2408 9832 2412
rect 9768 2308 9832 2312
rect 9768 2252 9772 2308
rect 9772 2252 9828 2308
rect 9828 2252 9832 2308
rect 9768 2248 9832 2252
rect 9768 2148 9832 2152
rect 9768 2092 9772 2148
rect 9772 2092 9828 2148
rect 9828 2092 9832 2148
rect 9768 2088 9832 2092
rect 9768 1988 9832 1992
rect 9768 1932 9772 1988
rect 9772 1932 9828 1988
rect 9828 1932 9832 1988
rect 9768 1928 9832 1932
rect 9768 1768 9832 1832
rect 9768 1668 9832 1672
rect 9768 1612 9772 1668
rect 9772 1612 9828 1668
rect 9828 1612 9832 1668
rect 9768 1608 9832 1612
rect 9768 1508 9832 1512
rect 9768 1452 9772 1508
rect 9772 1452 9828 1508
rect 9828 1452 9832 1508
rect 9768 1448 9832 1452
rect 9768 1348 9832 1352
rect 9768 1292 9772 1348
rect 9772 1292 9828 1348
rect 9828 1292 9832 1348
rect 9768 1288 9832 1292
rect 9768 1188 9832 1192
rect 9768 1132 9772 1188
rect 9772 1132 9828 1188
rect 9828 1132 9832 1188
rect 9768 1128 9832 1132
rect 9768 1028 9832 1032
rect 9768 972 9772 1028
rect 9772 972 9828 1028
rect 9828 972 9832 1028
rect 9768 968 9832 972
rect 9768 808 9832 872
rect 9768 648 9832 712
rect 9768 548 9832 552
rect 9768 492 9772 548
rect 9772 492 9828 548
rect 9828 492 9832 548
rect 9768 488 9832 492
rect 9768 388 9832 392
rect 9768 332 9772 388
rect 9772 332 9828 388
rect 9828 332 9832 388
rect 9768 328 9832 332
rect 9768 228 9832 232
rect 9768 172 9772 228
rect 9772 172 9828 228
rect 9828 172 9832 228
rect 9768 168 9832 172
rect 9768 68 9832 72
rect 9768 12 9772 68
rect 9772 12 9828 68
rect 9828 12 9832 68
rect 9768 8 9832 12
rect 9448 -1112 9512 -1048
rect 9448 -1192 9512 -1128
rect 9448 -1272 9512 -1208
rect 9448 -1352 9512 -1288
rect 9448 -1432 9512 -1368
rect 10088 31428 10152 31432
rect 10088 31372 10092 31428
rect 10092 31372 10148 31428
rect 10148 31372 10152 31428
rect 10088 31368 10152 31372
rect 10088 31268 10152 31272
rect 10088 31212 10092 31268
rect 10092 31212 10148 31268
rect 10148 31212 10152 31268
rect 10088 31208 10152 31212
rect 10088 31108 10152 31112
rect 10088 31052 10092 31108
rect 10092 31052 10148 31108
rect 10148 31052 10152 31108
rect 10088 31048 10152 31052
rect 10088 30948 10152 30952
rect 10088 30892 10092 30948
rect 10092 30892 10148 30948
rect 10148 30892 10152 30948
rect 10088 30888 10152 30892
rect 10088 30788 10152 30792
rect 10088 30732 10092 30788
rect 10092 30732 10148 30788
rect 10148 30732 10152 30788
rect 10088 30728 10152 30732
rect 10088 30628 10152 30632
rect 10088 30572 10092 30628
rect 10092 30572 10148 30628
rect 10148 30572 10152 30628
rect 10088 30568 10152 30572
rect 10088 30468 10152 30472
rect 10088 30412 10092 30468
rect 10092 30412 10148 30468
rect 10148 30412 10152 30468
rect 10088 30408 10152 30412
rect 10088 30308 10152 30312
rect 10088 30252 10092 30308
rect 10092 30252 10148 30308
rect 10148 30252 10152 30308
rect 10088 30248 10152 30252
rect 10088 30088 10152 30152
rect 10088 29988 10152 29992
rect 10088 29932 10092 29988
rect 10092 29932 10148 29988
rect 10148 29932 10152 29988
rect 10088 29928 10152 29932
rect 10088 29828 10152 29832
rect 10088 29772 10092 29828
rect 10092 29772 10148 29828
rect 10148 29772 10152 29828
rect 10088 29768 10152 29772
rect 10088 29668 10152 29672
rect 10088 29612 10092 29668
rect 10092 29612 10148 29668
rect 10148 29612 10152 29668
rect 10088 29608 10152 29612
rect 10088 29508 10152 29512
rect 10088 29452 10092 29508
rect 10092 29452 10148 29508
rect 10148 29452 10152 29508
rect 10088 29448 10152 29452
rect 10088 29348 10152 29352
rect 10088 29292 10092 29348
rect 10092 29292 10148 29348
rect 10148 29292 10152 29348
rect 10088 29288 10152 29292
rect 10088 29188 10152 29192
rect 10088 29132 10092 29188
rect 10092 29132 10148 29188
rect 10148 29132 10152 29188
rect 10088 29128 10152 29132
rect 10088 29028 10152 29032
rect 10088 28972 10092 29028
rect 10092 28972 10148 29028
rect 10148 28972 10152 29028
rect 10088 28968 10152 28972
rect 10088 28868 10152 28872
rect 10088 28812 10092 28868
rect 10092 28812 10148 28868
rect 10148 28812 10152 28868
rect 10088 28808 10152 28812
rect 10088 28648 10152 28712
rect 10088 28488 10152 28552
rect 10088 28328 10152 28392
rect 10088 28168 10152 28232
rect 10088 28068 10152 28072
rect 10088 28012 10092 28068
rect 10092 28012 10148 28068
rect 10148 28012 10152 28068
rect 10088 28008 10152 28012
rect 10088 27908 10152 27912
rect 10088 27852 10092 27908
rect 10092 27852 10148 27908
rect 10148 27852 10152 27908
rect 10088 27848 10152 27852
rect 10088 27748 10152 27752
rect 10088 27692 10092 27748
rect 10092 27692 10148 27748
rect 10148 27692 10152 27748
rect 10088 27688 10152 27692
rect 10088 27588 10152 27592
rect 10088 27532 10092 27588
rect 10092 27532 10148 27588
rect 10148 27532 10152 27588
rect 10088 27528 10152 27532
rect 10088 27428 10152 27432
rect 10088 27372 10092 27428
rect 10092 27372 10148 27428
rect 10148 27372 10152 27428
rect 10088 27368 10152 27372
rect 10088 27268 10152 27272
rect 10088 27212 10092 27268
rect 10092 27212 10148 27268
rect 10148 27212 10152 27268
rect 10088 27208 10152 27212
rect 10088 27108 10152 27112
rect 10088 27052 10092 27108
rect 10092 27052 10148 27108
rect 10148 27052 10152 27108
rect 10088 27048 10152 27052
rect 10088 26948 10152 26952
rect 10088 26892 10092 26948
rect 10092 26892 10148 26948
rect 10148 26892 10152 26948
rect 10088 26888 10152 26892
rect 10088 26728 10152 26792
rect 10088 26568 10152 26632
rect 10088 26408 10152 26472
rect 10088 26248 10152 26312
rect 10088 26148 10152 26152
rect 10088 26092 10092 26148
rect 10092 26092 10148 26148
rect 10148 26092 10152 26148
rect 10088 26088 10152 26092
rect 10088 25988 10152 25992
rect 10088 25932 10092 25988
rect 10092 25932 10148 25988
rect 10148 25932 10152 25988
rect 10088 25928 10152 25932
rect 10088 25828 10152 25832
rect 10088 25772 10092 25828
rect 10092 25772 10148 25828
rect 10148 25772 10152 25828
rect 10088 25768 10152 25772
rect 10088 25668 10152 25672
rect 10088 25612 10092 25668
rect 10092 25612 10148 25668
rect 10148 25612 10152 25668
rect 10088 25608 10152 25612
rect 10088 25508 10152 25512
rect 10088 25452 10092 25508
rect 10092 25452 10148 25508
rect 10148 25452 10152 25508
rect 10088 25448 10152 25452
rect 10088 25348 10152 25352
rect 10088 25292 10092 25348
rect 10092 25292 10148 25348
rect 10148 25292 10152 25348
rect 10088 25288 10152 25292
rect 10088 25188 10152 25192
rect 10088 25132 10092 25188
rect 10092 25132 10148 25188
rect 10148 25132 10152 25188
rect 10088 25128 10152 25132
rect 10088 25028 10152 25032
rect 10088 24972 10092 25028
rect 10092 24972 10148 25028
rect 10148 24972 10152 25028
rect 10088 24968 10152 24972
rect 10088 24808 10152 24872
rect 10088 24708 10152 24712
rect 10088 24652 10092 24708
rect 10092 24652 10148 24708
rect 10148 24652 10152 24708
rect 10088 24648 10152 24652
rect 10088 24548 10152 24552
rect 10088 24492 10092 24548
rect 10092 24492 10148 24548
rect 10148 24492 10152 24548
rect 10088 24488 10152 24492
rect 10088 24388 10152 24392
rect 10088 24332 10092 24388
rect 10092 24332 10148 24388
rect 10148 24332 10152 24388
rect 10088 24328 10152 24332
rect 10088 24228 10152 24232
rect 10088 24172 10092 24228
rect 10092 24172 10148 24228
rect 10148 24172 10152 24228
rect 10088 24168 10152 24172
rect 10088 24068 10152 24072
rect 10088 24012 10092 24068
rect 10092 24012 10148 24068
rect 10148 24012 10152 24068
rect 10088 24008 10152 24012
rect 10088 23908 10152 23912
rect 10088 23852 10092 23908
rect 10092 23852 10148 23908
rect 10148 23852 10152 23908
rect 10088 23848 10152 23852
rect 10088 23748 10152 23752
rect 10088 23692 10092 23748
rect 10092 23692 10148 23748
rect 10148 23692 10152 23748
rect 10088 23688 10152 23692
rect 10088 23588 10152 23592
rect 10088 23532 10092 23588
rect 10092 23532 10148 23588
rect 10148 23532 10152 23588
rect 10088 23528 10152 23532
rect 10088 23428 10152 23432
rect 10088 23372 10092 23428
rect 10092 23372 10148 23428
rect 10148 23372 10152 23428
rect 10088 23368 10152 23372
rect 10088 23268 10152 23272
rect 10088 23212 10092 23268
rect 10092 23212 10148 23268
rect 10148 23212 10152 23268
rect 10088 23208 10152 23212
rect 10088 23108 10152 23112
rect 10088 23052 10092 23108
rect 10092 23052 10148 23108
rect 10148 23052 10152 23108
rect 10088 23048 10152 23052
rect 10088 22948 10152 22952
rect 10088 22892 10092 22948
rect 10092 22892 10148 22948
rect 10148 22892 10152 22948
rect 10088 22888 10152 22892
rect 10088 22788 10152 22792
rect 10088 22732 10092 22788
rect 10092 22732 10148 22788
rect 10148 22732 10152 22788
rect 10088 22728 10152 22732
rect 10088 22628 10152 22632
rect 10088 22572 10092 22628
rect 10092 22572 10148 22628
rect 10148 22572 10152 22628
rect 10088 22568 10152 22572
rect 10088 22468 10152 22472
rect 10088 22412 10092 22468
rect 10092 22412 10148 22468
rect 10148 22412 10152 22468
rect 10088 22408 10152 22412
rect 10088 22308 10152 22312
rect 10088 22252 10092 22308
rect 10092 22252 10148 22308
rect 10148 22252 10152 22308
rect 10088 22248 10152 22252
rect 10088 22148 10152 22152
rect 10088 22092 10092 22148
rect 10092 22092 10148 22148
rect 10148 22092 10152 22148
rect 10088 22088 10152 22092
rect 10088 21928 10152 21992
rect 10088 21828 10152 21832
rect 10088 21772 10092 21828
rect 10092 21772 10148 21828
rect 10148 21772 10152 21828
rect 10088 21768 10152 21772
rect 10088 21668 10152 21672
rect 10088 21612 10092 21668
rect 10092 21612 10148 21668
rect 10148 21612 10152 21668
rect 10088 21608 10152 21612
rect 10088 21508 10152 21512
rect 10088 21452 10092 21508
rect 10092 21452 10148 21508
rect 10148 21452 10152 21508
rect 10088 21448 10152 21452
rect 10088 21348 10152 21352
rect 10088 21292 10092 21348
rect 10092 21292 10148 21348
rect 10148 21292 10152 21348
rect 10088 21288 10152 21292
rect 10088 21188 10152 21192
rect 10088 21132 10092 21188
rect 10092 21132 10148 21188
rect 10148 21132 10152 21188
rect 10088 21128 10152 21132
rect 10088 21028 10152 21032
rect 10088 20972 10092 21028
rect 10092 20972 10148 21028
rect 10148 20972 10152 21028
rect 10088 20968 10152 20972
rect 10088 20868 10152 20872
rect 10088 20812 10092 20868
rect 10092 20812 10148 20868
rect 10148 20812 10152 20868
rect 10088 20808 10152 20812
rect 10088 20708 10152 20712
rect 10088 20652 10092 20708
rect 10092 20652 10148 20708
rect 10148 20652 10152 20708
rect 10088 20648 10152 20652
rect 10088 20488 10152 20552
rect 10088 20328 10152 20392
rect 10088 20168 10152 20232
rect 10088 20008 10152 20072
rect 10088 19908 10152 19912
rect 10088 19852 10092 19908
rect 10092 19852 10148 19908
rect 10148 19852 10152 19908
rect 10088 19848 10152 19852
rect 10088 19748 10152 19752
rect 10088 19692 10092 19748
rect 10092 19692 10148 19748
rect 10148 19692 10152 19748
rect 10088 19688 10152 19692
rect 10088 19588 10152 19592
rect 10088 19532 10092 19588
rect 10092 19532 10148 19588
rect 10148 19532 10152 19588
rect 10088 19528 10152 19532
rect 10088 19428 10152 19432
rect 10088 19372 10092 19428
rect 10092 19372 10148 19428
rect 10148 19372 10152 19428
rect 10088 19368 10152 19372
rect 10088 19268 10152 19272
rect 10088 19212 10092 19268
rect 10092 19212 10148 19268
rect 10148 19212 10152 19268
rect 10088 19208 10152 19212
rect 10088 19108 10152 19112
rect 10088 19052 10092 19108
rect 10092 19052 10148 19108
rect 10148 19052 10152 19108
rect 10088 19048 10152 19052
rect 10088 18948 10152 18952
rect 10088 18892 10092 18948
rect 10092 18892 10148 18948
rect 10148 18892 10152 18948
rect 10088 18888 10152 18892
rect 10088 18788 10152 18792
rect 10088 18732 10092 18788
rect 10092 18732 10148 18788
rect 10148 18732 10152 18788
rect 10088 18728 10152 18732
rect 10088 18568 10152 18632
rect 10088 18408 10152 18472
rect 10088 18248 10152 18312
rect 10088 18088 10152 18152
rect 10088 17988 10152 17992
rect 10088 17932 10092 17988
rect 10092 17932 10148 17988
rect 10148 17932 10152 17988
rect 10088 17928 10152 17932
rect 10088 17828 10152 17832
rect 10088 17772 10092 17828
rect 10092 17772 10148 17828
rect 10148 17772 10152 17828
rect 10088 17768 10152 17772
rect 10088 17668 10152 17672
rect 10088 17612 10092 17668
rect 10092 17612 10148 17668
rect 10148 17612 10152 17668
rect 10088 17608 10152 17612
rect 10088 17508 10152 17512
rect 10088 17452 10092 17508
rect 10092 17452 10148 17508
rect 10148 17452 10152 17508
rect 10088 17448 10152 17452
rect 10088 17348 10152 17352
rect 10088 17292 10092 17348
rect 10092 17292 10148 17348
rect 10148 17292 10152 17348
rect 10088 17288 10152 17292
rect 10088 17188 10152 17192
rect 10088 17132 10092 17188
rect 10092 17132 10148 17188
rect 10148 17132 10152 17188
rect 10088 17128 10152 17132
rect 10088 17028 10152 17032
rect 10088 16972 10092 17028
rect 10092 16972 10148 17028
rect 10148 16972 10152 17028
rect 10088 16968 10152 16972
rect 10088 16868 10152 16872
rect 10088 16812 10092 16868
rect 10092 16812 10148 16868
rect 10148 16812 10152 16868
rect 10088 16808 10152 16812
rect 10088 16648 10152 16712
rect 10088 16548 10152 16552
rect 10088 16492 10092 16548
rect 10092 16492 10148 16548
rect 10148 16492 10152 16548
rect 10088 16488 10152 16492
rect 10088 16388 10152 16392
rect 10088 16332 10092 16388
rect 10092 16332 10148 16388
rect 10148 16332 10152 16388
rect 10088 16328 10152 16332
rect 10088 16228 10152 16232
rect 10088 16172 10092 16228
rect 10092 16172 10148 16228
rect 10148 16172 10152 16228
rect 10088 16168 10152 16172
rect 10088 16068 10152 16072
rect 10088 16012 10092 16068
rect 10092 16012 10148 16068
rect 10148 16012 10152 16068
rect 10088 16008 10152 16012
rect 10088 15908 10152 15912
rect 10088 15852 10092 15908
rect 10092 15852 10148 15908
rect 10148 15852 10152 15908
rect 10088 15848 10152 15852
rect 10088 15748 10152 15752
rect 10088 15692 10092 15748
rect 10092 15692 10148 15748
rect 10148 15692 10152 15748
rect 10088 15688 10152 15692
rect 10088 15588 10152 15592
rect 10088 15532 10092 15588
rect 10092 15532 10148 15588
rect 10148 15532 10152 15588
rect 10088 15528 10152 15532
rect 10088 15428 10152 15432
rect 10088 15372 10092 15428
rect 10092 15372 10148 15428
rect 10148 15372 10152 15428
rect 10088 15368 10152 15372
rect 10088 15268 10152 15272
rect 10088 15212 10092 15268
rect 10092 15212 10148 15268
rect 10148 15212 10152 15268
rect 10088 15208 10152 15212
rect 10088 15108 10152 15112
rect 10088 15052 10092 15108
rect 10092 15052 10148 15108
rect 10148 15052 10152 15108
rect 10088 15048 10152 15052
rect 10088 14948 10152 14952
rect 10088 14892 10092 14948
rect 10092 14892 10148 14948
rect 10148 14892 10152 14948
rect 10088 14888 10152 14892
rect 10088 14788 10152 14792
rect 10088 14732 10092 14788
rect 10092 14732 10148 14788
rect 10148 14732 10152 14788
rect 10088 14728 10152 14732
rect 10088 14628 10152 14632
rect 10088 14572 10092 14628
rect 10092 14572 10148 14628
rect 10148 14572 10152 14628
rect 10088 14568 10152 14572
rect 10088 14468 10152 14472
rect 10088 14412 10092 14468
rect 10092 14412 10148 14468
rect 10148 14412 10152 14468
rect 10088 14408 10152 14412
rect 10088 14308 10152 14312
rect 10088 14252 10092 14308
rect 10092 14252 10148 14308
rect 10148 14252 10152 14308
rect 10088 14248 10152 14252
rect 10088 14148 10152 14152
rect 10088 14092 10092 14148
rect 10092 14092 10148 14148
rect 10148 14092 10152 14148
rect 10088 14088 10152 14092
rect 10088 13988 10152 13992
rect 10088 13932 10092 13988
rect 10092 13932 10148 13988
rect 10148 13932 10152 13988
rect 10088 13928 10152 13932
rect 10088 13768 10152 13832
rect 10088 13668 10152 13672
rect 10088 13612 10092 13668
rect 10092 13612 10148 13668
rect 10148 13612 10152 13668
rect 10088 13608 10152 13612
rect 10088 13508 10152 13512
rect 10088 13452 10092 13508
rect 10092 13452 10148 13508
rect 10148 13452 10152 13508
rect 10088 13448 10152 13452
rect 10088 13348 10152 13352
rect 10088 13292 10092 13348
rect 10092 13292 10148 13348
rect 10148 13292 10152 13348
rect 10088 13288 10152 13292
rect 10088 13188 10152 13192
rect 10088 13132 10092 13188
rect 10092 13132 10148 13188
rect 10148 13132 10152 13188
rect 10088 13128 10152 13132
rect 10088 13028 10152 13032
rect 10088 12972 10092 13028
rect 10092 12972 10148 13028
rect 10148 12972 10152 13028
rect 10088 12968 10152 12972
rect 10088 12868 10152 12872
rect 10088 12812 10092 12868
rect 10092 12812 10148 12868
rect 10148 12812 10152 12868
rect 10088 12808 10152 12812
rect 10088 12708 10152 12712
rect 10088 12652 10092 12708
rect 10092 12652 10148 12708
rect 10148 12652 10152 12708
rect 10088 12648 10152 12652
rect 10088 12548 10152 12552
rect 10088 12492 10092 12548
rect 10092 12492 10148 12548
rect 10148 12492 10152 12548
rect 10088 12488 10152 12492
rect 10088 12328 10152 12392
rect 10088 12168 10152 12232
rect 10088 12008 10152 12072
rect 10088 11848 10152 11912
rect 10088 11748 10152 11752
rect 10088 11692 10092 11748
rect 10092 11692 10148 11748
rect 10148 11692 10152 11748
rect 10088 11688 10152 11692
rect 10088 11588 10152 11592
rect 10088 11532 10092 11588
rect 10092 11532 10148 11588
rect 10148 11532 10152 11588
rect 10088 11528 10152 11532
rect 10088 11428 10152 11432
rect 10088 11372 10092 11428
rect 10092 11372 10148 11428
rect 10148 11372 10152 11428
rect 10088 11368 10152 11372
rect 10088 11268 10152 11272
rect 10088 11212 10092 11268
rect 10092 11212 10148 11268
rect 10148 11212 10152 11268
rect 10088 11208 10152 11212
rect 10088 11108 10152 11112
rect 10088 11052 10092 11108
rect 10092 11052 10148 11108
rect 10148 11052 10152 11108
rect 10088 11048 10152 11052
rect 10088 10948 10152 10952
rect 10088 10892 10092 10948
rect 10092 10892 10148 10948
rect 10148 10892 10152 10948
rect 10088 10888 10152 10892
rect 10088 10788 10152 10792
rect 10088 10732 10092 10788
rect 10092 10732 10148 10788
rect 10148 10732 10152 10788
rect 10088 10728 10152 10732
rect 10088 10628 10152 10632
rect 10088 10572 10092 10628
rect 10092 10572 10148 10628
rect 10148 10572 10152 10628
rect 10088 10568 10152 10572
rect 10088 10468 10152 10472
rect 10088 10412 10092 10468
rect 10092 10412 10148 10468
rect 10148 10412 10152 10468
rect 10088 10408 10152 10412
rect 10088 10308 10152 10312
rect 10088 10252 10092 10308
rect 10092 10252 10148 10308
rect 10148 10252 10152 10308
rect 10088 10248 10152 10252
rect 10088 10148 10152 10152
rect 10088 10092 10092 10148
rect 10092 10092 10148 10148
rect 10148 10092 10152 10148
rect 10088 10088 10152 10092
rect 10088 9988 10152 9992
rect 10088 9932 10092 9988
rect 10092 9932 10148 9988
rect 10148 9932 10152 9988
rect 10088 9928 10152 9932
rect 10088 9828 10152 9832
rect 10088 9772 10092 9828
rect 10092 9772 10148 9828
rect 10148 9772 10152 9828
rect 10088 9768 10152 9772
rect 10088 9608 10152 9672
rect 10088 9508 10152 9512
rect 10088 9452 10092 9508
rect 10092 9452 10148 9508
rect 10148 9452 10152 9508
rect 10088 9448 10152 9452
rect 10088 9348 10152 9352
rect 10088 9292 10092 9348
rect 10092 9292 10148 9348
rect 10148 9292 10152 9348
rect 10088 9288 10152 9292
rect 10088 9128 10152 9192
rect 10088 9028 10152 9032
rect 10088 8972 10092 9028
rect 10092 8972 10148 9028
rect 10148 8972 10152 9028
rect 10088 8968 10152 8972
rect 10088 8868 10152 8872
rect 10088 8812 10092 8868
rect 10092 8812 10148 8868
rect 10148 8812 10152 8868
rect 10088 8808 10152 8812
rect 10088 8708 10152 8712
rect 10088 8652 10092 8708
rect 10092 8652 10148 8708
rect 10148 8652 10152 8708
rect 10088 8648 10152 8652
rect 10088 8548 10152 8552
rect 10088 8492 10092 8548
rect 10092 8492 10148 8548
rect 10148 8492 10152 8548
rect 10088 8488 10152 8492
rect 10088 8388 10152 8392
rect 10088 8332 10092 8388
rect 10092 8332 10148 8388
rect 10148 8332 10152 8388
rect 10088 8328 10152 8332
rect 10088 8228 10152 8232
rect 10088 8172 10092 8228
rect 10092 8172 10148 8228
rect 10148 8172 10152 8228
rect 10088 8168 10152 8172
rect 10088 8068 10152 8072
rect 10088 8012 10092 8068
rect 10092 8012 10148 8068
rect 10148 8012 10152 8068
rect 10088 8008 10152 8012
rect 10088 7908 10152 7912
rect 10088 7852 10092 7908
rect 10092 7852 10148 7908
rect 10148 7852 10152 7908
rect 10088 7848 10152 7852
rect 10088 7748 10152 7752
rect 10088 7692 10092 7748
rect 10092 7692 10148 7748
rect 10148 7692 10152 7748
rect 10088 7688 10152 7692
rect 10088 7528 10152 7592
rect 10088 7428 10152 7432
rect 10088 7372 10092 7428
rect 10092 7372 10148 7428
rect 10148 7372 10152 7428
rect 10088 7368 10152 7372
rect 10088 7268 10152 7272
rect 10088 7212 10092 7268
rect 10092 7212 10148 7268
rect 10148 7212 10152 7268
rect 10088 7208 10152 7212
rect 10088 7048 10152 7112
rect 10088 6948 10152 6952
rect 10088 6892 10092 6948
rect 10092 6892 10148 6948
rect 10148 6892 10152 6948
rect 10088 6888 10152 6892
rect 10088 6788 10152 6792
rect 10088 6732 10092 6788
rect 10092 6732 10148 6788
rect 10148 6732 10152 6788
rect 10088 6728 10152 6732
rect 10088 6568 10152 6632
rect 10088 6468 10152 6472
rect 10088 6412 10092 6468
rect 10092 6412 10148 6468
rect 10148 6412 10152 6468
rect 10088 6408 10152 6412
rect 10088 6308 10152 6312
rect 10088 6252 10092 6308
rect 10092 6252 10148 6308
rect 10148 6252 10152 6308
rect 10088 6248 10152 6252
rect 10088 6148 10152 6152
rect 10088 6092 10092 6148
rect 10092 6092 10148 6148
rect 10148 6092 10152 6148
rect 10088 6088 10152 6092
rect 10088 5988 10152 5992
rect 10088 5932 10092 5988
rect 10092 5932 10148 5988
rect 10148 5932 10152 5988
rect 10088 5928 10152 5932
rect 10088 5828 10152 5832
rect 10088 5772 10092 5828
rect 10092 5772 10148 5828
rect 10148 5772 10152 5828
rect 10088 5768 10152 5772
rect 10088 5668 10152 5672
rect 10088 5612 10092 5668
rect 10092 5612 10148 5668
rect 10148 5612 10152 5668
rect 10088 5608 10152 5612
rect 10088 5508 10152 5512
rect 10088 5452 10092 5508
rect 10092 5452 10148 5508
rect 10148 5452 10152 5508
rect 10088 5448 10152 5452
rect 10088 5348 10152 5352
rect 10088 5292 10092 5348
rect 10092 5292 10148 5348
rect 10148 5292 10152 5348
rect 10088 5288 10152 5292
rect 10088 5188 10152 5192
rect 10088 5132 10092 5188
rect 10092 5132 10148 5188
rect 10148 5132 10152 5188
rect 10088 5128 10152 5132
rect 10088 5028 10152 5032
rect 10088 4972 10092 5028
rect 10092 4972 10148 5028
rect 10148 4972 10152 5028
rect 10088 4968 10152 4972
rect 10088 4868 10152 4872
rect 10088 4812 10092 4868
rect 10092 4812 10148 4868
rect 10148 4812 10152 4868
rect 10088 4808 10152 4812
rect 10088 4708 10152 4712
rect 10088 4652 10092 4708
rect 10092 4652 10148 4708
rect 10148 4652 10152 4708
rect 10088 4648 10152 4652
rect 10088 4548 10152 4552
rect 10088 4492 10092 4548
rect 10092 4492 10148 4548
rect 10148 4492 10152 4548
rect 10088 4488 10152 4492
rect 10088 4388 10152 4392
rect 10088 4332 10092 4388
rect 10092 4332 10148 4388
rect 10148 4332 10152 4388
rect 10088 4328 10152 4332
rect 10088 4228 10152 4232
rect 10088 4172 10092 4228
rect 10092 4172 10148 4228
rect 10148 4172 10152 4228
rect 10088 4168 10152 4172
rect 10088 4068 10152 4072
rect 10088 4012 10092 4068
rect 10092 4012 10148 4068
rect 10148 4012 10152 4068
rect 10088 4008 10152 4012
rect 10088 3908 10152 3912
rect 10088 3852 10092 3908
rect 10092 3852 10148 3908
rect 10148 3852 10152 3908
rect 10088 3848 10152 3852
rect 10088 3688 10152 3752
rect 10088 3528 10152 3592
rect 10088 3428 10152 3432
rect 10088 3372 10092 3428
rect 10092 3372 10148 3428
rect 10148 3372 10152 3428
rect 10088 3368 10152 3372
rect 10088 3268 10152 3272
rect 10088 3212 10092 3268
rect 10092 3212 10148 3268
rect 10148 3212 10152 3268
rect 10088 3208 10152 3212
rect 10088 3108 10152 3112
rect 10088 3052 10092 3108
rect 10092 3052 10148 3108
rect 10148 3052 10152 3108
rect 10088 3048 10152 3052
rect 10088 2948 10152 2952
rect 10088 2892 10092 2948
rect 10092 2892 10148 2948
rect 10148 2892 10152 2948
rect 10088 2888 10152 2892
rect 10088 2788 10152 2792
rect 10088 2732 10092 2788
rect 10092 2732 10148 2788
rect 10148 2732 10152 2788
rect 10088 2728 10152 2732
rect 10088 2628 10152 2632
rect 10088 2572 10092 2628
rect 10092 2572 10148 2628
rect 10148 2572 10152 2628
rect 10088 2568 10152 2572
rect 10088 2468 10152 2472
rect 10088 2412 10092 2468
rect 10092 2412 10148 2468
rect 10148 2412 10152 2468
rect 10088 2408 10152 2412
rect 10088 2308 10152 2312
rect 10088 2252 10092 2308
rect 10092 2252 10148 2308
rect 10148 2252 10152 2308
rect 10088 2248 10152 2252
rect 10088 2148 10152 2152
rect 10088 2092 10092 2148
rect 10092 2092 10148 2148
rect 10148 2092 10152 2148
rect 10088 2088 10152 2092
rect 10088 1988 10152 1992
rect 10088 1932 10092 1988
rect 10092 1932 10148 1988
rect 10148 1932 10152 1988
rect 10088 1928 10152 1932
rect 10088 1768 10152 1832
rect 10088 1668 10152 1672
rect 10088 1612 10092 1668
rect 10092 1612 10148 1668
rect 10148 1612 10152 1668
rect 10088 1608 10152 1612
rect 10088 1508 10152 1512
rect 10088 1452 10092 1508
rect 10092 1452 10148 1508
rect 10148 1452 10152 1508
rect 10088 1448 10152 1452
rect 10088 1348 10152 1352
rect 10088 1292 10092 1348
rect 10092 1292 10148 1348
rect 10148 1292 10152 1348
rect 10088 1288 10152 1292
rect 10088 1188 10152 1192
rect 10088 1132 10092 1188
rect 10092 1132 10148 1188
rect 10148 1132 10152 1188
rect 10088 1128 10152 1132
rect 10088 1028 10152 1032
rect 10088 972 10092 1028
rect 10092 972 10148 1028
rect 10148 972 10152 1028
rect 10088 968 10152 972
rect 10088 808 10152 872
rect 10088 648 10152 712
rect 10088 548 10152 552
rect 10088 492 10092 548
rect 10092 492 10148 548
rect 10148 492 10152 548
rect 10088 488 10152 492
rect 10088 388 10152 392
rect 10088 332 10092 388
rect 10092 332 10148 388
rect 10148 332 10152 388
rect 10088 328 10152 332
rect 10088 228 10152 232
rect 10088 172 10092 228
rect 10092 172 10148 228
rect 10148 172 10152 228
rect 10088 168 10152 172
rect 10088 68 10152 72
rect 10088 12 10092 68
rect 10092 12 10148 68
rect 10148 12 10152 68
rect 10088 8 10152 12
rect 9768 -1112 9832 -1048
rect 9768 -1192 9832 -1128
rect 9768 -1272 9832 -1208
rect 9768 -1352 9832 -1288
rect 9768 -1432 9832 -1368
rect 10408 31428 10472 31432
rect 10408 31372 10412 31428
rect 10412 31372 10468 31428
rect 10468 31372 10472 31428
rect 10408 31368 10472 31372
rect 10408 31268 10472 31272
rect 10408 31212 10412 31268
rect 10412 31212 10468 31268
rect 10468 31212 10472 31268
rect 10408 31208 10472 31212
rect 10408 31108 10472 31112
rect 10408 31052 10412 31108
rect 10412 31052 10468 31108
rect 10468 31052 10472 31108
rect 10408 31048 10472 31052
rect 10408 30948 10472 30952
rect 10408 30892 10412 30948
rect 10412 30892 10468 30948
rect 10468 30892 10472 30948
rect 10408 30888 10472 30892
rect 10408 30788 10472 30792
rect 10408 30732 10412 30788
rect 10412 30732 10468 30788
rect 10468 30732 10472 30788
rect 10408 30728 10472 30732
rect 10408 30628 10472 30632
rect 10408 30572 10412 30628
rect 10412 30572 10468 30628
rect 10468 30572 10472 30628
rect 10408 30568 10472 30572
rect 10408 30468 10472 30472
rect 10408 30412 10412 30468
rect 10412 30412 10468 30468
rect 10468 30412 10472 30468
rect 10408 30408 10472 30412
rect 10408 30308 10472 30312
rect 10408 30252 10412 30308
rect 10412 30252 10468 30308
rect 10468 30252 10472 30308
rect 10408 30248 10472 30252
rect 10408 30088 10472 30152
rect 10408 29988 10472 29992
rect 10408 29932 10412 29988
rect 10412 29932 10468 29988
rect 10468 29932 10472 29988
rect 10408 29928 10472 29932
rect 10408 29828 10472 29832
rect 10408 29772 10412 29828
rect 10412 29772 10468 29828
rect 10468 29772 10472 29828
rect 10408 29768 10472 29772
rect 10408 29668 10472 29672
rect 10408 29612 10412 29668
rect 10412 29612 10468 29668
rect 10468 29612 10472 29668
rect 10408 29608 10472 29612
rect 10408 29508 10472 29512
rect 10408 29452 10412 29508
rect 10412 29452 10468 29508
rect 10468 29452 10472 29508
rect 10408 29448 10472 29452
rect 10408 29348 10472 29352
rect 10408 29292 10412 29348
rect 10412 29292 10468 29348
rect 10468 29292 10472 29348
rect 10408 29288 10472 29292
rect 10408 29188 10472 29192
rect 10408 29132 10412 29188
rect 10412 29132 10468 29188
rect 10468 29132 10472 29188
rect 10408 29128 10472 29132
rect 10408 29028 10472 29032
rect 10408 28972 10412 29028
rect 10412 28972 10468 29028
rect 10468 28972 10472 29028
rect 10408 28968 10472 28972
rect 10408 28868 10472 28872
rect 10408 28812 10412 28868
rect 10412 28812 10468 28868
rect 10468 28812 10472 28868
rect 10408 28808 10472 28812
rect 10408 28648 10472 28712
rect 10408 28488 10472 28552
rect 10408 28328 10472 28392
rect 10408 28168 10472 28232
rect 10408 28068 10472 28072
rect 10408 28012 10412 28068
rect 10412 28012 10468 28068
rect 10468 28012 10472 28068
rect 10408 28008 10472 28012
rect 10408 27908 10472 27912
rect 10408 27852 10412 27908
rect 10412 27852 10468 27908
rect 10468 27852 10472 27908
rect 10408 27848 10472 27852
rect 10408 27748 10472 27752
rect 10408 27692 10412 27748
rect 10412 27692 10468 27748
rect 10468 27692 10472 27748
rect 10408 27688 10472 27692
rect 10408 27588 10472 27592
rect 10408 27532 10412 27588
rect 10412 27532 10468 27588
rect 10468 27532 10472 27588
rect 10408 27528 10472 27532
rect 10408 27428 10472 27432
rect 10408 27372 10412 27428
rect 10412 27372 10468 27428
rect 10468 27372 10472 27428
rect 10408 27368 10472 27372
rect 10408 27268 10472 27272
rect 10408 27212 10412 27268
rect 10412 27212 10468 27268
rect 10468 27212 10472 27268
rect 10408 27208 10472 27212
rect 10408 27108 10472 27112
rect 10408 27052 10412 27108
rect 10412 27052 10468 27108
rect 10468 27052 10472 27108
rect 10408 27048 10472 27052
rect 10408 26948 10472 26952
rect 10408 26892 10412 26948
rect 10412 26892 10468 26948
rect 10468 26892 10472 26948
rect 10408 26888 10472 26892
rect 10408 26728 10472 26792
rect 10408 26568 10472 26632
rect 10408 26408 10472 26472
rect 10408 26248 10472 26312
rect 10408 26148 10472 26152
rect 10408 26092 10412 26148
rect 10412 26092 10468 26148
rect 10468 26092 10472 26148
rect 10408 26088 10472 26092
rect 10408 25988 10472 25992
rect 10408 25932 10412 25988
rect 10412 25932 10468 25988
rect 10468 25932 10472 25988
rect 10408 25928 10472 25932
rect 10408 25828 10472 25832
rect 10408 25772 10412 25828
rect 10412 25772 10468 25828
rect 10468 25772 10472 25828
rect 10408 25768 10472 25772
rect 10408 25668 10472 25672
rect 10408 25612 10412 25668
rect 10412 25612 10468 25668
rect 10468 25612 10472 25668
rect 10408 25608 10472 25612
rect 10408 25508 10472 25512
rect 10408 25452 10412 25508
rect 10412 25452 10468 25508
rect 10468 25452 10472 25508
rect 10408 25448 10472 25452
rect 10408 25348 10472 25352
rect 10408 25292 10412 25348
rect 10412 25292 10468 25348
rect 10468 25292 10472 25348
rect 10408 25288 10472 25292
rect 10408 25188 10472 25192
rect 10408 25132 10412 25188
rect 10412 25132 10468 25188
rect 10468 25132 10472 25188
rect 10408 25128 10472 25132
rect 10408 25028 10472 25032
rect 10408 24972 10412 25028
rect 10412 24972 10468 25028
rect 10468 24972 10472 25028
rect 10408 24968 10472 24972
rect 10408 24808 10472 24872
rect 10408 24708 10472 24712
rect 10408 24652 10412 24708
rect 10412 24652 10468 24708
rect 10468 24652 10472 24708
rect 10408 24648 10472 24652
rect 10408 24548 10472 24552
rect 10408 24492 10412 24548
rect 10412 24492 10468 24548
rect 10468 24492 10472 24548
rect 10408 24488 10472 24492
rect 10408 24388 10472 24392
rect 10408 24332 10412 24388
rect 10412 24332 10468 24388
rect 10468 24332 10472 24388
rect 10408 24328 10472 24332
rect 10408 24228 10472 24232
rect 10408 24172 10412 24228
rect 10412 24172 10468 24228
rect 10468 24172 10472 24228
rect 10408 24168 10472 24172
rect 10408 24068 10472 24072
rect 10408 24012 10412 24068
rect 10412 24012 10468 24068
rect 10468 24012 10472 24068
rect 10408 24008 10472 24012
rect 10408 23908 10472 23912
rect 10408 23852 10412 23908
rect 10412 23852 10468 23908
rect 10468 23852 10472 23908
rect 10408 23848 10472 23852
rect 10408 23748 10472 23752
rect 10408 23692 10412 23748
rect 10412 23692 10468 23748
rect 10468 23692 10472 23748
rect 10408 23688 10472 23692
rect 10408 23588 10472 23592
rect 10408 23532 10412 23588
rect 10412 23532 10468 23588
rect 10468 23532 10472 23588
rect 10408 23528 10472 23532
rect 10408 23428 10472 23432
rect 10408 23372 10412 23428
rect 10412 23372 10468 23428
rect 10468 23372 10472 23428
rect 10408 23368 10472 23372
rect 10408 23268 10472 23272
rect 10408 23212 10412 23268
rect 10412 23212 10468 23268
rect 10468 23212 10472 23268
rect 10408 23208 10472 23212
rect 10408 23108 10472 23112
rect 10408 23052 10412 23108
rect 10412 23052 10468 23108
rect 10468 23052 10472 23108
rect 10408 23048 10472 23052
rect 10408 22948 10472 22952
rect 10408 22892 10412 22948
rect 10412 22892 10468 22948
rect 10468 22892 10472 22948
rect 10408 22888 10472 22892
rect 10408 22788 10472 22792
rect 10408 22732 10412 22788
rect 10412 22732 10468 22788
rect 10468 22732 10472 22788
rect 10408 22728 10472 22732
rect 10408 22628 10472 22632
rect 10408 22572 10412 22628
rect 10412 22572 10468 22628
rect 10468 22572 10472 22628
rect 10408 22568 10472 22572
rect 10408 22468 10472 22472
rect 10408 22412 10412 22468
rect 10412 22412 10468 22468
rect 10468 22412 10472 22468
rect 10408 22408 10472 22412
rect 10408 22308 10472 22312
rect 10408 22252 10412 22308
rect 10412 22252 10468 22308
rect 10468 22252 10472 22308
rect 10408 22248 10472 22252
rect 10408 22148 10472 22152
rect 10408 22092 10412 22148
rect 10412 22092 10468 22148
rect 10468 22092 10472 22148
rect 10408 22088 10472 22092
rect 10408 21928 10472 21992
rect 10408 21828 10472 21832
rect 10408 21772 10412 21828
rect 10412 21772 10468 21828
rect 10468 21772 10472 21828
rect 10408 21768 10472 21772
rect 10408 21668 10472 21672
rect 10408 21612 10412 21668
rect 10412 21612 10468 21668
rect 10468 21612 10472 21668
rect 10408 21608 10472 21612
rect 10408 21508 10472 21512
rect 10408 21452 10412 21508
rect 10412 21452 10468 21508
rect 10468 21452 10472 21508
rect 10408 21448 10472 21452
rect 10408 21348 10472 21352
rect 10408 21292 10412 21348
rect 10412 21292 10468 21348
rect 10468 21292 10472 21348
rect 10408 21288 10472 21292
rect 10408 21188 10472 21192
rect 10408 21132 10412 21188
rect 10412 21132 10468 21188
rect 10468 21132 10472 21188
rect 10408 21128 10472 21132
rect 10408 21028 10472 21032
rect 10408 20972 10412 21028
rect 10412 20972 10468 21028
rect 10468 20972 10472 21028
rect 10408 20968 10472 20972
rect 10408 20868 10472 20872
rect 10408 20812 10412 20868
rect 10412 20812 10468 20868
rect 10468 20812 10472 20868
rect 10408 20808 10472 20812
rect 10408 20708 10472 20712
rect 10408 20652 10412 20708
rect 10412 20652 10468 20708
rect 10468 20652 10472 20708
rect 10408 20648 10472 20652
rect 10408 20488 10472 20552
rect 10408 20328 10472 20392
rect 10408 20168 10472 20232
rect 10408 20008 10472 20072
rect 10408 19908 10472 19912
rect 10408 19852 10412 19908
rect 10412 19852 10468 19908
rect 10468 19852 10472 19908
rect 10408 19848 10472 19852
rect 10408 19748 10472 19752
rect 10408 19692 10412 19748
rect 10412 19692 10468 19748
rect 10468 19692 10472 19748
rect 10408 19688 10472 19692
rect 10408 19588 10472 19592
rect 10408 19532 10412 19588
rect 10412 19532 10468 19588
rect 10468 19532 10472 19588
rect 10408 19528 10472 19532
rect 10408 19428 10472 19432
rect 10408 19372 10412 19428
rect 10412 19372 10468 19428
rect 10468 19372 10472 19428
rect 10408 19368 10472 19372
rect 10408 19268 10472 19272
rect 10408 19212 10412 19268
rect 10412 19212 10468 19268
rect 10468 19212 10472 19268
rect 10408 19208 10472 19212
rect 10408 19108 10472 19112
rect 10408 19052 10412 19108
rect 10412 19052 10468 19108
rect 10468 19052 10472 19108
rect 10408 19048 10472 19052
rect 10408 18948 10472 18952
rect 10408 18892 10412 18948
rect 10412 18892 10468 18948
rect 10468 18892 10472 18948
rect 10408 18888 10472 18892
rect 10408 18788 10472 18792
rect 10408 18732 10412 18788
rect 10412 18732 10468 18788
rect 10468 18732 10472 18788
rect 10408 18728 10472 18732
rect 10408 18568 10472 18632
rect 10408 18408 10472 18472
rect 10408 18248 10472 18312
rect 10408 18088 10472 18152
rect 10408 17988 10472 17992
rect 10408 17932 10412 17988
rect 10412 17932 10468 17988
rect 10468 17932 10472 17988
rect 10408 17928 10472 17932
rect 10408 17828 10472 17832
rect 10408 17772 10412 17828
rect 10412 17772 10468 17828
rect 10468 17772 10472 17828
rect 10408 17768 10472 17772
rect 10408 17668 10472 17672
rect 10408 17612 10412 17668
rect 10412 17612 10468 17668
rect 10468 17612 10472 17668
rect 10408 17608 10472 17612
rect 10408 17508 10472 17512
rect 10408 17452 10412 17508
rect 10412 17452 10468 17508
rect 10468 17452 10472 17508
rect 10408 17448 10472 17452
rect 10408 17348 10472 17352
rect 10408 17292 10412 17348
rect 10412 17292 10468 17348
rect 10468 17292 10472 17348
rect 10408 17288 10472 17292
rect 10408 17188 10472 17192
rect 10408 17132 10412 17188
rect 10412 17132 10468 17188
rect 10468 17132 10472 17188
rect 10408 17128 10472 17132
rect 10408 17028 10472 17032
rect 10408 16972 10412 17028
rect 10412 16972 10468 17028
rect 10468 16972 10472 17028
rect 10408 16968 10472 16972
rect 10408 16868 10472 16872
rect 10408 16812 10412 16868
rect 10412 16812 10468 16868
rect 10468 16812 10472 16868
rect 10408 16808 10472 16812
rect 10408 16648 10472 16712
rect 10408 16548 10472 16552
rect 10408 16492 10412 16548
rect 10412 16492 10468 16548
rect 10468 16492 10472 16548
rect 10408 16488 10472 16492
rect 10408 16388 10472 16392
rect 10408 16332 10412 16388
rect 10412 16332 10468 16388
rect 10468 16332 10472 16388
rect 10408 16328 10472 16332
rect 10408 16228 10472 16232
rect 10408 16172 10412 16228
rect 10412 16172 10468 16228
rect 10468 16172 10472 16228
rect 10408 16168 10472 16172
rect 10408 16068 10472 16072
rect 10408 16012 10412 16068
rect 10412 16012 10468 16068
rect 10468 16012 10472 16068
rect 10408 16008 10472 16012
rect 10408 15908 10472 15912
rect 10408 15852 10412 15908
rect 10412 15852 10468 15908
rect 10468 15852 10472 15908
rect 10408 15848 10472 15852
rect 10408 15748 10472 15752
rect 10408 15692 10412 15748
rect 10412 15692 10468 15748
rect 10468 15692 10472 15748
rect 10408 15688 10472 15692
rect 10408 15588 10472 15592
rect 10408 15532 10412 15588
rect 10412 15532 10468 15588
rect 10468 15532 10472 15588
rect 10408 15528 10472 15532
rect 10408 15428 10472 15432
rect 10408 15372 10412 15428
rect 10412 15372 10468 15428
rect 10468 15372 10472 15428
rect 10408 15368 10472 15372
rect 10408 15268 10472 15272
rect 10408 15212 10412 15268
rect 10412 15212 10468 15268
rect 10468 15212 10472 15268
rect 10408 15208 10472 15212
rect 10408 15108 10472 15112
rect 10408 15052 10412 15108
rect 10412 15052 10468 15108
rect 10468 15052 10472 15108
rect 10408 15048 10472 15052
rect 10408 14948 10472 14952
rect 10408 14892 10412 14948
rect 10412 14892 10468 14948
rect 10468 14892 10472 14948
rect 10408 14888 10472 14892
rect 10408 14788 10472 14792
rect 10408 14732 10412 14788
rect 10412 14732 10468 14788
rect 10468 14732 10472 14788
rect 10408 14728 10472 14732
rect 10408 14628 10472 14632
rect 10408 14572 10412 14628
rect 10412 14572 10468 14628
rect 10468 14572 10472 14628
rect 10408 14568 10472 14572
rect 10408 14468 10472 14472
rect 10408 14412 10412 14468
rect 10412 14412 10468 14468
rect 10468 14412 10472 14468
rect 10408 14408 10472 14412
rect 10408 14308 10472 14312
rect 10408 14252 10412 14308
rect 10412 14252 10468 14308
rect 10468 14252 10472 14308
rect 10408 14248 10472 14252
rect 10408 14148 10472 14152
rect 10408 14092 10412 14148
rect 10412 14092 10468 14148
rect 10468 14092 10472 14148
rect 10408 14088 10472 14092
rect 10408 13988 10472 13992
rect 10408 13932 10412 13988
rect 10412 13932 10468 13988
rect 10468 13932 10472 13988
rect 10408 13928 10472 13932
rect 10408 13768 10472 13832
rect 10408 13668 10472 13672
rect 10408 13612 10412 13668
rect 10412 13612 10468 13668
rect 10468 13612 10472 13668
rect 10408 13608 10472 13612
rect 10408 13508 10472 13512
rect 10408 13452 10412 13508
rect 10412 13452 10468 13508
rect 10468 13452 10472 13508
rect 10408 13448 10472 13452
rect 10408 13348 10472 13352
rect 10408 13292 10412 13348
rect 10412 13292 10468 13348
rect 10468 13292 10472 13348
rect 10408 13288 10472 13292
rect 10408 13188 10472 13192
rect 10408 13132 10412 13188
rect 10412 13132 10468 13188
rect 10468 13132 10472 13188
rect 10408 13128 10472 13132
rect 10408 13028 10472 13032
rect 10408 12972 10412 13028
rect 10412 12972 10468 13028
rect 10468 12972 10472 13028
rect 10408 12968 10472 12972
rect 10408 12868 10472 12872
rect 10408 12812 10412 12868
rect 10412 12812 10468 12868
rect 10468 12812 10472 12868
rect 10408 12808 10472 12812
rect 10408 12708 10472 12712
rect 10408 12652 10412 12708
rect 10412 12652 10468 12708
rect 10468 12652 10472 12708
rect 10408 12648 10472 12652
rect 10408 12548 10472 12552
rect 10408 12492 10412 12548
rect 10412 12492 10468 12548
rect 10468 12492 10472 12548
rect 10408 12488 10472 12492
rect 10408 12328 10472 12392
rect 10408 12168 10472 12232
rect 10408 12008 10472 12072
rect 10408 11848 10472 11912
rect 10408 11748 10472 11752
rect 10408 11692 10412 11748
rect 10412 11692 10468 11748
rect 10468 11692 10472 11748
rect 10408 11688 10472 11692
rect 10408 11588 10472 11592
rect 10408 11532 10412 11588
rect 10412 11532 10468 11588
rect 10468 11532 10472 11588
rect 10408 11528 10472 11532
rect 10408 11428 10472 11432
rect 10408 11372 10412 11428
rect 10412 11372 10468 11428
rect 10468 11372 10472 11428
rect 10408 11368 10472 11372
rect 10408 11268 10472 11272
rect 10408 11212 10412 11268
rect 10412 11212 10468 11268
rect 10468 11212 10472 11268
rect 10408 11208 10472 11212
rect 10408 11108 10472 11112
rect 10408 11052 10412 11108
rect 10412 11052 10468 11108
rect 10468 11052 10472 11108
rect 10408 11048 10472 11052
rect 10408 10948 10472 10952
rect 10408 10892 10412 10948
rect 10412 10892 10468 10948
rect 10468 10892 10472 10948
rect 10408 10888 10472 10892
rect 10408 10788 10472 10792
rect 10408 10732 10412 10788
rect 10412 10732 10468 10788
rect 10468 10732 10472 10788
rect 10408 10728 10472 10732
rect 10408 10628 10472 10632
rect 10408 10572 10412 10628
rect 10412 10572 10468 10628
rect 10468 10572 10472 10628
rect 10408 10568 10472 10572
rect 10408 10468 10472 10472
rect 10408 10412 10412 10468
rect 10412 10412 10468 10468
rect 10468 10412 10472 10468
rect 10408 10408 10472 10412
rect 10408 10308 10472 10312
rect 10408 10252 10412 10308
rect 10412 10252 10468 10308
rect 10468 10252 10472 10308
rect 10408 10248 10472 10252
rect 10408 10148 10472 10152
rect 10408 10092 10412 10148
rect 10412 10092 10468 10148
rect 10468 10092 10472 10148
rect 10408 10088 10472 10092
rect 10408 9988 10472 9992
rect 10408 9932 10412 9988
rect 10412 9932 10468 9988
rect 10468 9932 10472 9988
rect 10408 9928 10472 9932
rect 10408 9828 10472 9832
rect 10408 9772 10412 9828
rect 10412 9772 10468 9828
rect 10468 9772 10472 9828
rect 10408 9768 10472 9772
rect 10408 9608 10472 9672
rect 10408 9508 10472 9512
rect 10408 9452 10412 9508
rect 10412 9452 10468 9508
rect 10468 9452 10472 9508
rect 10408 9448 10472 9452
rect 10408 9348 10472 9352
rect 10408 9292 10412 9348
rect 10412 9292 10468 9348
rect 10468 9292 10472 9348
rect 10408 9288 10472 9292
rect 10408 9128 10472 9192
rect 10408 9028 10472 9032
rect 10408 8972 10412 9028
rect 10412 8972 10468 9028
rect 10468 8972 10472 9028
rect 10408 8968 10472 8972
rect 10408 8868 10472 8872
rect 10408 8812 10412 8868
rect 10412 8812 10468 8868
rect 10468 8812 10472 8868
rect 10408 8808 10472 8812
rect 10408 8708 10472 8712
rect 10408 8652 10412 8708
rect 10412 8652 10468 8708
rect 10468 8652 10472 8708
rect 10408 8648 10472 8652
rect 10408 8548 10472 8552
rect 10408 8492 10412 8548
rect 10412 8492 10468 8548
rect 10468 8492 10472 8548
rect 10408 8488 10472 8492
rect 10408 8388 10472 8392
rect 10408 8332 10412 8388
rect 10412 8332 10468 8388
rect 10468 8332 10472 8388
rect 10408 8328 10472 8332
rect 10408 8228 10472 8232
rect 10408 8172 10412 8228
rect 10412 8172 10468 8228
rect 10468 8172 10472 8228
rect 10408 8168 10472 8172
rect 10408 8068 10472 8072
rect 10408 8012 10412 8068
rect 10412 8012 10468 8068
rect 10468 8012 10472 8068
rect 10408 8008 10472 8012
rect 10408 7908 10472 7912
rect 10408 7852 10412 7908
rect 10412 7852 10468 7908
rect 10468 7852 10472 7908
rect 10408 7848 10472 7852
rect 10408 7748 10472 7752
rect 10408 7692 10412 7748
rect 10412 7692 10468 7748
rect 10468 7692 10472 7748
rect 10408 7688 10472 7692
rect 10408 7528 10472 7592
rect 10408 7428 10472 7432
rect 10408 7372 10412 7428
rect 10412 7372 10468 7428
rect 10468 7372 10472 7428
rect 10408 7368 10472 7372
rect 10408 7268 10472 7272
rect 10408 7212 10412 7268
rect 10412 7212 10468 7268
rect 10468 7212 10472 7268
rect 10408 7208 10472 7212
rect 10408 7048 10472 7112
rect 10408 6948 10472 6952
rect 10408 6892 10412 6948
rect 10412 6892 10468 6948
rect 10468 6892 10472 6948
rect 10408 6888 10472 6892
rect 10408 6788 10472 6792
rect 10408 6732 10412 6788
rect 10412 6732 10468 6788
rect 10468 6732 10472 6788
rect 10408 6728 10472 6732
rect 10408 6568 10472 6632
rect 10408 6468 10472 6472
rect 10408 6412 10412 6468
rect 10412 6412 10468 6468
rect 10468 6412 10472 6468
rect 10408 6408 10472 6412
rect 10408 6308 10472 6312
rect 10408 6252 10412 6308
rect 10412 6252 10468 6308
rect 10468 6252 10472 6308
rect 10408 6248 10472 6252
rect 10408 6148 10472 6152
rect 10408 6092 10412 6148
rect 10412 6092 10468 6148
rect 10468 6092 10472 6148
rect 10408 6088 10472 6092
rect 10408 5988 10472 5992
rect 10408 5932 10412 5988
rect 10412 5932 10468 5988
rect 10468 5932 10472 5988
rect 10408 5928 10472 5932
rect 10408 5828 10472 5832
rect 10408 5772 10412 5828
rect 10412 5772 10468 5828
rect 10468 5772 10472 5828
rect 10408 5768 10472 5772
rect 10408 5668 10472 5672
rect 10408 5612 10412 5668
rect 10412 5612 10468 5668
rect 10468 5612 10472 5668
rect 10408 5608 10472 5612
rect 10408 5508 10472 5512
rect 10408 5452 10412 5508
rect 10412 5452 10468 5508
rect 10468 5452 10472 5508
rect 10408 5448 10472 5452
rect 10408 5348 10472 5352
rect 10408 5292 10412 5348
rect 10412 5292 10468 5348
rect 10468 5292 10472 5348
rect 10408 5288 10472 5292
rect 10408 5188 10472 5192
rect 10408 5132 10412 5188
rect 10412 5132 10468 5188
rect 10468 5132 10472 5188
rect 10408 5128 10472 5132
rect 10408 5028 10472 5032
rect 10408 4972 10412 5028
rect 10412 4972 10468 5028
rect 10468 4972 10472 5028
rect 10408 4968 10472 4972
rect 10408 4868 10472 4872
rect 10408 4812 10412 4868
rect 10412 4812 10468 4868
rect 10468 4812 10472 4868
rect 10408 4808 10472 4812
rect 10408 4708 10472 4712
rect 10408 4652 10412 4708
rect 10412 4652 10468 4708
rect 10468 4652 10472 4708
rect 10408 4648 10472 4652
rect 10408 4548 10472 4552
rect 10408 4492 10412 4548
rect 10412 4492 10468 4548
rect 10468 4492 10472 4548
rect 10408 4488 10472 4492
rect 10408 4388 10472 4392
rect 10408 4332 10412 4388
rect 10412 4332 10468 4388
rect 10468 4332 10472 4388
rect 10408 4328 10472 4332
rect 10408 4228 10472 4232
rect 10408 4172 10412 4228
rect 10412 4172 10468 4228
rect 10468 4172 10472 4228
rect 10408 4168 10472 4172
rect 10408 4068 10472 4072
rect 10408 4012 10412 4068
rect 10412 4012 10468 4068
rect 10468 4012 10472 4068
rect 10408 4008 10472 4012
rect 10408 3908 10472 3912
rect 10408 3852 10412 3908
rect 10412 3852 10468 3908
rect 10468 3852 10472 3908
rect 10408 3848 10472 3852
rect 10408 3688 10472 3752
rect 10408 3528 10472 3592
rect 10408 3428 10472 3432
rect 10408 3372 10412 3428
rect 10412 3372 10468 3428
rect 10468 3372 10472 3428
rect 10408 3368 10472 3372
rect 10408 3268 10472 3272
rect 10408 3212 10412 3268
rect 10412 3212 10468 3268
rect 10468 3212 10472 3268
rect 10408 3208 10472 3212
rect 10408 3108 10472 3112
rect 10408 3052 10412 3108
rect 10412 3052 10468 3108
rect 10468 3052 10472 3108
rect 10408 3048 10472 3052
rect 10408 2948 10472 2952
rect 10408 2892 10412 2948
rect 10412 2892 10468 2948
rect 10468 2892 10472 2948
rect 10408 2888 10472 2892
rect 10408 2788 10472 2792
rect 10408 2732 10412 2788
rect 10412 2732 10468 2788
rect 10468 2732 10472 2788
rect 10408 2728 10472 2732
rect 10408 2628 10472 2632
rect 10408 2572 10412 2628
rect 10412 2572 10468 2628
rect 10468 2572 10472 2628
rect 10408 2568 10472 2572
rect 10408 2468 10472 2472
rect 10408 2412 10412 2468
rect 10412 2412 10468 2468
rect 10468 2412 10472 2468
rect 10408 2408 10472 2412
rect 10408 2308 10472 2312
rect 10408 2252 10412 2308
rect 10412 2252 10468 2308
rect 10468 2252 10472 2308
rect 10408 2248 10472 2252
rect 10408 2148 10472 2152
rect 10408 2092 10412 2148
rect 10412 2092 10468 2148
rect 10468 2092 10472 2148
rect 10408 2088 10472 2092
rect 10408 1988 10472 1992
rect 10408 1932 10412 1988
rect 10412 1932 10468 1988
rect 10468 1932 10472 1988
rect 10408 1928 10472 1932
rect 10408 1768 10472 1832
rect 10408 1668 10472 1672
rect 10408 1612 10412 1668
rect 10412 1612 10468 1668
rect 10468 1612 10472 1668
rect 10408 1608 10472 1612
rect 10408 1508 10472 1512
rect 10408 1452 10412 1508
rect 10412 1452 10468 1508
rect 10468 1452 10472 1508
rect 10408 1448 10472 1452
rect 10408 1348 10472 1352
rect 10408 1292 10412 1348
rect 10412 1292 10468 1348
rect 10468 1292 10472 1348
rect 10408 1288 10472 1292
rect 10408 1188 10472 1192
rect 10408 1132 10412 1188
rect 10412 1132 10468 1188
rect 10468 1132 10472 1188
rect 10408 1128 10472 1132
rect 10408 1028 10472 1032
rect 10408 972 10412 1028
rect 10412 972 10468 1028
rect 10468 972 10472 1028
rect 10408 968 10472 972
rect 10408 808 10472 872
rect 10408 648 10472 712
rect 10408 548 10472 552
rect 10408 492 10412 548
rect 10412 492 10468 548
rect 10468 492 10472 548
rect 10408 488 10472 492
rect 10408 388 10472 392
rect 10408 332 10412 388
rect 10412 332 10468 388
rect 10468 332 10472 388
rect 10408 328 10472 332
rect 10408 228 10472 232
rect 10408 172 10412 228
rect 10412 172 10468 228
rect 10468 172 10472 228
rect 10408 168 10472 172
rect 10408 68 10472 72
rect 10408 12 10412 68
rect 10412 12 10468 68
rect 10468 12 10472 68
rect 10408 8 10472 12
rect 10088 -1112 10152 -1048
rect 10088 -1192 10152 -1128
rect 10088 -1272 10152 -1208
rect 10088 -1352 10152 -1288
rect 10088 -1432 10152 -1368
rect 10728 31428 10792 31432
rect 10728 31372 10732 31428
rect 10732 31372 10788 31428
rect 10788 31372 10792 31428
rect 10728 31368 10792 31372
rect 10728 31268 10792 31272
rect 10728 31212 10732 31268
rect 10732 31212 10788 31268
rect 10788 31212 10792 31268
rect 10728 31208 10792 31212
rect 10728 31108 10792 31112
rect 10728 31052 10732 31108
rect 10732 31052 10788 31108
rect 10788 31052 10792 31108
rect 10728 31048 10792 31052
rect 10728 30948 10792 30952
rect 10728 30892 10732 30948
rect 10732 30892 10788 30948
rect 10788 30892 10792 30948
rect 10728 30888 10792 30892
rect 10728 30788 10792 30792
rect 10728 30732 10732 30788
rect 10732 30732 10788 30788
rect 10788 30732 10792 30788
rect 10728 30728 10792 30732
rect 10728 30628 10792 30632
rect 10728 30572 10732 30628
rect 10732 30572 10788 30628
rect 10788 30572 10792 30628
rect 10728 30568 10792 30572
rect 10728 30468 10792 30472
rect 10728 30412 10732 30468
rect 10732 30412 10788 30468
rect 10788 30412 10792 30468
rect 10728 30408 10792 30412
rect 10728 30308 10792 30312
rect 10728 30252 10732 30308
rect 10732 30252 10788 30308
rect 10788 30252 10792 30308
rect 10728 30248 10792 30252
rect 10728 30088 10792 30152
rect 10728 29988 10792 29992
rect 10728 29932 10732 29988
rect 10732 29932 10788 29988
rect 10788 29932 10792 29988
rect 10728 29928 10792 29932
rect 10728 29828 10792 29832
rect 10728 29772 10732 29828
rect 10732 29772 10788 29828
rect 10788 29772 10792 29828
rect 10728 29768 10792 29772
rect 10728 29668 10792 29672
rect 10728 29612 10732 29668
rect 10732 29612 10788 29668
rect 10788 29612 10792 29668
rect 10728 29608 10792 29612
rect 10728 29508 10792 29512
rect 10728 29452 10732 29508
rect 10732 29452 10788 29508
rect 10788 29452 10792 29508
rect 10728 29448 10792 29452
rect 10728 29348 10792 29352
rect 10728 29292 10732 29348
rect 10732 29292 10788 29348
rect 10788 29292 10792 29348
rect 10728 29288 10792 29292
rect 10728 29188 10792 29192
rect 10728 29132 10732 29188
rect 10732 29132 10788 29188
rect 10788 29132 10792 29188
rect 10728 29128 10792 29132
rect 10728 29028 10792 29032
rect 10728 28972 10732 29028
rect 10732 28972 10788 29028
rect 10788 28972 10792 29028
rect 10728 28968 10792 28972
rect 10728 28868 10792 28872
rect 10728 28812 10732 28868
rect 10732 28812 10788 28868
rect 10788 28812 10792 28868
rect 10728 28808 10792 28812
rect 10728 28648 10792 28712
rect 10728 28488 10792 28552
rect 10728 28328 10792 28392
rect 10728 28168 10792 28232
rect 10728 28068 10792 28072
rect 10728 28012 10732 28068
rect 10732 28012 10788 28068
rect 10788 28012 10792 28068
rect 10728 28008 10792 28012
rect 10728 27908 10792 27912
rect 10728 27852 10732 27908
rect 10732 27852 10788 27908
rect 10788 27852 10792 27908
rect 10728 27848 10792 27852
rect 10728 27748 10792 27752
rect 10728 27692 10732 27748
rect 10732 27692 10788 27748
rect 10788 27692 10792 27748
rect 10728 27688 10792 27692
rect 10728 27588 10792 27592
rect 10728 27532 10732 27588
rect 10732 27532 10788 27588
rect 10788 27532 10792 27588
rect 10728 27528 10792 27532
rect 10728 27428 10792 27432
rect 10728 27372 10732 27428
rect 10732 27372 10788 27428
rect 10788 27372 10792 27428
rect 10728 27368 10792 27372
rect 10728 27268 10792 27272
rect 10728 27212 10732 27268
rect 10732 27212 10788 27268
rect 10788 27212 10792 27268
rect 10728 27208 10792 27212
rect 10728 27108 10792 27112
rect 10728 27052 10732 27108
rect 10732 27052 10788 27108
rect 10788 27052 10792 27108
rect 10728 27048 10792 27052
rect 10728 26948 10792 26952
rect 10728 26892 10732 26948
rect 10732 26892 10788 26948
rect 10788 26892 10792 26948
rect 10728 26888 10792 26892
rect 10728 26728 10792 26792
rect 10728 26568 10792 26632
rect 10728 26408 10792 26472
rect 10728 26248 10792 26312
rect 10728 26148 10792 26152
rect 10728 26092 10732 26148
rect 10732 26092 10788 26148
rect 10788 26092 10792 26148
rect 10728 26088 10792 26092
rect 10728 25988 10792 25992
rect 10728 25932 10732 25988
rect 10732 25932 10788 25988
rect 10788 25932 10792 25988
rect 10728 25928 10792 25932
rect 10728 25828 10792 25832
rect 10728 25772 10732 25828
rect 10732 25772 10788 25828
rect 10788 25772 10792 25828
rect 10728 25768 10792 25772
rect 10728 25668 10792 25672
rect 10728 25612 10732 25668
rect 10732 25612 10788 25668
rect 10788 25612 10792 25668
rect 10728 25608 10792 25612
rect 10728 25508 10792 25512
rect 10728 25452 10732 25508
rect 10732 25452 10788 25508
rect 10788 25452 10792 25508
rect 10728 25448 10792 25452
rect 10728 25348 10792 25352
rect 10728 25292 10732 25348
rect 10732 25292 10788 25348
rect 10788 25292 10792 25348
rect 10728 25288 10792 25292
rect 10728 25188 10792 25192
rect 10728 25132 10732 25188
rect 10732 25132 10788 25188
rect 10788 25132 10792 25188
rect 10728 25128 10792 25132
rect 10728 25028 10792 25032
rect 10728 24972 10732 25028
rect 10732 24972 10788 25028
rect 10788 24972 10792 25028
rect 10728 24968 10792 24972
rect 10728 24808 10792 24872
rect 10728 24708 10792 24712
rect 10728 24652 10732 24708
rect 10732 24652 10788 24708
rect 10788 24652 10792 24708
rect 10728 24648 10792 24652
rect 10728 24548 10792 24552
rect 10728 24492 10732 24548
rect 10732 24492 10788 24548
rect 10788 24492 10792 24548
rect 10728 24488 10792 24492
rect 10728 24388 10792 24392
rect 10728 24332 10732 24388
rect 10732 24332 10788 24388
rect 10788 24332 10792 24388
rect 10728 24328 10792 24332
rect 10728 24228 10792 24232
rect 10728 24172 10732 24228
rect 10732 24172 10788 24228
rect 10788 24172 10792 24228
rect 10728 24168 10792 24172
rect 10728 24068 10792 24072
rect 10728 24012 10732 24068
rect 10732 24012 10788 24068
rect 10788 24012 10792 24068
rect 10728 24008 10792 24012
rect 10728 23908 10792 23912
rect 10728 23852 10732 23908
rect 10732 23852 10788 23908
rect 10788 23852 10792 23908
rect 10728 23848 10792 23852
rect 10728 23748 10792 23752
rect 10728 23692 10732 23748
rect 10732 23692 10788 23748
rect 10788 23692 10792 23748
rect 10728 23688 10792 23692
rect 10728 23588 10792 23592
rect 10728 23532 10732 23588
rect 10732 23532 10788 23588
rect 10788 23532 10792 23588
rect 10728 23528 10792 23532
rect 10728 23428 10792 23432
rect 10728 23372 10732 23428
rect 10732 23372 10788 23428
rect 10788 23372 10792 23428
rect 10728 23368 10792 23372
rect 10728 23268 10792 23272
rect 10728 23212 10732 23268
rect 10732 23212 10788 23268
rect 10788 23212 10792 23268
rect 10728 23208 10792 23212
rect 10728 23108 10792 23112
rect 10728 23052 10732 23108
rect 10732 23052 10788 23108
rect 10788 23052 10792 23108
rect 10728 23048 10792 23052
rect 10728 22948 10792 22952
rect 10728 22892 10732 22948
rect 10732 22892 10788 22948
rect 10788 22892 10792 22948
rect 10728 22888 10792 22892
rect 10728 22788 10792 22792
rect 10728 22732 10732 22788
rect 10732 22732 10788 22788
rect 10788 22732 10792 22788
rect 10728 22728 10792 22732
rect 10728 22628 10792 22632
rect 10728 22572 10732 22628
rect 10732 22572 10788 22628
rect 10788 22572 10792 22628
rect 10728 22568 10792 22572
rect 10728 22468 10792 22472
rect 10728 22412 10732 22468
rect 10732 22412 10788 22468
rect 10788 22412 10792 22468
rect 10728 22408 10792 22412
rect 10728 22308 10792 22312
rect 10728 22252 10732 22308
rect 10732 22252 10788 22308
rect 10788 22252 10792 22308
rect 10728 22248 10792 22252
rect 10728 22148 10792 22152
rect 10728 22092 10732 22148
rect 10732 22092 10788 22148
rect 10788 22092 10792 22148
rect 10728 22088 10792 22092
rect 10728 21928 10792 21992
rect 10728 21828 10792 21832
rect 10728 21772 10732 21828
rect 10732 21772 10788 21828
rect 10788 21772 10792 21828
rect 10728 21768 10792 21772
rect 10728 21668 10792 21672
rect 10728 21612 10732 21668
rect 10732 21612 10788 21668
rect 10788 21612 10792 21668
rect 10728 21608 10792 21612
rect 10728 21508 10792 21512
rect 10728 21452 10732 21508
rect 10732 21452 10788 21508
rect 10788 21452 10792 21508
rect 10728 21448 10792 21452
rect 10728 21348 10792 21352
rect 10728 21292 10732 21348
rect 10732 21292 10788 21348
rect 10788 21292 10792 21348
rect 10728 21288 10792 21292
rect 10728 21188 10792 21192
rect 10728 21132 10732 21188
rect 10732 21132 10788 21188
rect 10788 21132 10792 21188
rect 10728 21128 10792 21132
rect 10728 21028 10792 21032
rect 10728 20972 10732 21028
rect 10732 20972 10788 21028
rect 10788 20972 10792 21028
rect 10728 20968 10792 20972
rect 10728 20868 10792 20872
rect 10728 20812 10732 20868
rect 10732 20812 10788 20868
rect 10788 20812 10792 20868
rect 10728 20808 10792 20812
rect 10728 20708 10792 20712
rect 10728 20652 10732 20708
rect 10732 20652 10788 20708
rect 10788 20652 10792 20708
rect 10728 20648 10792 20652
rect 10728 20488 10792 20552
rect 10728 20328 10792 20392
rect 10728 20168 10792 20232
rect 10728 20008 10792 20072
rect 10728 19908 10792 19912
rect 10728 19852 10732 19908
rect 10732 19852 10788 19908
rect 10788 19852 10792 19908
rect 10728 19848 10792 19852
rect 10728 19748 10792 19752
rect 10728 19692 10732 19748
rect 10732 19692 10788 19748
rect 10788 19692 10792 19748
rect 10728 19688 10792 19692
rect 10728 19588 10792 19592
rect 10728 19532 10732 19588
rect 10732 19532 10788 19588
rect 10788 19532 10792 19588
rect 10728 19528 10792 19532
rect 10728 19428 10792 19432
rect 10728 19372 10732 19428
rect 10732 19372 10788 19428
rect 10788 19372 10792 19428
rect 10728 19368 10792 19372
rect 10728 19268 10792 19272
rect 10728 19212 10732 19268
rect 10732 19212 10788 19268
rect 10788 19212 10792 19268
rect 10728 19208 10792 19212
rect 10728 19108 10792 19112
rect 10728 19052 10732 19108
rect 10732 19052 10788 19108
rect 10788 19052 10792 19108
rect 10728 19048 10792 19052
rect 10728 18948 10792 18952
rect 10728 18892 10732 18948
rect 10732 18892 10788 18948
rect 10788 18892 10792 18948
rect 10728 18888 10792 18892
rect 10728 18788 10792 18792
rect 10728 18732 10732 18788
rect 10732 18732 10788 18788
rect 10788 18732 10792 18788
rect 10728 18728 10792 18732
rect 10728 18568 10792 18632
rect 10728 18408 10792 18472
rect 10728 18248 10792 18312
rect 10728 18088 10792 18152
rect 10728 17988 10792 17992
rect 10728 17932 10732 17988
rect 10732 17932 10788 17988
rect 10788 17932 10792 17988
rect 10728 17928 10792 17932
rect 10728 17828 10792 17832
rect 10728 17772 10732 17828
rect 10732 17772 10788 17828
rect 10788 17772 10792 17828
rect 10728 17768 10792 17772
rect 10728 17668 10792 17672
rect 10728 17612 10732 17668
rect 10732 17612 10788 17668
rect 10788 17612 10792 17668
rect 10728 17608 10792 17612
rect 10728 17508 10792 17512
rect 10728 17452 10732 17508
rect 10732 17452 10788 17508
rect 10788 17452 10792 17508
rect 10728 17448 10792 17452
rect 10728 17348 10792 17352
rect 10728 17292 10732 17348
rect 10732 17292 10788 17348
rect 10788 17292 10792 17348
rect 10728 17288 10792 17292
rect 10728 17188 10792 17192
rect 10728 17132 10732 17188
rect 10732 17132 10788 17188
rect 10788 17132 10792 17188
rect 10728 17128 10792 17132
rect 10728 17028 10792 17032
rect 10728 16972 10732 17028
rect 10732 16972 10788 17028
rect 10788 16972 10792 17028
rect 10728 16968 10792 16972
rect 10728 16868 10792 16872
rect 10728 16812 10732 16868
rect 10732 16812 10788 16868
rect 10788 16812 10792 16868
rect 10728 16808 10792 16812
rect 10728 16648 10792 16712
rect 10728 16548 10792 16552
rect 10728 16492 10732 16548
rect 10732 16492 10788 16548
rect 10788 16492 10792 16548
rect 10728 16488 10792 16492
rect 10728 16388 10792 16392
rect 10728 16332 10732 16388
rect 10732 16332 10788 16388
rect 10788 16332 10792 16388
rect 10728 16328 10792 16332
rect 10728 16228 10792 16232
rect 10728 16172 10732 16228
rect 10732 16172 10788 16228
rect 10788 16172 10792 16228
rect 10728 16168 10792 16172
rect 10728 16068 10792 16072
rect 10728 16012 10732 16068
rect 10732 16012 10788 16068
rect 10788 16012 10792 16068
rect 10728 16008 10792 16012
rect 10728 15908 10792 15912
rect 10728 15852 10732 15908
rect 10732 15852 10788 15908
rect 10788 15852 10792 15908
rect 10728 15848 10792 15852
rect 10728 15748 10792 15752
rect 10728 15692 10732 15748
rect 10732 15692 10788 15748
rect 10788 15692 10792 15748
rect 10728 15688 10792 15692
rect 10728 15588 10792 15592
rect 10728 15532 10732 15588
rect 10732 15532 10788 15588
rect 10788 15532 10792 15588
rect 10728 15528 10792 15532
rect 10728 15428 10792 15432
rect 10728 15372 10732 15428
rect 10732 15372 10788 15428
rect 10788 15372 10792 15428
rect 10728 15368 10792 15372
rect 10728 15268 10792 15272
rect 10728 15212 10732 15268
rect 10732 15212 10788 15268
rect 10788 15212 10792 15268
rect 10728 15208 10792 15212
rect 10728 15108 10792 15112
rect 10728 15052 10732 15108
rect 10732 15052 10788 15108
rect 10788 15052 10792 15108
rect 10728 15048 10792 15052
rect 10728 14948 10792 14952
rect 10728 14892 10732 14948
rect 10732 14892 10788 14948
rect 10788 14892 10792 14948
rect 10728 14888 10792 14892
rect 10728 14788 10792 14792
rect 10728 14732 10732 14788
rect 10732 14732 10788 14788
rect 10788 14732 10792 14788
rect 10728 14728 10792 14732
rect 10728 14628 10792 14632
rect 10728 14572 10732 14628
rect 10732 14572 10788 14628
rect 10788 14572 10792 14628
rect 10728 14568 10792 14572
rect 10728 14468 10792 14472
rect 10728 14412 10732 14468
rect 10732 14412 10788 14468
rect 10788 14412 10792 14468
rect 10728 14408 10792 14412
rect 10728 14308 10792 14312
rect 10728 14252 10732 14308
rect 10732 14252 10788 14308
rect 10788 14252 10792 14308
rect 10728 14248 10792 14252
rect 10728 14148 10792 14152
rect 10728 14092 10732 14148
rect 10732 14092 10788 14148
rect 10788 14092 10792 14148
rect 10728 14088 10792 14092
rect 10728 13988 10792 13992
rect 10728 13932 10732 13988
rect 10732 13932 10788 13988
rect 10788 13932 10792 13988
rect 10728 13928 10792 13932
rect 10728 13768 10792 13832
rect 10728 13668 10792 13672
rect 10728 13612 10732 13668
rect 10732 13612 10788 13668
rect 10788 13612 10792 13668
rect 10728 13608 10792 13612
rect 10728 13508 10792 13512
rect 10728 13452 10732 13508
rect 10732 13452 10788 13508
rect 10788 13452 10792 13508
rect 10728 13448 10792 13452
rect 10728 13348 10792 13352
rect 10728 13292 10732 13348
rect 10732 13292 10788 13348
rect 10788 13292 10792 13348
rect 10728 13288 10792 13292
rect 10728 13188 10792 13192
rect 10728 13132 10732 13188
rect 10732 13132 10788 13188
rect 10788 13132 10792 13188
rect 10728 13128 10792 13132
rect 10728 13028 10792 13032
rect 10728 12972 10732 13028
rect 10732 12972 10788 13028
rect 10788 12972 10792 13028
rect 10728 12968 10792 12972
rect 10728 12868 10792 12872
rect 10728 12812 10732 12868
rect 10732 12812 10788 12868
rect 10788 12812 10792 12868
rect 10728 12808 10792 12812
rect 10728 12708 10792 12712
rect 10728 12652 10732 12708
rect 10732 12652 10788 12708
rect 10788 12652 10792 12708
rect 10728 12648 10792 12652
rect 10728 12548 10792 12552
rect 10728 12492 10732 12548
rect 10732 12492 10788 12548
rect 10788 12492 10792 12548
rect 10728 12488 10792 12492
rect 10728 12328 10792 12392
rect 10728 12168 10792 12232
rect 10728 12008 10792 12072
rect 10728 11848 10792 11912
rect 10728 11748 10792 11752
rect 10728 11692 10732 11748
rect 10732 11692 10788 11748
rect 10788 11692 10792 11748
rect 10728 11688 10792 11692
rect 10728 11588 10792 11592
rect 10728 11532 10732 11588
rect 10732 11532 10788 11588
rect 10788 11532 10792 11588
rect 10728 11528 10792 11532
rect 10728 11428 10792 11432
rect 10728 11372 10732 11428
rect 10732 11372 10788 11428
rect 10788 11372 10792 11428
rect 10728 11368 10792 11372
rect 10728 11268 10792 11272
rect 10728 11212 10732 11268
rect 10732 11212 10788 11268
rect 10788 11212 10792 11268
rect 10728 11208 10792 11212
rect 10728 11108 10792 11112
rect 10728 11052 10732 11108
rect 10732 11052 10788 11108
rect 10788 11052 10792 11108
rect 10728 11048 10792 11052
rect 10728 10948 10792 10952
rect 10728 10892 10732 10948
rect 10732 10892 10788 10948
rect 10788 10892 10792 10948
rect 10728 10888 10792 10892
rect 10728 10788 10792 10792
rect 10728 10732 10732 10788
rect 10732 10732 10788 10788
rect 10788 10732 10792 10788
rect 10728 10728 10792 10732
rect 10728 10628 10792 10632
rect 10728 10572 10732 10628
rect 10732 10572 10788 10628
rect 10788 10572 10792 10628
rect 10728 10568 10792 10572
rect 10728 10468 10792 10472
rect 10728 10412 10732 10468
rect 10732 10412 10788 10468
rect 10788 10412 10792 10468
rect 10728 10408 10792 10412
rect 10728 10308 10792 10312
rect 10728 10252 10732 10308
rect 10732 10252 10788 10308
rect 10788 10252 10792 10308
rect 10728 10248 10792 10252
rect 10728 10148 10792 10152
rect 10728 10092 10732 10148
rect 10732 10092 10788 10148
rect 10788 10092 10792 10148
rect 10728 10088 10792 10092
rect 10728 9988 10792 9992
rect 10728 9932 10732 9988
rect 10732 9932 10788 9988
rect 10788 9932 10792 9988
rect 10728 9928 10792 9932
rect 10728 9828 10792 9832
rect 10728 9772 10732 9828
rect 10732 9772 10788 9828
rect 10788 9772 10792 9828
rect 10728 9768 10792 9772
rect 10728 9608 10792 9672
rect 10728 9508 10792 9512
rect 10728 9452 10732 9508
rect 10732 9452 10788 9508
rect 10788 9452 10792 9508
rect 10728 9448 10792 9452
rect 10728 9348 10792 9352
rect 10728 9292 10732 9348
rect 10732 9292 10788 9348
rect 10788 9292 10792 9348
rect 10728 9288 10792 9292
rect 10728 9128 10792 9192
rect 10728 9028 10792 9032
rect 10728 8972 10732 9028
rect 10732 8972 10788 9028
rect 10788 8972 10792 9028
rect 10728 8968 10792 8972
rect 10728 8868 10792 8872
rect 10728 8812 10732 8868
rect 10732 8812 10788 8868
rect 10788 8812 10792 8868
rect 10728 8808 10792 8812
rect 10728 8708 10792 8712
rect 10728 8652 10732 8708
rect 10732 8652 10788 8708
rect 10788 8652 10792 8708
rect 10728 8648 10792 8652
rect 10728 8548 10792 8552
rect 10728 8492 10732 8548
rect 10732 8492 10788 8548
rect 10788 8492 10792 8548
rect 10728 8488 10792 8492
rect 10728 8388 10792 8392
rect 10728 8332 10732 8388
rect 10732 8332 10788 8388
rect 10788 8332 10792 8388
rect 10728 8328 10792 8332
rect 10728 8228 10792 8232
rect 10728 8172 10732 8228
rect 10732 8172 10788 8228
rect 10788 8172 10792 8228
rect 10728 8168 10792 8172
rect 10728 8068 10792 8072
rect 10728 8012 10732 8068
rect 10732 8012 10788 8068
rect 10788 8012 10792 8068
rect 10728 8008 10792 8012
rect 10728 7908 10792 7912
rect 10728 7852 10732 7908
rect 10732 7852 10788 7908
rect 10788 7852 10792 7908
rect 10728 7848 10792 7852
rect 10728 7748 10792 7752
rect 10728 7692 10732 7748
rect 10732 7692 10788 7748
rect 10788 7692 10792 7748
rect 10728 7688 10792 7692
rect 10728 7528 10792 7592
rect 10728 7428 10792 7432
rect 10728 7372 10732 7428
rect 10732 7372 10788 7428
rect 10788 7372 10792 7428
rect 10728 7368 10792 7372
rect 10728 7268 10792 7272
rect 10728 7212 10732 7268
rect 10732 7212 10788 7268
rect 10788 7212 10792 7268
rect 10728 7208 10792 7212
rect 10728 7048 10792 7112
rect 10728 6948 10792 6952
rect 10728 6892 10732 6948
rect 10732 6892 10788 6948
rect 10788 6892 10792 6948
rect 10728 6888 10792 6892
rect 10728 6788 10792 6792
rect 10728 6732 10732 6788
rect 10732 6732 10788 6788
rect 10788 6732 10792 6788
rect 10728 6728 10792 6732
rect 10728 6568 10792 6632
rect 10728 6468 10792 6472
rect 10728 6412 10732 6468
rect 10732 6412 10788 6468
rect 10788 6412 10792 6468
rect 10728 6408 10792 6412
rect 10728 6308 10792 6312
rect 10728 6252 10732 6308
rect 10732 6252 10788 6308
rect 10788 6252 10792 6308
rect 10728 6248 10792 6252
rect 10728 6148 10792 6152
rect 10728 6092 10732 6148
rect 10732 6092 10788 6148
rect 10788 6092 10792 6148
rect 10728 6088 10792 6092
rect 10728 5988 10792 5992
rect 10728 5932 10732 5988
rect 10732 5932 10788 5988
rect 10788 5932 10792 5988
rect 10728 5928 10792 5932
rect 10728 5828 10792 5832
rect 10728 5772 10732 5828
rect 10732 5772 10788 5828
rect 10788 5772 10792 5828
rect 10728 5768 10792 5772
rect 10728 5668 10792 5672
rect 10728 5612 10732 5668
rect 10732 5612 10788 5668
rect 10788 5612 10792 5668
rect 10728 5608 10792 5612
rect 10728 5508 10792 5512
rect 10728 5452 10732 5508
rect 10732 5452 10788 5508
rect 10788 5452 10792 5508
rect 10728 5448 10792 5452
rect 10728 5348 10792 5352
rect 10728 5292 10732 5348
rect 10732 5292 10788 5348
rect 10788 5292 10792 5348
rect 10728 5288 10792 5292
rect 10728 5188 10792 5192
rect 10728 5132 10732 5188
rect 10732 5132 10788 5188
rect 10788 5132 10792 5188
rect 10728 5128 10792 5132
rect 10728 5028 10792 5032
rect 10728 4972 10732 5028
rect 10732 4972 10788 5028
rect 10788 4972 10792 5028
rect 10728 4968 10792 4972
rect 10728 4868 10792 4872
rect 10728 4812 10732 4868
rect 10732 4812 10788 4868
rect 10788 4812 10792 4868
rect 10728 4808 10792 4812
rect 10728 4708 10792 4712
rect 10728 4652 10732 4708
rect 10732 4652 10788 4708
rect 10788 4652 10792 4708
rect 10728 4648 10792 4652
rect 10728 4548 10792 4552
rect 10728 4492 10732 4548
rect 10732 4492 10788 4548
rect 10788 4492 10792 4548
rect 10728 4488 10792 4492
rect 10728 4388 10792 4392
rect 10728 4332 10732 4388
rect 10732 4332 10788 4388
rect 10788 4332 10792 4388
rect 10728 4328 10792 4332
rect 10728 4228 10792 4232
rect 10728 4172 10732 4228
rect 10732 4172 10788 4228
rect 10788 4172 10792 4228
rect 10728 4168 10792 4172
rect 10728 4068 10792 4072
rect 10728 4012 10732 4068
rect 10732 4012 10788 4068
rect 10788 4012 10792 4068
rect 10728 4008 10792 4012
rect 10728 3908 10792 3912
rect 10728 3852 10732 3908
rect 10732 3852 10788 3908
rect 10788 3852 10792 3908
rect 10728 3848 10792 3852
rect 10728 3688 10792 3752
rect 10728 3528 10792 3592
rect 10728 3428 10792 3432
rect 10728 3372 10732 3428
rect 10732 3372 10788 3428
rect 10788 3372 10792 3428
rect 10728 3368 10792 3372
rect 10728 3268 10792 3272
rect 10728 3212 10732 3268
rect 10732 3212 10788 3268
rect 10788 3212 10792 3268
rect 10728 3208 10792 3212
rect 10728 3108 10792 3112
rect 10728 3052 10732 3108
rect 10732 3052 10788 3108
rect 10788 3052 10792 3108
rect 10728 3048 10792 3052
rect 10728 2948 10792 2952
rect 10728 2892 10732 2948
rect 10732 2892 10788 2948
rect 10788 2892 10792 2948
rect 10728 2888 10792 2892
rect 10728 2788 10792 2792
rect 10728 2732 10732 2788
rect 10732 2732 10788 2788
rect 10788 2732 10792 2788
rect 10728 2728 10792 2732
rect 10728 2628 10792 2632
rect 10728 2572 10732 2628
rect 10732 2572 10788 2628
rect 10788 2572 10792 2628
rect 10728 2568 10792 2572
rect 10728 2468 10792 2472
rect 10728 2412 10732 2468
rect 10732 2412 10788 2468
rect 10788 2412 10792 2468
rect 10728 2408 10792 2412
rect 10728 2308 10792 2312
rect 10728 2252 10732 2308
rect 10732 2252 10788 2308
rect 10788 2252 10792 2308
rect 10728 2248 10792 2252
rect 10728 2148 10792 2152
rect 10728 2092 10732 2148
rect 10732 2092 10788 2148
rect 10788 2092 10792 2148
rect 10728 2088 10792 2092
rect 10728 1988 10792 1992
rect 10728 1932 10732 1988
rect 10732 1932 10788 1988
rect 10788 1932 10792 1988
rect 10728 1928 10792 1932
rect 10728 1768 10792 1832
rect 10728 1668 10792 1672
rect 10728 1612 10732 1668
rect 10732 1612 10788 1668
rect 10788 1612 10792 1668
rect 10728 1608 10792 1612
rect 10728 1508 10792 1512
rect 10728 1452 10732 1508
rect 10732 1452 10788 1508
rect 10788 1452 10792 1508
rect 10728 1448 10792 1452
rect 10728 1348 10792 1352
rect 10728 1292 10732 1348
rect 10732 1292 10788 1348
rect 10788 1292 10792 1348
rect 10728 1288 10792 1292
rect 10728 1188 10792 1192
rect 10728 1132 10732 1188
rect 10732 1132 10788 1188
rect 10788 1132 10792 1188
rect 10728 1128 10792 1132
rect 10728 1028 10792 1032
rect 10728 972 10732 1028
rect 10732 972 10788 1028
rect 10788 972 10792 1028
rect 10728 968 10792 972
rect 10728 808 10792 872
rect 10728 648 10792 712
rect 10728 548 10792 552
rect 10728 492 10732 548
rect 10732 492 10788 548
rect 10788 492 10792 548
rect 10728 488 10792 492
rect 10728 388 10792 392
rect 10728 332 10732 388
rect 10732 332 10788 388
rect 10788 332 10792 388
rect 10728 328 10792 332
rect 10728 228 10792 232
rect 10728 172 10732 228
rect 10732 172 10788 228
rect 10788 172 10792 228
rect 10728 168 10792 172
rect 10728 68 10792 72
rect 10728 12 10732 68
rect 10732 12 10788 68
rect 10788 12 10792 68
rect 10728 8 10792 12
rect 10408 -1112 10472 -1048
rect 10408 -1192 10472 -1128
rect 10408 -1272 10472 -1208
rect 10408 -1352 10472 -1288
rect 10408 -1432 10472 -1368
rect 11048 31428 11112 31432
rect 11048 31372 11052 31428
rect 11052 31372 11108 31428
rect 11108 31372 11112 31428
rect 11048 31368 11112 31372
rect 11048 31268 11112 31272
rect 11048 31212 11052 31268
rect 11052 31212 11108 31268
rect 11108 31212 11112 31268
rect 11048 31208 11112 31212
rect 11048 31108 11112 31112
rect 11048 31052 11052 31108
rect 11052 31052 11108 31108
rect 11108 31052 11112 31108
rect 11048 31048 11112 31052
rect 11048 30948 11112 30952
rect 11048 30892 11052 30948
rect 11052 30892 11108 30948
rect 11108 30892 11112 30948
rect 11048 30888 11112 30892
rect 11048 30788 11112 30792
rect 11048 30732 11052 30788
rect 11052 30732 11108 30788
rect 11108 30732 11112 30788
rect 11048 30728 11112 30732
rect 11048 30628 11112 30632
rect 11048 30572 11052 30628
rect 11052 30572 11108 30628
rect 11108 30572 11112 30628
rect 11048 30568 11112 30572
rect 11048 30468 11112 30472
rect 11048 30412 11052 30468
rect 11052 30412 11108 30468
rect 11108 30412 11112 30468
rect 11048 30408 11112 30412
rect 11048 30308 11112 30312
rect 11048 30252 11052 30308
rect 11052 30252 11108 30308
rect 11108 30252 11112 30308
rect 11048 30248 11112 30252
rect 11048 30088 11112 30152
rect 11048 29988 11112 29992
rect 11048 29932 11052 29988
rect 11052 29932 11108 29988
rect 11108 29932 11112 29988
rect 11048 29928 11112 29932
rect 11048 29828 11112 29832
rect 11048 29772 11052 29828
rect 11052 29772 11108 29828
rect 11108 29772 11112 29828
rect 11048 29768 11112 29772
rect 11048 29668 11112 29672
rect 11048 29612 11052 29668
rect 11052 29612 11108 29668
rect 11108 29612 11112 29668
rect 11048 29608 11112 29612
rect 11048 29508 11112 29512
rect 11048 29452 11052 29508
rect 11052 29452 11108 29508
rect 11108 29452 11112 29508
rect 11048 29448 11112 29452
rect 11048 29348 11112 29352
rect 11048 29292 11052 29348
rect 11052 29292 11108 29348
rect 11108 29292 11112 29348
rect 11048 29288 11112 29292
rect 11048 29188 11112 29192
rect 11048 29132 11052 29188
rect 11052 29132 11108 29188
rect 11108 29132 11112 29188
rect 11048 29128 11112 29132
rect 11048 29028 11112 29032
rect 11048 28972 11052 29028
rect 11052 28972 11108 29028
rect 11108 28972 11112 29028
rect 11048 28968 11112 28972
rect 11048 28868 11112 28872
rect 11048 28812 11052 28868
rect 11052 28812 11108 28868
rect 11108 28812 11112 28868
rect 11048 28808 11112 28812
rect 11048 28648 11112 28712
rect 11048 28488 11112 28552
rect 11048 28328 11112 28392
rect 11048 28168 11112 28232
rect 11048 28068 11112 28072
rect 11048 28012 11052 28068
rect 11052 28012 11108 28068
rect 11108 28012 11112 28068
rect 11048 28008 11112 28012
rect 11048 27908 11112 27912
rect 11048 27852 11052 27908
rect 11052 27852 11108 27908
rect 11108 27852 11112 27908
rect 11048 27848 11112 27852
rect 11048 27748 11112 27752
rect 11048 27692 11052 27748
rect 11052 27692 11108 27748
rect 11108 27692 11112 27748
rect 11048 27688 11112 27692
rect 11048 27588 11112 27592
rect 11048 27532 11052 27588
rect 11052 27532 11108 27588
rect 11108 27532 11112 27588
rect 11048 27528 11112 27532
rect 11048 27428 11112 27432
rect 11048 27372 11052 27428
rect 11052 27372 11108 27428
rect 11108 27372 11112 27428
rect 11048 27368 11112 27372
rect 11048 27268 11112 27272
rect 11048 27212 11052 27268
rect 11052 27212 11108 27268
rect 11108 27212 11112 27268
rect 11048 27208 11112 27212
rect 11048 27108 11112 27112
rect 11048 27052 11052 27108
rect 11052 27052 11108 27108
rect 11108 27052 11112 27108
rect 11048 27048 11112 27052
rect 11048 26948 11112 26952
rect 11048 26892 11052 26948
rect 11052 26892 11108 26948
rect 11108 26892 11112 26948
rect 11048 26888 11112 26892
rect 11048 26728 11112 26792
rect 11048 26568 11112 26632
rect 11048 26408 11112 26472
rect 11048 26248 11112 26312
rect 11048 26148 11112 26152
rect 11048 26092 11052 26148
rect 11052 26092 11108 26148
rect 11108 26092 11112 26148
rect 11048 26088 11112 26092
rect 11048 25988 11112 25992
rect 11048 25932 11052 25988
rect 11052 25932 11108 25988
rect 11108 25932 11112 25988
rect 11048 25928 11112 25932
rect 11048 25828 11112 25832
rect 11048 25772 11052 25828
rect 11052 25772 11108 25828
rect 11108 25772 11112 25828
rect 11048 25768 11112 25772
rect 11048 25668 11112 25672
rect 11048 25612 11052 25668
rect 11052 25612 11108 25668
rect 11108 25612 11112 25668
rect 11048 25608 11112 25612
rect 11048 25508 11112 25512
rect 11048 25452 11052 25508
rect 11052 25452 11108 25508
rect 11108 25452 11112 25508
rect 11048 25448 11112 25452
rect 11048 25348 11112 25352
rect 11048 25292 11052 25348
rect 11052 25292 11108 25348
rect 11108 25292 11112 25348
rect 11048 25288 11112 25292
rect 11048 25188 11112 25192
rect 11048 25132 11052 25188
rect 11052 25132 11108 25188
rect 11108 25132 11112 25188
rect 11048 25128 11112 25132
rect 11048 25028 11112 25032
rect 11048 24972 11052 25028
rect 11052 24972 11108 25028
rect 11108 24972 11112 25028
rect 11048 24968 11112 24972
rect 11048 24808 11112 24872
rect 11048 24708 11112 24712
rect 11048 24652 11052 24708
rect 11052 24652 11108 24708
rect 11108 24652 11112 24708
rect 11048 24648 11112 24652
rect 11048 24548 11112 24552
rect 11048 24492 11052 24548
rect 11052 24492 11108 24548
rect 11108 24492 11112 24548
rect 11048 24488 11112 24492
rect 11048 24388 11112 24392
rect 11048 24332 11052 24388
rect 11052 24332 11108 24388
rect 11108 24332 11112 24388
rect 11048 24328 11112 24332
rect 11048 24228 11112 24232
rect 11048 24172 11052 24228
rect 11052 24172 11108 24228
rect 11108 24172 11112 24228
rect 11048 24168 11112 24172
rect 11048 24068 11112 24072
rect 11048 24012 11052 24068
rect 11052 24012 11108 24068
rect 11108 24012 11112 24068
rect 11048 24008 11112 24012
rect 11048 23908 11112 23912
rect 11048 23852 11052 23908
rect 11052 23852 11108 23908
rect 11108 23852 11112 23908
rect 11048 23848 11112 23852
rect 11048 23748 11112 23752
rect 11048 23692 11052 23748
rect 11052 23692 11108 23748
rect 11108 23692 11112 23748
rect 11048 23688 11112 23692
rect 11048 23588 11112 23592
rect 11048 23532 11052 23588
rect 11052 23532 11108 23588
rect 11108 23532 11112 23588
rect 11048 23528 11112 23532
rect 11048 23428 11112 23432
rect 11048 23372 11052 23428
rect 11052 23372 11108 23428
rect 11108 23372 11112 23428
rect 11048 23368 11112 23372
rect 11048 23268 11112 23272
rect 11048 23212 11052 23268
rect 11052 23212 11108 23268
rect 11108 23212 11112 23268
rect 11048 23208 11112 23212
rect 11048 23108 11112 23112
rect 11048 23052 11052 23108
rect 11052 23052 11108 23108
rect 11108 23052 11112 23108
rect 11048 23048 11112 23052
rect 11048 22948 11112 22952
rect 11048 22892 11052 22948
rect 11052 22892 11108 22948
rect 11108 22892 11112 22948
rect 11048 22888 11112 22892
rect 11048 22788 11112 22792
rect 11048 22732 11052 22788
rect 11052 22732 11108 22788
rect 11108 22732 11112 22788
rect 11048 22728 11112 22732
rect 11048 22628 11112 22632
rect 11048 22572 11052 22628
rect 11052 22572 11108 22628
rect 11108 22572 11112 22628
rect 11048 22568 11112 22572
rect 11048 22468 11112 22472
rect 11048 22412 11052 22468
rect 11052 22412 11108 22468
rect 11108 22412 11112 22468
rect 11048 22408 11112 22412
rect 11048 22308 11112 22312
rect 11048 22252 11052 22308
rect 11052 22252 11108 22308
rect 11108 22252 11112 22308
rect 11048 22248 11112 22252
rect 11048 22148 11112 22152
rect 11048 22092 11052 22148
rect 11052 22092 11108 22148
rect 11108 22092 11112 22148
rect 11048 22088 11112 22092
rect 11048 21928 11112 21992
rect 11048 21828 11112 21832
rect 11048 21772 11052 21828
rect 11052 21772 11108 21828
rect 11108 21772 11112 21828
rect 11048 21768 11112 21772
rect 11048 21668 11112 21672
rect 11048 21612 11052 21668
rect 11052 21612 11108 21668
rect 11108 21612 11112 21668
rect 11048 21608 11112 21612
rect 11048 21508 11112 21512
rect 11048 21452 11052 21508
rect 11052 21452 11108 21508
rect 11108 21452 11112 21508
rect 11048 21448 11112 21452
rect 11048 21348 11112 21352
rect 11048 21292 11052 21348
rect 11052 21292 11108 21348
rect 11108 21292 11112 21348
rect 11048 21288 11112 21292
rect 11048 21188 11112 21192
rect 11048 21132 11052 21188
rect 11052 21132 11108 21188
rect 11108 21132 11112 21188
rect 11048 21128 11112 21132
rect 11048 21028 11112 21032
rect 11048 20972 11052 21028
rect 11052 20972 11108 21028
rect 11108 20972 11112 21028
rect 11048 20968 11112 20972
rect 11048 20868 11112 20872
rect 11048 20812 11052 20868
rect 11052 20812 11108 20868
rect 11108 20812 11112 20868
rect 11048 20808 11112 20812
rect 11048 20708 11112 20712
rect 11048 20652 11052 20708
rect 11052 20652 11108 20708
rect 11108 20652 11112 20708
rect 11048 20648 11112 20652
rect 11048 20488 11112 20552
rect 11048 20328 11112 20392
rect 11048 20168 11112 20232
rect 11048 20008 11112 20072
rect 11048 19908 11112 19912
rect 11048 19852 11052 19908
rect 11052 19852 11108 19908
rect 11108 19852 11112 19908
rect 11048 19848 11112 19852
rect 11048 19748 11112 19752
rect 11048 19692 11052 19748
rect 11052 19692 11108 19748
rect 11108 19692 11112 19748
rect 11048 19688 11112 19692
rect 11048 19588 11112 19592
rect 11048 19532 11052 19588
rect 11052 19532 11108 19588
rect 11108 19532 11112 19588
rect 11048 19528 11112 19532
rect 11048 19428 11112 19432
rect 11048 19372 11052 19428
rect 11052 19372 11108 19428
rect 11108 19372 11112 19428
rect 11048 19368 11112 19372
rect 11048 19268 11112 19272
rect 11048 19212 11052 19268
rect 11052 19212 11108 19268
rect 11108 19212 11112 19268
rect 11048 19208 11112 19212
rect 11048 19108 11112 19112
rect 11048 19052 11052 19108
rect 11052 19052 11108 19108
rect 11108 19052 11112 19108
rect 11048 19048 11112 19052
rect 11048 18948 11112 18952
rect 11048 18892 11052 18948
rect 11052 18892 11108 18948
rect 11108 18892 11112 18948
rect 11048 18888 11112 18892
rect 11048 18788 11112 18792
rect 11048 18732 11052 18788
rect 11052 18732 11108 18788
rect 11108 18732 11112 18788
rect 11048 18728 11112 18732
rect 11048 18568 11112 18632
rect 11048 18408 11112 18472
rect 11048 18248 11112 18312
rect 11048 18088 11112 18152
rect 11048 17988 11112 17992
rect 11048 17932 11052 17988
rect 11052 17932 11108 17988
rect 11108 17932 11112 17988
rect 11048 17928 11112 17932
rect 11048 17828 11112 17832
rect 11048 17772 11052 17828
rect 11052 17772 11108 17828
rect 11108 17772 11112 17828
rect 11048 17768 11112 17772
rect 11048 17668 11112 17672
rect 11048 17612 11052 17668
rect 11052 17612 11108 17668
rect 11108 17612 11112 17668
rect 11048 17608 11112 17612
rect 11048 17508 11112 17512
rect 11048 17452 11052 17508
rect 11052 17452 11108 17508
rect 11108 17452 11112 17508
rect 11048 17448 11112 17452
rect 11048 17348 11112 17352
rect 11048 17292 11052 17348
rect 11052 17292 11108 17348
rect 11108 17292 11112 17348
rect 11048 17288 11112 17292
rect 11048 17188 11112 17192
rect 11048 17132 11052 17188
rect 11052 17132 11108 17188
rect 11108 17132 11112 17188
rect 11048 17128 11112 17132
rect 11048 17028 11112 17032
rect 11048 16972 11052 17028
rect 11052 16972 11108 17028
rect 11108 16972 11112 17028
rect 11048 16968 11112 16972
rect 11048 16868 11112 16872
rect 11048 16812 11052 16868
rect 11052 16812 11108 16868
rect 11108 16812 11112 16868
rect 11048 16808 11112 16812
rect 11048 16648 11112 16712
rect 11048 16548 11112 16552
rect 11048 16492 11052 16548
rect 11052 16492 11108 16548
rect 11108 16492 11112 16548
rect 11048 16488 11112 16492
rect 11048 16388 11112 16392
rect 11048 16332 11052 16388
rect 11052 16332 11108 16388
rect 11108 16332 11112 16388
rect 11048 16328 11112 16332
rect 11048 16228 11112 16232
rect 11048 16172 11052 16228
rect 11052 16172 11108 16228
rect 11108 16172 11112 16228
rect 11048 16168 11112 16172
rect 11048 16068 11112 16072
rect 11048 16012 11052 16068
rect 11052 16012 11108 16068
rect 11108 16012 11112 16068
rect 11048 16008 11112 16012
rect 11048 15908 11112 15912
rect 11048 15852 11052 15908
rect 11052 15852 11108 15908
rect 11108 15852 11112 15908
rect 11048 15848 11112 15852
rect 11048 15748 11112 15752
rect 11048 15692 11052 15748
rect 11052 15692 11108 15748
rect 11108 15692 11112 15748
rect 11048 15688 11112 15692
rect 11048 15588 11112 15592
rect 11048 15532 11052 15588
rect 11052 15532 11108 15588
rect 11108 15532 11112 15588
rect 11048 15528 11112 15532
rect 11048 15428 11112 15432
rect 11048 15372 11052 15428
rect 11052 15372 11108 15428
rect 11108 15372 11112 15428
rect 11048 15368 11112 15372
rect 11048 15268 11112 15272
rect 11048 15212 11052 15268
rect 11052 15212 11108 15268
rect 11108 15212 11112 15268
rect 11048 15208 11112 15212
rect 11048 15108 11112 15112
rect 11048 15052 11052 15108
rect 11052 15052 11108 15108
rect 11108 15052 11112 15108
rect 11048 15048 11112 15052
rect 11048 14948 11112 14952
rect 11048 14892 11052 14948
rect 11052 14892 11108 14948
rect 11108 14892 11112 14948
rect 11048 14888 11112 14892
rect 11048 14788 11112 14792
rect 11048 14732 11052 14788
rect 11052 14732 11108 14788
rect 11108 14732 11112 14788
rect 11048 14728 11112 14732
rect 11048 14628 11112 14632
rect 11048 14572 11052 14628
rect 11052 14572 11108 14628
rect 11108 14572 11112 14628
rect 11048 14568 11112 14572
rect 11048 14468 11112 14472
rect 11048 14412 11052 14468
rect 11052 14412 11108 14468
rect 11108 14412 11112 14468
rect 11048 14408 11112 14412
rect 11048 14308 11112 14312
rect 11048 14252 11052 14308
rect 11052 14252 11108 14308
rect 11108 14252 11112 14308
rect 11048 14248 11112 14252
rect 11048 14148 11112 14152
rect 11048 14092 11052 14148
rect 11052 14092 11108 14148
rect 11108 14092 11112 14148
rect 11048 14088 11112 14092
rect 11048 13988 11112 13992
rect 11048 13932 11052 13988
rect 11052 13932 11108 13988
rect 11108 13932 11112 13988
rect 11048 13928 11112 13932
rect 11048 13768 11112 13832
rect 11048 13668 11112 13672
rect 11048 13612 11052 13668
rect 11052 13612 11108 13668
rect 11108 13612 11112 13668
rect 11048 13608 11112 13612
rect 11048 13508 11112 13512
rect 11048 13452 11052 13508
rect 11052 13452 11108 13508
rect 11108 13452 11112 13508
rect 11048 13448 11112 13452
rect 11048 13348 11112 13352
rect 11048 13292 11052 13348
rect 11052 13292 11108 13348
rect 11108 13292 11112 13348
rect 11048 13288 11112 13292
rect 11048 13188 11112 13192
rect 11048 13132 11052 13188
rect 11052 13132 11108 13188
rect 11108 13132 11112 13188
rect 11048 13128 11112 13132
rect 11048 13028 11112 13032
rect 11048 12972 11052 13028
rect 11052 12972 11108 13028
rect 11108 12972 11112 13028
rect 11048 12968 11112 12972
rect 11048 12868 11112 12872
rect 11048 12812 11052 12868
rect 11052 12812 11108 12868
rect 11108 12812 11112 12868
rect 11048 12808 11112 12812
rect 11048 12708 11112 12712
rect 11048 12652 11052 12708
rect 11052 12652 11108 12708
rect 11108 12652 11112 12708
rect 11048 12648 11112 12652
rect 11048 12548 11112 12552
rect 11048 12492 11052 12548
rect 11052 12492 11108 12548
rect 11108 12492 11112 12548
rect 11048 12488 11112 12492
rect 11048 12328 11112 12392
rect 11048 12168 11112 12232
rect 11048 12008 11112 12072
rect 11048 11848 11112 11912
rect 11048 11748 11112 11752
rect 11048 11692 11052 11748
rect 11052 11692 11108 11748
rect 11108 11692 11112 11748
rect 11048 11688 11112 11692
rect 11048 11588 11112 11592
rect 11048 11532 11052 11588
rect 11052 11532 11108 11588
rect 11108 11532 11112 11588
rect 11048 11528 11112 11532
rect 11048 11428 11112 11432
rect 11048 11372 11052 11428
rect 11052 11372 11108 11428
rect 11108 11372 11112 11428
rect 11048 11368 11112 11372
rect 11048 11268 11112 11272
rect 11048 11212 11052 11268
rect 11052 11212 11108 11268
rect 11108 11212 11112 11268
rect 11048 11208 11112 11212
rect 11048 11108 11112 11112
rect 11048 11052 11052 11108
rect 11052 11052 11108 11108
rect 11108 11052 11112 11108
rect 11048 11048 11112 11052
rect 11048 10948 11112 10952
rect 11048 10892 11052 10948
rect 11052 10892 11108 10948
rect 11108 10892 11112 10948
rect 11048 10888 11112 10892
rect 11048 10788 11112 10792
rect 11048 10732 11052 10788
rect 11052 10732 11108 10788
rect 11108 10732 11112 10788
rect 11048 10728 11112 10732
rect 11048 10628 11112 10632
rect 11048 10572 11052 10628
rect 11052 10572 11108 10628
rect 11108 10572 11112 10628
rect 11048 10568 11112 10572
rect 11048 10468 11112 10472
rect 11048 10412 11052 10468
rect 11052 10412 11108 10468
rect 11108 10412 11112 10468
rect 11048 10408 11112 10412
rect 11048 10308 11112 10312
rect 11048 10252 11052 10308
rect 11052 10252 11108 10308
rect 11108 10252 11112 10308
rect 11048 10248 11112 10252
rect 11048 10148 11112 10152
rect 11048 10092 11052 10148
rect 11052 10092 11108 10148
rect 11108 10092 11112 10148
rect 11048 10088 11112 10092
rect 11048 9988 11112 9992
rect 11048 9932 11052 9988
rect 11052 9932 11108 9988
rect 11108 9932 11112 9988
rect 11048 9928 11112 9932
rect 11048 9828 11112 9832
rect 11048 9772 11052 9828
rect 11052 9772 11108 9828
rect 11108 9772 11112 9828
rect 11048 9768 11112 9772
rect 11048 9608 11112 9672
rect 11048 9508 11112 9512
rect 11048 9452 11052 9508
rect 11052 9452 11108 9508
rect 11108 9452 11112 9508
rect 11048 9448 11112 9452
rect 11048 9348 11112 9352
rect 11048 9292 11052 9348
rect 11052 9292 11108 9348
rect 11108 9292 11112 9348
rect 11048 9288 11112 9292
rect 11048 9128 11112 9192
rect 11048 9028 11112 9032
rect 11048 8972 11052 9028
rect 11052 8972 11108 9028
rect 11108 8972 11112 9028
rect 11048 8968 11112 8972
rect 11048 8868 11112 8872
rect 11048 8812 11052 8868
rect 11052 8812 11108 8868
rect 11108 8812 11112 8868
rect 11048 8808 11112 8812
rect 11048 8708 11112 8712
rect 11048 8652 11052 8708
rect 11052 8652 11108 8708
rect 11108 8652 11112 8708
rect 11048 8648 11112 8652
rect 11048 8548 11112 8552
rect 11048 8492 11052 8548
rect 11052 8492 11108 8548
rect 11108 8492 11112 8548
rect 11048 8488 11112 8492
rect 11048 8388 11112 8392
rect 11048 8332 11052 8388
rect 11052 8332 11108 8388
rect 11108 8332 11112 8388
rect 11048 8328 11112 8332
rect 11048 8228 11112 8232
rect 11048 8172 11052 8228
rect 11052 8172 11108 8228
rect 11108 8172 11112 8228
rect 11048 8168 11112 8172
rect 11048 8068 11112 8072
rect 11048 8012 11052 8068
rect 11052 8012 11108 8068
rect 11108 8012 11112 8068
rect 11048 8008 11112 8012
rect 11048 7908 11112 7912
rect 11048 7852 11052 7908
rect 11052 7852 11108 7908
rect 11108 7852 11112 7908
rect 11048 7848 11112 7852
rect 11048 7748 11112 7752
rect 11048 7692 11052 7748
rect 11052 7692 11108 7748
rect 11108 7692 11112 7748
rect 11048 7688 11112 7692
rect 11048 7528 11112 7592
rect 11048 7428 11112 7432
rect 11048 7372 11052 7428
rect 11052 7372 11108 7428
rect 11108 7372 11112 7428
rect 11048 7368 11112 7372
rect 11048 7268 11112 7272
rect 11048 7212 11052 7268
rect 11052 7212 11108 7268
rect 11108 7212 11112 7268
rect 11048 7208 11112 7212
rect 11048 7048 11112 7112
rect 11048 6948 11112 6952
rect 11048 6892 11052 6948
rect 11052 6892 11108 6948
rect 11108 6892 11112 6948
rect 11048 6888 11112 6892
rect 11048 6788 11112 6792
rect 11048 6732 11052 6788
rect 11052 6732 11108 6788
rect 11108 6732 11112 6788
rect 11048 6728 11112 6732
rect 11048 6568 11112 6632
rect 11048 6468 11112 6472
rect 11048 6412 11052 6468
rect 11052 6412 11108 6468
rect 11108 6412 11112 6468
rect 11048 6408 11112 6412
rect 11048 6308 11112 6312
rect 11048 6252 11052 6308
rect 11052 6252 11108 6308
rect 11108 6252 11112 6308
rect 11048 6248 11112 6252
rect 11048 6148 11112 6152
rect 11048 6092 11052 6148
rect 11052 6092 11108 6148
rect 11108 6092 11112 6148
rect 11048 6088 11112 6092
rect 11048 5988 11112 5992
rect 11048 5932 11052 5988
rect 11052 5932 11108 5988
rect 11108 5932 11112 5988
rect 11048 5928 11112 5932
rect 11048 5828 11112 5832
rect 11048 5772 11052 5828
rect 11052 5772 11108 5828
rect 11108 5772 11112 5828
rect 11048 5768 11112 5772
rect 11048 5668 11112 5672
rect 11048 5612 11052 5668
rect 11052 5612 11108 5668
rect 11108 5612 11112 5668
rect 11048 5608 11112 5612
rect 11048 5508 11112 5512
rect 11048 5452 11052 5508
rect 11052 5452 11108 5508
rect 11108 5452 11112 5508
rect 11048 5448 11112 5452
rect 11048 5348 11112 5352
rect 11048 5292 11052 5348
rect 11052 5292 11108 5348
rect 11108 5292 11112 5348
rect 11048 5288 11112 5292
rect 11048 5188 11112 5192
rect 11048 5132 11052 5188
rect 11052 5132 11108 5188
rect 11108 5132 11112 5188
rect 11048 5128 11112 5132
rect 11048 5028 11112 5032
rect 11048 4972 11052 5028
rect 11052 4972 11108 5028
rect 11108 4972 11112 5028
rect 11048 4968 11112 4972
rect 11048 4868 11112 4872
rect 11048 4812 11052 4868
rect 11052 4812 11108 4868
rect 11108 4812 11112 4868
rect 11048 4808 11112 4812
rect 11048 4708 11112 4712
rect 11048 4652 11052 4708
rect 11052 4652 11108 4708
rect 11108 4652 11112 4708
rect 11048 4648 11112 4652
rect 11048 4548 11112 4552
rect 11048 4492 11052 4548
rect 11052 4492 11108 4548
rect 11108 4492 11112 4548
rect 11048 4488 11112 4492
rect 11048 4388 11112 4392
rect 11048 4332 11052 4388
rect 11052 4332 11108 4388
rect 11108 4332 11112 4388
rect 11048 4328 11112 4332
rect 11048 4228 11112 4232
rect 11048 4172 11052 4228
rect 11052 4172 11108 4228
rect 11108 4172 11112 4228
rect 11048 4168 11112 4172
rect 11048 4068 11112 4072
rect 11048 4012 11052 4068
rect 11052 4012 11108 4068
rect 11108 4012 11112 4068
rect 11048 4008 11112 4012
rect 11048 3908 11112 3912
rect 11048 3852 11052 3908
rect 11052 3852 11108 3908
rect 11108 3852 11112 3908
rect 11048 3848 11112 3852
rect 11048 3688 11112 3752
rect 11048 3528 11112 3592
rect 11048 3428 11112 3432
rect 11048 3372 11052 3428
rect 11052 3372 11108 3428
rect 11108 3372 11112 3428
rect 11048 3368 11112 3372
rect 11048 3268 11112 3272
rect 11048 3212 11052 3268
rect 11052 3212 11108 3268
rect 11108 3212 11112 3268
rect 11048 3208 11112 3212
rect 11048 3108 11112 3112
rect 11048 3052 11052 3108
rect 11052 3052 11108 3108
rect 11108 3052 11112 3108
rect 11048 3048 11112 3052
rect 11048 2948 11112 2952
rect 11048 2892 11052 2948
rect 11052 2892 11108 2948
rect 11108 2892 11112 2948
rect 11048 2888 11112 2892
rect 11048 2788 11112 2792
rect 11048 2732 11052 2788
rect 11052 2732 11108 2788
rect 11108 2732 11112 2788
rect 11048 2728 11112 2732
rect 11048 2628 11112 2632
rect 11048 2572 11052 2628
rect 11052 2572 11108 2628
rect 11108 2572 11112 2628
rect 11048 2568 11112 2572
rect 11048 2468 11112 2472
rect 11048 2412 11052 2468
rect 11052 2412 11108 2468
rect 11108 2412 11112 2468
rect 11048 2408 11112 2412
rect 11048 2308 11112 2312
rect 11048 2252 11052 2308
rect 11052 2252 11108 2308
rect 11108 2252 11112 2308
rect 11048 2248 11112 2252
rect 11048 2148 11112 2152
rect 11048 2092 11052 2148
rect 11052 2092 11108 2148
rect 11108 2092 11112 2148
rect 11048 2088 11112 2092
rect 11048 1988 11112 1992
rect 11048 1932 11052 1988
rect 11052 1932 11108 1988
rect 11108 1932 11112 1988
rect 11048 1928 11112 1932
rect 11048 1768 11112 1832
rect 11048 1668 11112 1672
rect 11048 1612 11052 1668
rect 11052 1612 11108 1668
rect 11108 1612 11112 1668
rect 11048 1608 11112 1612
rect 11048 1508 11112 1512
rect 11048 1452 11052 1508
rect 11052 1452 11108 1508
rect 11108 1452 11112 1508
rect 11048 1448 11112 1452
rect 11048 1348 11112 1352
rect 11048 1292 11052 1348
rect 11052 1292 11108 1348
rect 11108 1292 11112 1348
rect 11048 1288 11112 1292
rect 11048 1188 11112 1192
rect 11048 1132 11052 1188
rect 11052 1132 11108 1188
rect 11108 1132 11112 1188
rect 11048 1128 11112 1132
rect 11048 1028 11112 1032
rect 11048 972 11052 1028
rect 11052 972 11108 1028
rect 11108 972 11112 1028
rect 11048 968 11112 972
rect 11048 808 11112 872
rect 11048 648 11112 712
rect 11048 548 11112 552
rect 11048 492 11052 548
rect 11052 492 11108 548
rect 11108 492 11112 548
rect 11048 488 11112 492
rect 11048 388 11112 392
rect 11048 332 11052 388
rect 11052 332 11108 388
rect 11108 332 11112 388
rect 11048 328 11112 332
rect 11048 228 11112 232
rect 11048 172 11052 228
rect 11052 172 11108 228
rect 11108 172 11112 228
rect 11048 168 11112 172
rect 11048 68 11112 72
rect 11048 12 11052 68
rect 11052 12 11108 68
rect 11108 12 11112 68
rect 11048 8 11112 12
rect 10728 -1112 10792 -1048
rect 10728 -1192 10792 -1128
rect 10728 -1272 10792 -1208
rect 10728 -1352 10792 -1288
rect 10728 -1432 10792 -1368
rect 11368 31428 11432 31432
rect 11368 31372 11372 31428
rect 11372 31372 11428 31428
rect 11428 31372 11432 31428
rect 11368 31368 11432 31372
rect 11368 31268 11432 31272
rect 11368 31212 11372 31268
rect 11372 31212 11428 31268
rect 11428 31212 11432 31268
rect 11368 31208 11432 31212
rect 11368 31108 11432 31112
rect 11368 31052 11372 31108
rect 11372 31052 11428 31108
rect 11428 31052 11432 31108
rect 11368 31048 11432 31052
rect 11368 30948 11432 30952
rect 11368 30892 11372 30948
rect 11372 30892 11428 30948
rect 11428 30892 11432 30948
rect 11368 30888 11432 30892
rect 11368 30788 11432 30792
rect 11368 30732 11372 30788
rect 11372 30732 11428 30788
rect 11428 30732 11432 30788
rect 11368 30728 11432 30732
rect 11368 30628 11432 30632
rect 11368 30572 11372 30628
rect 11372 30572 11428 30628
rect 11428 30572 11432 30628
rect 11368 30568 11432 30572
rect 11368 30468 11432 30472
rect 11368 30412 11372 30468
rect 11372 30412 11428 30468
rect 11428 30412 11432 30468
rect 11368 30408 11432 30412
rect 11368 30308 11432 30312
rect 11368 30252 11372 30308
rect 11372 30252 11428 30308
rect 11428 30252 11432 30308
rect 11368 30248 11432 30252
rect 11368 30088 11432 30152
rect 11368 29988 11432 29992
rect 11368 29932 11372 29988
rect 11372 29932 11428 29988
rect 11428 29932 11432 29988
rect 11368 29928 11432 29932
rect 11368 29828 11432 29832
rect 11368 29772 11372 29828
rect 11372 29772 11428 29828
rect 11428 29772 11432 29828
rect 11368 29768 11432 29772
rect 11368 29668 11432 29672
rect 11368 29612 11372 29668
rect 11372 29612 11428 29668
rect 11428 29612 11432 29668
rect 11368 29608 11432 29612
rect 11368 29508 11432 29512
rect 11368 29452 11372 29508
rect 11372 29452 11428 29508
rect 11428 29452 11432 29508
rect 11368 29448 11432 29452
rect 11368 29348 11432 29352
rect 11368 29292 11372 29348
rect 11372 29292 11428 29348
rect 11428 29292 11432 29348
rect 11368 29288 11432 29292
rect 11368 29188 11432 29192
rect 11368 29132 11372 29188
rect 11372 29132 11428 29188
rect 11428 29132 11432 29188
rect 11368 29128 11432 29132
rect 11368 29028 11432 29032
rect 11368 28972 11372 29028
rect 11372 28972 11428 29028
rect 11428 28972 11432 29028
rect 11368 28968 11432 28972
rect 11368 28868 11432 28872
rect 11368 28812 11372 28868
rect 11372 28812 11428 28868
rect 11428 28812 11432 28868
rect 11368 28808 11432 28812
rect 11368 28648 11432 28712
rect 11368 28488 11432 28552
rect 11368 28328 11432 28392
rect 11368 28168 11432 28232
rect 11368 28068 11432 28072
rect 11368 28012 11372 28068
rect 11372 28012 11428 28068
rect 11428 28012 11432 28068
rect 11368 28008 11432 28012
rect 11368 27908 11432 27912
rect 11368 27852 11372 27908
rect 11372 27852 11428 27908
rect 11428 27852 11432 27908
rect 11368 27848 11432 27852
rect 11368 27748 11432 27752
rect 11368 27692 11372 27748
rect 11372 27692 11428 27748
rect 11428 27692 11432 27748
rect 11368 27688 11432 27692
rect 11368 27588 11432 27592
rect 11368 27532 11372 27588
rect 11372 27532 11428 27588
rect 11428 27532 11432 27588
rect 11368 27528 11432 27532
rect 11368 27428 11432 27432
rect 11368 27372 11372 27428
rect 11372 27372 11428 27428
rect 11428 27372 11432 27428
rect 11368 27368 11432 27372
rect 11368 27268 11432 27272
rect 11368 27212 11372 27268
rect 11372 27212 11428 27268
rect 11428 27212 11432 27268
rect 11368 27208 11432 27212
rect 11368 27108 11432 27112
rect 11368 27052 11372 27108
rect 11372 27052 11428 27108
rect 11428 27052 11432 27108
rect 11368 27048 11432 27052
rect 11368 26948 11432 26952
rect 11368 26892 11372 26948
rect 11372 26892 11428 26948
rect 11428 26892 11432 26948
rect 11368 26888 11432 26892
rect 11368 26728 11432 26792
rect 11368 26568 11432 26632
rect 11368 26408 11432 26472
rect 11368 26248 11432 26312
rect 11368 26148 11432 26152
rect 11368 26092 11372 26148
rect 11372 26092 11428 26148
rect 11428 26092 11432 26148
rect 11368 26088 11432 26092
rect 11368 25988 11432 25992
rect 11368 25932 11372 25988
rect 11372 25932 11428 25988
rect 11428 25932 11432 25988
rect 11368 25928 11432 25932
rect 11368 25828 11432 25832
rect 11368 25772 11372 25828
rect 11372 25772 11428 25828
rect 11428 25772 11432 25828
rect 11368 25768 11432 25772
rect 11368 25668 11432 25672
rect 11368 25612 11372 25668
rect 11372 25612 11428 25668
rect 11428 25612 11432 25668
rect 11368 25608 11432 25612
rect 11368 25508 11432 25512
rect 11368 25452 11372 25508
rect 11372 25452 11428 25508
rect 11428 25452 11432 25508
rect 11368 25448 11432 25452
rect 11368 25348 11432 25352
rect 11368 25292 11372 25348
rect 11372 25292 11428 25348
rect 11428 25292 11432 25348
rect 11368 25288 11432 25292
rect 11368 25188 11432 25192
rect 11368 25132 11372 25188
rect 11372 25132 11428 25188
rect 11428 25132 11432 25188
rect 11368 25128 11432 25132
rect 11368 25028 11432 25032
rect 11368 24972 11372 25028
rect 11372 24972 11428 25028
rect 11428 24972 11432 25028
rect 11368 24968 11432 24972
rect 11368 24808 11432 24872
rect 11368 24708 11432 24712
rect 11368 24652 11372 24708
rect 11372 24652 11428 24708
rect 11428 24652 11432 24708
rect 11368 24648 11432 24652
rect 11368 24548 11432 24552
rect 11368 24492 11372 24548
rect 11372 24492 11428 24548
rect 11428 24492 11432 24548
rect 11368 24488 11432 24492
rect 11368 24388 11432 24392
rect 11368 24332 11372 24388
rect 11372 24332 11428 24388
rect 11428 24332 11432 24388
rect 11368 24328 11432 24332
rect 11368 24228 11432 24232
rect 11368 24172 11372 24228
rect 11372 24172 11428 24228
rect 11428 24172 11432 24228
rect 11368 24168 11432 24172
rect 11368 24068 11432 24072
rect 11368 24012 11372 24068
rect 11372 24012 11428 24068
rect 11428 24012 11432 24068
rect 11368 24008 11432 24012
rect 11368 23908 11432 23912
rect 11368 23852 11372 23908
rect 11372 23852 11428 23908
rect 11428 23852 11432 23908
rect 11368 23848 11432 23852
rect 11368 23748 11432 23752
rect 11368 23692 11372 23748
rect 11372 23692 11428 23748
rect 11428 23692 11432 23748
rect 11368 23688 11432 23692
rect 11368 23588 11432 23592
rect 11368 23532 11372 23588
rect 11372 23532 11428 23588
rect 11428 23532 11432 23588
rect 11368 23528 11432 23532
rect 11368 23428 11432 23432
rect 11368 23372 11372 23428
rect 11372 23372 11428 23428
rect 11428 23372 11432 23428
rect 11368 23368 11432 23372
rect 11368 23268 11432 23272
rect 11368 23212 11372 23268
rect 11372 23212 11428 23268
rect 11428 23212 11432 23268
rect 11368 23208 11432 23212
rect 11368 23108 11432 23112
rect 11368 23052 11372 23108
rect 11372 23052 11428 23108
rect 11428 23052 11432 23108
rect 11368 23048 11432 23052
rect 11368 22948 11432 22952
rect 11368 22892 11372 22948
rect 11372 22892 11428 22948
rect 11428 22892 11432 22948
rect 11368 22888 11432 22892
rect 11368 22788 11432 22792
rect 11368 22732 11372 22788
rect 11372 22732 11428 22788
rect 11428 22732 11432 22788
rect 11368 22728 11432 22732
rect 11368 22628 11432 22632
rect 11368 22572 11372 22628
rect 11372 22572 11428 22628
rect 11428 22572 11432 22628
rect 11368 22568 11432 22572
rect 11368 22468 11432 22472
rect 11368 22412 11372 22468
rect 11372 22412 11428 22468
rect 11428 22412 11432 22468
rect 11368 22408 11432 22412
rect 11368 22308 11432 22312
rect 11368 22252 11372 22308
rect 11372 22252 11428 22308
rect 11428 22252 11432 22308
rect 11368 22248 11432 22252
rect 11368 22148 11432 22152
rect 11368 22092 11372 22148
rect 11372 22092 11428 22148
rect 11428 22092 11432 22148
rect 11368 22088 11432 22092
rect 11368 21928 11432 21992
rect 11368 21828 11432 21832
rect 11368 21772 11372 21828
rect 11372 21772 11428 21828
rect 11428 21772 11432 21828
rect 11368 21768 11432 21772
rect 11368 21668 11432 21672
rect 11368 21612 11372 21668
rect 11372 21612 11428 21668
rect 11428 21612 11432 21668
rect 11368 21608 11432 21612
rect 11368 21508 11432 21512
rect 11368 21452 11372 21508
rect 11372 21452 11428 21508
rect 11428 21452 11432 21508
rect 11368 21448 11432 21452
rect 11368 21348 11432 21352
rect 11368 21292 11372 21348
rect 11372 21292 11428 21348
rect 11428 21292 11432 21348
rect 11368 21288 11432 21292
rect 11368 21188 11432 21192
rect 11368 21132 11372 21188
rect 11372 21132 11428 21188
rect 11428 21132 11432 21188
rect 11368 21128 11432 21132
rect 11368 21028 11432 21032
rect 11368 20972 11372 21028
rect 11372 20972 11428 21028
rect 11428 20972 11432 21028
rect 11368 20968 11432 20972
rect 11368 20868 11432 20872
rect 11368 20812 11372 20868
rect 11372 20812 11428 20868
rect 11428 20812 11432 20868
rect 11368 20808 11432 20812
rect 11368 20708 11432 20712
rect 11368 20652 11372 20708
rect 11372 20652 11428 20708
rect 11428 20652 11432 20708
rect 11368 20648 11432 20652
rect 11368 20488 11432 20552
rect 11368 20328 11432 20392
rect 11368 20168 11432 20232
rect 11368 20008 11432 20072
rect 11368 19908 11432 19912
rect 11368 19852 11372 19908
rect 11372 19852 11428 19908
rect 11428 19852 11432 19908
rect 11368 19848 11432 19852
rect 11368 19748 11432 19752
rect 11368 19692 11372 19748
rect 11372 19692 11428 19748
rect 11428 19692 11432 19748
rect 11368 19688 11432 19692
rect 11368 19588 11432 19592
rect 11368 19532 11372 19588
rect 11372 19532 11428 19588
rect 11428 19532 11432 19588
rect 11368 19528 11432 19532
rect 11368 19428 11432 19432
rect 11368 19372 11372 19428
rect 11372 19372 11428 19428
rect 11428 19372 11432 19428
rect 11368 19368 11432 19372
rect 11368 19268 11432 19272
rect 11368 19212 11372 19268
rect 11372 19212 11428 19268
rect 11428 19212 11432 19268
rect 11368 19208 11432 19212
rect 11368 19108 11432 19112
rect 11368 19052 11372 19108
rect 11372 19052 11428 19108
rect 11428 19052 11432 19108
rect 11368 19048 11432 19052
rect 11368 18948 11432 18952
rect 11368 18892 11372 18948
rect 11372 18892 11428 18948
rect 11428 18892 11432 18948
rect 11368 18888 11432 18892
rect 11368 18788 11432 18792
rect 11368 18732 11372 18788
rect 11372 18732 11428 18788
rect 11428 18732 11432 18788
rect 11368 18728 11432 18732
rect 11368 18568 11432 18632
rect 11368 18408 11432 18472
rect 11368 18248 11432 18312
rect 11368 18088 11432 18152
rect 11368 17988 11432 17992
rect 11368 17932 11372 17988
rect 11372 17932 11428 17988
rect 11428 17932 11432 17988
rect 11368 17928 11432 17932
rect 11368 17828 11432 17832
rect 11368 17772 11372 17828
rect 11372 17772 11428 17828
rect 11428 17772 11432 17828
rect 11368 17768 11432 17772
rect 11368 17668 11432 17672
rect 11368 17612 11372 17668
rect 11372 17612 11428 17668
rect 11428 17612 11432 17668
rect 11368 17608 11432 17612
rect 11368 17508 11432 17512
rect 11368 17452 11372 17508
rect 11372 17452 11428 17508
rect 11428 17452 11432 17508
rect 11368 17448 11432 17452
rect 11368 17348 11432 17352
rect 11368 17292 11372 17348
rect 11372 17292 11428 17348
rect 11428 17292 11432 17348
rect 11368 17288 11432 17292
rect 11368 17188 11432 17192
rect 11368 17132 11372 17188
rect 11372 17132 11428 17188
rect 11428 17132 11432 17188
rect 11368 17128 11432 17132
rect 11368 17028 11432 17032
rect 11368 16972 11372 17028
rect 11372 16972 11428 17028
rect 11428 16972 11432 17028
rect 11368 16968 11432 16972
rect 11368 16868 11432 16872
rect 11368 16812 11372 16868
rect 11372 16812 11428 16868
rect 11428 16812 11432 16868
rect 11368 16808 11432 16812
rect 11368 16648 11432 16712
rect 11368 16548 11432 16552
rect 11368 16492 11372 16548
rect 11372 16492 11428 16548
rect 11428 16492 11432 16548
rect 11368 16488 11432 16492
rect 11368 16388 11432 16392
rect 11368 16332 11372 16388
rect 11372 16332 11428 16388
rect 11428 16332 11432 16388
rect 11368 16328 11432 16332
rect 11368 16228 11432 16232
rect 11368 16172 11372 16228
rect 11372 16172 11428 16228
rect 11428 16172 11432 16228
rect 11368 16168 11432 16172
rect 11368 16068 11432 16072
rect 11368 16012 11372 16068
rect 11372 16012 11428 16068
rect 11428 16012 11432 16068
rect 11368 16008 11432 16012
rect 11368 15908 11432 15912
rect 11368 15852 11372 15908
rect 11372 15852 11428 15908
rect 11428 15852 11432 15908
rect 11368 15848 11432 15852
rect 11368 15748 11432 15752
rect 11368 15692 11372 15748
rect 11372 15692 11428 15748
rect 11428 15692 11432 15748
rect 11368 15688 11432 15692
rect 11368 15588 11432 15592
rect 11368 15532 11372 15588
rect 11372 15532 11428 15588
rect 11428 15532 11432 15588
rect 11368 15528 11432 15532
rect 11368 15428 11432 15432
rect 11368 15372 11372 15428
rect 11372 15372 11428 15428
rect 11428 15372 11432 15428
rect 11368 15368 11432 15372
rect 11368 15268 11432 15272
rect 11368 15212 11372 15268
rect 11372 15212 11428 15268
rect 11428 15212 11432 15268
rect 11368 15208 11432 15212
rect 11368 15108 11432 15112
rect 11368 15052 11372 15108
rect 11372 15052 11428 15108
rect 11428 15052 11432 15108
rect 11368 15048 11432 15052
rect 11368 14948 11432 14952
rect 11368 14892 11372 14948
rect 11372 14892 11428 14948
rect 11428 14892 11432 14948
rect 11368 14888 11432 14892
rect 11368 14788 11432 14792
rect 11368 14732 11372 14788
rect 11372 14732 11428 14788
rect 11428 14732 11432 14788
rect 11368 14728 11432 14732
rect 11368 14628 11432 14632
rect 11368 14572 11372 14628
rect 11372 14572 11428 14628
rect 11428 14572 11432 14628
rect 11368 14568 11432 14572
rect 11368 14468 11432 14472
rect 11368 14412 11372 14468
rect 11372 14412 11428 14468
rect 11428 14412 11432 14468
rect 11368 14408 11432 14412
rect 11368 14308 11432 14312
rect 11368 14252 11372 14308
rect 11372 14252 11428 14308
rect 11428 14252 11432 14308
rect 11368 14248 11432 14252
rect 11368 14148 11432 14152
rect 11368 14092 11372 14148
rect 11372 14092 11428 14148
rect 11428 14092 11432 14148
rect 11368 14088 11432 14092
rect 11368 13988 11432 13992
rect 11368 13932 11372 13988
rect 11372 13932 11428 13988
rect 11428 13932 11432 13988
rect 11368 13928 11432 13932
rect 11368 13768 11432 13832
rect 11368 13668 11432 13672
rect 11368 13612 11372 13668
rect 11372 13612 11428 13668
rect 11428 13612 11432 13668
rect 11368 13608 11432 13612
rect 11368 13508 11432 13512
rect 11368 13452 11372 13508
rect 11372 13452 11428 13508
rect 11428 13452 11432 13508
rect 11368 13448 11432 13452
rect 11368 13348 11432 13352
rect 11368 13292 11372 13348
rect 11372 13292 11428 13348
rect 11428 13292 11432 13348
rect 11368 13288 11432 13292
rect 11368 13188 11432 13192
rect 11368 13132 11372 13188
rect 11372 13132 11428 13188
rect 11428 13132 11432 13188
rect 11368 13128 11432 13132
rect 11368 13028 11432 13032
rect 11368 12972 11372 13028
rect 11372 12972 11428 13028
rect 11428 12972 11432 13028
rect 11368 12968 11432 12972
rect 11368 12868 11432 12872
rect 11368 12812 11372 12868
rect 11372 12812 11428 12868
rect 11428 12812 11432 12868
rect 11368 12808 11432 12812
rect 11368 12708 11432 12712
rect 11368 12652 11372 12708
rect 11372 12652 11428 12708
rect 11428 12652 11432 12708
rect 11368 12648 11432 12652
rect 11368 12548 11432 12552
rect 11368 12492 11372 12548
rect 11372 12492 11428 12548
rect 11428 12492 11432 12548
rect 11368 12488 11432 12492
rect 11368 12328 11432 12392
rect 11368 12168 11432 12232
rect 11368 12008 11432 12072
rect 11368 11848 11432 11912
rect 11368 11748 11432 11752
rect 11368 11692 11372 11748
rect 11372 11692 11428 11748
rect 11428 11692 11432 11748
rect 11368 11688 11432 11692
rect 11368 11588 11432 11592
rect 11368 11532 11372 11588
rect 11372 11532 11428 11588
rect 11428 11532 11432 11588
rect 11368 11528 11432 11532
rect 11368 11428 11432 11432
rect 11368 11372 11372 11428
rect 11372 11372 11428 11428
rect 11428 11372 11432 11428
rect 11368 11368 11432 11372
rect 11368 11268 11432 11272
rect 11368 11212 11372 11268
rect 11372 11212 11428 11268
rect 11428 11212 11432 11268
rect 11368 11208 11432 11212
rect 11368 11108 11432 11112
rect 11368 11052 11372 11108
rect 11372 11052 11428 11108
rect 11428 11052 11432 11108
rect 11368 11048 11432 11052
rect 11368 10948 11432 10952
rect 11368 10892 11372 10948
rect 11372 10892 11428 10948
rect 11428 10892 11432 10948
rect 11368 10888 11432 10892
rect 11368 10788 11432 10792
rect 11368 10732 11372 10788
rect 11372 10732 11428 10788
rect 11428 10732 11432 10788
rect 11368 10728 11432 10732
rect 11368 10628 11432 10632
rect 11368 10572 11372 10628
rect 11372 10572 11428 10628
rect 11428 10572 11432 10628
rect 11368 10568 11432 10572
rect 11368 10468 11432 10472
rect 11368 10412 11372 10468
rect 11372 10412 11428 10468
rect 11428 10412 11432 10468
rect 11368 10408 11432 10412
rect 11368 10308 11432 10312
rect 11368 10252 11372 10308
rect 11372 10252 11428 10308
rect 11428 10252 11432 10308
rect 11368 10248 11432 10252
rect 11368 10148 11432 10152
rect 11368 10092 11372 10148
rect 11372 10092 11428 10148
rect 11428 10092 11432 10148
rect 11368 10088 11432 10092
rect 11368 9988 11432 9992
rect 11368 9932 11372 9988
rect 11372 9932 11428 9988
rect 11428 9932 11432 9988
rect 11368 9928 11432 9932
rect 11368 9828 11432 9832
rect 11368 9772 11372 9828
rect 11372 9772 11428 9828
rect 11428 9772 11432 9828
rect 11368 9768 11432 9772
rect 11368 9608 11432 9672
rect 11368 9508 11432 9512
rect 11368 9452 11372 9508
rect 11372 9452 11428 9508
rect 11428 9452 11432 9508
rect 11368 9448 11432 9452
rect 11368 9348 11432 9352
rect 11368 9292 11372 9348
rect 11372 9292 11428 9348
rect 11428 9292 11432 9348
rect 11368 9288 11432 9292
rect 11368 9128 11432 9192
rect 11368 9028 11432 9032
rect 11368 8972 11372 9028
rect 11372 8972 11428 9028
rect 11428 8972 11432 9028
rect 11368 8968 11432 8972
rect 11368 8868 11432 8872
rect 11368 8812 11372 8868
rect 11372 8812 11428 8868
rect 11428 8812 11432 8868
rect 11368 8808 11432 8812
rect 11368 8708 11432 8712
rect 11368 8652 11372 8708
rect 11372 8652 11428 8708
rect 11428 8652 11432 8708
rect 11368 8648 11432 8652
rect 11368 8548 11432 8552
rect 11368 8492 11372 8548
rect 11372 8492 11428 8548
rect 11428 8492 11432 8548
rect 11368 8488 11432 8492
rect 11368 8388 11432 8392
rect 11368 8332 11372 8388
rect 11372 8332 11428 8388
rect 11428 8332 11432 8388
rect 11368 8328 11432 8332
rect 11368 8228 11432 8232
rect 11368 8172 11372 8228
rect 11372 8172 11428 8228
rect 11428 8172 11432 8228
rect 11368 8168 11432 8172
rect 11368 8068 11432 8072
rect 11368 8012 11372 8068
rect 11372 8012 11428 8068
rect 11428 8012 11432 8068
rect 11368 8008 11432 8012
rect 11368 7908 11432 7912
rect 11368 7852 11372 7908
rect 11372 7852 11428 7908
rect 11428 7852 11432 7908
rect 11368 7848 11432 7852
rect 11368 7748 11432 7752
rect 11368 7692 11372 7748
rect 11372 7692 11428 7748
rect 11428 7692 11432 7748
rect 11368 7688 11432 7692
rect 11368 7528 11432 7592
rect 11368 7428 11432 7432
rect 11368 7372 11372 7428
rect 11372 7372 11428 7428
rect 11428 7372 11432 7428
rect 11368 7368 11432 7372
rect 11368 7268 11432 7272
rect 11368 7212 11372 7268
rect 11372 7212 11428 7268
rect 11428 7212 11432 7268
rect 11368 7208 11432 7212
rect 11368 7048 11432 7112
rect 11368 6948 11432 6952
rect 11368 6892 11372 6948
rect 11372 6892 11428 6948
rect 11428 6892 11432 6948
rect 11368 6888 11432 6892
rect 11368 6788 11432 6792
rect 11368 6732 11372 6788
rect 11372 6732 11428 6788
rect 11428 6732 11432 6788
rect 11368 6728 11432 6732
rect 11368 6568 11432 6632
rect 11368 6468 11432 6472
rect 11368 6412 11372 6468
rect 11372 6412 11428 6468
rect 11428 6412 11432 6468
rect 11368 6408 11432 6412
rect 11368 6308 11432 6312
rect 11368 6252 11372 6308
rect 11372 6252 11428 6308
rect 11428 6252 11432 6308
rect 11368 6248 11432 6252
rect 11368 6148 11432 6152
rect 11368 6092 11372 6148
rect 11372 6092 11428 6148
rect 11428 6092 11432 6148
rect 11368 6088 11432 6092
rect 11368 5988 11432 5992
rect 11368 5932 11372 5988
rect 11372 5932 11428 5988
rect 11428 5932 11432 5988
rect 11368 5928 11432 5932
rect 11368 5828 11432 5832
rect 11368 5772 11372 5828
rect 11372 5772 11428 5828
rect 11428 5772 11432 5828
rect 11368 5768 11432 5772
rect 11368 5668 11432 5672
rect 11368 5612 11372 5668
rect 11372 5612 11428 5668
rect 11428 5612 11432 5668
rect 11368 5608 11432 5612
rect 11368 5508 11432 5512
rect 11368 5452 11372 5508
rect 11372 5452 11428 5508
rect 11428 5452 11432 5508
rect 11368 5448 11432 5452
rect 11368 5348 11432 5352
rect 11368 5292 11372 5348
rect 11372 5292 11428 5348
rect 11428 5292 11432 5348
rect 11368 5288 11432 5292
rect 11368 5188 11432 5192
rect 11368 5132 11372 5188
rect 11372 5132 11428 5188
rect 11428 5132 11432 5188
rect 11368 5128 11432 5132
rect 11368 5028 11432 5032
rect 11368 4972 11372 5028
rect 11372 4972 11428 5028
rect 11428 4972 11432 5028
rect 11368 4968 11432 4972
rect 11368 4868 11432 4872
rect 11368 4812 11372 4868
rect 11372 4812 11428 4868
rect 11428 4812 11432 4868
rect 11368 4808 11432 4812
rect 11368 4708 11432 4712
rect 11368 4652 11372 4708
rect 11372 4652 11428 4708
rect 11428 4652 11432 4708
rect 11368 4648 11432 4652
rect 11368 4548 11432 4552
rect 11368 4492 11372 4548
rect 11372 4492 11428 4548
rect 11428 4492 11432 4548
rect 11368 4488 11432 4492
rect 11368 4388 11432 4392
rect 11368 4332 11372 4388
rect 11372 4332 11428 4388
rect 11428 4332 11432 4388
rect 11368 4328 11432 4332
rect 11368 4228 11432 4232
rect 11368 4172 11372 4228
rect 11372 4172 11428 4228
rect 11428 4172 11432 4228
rect 11368 4168 11432 4172
rect 11368 4068 11432 4072
rect 11368 4012 11372 4068
rect 11372 4012 11428 4068
rect 11428 4012 11432 4068
rect 11368 4008 11432 4012
rect 11368 3908 11432 3912
rect 11368 3852 11372 3908
rect 11372 3852 11428 3908
rect 11428 3852 11432 3908
rect 11368 3848 11432 3852
rect 11368 3688 11432 3752
rect 11368 3528 11432 3592
rect 11368 3428 11432 3432
rect 11368 3372 11372 3428
rect 11372 3372 11428 3428
rect 11428 3372 11432 3428
rect 11368 3368 11432 3372
rect 11368 3268 11432 3272
rect 11368 3212 11372 3268
rect 11372 3212 11428 3268
rect 11428 3212 11432 3268
rect 11368 3208 11432 3212
rect 11368 3108 11432 3112
rect 11368 3052 11372 3108
rect 11372 3052 11428 3108
rect 11428 3052 11432 3108
rect 11368 3048 11432 3052
rect 11368 2948 11432 2952
rect 11368 2892 11372 2948
rect 11372 2892 11428 2948
rect 11428 2892 11432 2948
rect 11368 2888 11432 2892
rect 11368 2788 11432 2792
rect 11368 2732 11372 2788
rect 11372 2732 11428 2788
rect 11428 2732 11432 2788
rect 11368 2728 11432 2732
rect 11368 2628 11432 2632
rect 11368 2572 11372 2628
rect 11372 2572 11428 2628
rect 11428 2572 11432 2628
rect 11368 2568 11432 2572
rect 11368 2468 11432 2472
rect 11368 2412 11372 2468
rect 11372 2412 11428 2468
rect 11428 2412 11432 2468
rect 11368 2408 11432 2412
rect 11368 2308 11432 2312
rect 11368 2252 11372 2308
rect 11372 2252 11428 2308
rect 11428 2252 11432 2308
rect 11368 2248 11432 2252
rect 11368 2148 11432 2152
rect 11368 2092 11372 2148
rect 11372 2092 11428 2148
rect 11428 2092 11432 2148
rect 11368 2088 11432 2092
rect 11368 1988 11432 1992
rect 11368 1932 11372 1988
rect 11372 1932 11428 1988
rect 11428 1932 11432 1988
rect 11368 1928 11432 1932
rect 11368 1768 11432 1832
rect 11368 1668 11432 1672
rect 11368 1612 11372 1668
rect 11372 1612 11428 1668
rect 11428 1612 11432 1668
rect 11368 1608 11432 1612
rect 11368 1508 11432 1512
rect 11368 1452 11372 1508
rect 11372 1452 11428 1508
rect 11428 1452 11432 1508
rect 11368 1448 11432 1452
rect 11368 1348 11432 1352
rect 11368 1292 11372 1348
rect 11372 1292 11428 1348
rect 11428 1292 11432 1348
rect 11368 1288 11432 1292
rect 11368 1188 11432 1192
rect 11368 1132 11372 1188
rect 11372 1132 11428 1188
rect 11428 1132 11432 1188
rect 11368 1128 11432 1132
rect 11368 1028 11432 1032
rect 11368 972 11372 1028
rect 11372 972 11428 1028
rect 11428 972 11432 1028
rect 11368 968 11432 972
rect 11368 808 11432 872
rect 11368 648 11432 712
rect 11368 548 11432 552
rect 11368 492 11372 548
rect 11372 492 11428 548
rect 11428 492 11432 548
rect 11368 488 11432 492
rect 11368 388 11432 392
rect 11368 332 11372 388
rect 11372 332 11428 388
rect 11428 332 11432 388
rect 11368 328 11432 332
rect 11368 228 11432 232
rect 11368 172 11372 228
rect 11372 172 11428 228
rect 11428 172 11432 228
rect 11368 168 11432 172
rect 11368 68 11432 72
rect 11368 12 11372 68
rect 11372 12 11428 68
rect 11428 12 11432 68
rect 11368 8 11432 12
rect 11048 -1112 11112 -1048
rect 11048 -1192 11112 -1128
rect 11048 -1272 11112 -1208
rect 11048 -1352 11112 -1288
rect 11048 -1432 11112 -1368
rect 11368 -1112 11432 -1048
rect 11368 -1192 11432 -1128
rect 11368 -1272 11432 -1208
rect 11368 -1352 11432 -1288
rect 11368 -1432 11432 -1368
rect 11528 31428 11592 31432
rect 11528 31372 11532 31428
rect 11532 31372 11588 31428
rect 11588 31372 11592 31428
rect 11528 31368 11592 31372
rect 11528 31268 11592 31272
rect 11528 31212 11532 31268
rect 11532 31212 11588 31268
rect 11588 31212 11592 31268
rect 11528 31208 11592 31212
rect 11528 31108 11592 31112
rect 11528 31052 11532 31108
rect 11532 31052 11588 31108
rect 11588 31052 11592 31108
rect 11528 31048 11592 31052
rect 11528 30948 11592 30952
rect 11528 30892 11532 30948
rect 11532 30892 11588 30948
rect 11588 30892 11592 30948
rect 11528 30888 11592 30892
rect 11528 30788 11592 30792
rect 11528 30732 11532 30788
rect 11532 30732 11588 30788
rect 11588 30732 11592 30788
rect 11528 30728 11592 30732
rect 11528 30628 11592 30632
rect 11528 30572 11532 30628
rect 11532 30572 11588 30628
rect 11588 30572 11592 30628
rect 11528 30568 11592 30572
rect 11528 30468 11592 30472
rect 11528 30412 11532 30468
rect 11532 30412 11588 30468
rect 11588 30412 11592 30468
rect 11528 30408 11592 30412
rect 11528 30308 11592 30312
rect 11528 30252 11532 30308
rect 11532 30252 11588 30308
rect 11588 30252 11592 30308
rect 11528 30248 11592 30252
rect 11528 30088 11592 30152
rect 11528 29988 11592 29992
rect 11528 29932 11532 29988
rect 11532 29932 11588 29988
rect 11588 29932 11592 29988
rect 11528 29928 11592 29932
rect 11528 29828 11592 29832
rect 11528 29772 11532 29828
rect 11532 29772 11588 29828
rect 11588 29772 11592 29828
rect 11528 29768 11592 29772
rect 11528 29668 11592 29672
rect 11528 29612 11532 29668
rect 11532 29612 11588 29668
rect 11588 29612 11592 29668
rect 11528 29608 11592 29612
rect 11528 29508 11592 29512
rect 11528 29452 11532 29508
rect 11532 29452 11588 29508
rect 11588 29452 11592 29508
rect 11528 29448 11592 29452
rect 11528 29348 11592 29352
rect 11528 29292 11532 29348
rect 11532 29292 11588 29348
rect 11588 29292 11592 29348
rect 11528 29288 11592 29292
rect 11528 29188 11592 29192
rect 11528 29132 11532 29188
rect 11532 29132 11588 29188
rect 11588 29132 11592 29188
rect 11528 29128 11592 29132
rect 11528 29028 11592 29032
rect 11528 28972 11532 29028
rect 11532 28972 11588 29028
rect 11588 28972 11592 29028
rect 11528 28968 11592 28972
rect 11528 28868 11592 28872
rect 11528 28812 11532 28868
rect 11532 28812 11588 28868
rect 11588 28812 11592 28868
rect 11528 28808 11592 28812
rect 11528 28648 11592 28712
rect 11528 28488 11592 28552
rect 11528 28328 11592 28392
rect 11528 28168 11592 28232
rect 11528 28068 11592 28072
rect 11528 28012 11532 28068
rect 11532 28012 11588 28068
rect 11588 28012 11592 28068
rect 11528 28008 11592 28012
rect 11528 27908 11592 27912
rect 11528 27852 11532 27908
rect 11532 27852 11588 27908
rect 11588 27852 11592 27908
rect 11528 27848 11592 27852
rect 11528 27748 11592 27752
rect 11528 27692 11532 27748
rect 11532 27692 11588 27748
rect 11588 27692 11592 27748
rect 11528 27688 11592 27692
rect 11528 27588 11592 27592
rect 11528 27532 11532 27588
rect 11532 27532 11588 27588
rect 11588 27532 11592 27588
rect 11528 27528 11592 27532
rect 11528 27428 11592 27432
rect 11528 27372 11532 27428
rect 11532 27372 11588 27428
rect 11588 27372 11592 27428
rect 11528 27368 11592 27372
rect 11528 27268 11592 27272
rect 11528 27212 11532 27268
rect 11532 27212 11588 27268
rect 11588 27212 11592 27268
rect 11528 27208 11592 27212
rect 11528 27108 11592 27112
rect 11528 27052 11532 27108
rect 11532 27052 11588 27108
rect 11588 27052 11592 27108
rect 11528 27048 11592 27052
rect 11528 26948 11592 26952
rect 11528 26892 11532 26948
rect 11532 26892 11588 26948
rect 11588 26892 11592 26948
rect 11528 26888 11592 26892
rect 11528 26728 11592 26792
rect 11528 26568 11592 26632
rect 11528 26408 11592 26472
rect 11528 26248 11592 26312
rect 11528 26148 11592 26152
rect 11528 26092 11532 26148
rect 11532 26092 11588 26148
rect 11588 26092 11592 26148
rect 11528 26088 11592 26092
rect 11528 25988 11592 25992
rect 11528 25932 11532 25988
rect 11532 25932 11588 25988
rect 11588 25932 11592 25988
rect 11528 25928 11592 25932
rect 11528 25828 11592 25832
rect 11528 25772 11532 25828
rect 11532 25772 11588 25828
rect 11588 25772 11592 25828
rect 11528 25768 11592 25772
rect 11528 25668 11592 25672
rect 11528 25612 11532 25668
rect 11532 25612 11588 25668
rect 11588 25612 11592 25668
rect 11528 25608 11592 25612
rect 11528 25508 11592 25512
rect 11528 25452 11532 25508
rect 11532 25452 11588 25508
rect 11588 25452 11592 25508
rect 11528 25448 11592 25452
rect 11528 25348 11592 25352
rect 11528 25292 11532 25348
rect 11532 25292 11588 25348
rect 11588 25292 11592 25348
rect 11528 25288 11592 25292
rect 11528 25188 11592 25192
rect 11528 25132 11532 25188
rect 11532 25132 11588 25188
rect 11588 25132 11592 25188
rect 11528 25128 11592 25132
rect 11528 25028 11592 25032
rect 11528 24972 11532 25028
rect 11532 24972 11588 25028
rect 11588 24972 11592 25028
rect 11528 24968 11592 24972
rect 11528 24808 11592 24872
rect 11528 24708 11592 24712
rect 11528 24652 11532 24708
rect 11532 24652 11588 24708
rect 11588 24652 11592 24708
rect 11528 24648 11592 24652
rect 11528 24548 11592 24552
rect 11528 24492 11532 24548
rect 11532 24492 11588 24548
rect 11588 24492 11592 24548
rect 11528 24488 11592 24492
rect 11528 24388 11592 24392
rect 11528 24332 11532 24388
rect 11532 24332 11588 24388
rect 11588 24332 11592 24388
rect 11528 24328 11592 24332
rect 11528 24228 11592 24232
rect 11528 24172 11532 24228
rect 11532 24172 11588 24228
rect 11588 24172 11592 24228
rect 11528 24168 11592 24172
rect 11528 24068 11592 24072
rect 11528 24012 11532 24068
rect 11532 24012 11588 24068
rect 11588 24012 11592 24068
rect 11528 24008 11592 24012
rect 11528 23908 11592 23912
rect 11528 23852 11532 23908
rect 11532 23852 11588 23908
rect 11588 23852 11592 23908
rect 11528 23848 11592 23852
rect 11528 23748 11592 23752
rect 11528 23692 11532 23748
rect 11532 23692 11588 23748
rect 11588 23692 11592 23748
rect 11528 23688 11592 23692
rect 11528 23588 11592 23592
rect 11528 23532 11532 23588
rect 11532 23532 11588 23588
rect 11588 23532 11592 23588
rect 11528 23528 11592 23532
rect 11528 23428 11592 23432
rect 11528 23372 11532 23428
rect 11532 23372 11588 23428
rect 11588 23372 11592 23428
rect 11528 23368 11592 23372
rect 11528 23268 11592 23272
rect 11528 23212 11532 23268
rect 11532 23212 11588 23268
rect 11588 23212 11592 23268
rect 11528 23208 11592 23212
rect 11528 23108 11592 23112
rect 11528 23052 11532 23108
rect 11532 23052 11588 23108
rect 11588 23052 11592 23108
rect 11528 23048 11592 23052
rect 11528 22948 11592 22952
rect 11528 22892 11532 22948
rect 11532 22892 11588 22948
rect 11588 22892 11592 22948
rect 11528 22888 11592 22892
rect 11528 22788 11592 22792
rect 11528 22732 11532 22788
rect 11532 22732 11588 22788
rect 11588 22732 11592 22788
rect 11528 22728 11592 22732
rect 11528 22628 11592 22632
rect 11528 22572 11532 22628
rect 11532 22572 11588 22628
rect 11588 22572 11592 22628
rect 11528 22568 11592 22572
rect 11528 22468 11592 22472
rect 11528 22412 11532 22468
rect 11532 22412 11588 22468
rect 11588 22412 11592 22468
rect 11528 22408 11592 22412
rect 11528 22308 11592 22312
rect 11528 22252 11532 22308
rect 11532 22252 11588 22308
rect 11588 22252 11592 22308
rect 11528 22248 11592 22252
rect 11528 22148 11592 22152
rect 11528 22092 11532 22148
rect 11532 22092 11588 22148
rect 11588 22092 11592 22148
rect 11528 22088 11592 22092
rect 11528 21928 11592 21992
rect 11528 21828 11592 21832
rect 11528 21772 11532 21828
rect 11532 21772 11588 21828
rect 11588 21772 11592 21828
rect 11528 21768 11592 21772
rect 11528 21668 11592 21672
rect 11528 21612 11532 21668
rect 11532 21612 11588 21668
rect 11588 21612 11592 21668
rect 11528 21608 11592 21612
rect 11528 21508 11592 21512
rect 11528 21452 11532 21508
rect 11532 21452 11588 21508
rect 11588 21452 11592 21508
rect 11528 21448 11592 21452
rect 11528 21348 11592 21352
rect 11528 21292 11532 21348
rect 11532 21292 11588 21348
rect 11588 21292 11592 21348
rect 11528 21288 11592 21292
rect 11528 21188 11592 21192
rect 11528 21132 11532 21188
rect 11532 21132 11588 21188
rect 11588 21132 11592 21188
rect 11528 21128 11592 21132
rect 11528 21028 11592 21032
rect 11528 20972 11532 21028
rect 11532 20972 11588 21028
rect 11588 20972 11592 21028
rect 11528 20968 11592 20972
rect 11528 20868 11592 20872
rect 11528 20812 11532 20868
rect 11532 20812 11588 20868
rect 11588 20812 11592 20868
rect 11528 20808 11592 20812
rect 11528 20708 11592 20712
rect 11528 20652 11532 20708
rect 11532 20652 11588 20708
rect 11588 20652 11592 20708
rect 11528 20648 11592 20652
rect 11528 20488 11592 20552
rect 11528 20328 11592 20392
rect 11528 20168 11592 20232
rect 11528 20008 11592 20072
rect 11528 19908 11592 19912
rect 11528 19852 11532 19908
rect 11532 19852 11588 19908
rect 11588 19852 11592 19908
rect 11528 19848 11592 19852
rect 11528 19748 11592 19752
rect 11528 19692 11532 19748
rect 11532 19692 11588 19748
rect 11588 19692 11592 19748
rect 11528 19688 11592 19692
rect 11528 19588 11592 19592
rect 11528 19532 11532 19588
rect 11532 19532 11588 19588
rect 11588 19532 11592 19588
rect 11528 19528 11592 19532
rect 11528 19428 11592 19432
rect 11528 19372 11532 19428
rect 11532 19372 11588 19428
rect 11588 19372 11592 19428
rect 11528 19368 11592 19372
rect 11528 19268 11592 19272
rect 11528 19212 11532 19268
rect 11532 19212 11588 19268
rect 11588 19212 11592 19268
rect 11528 19208 11592 19212
rect 11528 19108 11592 19112
rect 11528 19052 11532 19108
rect 11532 19052 11588 19108
rect 11588 19052 11592 19108
rect 11528 19048 11592 19052
rect 11528 18948 11592 18952
rect 11528 18892 11532 18948
rect 11532 18892 11588 18948
rect 11588 18892 11592 18948
rect 11528 18888 11592 18892
rect 11528 18788 11592 18792
rect 11528 18732 11532 18788
rect 11532 18732 11588 18788
rect 11588 18732 11592 18788
rect 11528 18728 11592 18732
rect 11528 18568 11592 18632
rect 11528 18408 11592 18472
rect 11528 18248 11592 18312
rect 11528 18088 11592 18152
rect 11528 17988 11592 17992
rect 11528 17932 11532 17988
rect 11532 17932 11588 17988
rect 11588 17932 11592 17988
rect 11528 17928 11592 17932
rect 11528 17828 11592 17832
rect 11528 17772 11532 17828
rect 11532 17772 11588 17828
rect 11588 17772 11592 17828
rect 11528 17768 11592 17772
rect 11528 17668 11592 17672
rect 11528 17612 11532 17668
rect 11532 17612 11588 17668
rect 11588 17612 11592 17668
rect 11528 17608 11592 17612
rect 11528 17508 11592 17512
rect 11528 17452 11532 17508
rect 11532 17452 11588 17508
rect 11588 17452 11592 17508
rect 11528 17448 11592 17452
rect 11528 17348 11592 17352
rect 11528 17292 11532 17348
rect 11532 17292 11588 17348
rect 11588 17292 11592 17348
rect 11528 17288 11592 17292
rect 11528 17188 11592 17192
rect 11528 17132 11532 17188
rect 11532 17132 11588 17188
rect 11588 17132 11592 17188
rect 11528 17128 11592 17132
rect 11528 17028 11592 17032
rect 11528 16972 11532 17028
rect 11532 16972 11588 17028
rect 11588 16972 11592 17028
rect 11528 16968 11592 16972
rect 11528 16868 11592 16872
rect 11528 16812 11532 16868
rect 11532 16812 11588 16868
rect 11588 16812 11592 16868
rect 11528 16808 11592 16812
rect 11528 16648 11592 16712
rect 11528 16548 11592 16552
rect 11528 16492 11532 16548
rect 11532 16492 11588 16548
rect 11588 16492 11592 16548
rect 11528 16488 11592 16492
rect 11528 16388 11592 16392
rect 11528 16332 11532 16388
rect 11532 16332 11588 16388
rect 11588 16332 11592 16388
rect 11528 16328 11592 16332
rect 11528 16228 11592 16232
rect 11528 16172 11532 16228
rect 11532 16172 11588 16228
rect 11588 16172 11592 16228
rect 11528 16168 11592 16172
rect 11528 16068 11592 16072
rect 11528 16012 11532 16068
rect 11532 16012 11588 16068
rect 11588 16012 11592 16068
rect 11528 16008 11592 16012
rect 11528 15908 11592 15912
rect 11528 15852 11532 15908
rect 11532 15852 11588 15908
rect 11588 15852 11592 15908
rect 11528 15848 11592 15852
rect 11528 15748 11592 15752
rect 11528 15692 11532 15748
rect 11532 15692 11588 15748
rect 11588 15692 11592 15748
rect 11528 15688 11592 15692
rect 11528 15588 11592 15592
rect 11528 15532 11532 15588
rect 11532 15532 11588 15588
rect 11588 15532 11592 15588
rect 11528 15528 11592 15532
rect 11528 15428 11592 15432
rect 11528 15372 11532 15428
rect 11532 15372 11588 15428
rect 11588 15372 11592 15428
rect 11528 15368 11592 15372
rect 11528 15268 11592 15272
rect 11528 15212 11532 15268
rect 11532 15212 11588 15268
rect 11588 15212 11592 15268
rect 11528 15208 11592 15212
rect 11528 15108 11592 15112
rect 11528 15052 11532 15108
rect 11532 15052 11588 15108
rect 11588 15052 11592 15108
rect 11528 15048 11592 15052
rect 11528 14948 11592 14952
rect 11528 14892 11532 14948
rect 11532 14892 11588 14948
rect 11588 14892 11592 14948
rect 11528 14888 11592 14892
rect 11528 14788 11592 14792
rect 11528 14732 11532 14788
rect 11532 14732 11588 14788
rect 11588 14732 11592 14788
rect 11528 14728 11592 14732
rect 11528 14628 11592 14632
rect 11528 14572 11532 14628
rect 11532 14572 11588 14628
rect 11588 14572 11592 14628
rect 11528 14568 11592 14572
rect 11528 14468 11592 14472
rect 11528 14412 11532 14468
rect 11532 14412 11588 14468
rect 11588 14412 11592 14468
rect 11528 14408 11592 14412
rect 11528 14308 11592 14312
rect 11528 14252 11532 14308
rect 11532 14252 11588 14308
rect 11588 14252 11592 14308
rect 11528 14248 11592 14252
rect 11528 14148 11592 14152
rect 11528 14092 11532 14148
rect 11532 14092 11588 14148
rect 11588 14092 11592 14148
rect 11528 14088 11592 14092
rect 11528 13988 11592 13992
rect 11528 13932 11532 13988
rect 11532 13932 11588 13988
rect 11588 13932 11592 13988
rect 11528 13928 11592 13932
rect 11528 13768 11592 13832
rect 11528 13668 11592 13672
rect 11528 13612 11532 13668
rect 11532 13612 11588 13668
rect 11588 13612 11592 13668
rect 11528 13608 11592 13612
rect 11528 13508 11592 13512
rect 11528 13452 11532 13508
rect 11532 13452 11588 13508
rect 11588 13452 11592 13508
rect 11528 13448 11592 13452
rect 11528 13348 11592 13352
rect 11528 13292 11532 13348
rect 11532 13292 11588 13348
rect 11588 13292 11592 13348
rect 11528 13288 11592 13292
rect 11528 13188 11592 13192
rect 11528 13132 11532 13188
rect 11532 13132 11588 13188
rect 11588 13132 11592 13188
rect 11528 13128 11592 13132
rect 11528 13028 11592 13032
rect 11528 12972 11532 13028
rect 11532 12972 11588 13028
rect 11588 12972 11592 13028
rect 11528 12968 11592 12972
rect 11528 12868 11592 12872
rect 11528 12812 11532 12868
rect 11532 12812 11588 12868
rect 11588 12812 11592 12868
rect 11528 12808 11592 12812
rect 11528 12708 11592 12712
rect 11528 12652 11532 12708
rect 11532 12652 11588 12708
rect 11588 12652 11592 12708
rect 11528 12648 11592 12652
rect 11528 12548 11592 12552
rect 11528 12492 11532 12548
rect 11532 12492 11588 12548
rect 11588 12492 11592 12548
rect 11528 12488 11592 12492
rect 11528 12328 11592 12392
rect 11528 12168 11592 12232
rect 11528 12008 11592 12072
rect 11528 11848 11592 11912
rect 11528 11748 11592 11752
rect 11528 11692 11532 11748
rect 11532 11692 11588 11748
rect 11588 11692 11592 11748
rect 11528 11688 11592 11692
rect 11528 11588 11592 11592
rect 11528 11532 11532 11588
rect 11532 11532 11588 11588
rect 11588 11532 11592 11588
rect 11528 11528 11592 11532
rect 11528 11428 11592 11432
rect 11528 11372 11532 11428
rect 11532 11372 11588 11428
rect 11588 11372 11592 11428
rect 11528 11368 11592 11372
rect 11528 11268 11592 11272
rect 11528 11212 11532 11268
rect 11532 11212 11588 11268
rect 11588 11212 11592 11268
rect 11528 11208 11592 11212
rect 11528 11108 11592 11112
rect 11528 11052 11532 11108
rect 11532 11052 11588 11108
rect 11588 11052 11592 11108
rect 11528 11048 11592 11052
rect 11528 10948 11592 10952
rect 11528 10892 11532 10948
rect 11532 10892 11588 10948
rect 11588 10892 11592 10948
rect 11528 10888 11592 10892
rect 11528 10788 11592 10792
rect 11528 10732 11532 10788
rect 11532 10732 11588 10788
rect 11588 10732 11592 10788
rect 11528 10728 11592 10732
rect 11528 10628 11592 10632
rect 11528 10572 11532 10628
rect 11532 10572 11588 10628
rect 11588 10572 11592 10628
rect 11528 10568 11592 10572
rect 11528 10468 11592 10472
rect 11528 10412 11532 10468
rect 11532 10412 11588 10468
rect 11588 10412 11592 10468
rect 11528 10408 11592 10412
rect 11528 10308 11592 10312
rect 11528 10252 11532 10308
rect 11532 10252 11588 10308
rect 11588 10252 11592 10308
rect 11528 10248 11592 10252
rect 11528 10148 11592 10152
rect 11528 10092 11532 10148
rect 11532 10092 11588 10148
rect 11588 10092 11592 10148
rect 11528 10088 11592 10092
rect 11528 9988 11592 9992
rect 11528 9932 11532 9988
rect 11532 9932 11588 9988
rect 11588 9932 11592 9988
rect 11528 9928 11592 9932
rect 11528 9828 11592 9832
rect 11528 9772 11532 9828
rect 11532 9772 11588 9828
rect 11588 9772 11592 9828
rect 11528 9768 11592 9772
rect 11528 9608 11592 9672
rect 11528 9508 11592 9512
rect 11528 9452 11532 9508
rect 11532 9452 11588 9508
rect 11588 9452 11592 9508
rect 11528 9448 11592 9452
rect 11528 9348 11592 9352
rect 11528 9292 11532 9348
rect 11532 9292 11588 9348
rect 11588 9292 11592 9348
rect 11528 9288 11592 9292
rect 11528 9128 11592 9192
rect 11528 9028 11592 9032
rect 11528 8972 11532 9028
rect 11532 8972 11588 9028
rect 11588 8972 11592 9028
rect 11528 8968 11592 8972
rect 11528 8868 11592 8872
rect 11528 8812 11532 8868
rect 11532 8812 11588 8868
rect 11588 8812 11592 8868
rect 11528 8808 11592 8812
rect 11528 8708 11592 8712
rect 11528 8652 11532 8708
rect 11532 8652 11588 8708
rect 11588 8652 11592 8708
rect 11528 8648 11592 8652
rect 11528 8548 11592 8552
rect 11528 8492 11532 8548
rect 11532 8492 11588 8548
rect 11588 8492 11592 8548
rect 11528 8488 11592 8492
rect 11528 8388 11592 8392
rect 11528 8332 11532 8388
rect 11532 8332 11588 8388
rect 11588 8332 11592 8388
rect 11528 8328 11592 8332
rect 11528 8228 11592 8232
rect 11528 8172 11532 8228
rect 11532 8172 11588 8228
rect 11588 8172 11592 8228
rect 11528 8168 11592 8172
rect 11528 8068 11592 8072
rect 11528 8012 11532 8068
rect 11532 8012 11588 8068
rect 11588 8012 11592 8068
rect 11528 8008 11592 8012
rect 11528 7908 11592 7912
rect 11528 7852 11532 7908
rect 11532 7852 11588 7908
rect 11588 7852 11592 7908
rect 11528 7848 11592 7852
rect 11528 7748 11592 7752
rect 11528 7692 11532 7748
rect 11532 7692 11588 7748
rect 11588 7692 11592 7748
rect 11528 7688 11592 7692
rect 11528 7528 11592 7592
rect 11528 7428 11592 7432
rect 11528 7372 11532 7428
rect 11532 7372 11588 7428
rect 11588 7372 11592 7428
rect 11528 7368 11592 7372
rect 11528 7268 11592 7272
rect 11528 7212 11532 7268
rect 11532 7212 11588 7268
rect 11588 7212 11592 7268
rect 11528 7208 11592 7212
rect 11528 7048 11592 7112
rect 11528 6948 11592 6952
rect 11528 6892 11532 6948
rect 11532 6892 11588 6948
rect 11588 6892 11592 6948
rect 11528 6888 11592 6892
rect 11528 6788 11592 6792
rect 11528 6732 11532 6788
rect 11532 6732 11588 6788
rect 11588 6732 11592 6788
rect 11528 6728 11592 6732
rect 11528 6568 11592 6632
rect 11528 6468 11592 6472
rect 11528 6412 11532 6468
rect 11532 6412 11588 6468
rect 11588 6412 11592 6468
rect 11528 6408 11592 6412
rect 11528 6308 11592 6312
rect 11528 6252 11532 6308
rect 11532 6252 11588 6308
rect 11588 6252 11592 6308
rect 11528 6248 11592 6252
rect 11528 6148 11592 6152
rect 11528 6092 11532 6148
rect 11532 6092 11588 6148
rect 11588 6092 11592 6148
rect 11528 6088 11592 6092
rect 11528 5988 11592 5992
rect 11528 5932 11532 5988
rect 11532 5932 11588 5988
rect 11588 5932 11592 5988
rect 11528 5928 11592 5932
rect 11528 5828 11592 5832
rect 11528 5772 11532 5828
rect 11532 5772 11588 5828
rect 11588 5772 11592 5828
rect 11528 5768 11592 5772
rect 11528 5668 11592 5672
rect 11528 5612 11532 5668
rect 11532 5612 11588 5668
rect 11588 5612 11592 5668
rect 11528 5608 11592 5612
rect 11528 5508 11592 5512
rect 11528 5452 11532 5508
rect 11532 5452 11588 5508
rect 11588 5452 11592 5508
rect 11528 5448 11592 5452
rect 11528 5348 11592 5352
rect 11528 5292 11532 5348
rect 11532 5292 11588 5348
rect 11588 5292 11592 5348
rect 11528 5288 11592 5292
rect 11528 5188 11592 5192
rect 11528 5132 11532 5188
rect 11532 5132 11588 5188
rect 11588 5132 11592 5188
rect 11528 5128 11592 5132
rect 11528 5028 11592 5032
rect 11528 4972 11532 5028
rect 11532 4972 11588 5028
rect 11588 4972 11592 5028
rect 11528 4968 11592 4972
rect 11528 4868 11592 4872
rect 11528 4812 11532 4868
rect 11532 4812 11588 4868
rect 11588 4812 11592 4868
rect 11528 4808 11592 4812
rect 11528 4708 11592 4712
rect 11528 4652 11532 4708
rect 11532 4652 11588 4708
rect 11588 4652 11592 4708
rect 11528 4648 11592 4652
rect 11528 4548 11592 4552
rect 11528 4492 11532 4548
rect 11532 4492 11588 4548
rect 11588 4492 11592 4548
rect 11528 4488 11592 4492
rect 11528 4388 11592 4392
rect 11528 4332 11532 4388
rect 11532 4332 11588 4388
rect 11588 4332 11592 4388
rect 11528 4328 11592 4332
rect 11528 4228 11592 4232
rect 11528 4172 11532 4228
rect 11532 4172 11588 4228
rect 11588 4172 11592 4228
rect 11528 4168 11592 4172
rect 11528 4068 11592 4072
rect 11528 4012 11532 4068
rect 11532 4012 11588 4068
rect 11588 4012 11592 4068
rect 11528 4008 11592 4012
rect 11528 3908 11592 3912
rect 11528 3852 11532 3908
rect 11532 3852 11588 3908
rect 11588 3852 11592 3908
rect 11528 3848 11592 3852
rect 11528 3688 11592 3752
rect 11528 3528 11592 3592
rect 11528 3428 11592 3432
rect 11528 3372 11532 3428
rect 11532 3372 11588 3428
rect 11588 3372 11592 3428
rect 11528 3368 11592 3372
rect 11528 3268 11592 3272
rect 11528 3212 11532 3268
rect 11532 3212 11588 3268
rect 11588 3212 11592 3268
rect 11528 3208 11592 3212
rect 11528 3108 11592 3112
rect 11528 3052 11532 3108
rect 11532 3052 11588 3108
rect 11588 3052 11592 3108
rect 11528 3048 11592 3052
rect 11528 2948 11592 2952
rect 11528 2892 11532 2948
rect 11532 2892 11588 2948
rect 11588 2892 11592 2948
rect 11528 2888 11592 2892
rect 11528 2788 11592 2792
rect 11528 2732 11532 2788
rect 11532 2732 11588 2788
rect 11588 2732 11592 2788
rect 11528 2728 11592 2732
rect 11528 2628 11592 2632
rect 11528 2572 11532 2628
rect 11532 2572 11588 2628
rect 11588 2572 11592 2628
rect 11528 2568 11592 2572
rect 11528 2468 11592 2472
rect 11528 2412 11532 2468
rect 11532 2412 11588 2468
rect 11588 2412 11592 2468
rect 11528 2408 11592 2412
rect 11528 2308 11592 2312
rect 11528 2252 11532 2308
rect 11532 2252 11588 2308
rect 11588 2252 11592 2308
rect 11528 2248 11592 2252
rect 11528 2148 11592 2152
rect 11528 2092 11532 2148
rect 11532 2092 11588 2148
rect 11588 2092 11592 2148
rect 11528 2088 11592 2092
rect 11528 1988 11592 1992
rect 11528 1932 11532 1988
rect 11532 1932 11588 1988
rect 11588 1932 11592 1988
rect 11528 1928 11592 1932
rect 11528 1768 11592 1832
rect 11528 1668 11592 1672
rect 11528 1612 11532 1668
rect 11532 1612 11588 1668
rect 11588 1612 11592 1668
rect 11528 1608 11592 1612
rect 11528 1508 11592 1512
rect 11528 1452 11532 1508
rect 11532 1452 11588 1508
rect 11588 1452 11592 1508
rect 11528 1448 11592 1452
rect 11528 1348 11592 1352
rect 11528 1292 11532 1348
rect 11532 1292 11588 1348
rect 11588 1292 11592 1348
rect 11528 1288 11592 1292
rect 11528 1188 11592 1192
rect 11528 1132 11532 1188
rect 11532 1132 11588 1188
rect 11588 1132 11592 1188
rect 11528 1128 11592 1132
rect 11528 1028 11592 1032
rect 11528 972 11532 1028
rect 11532 972 11588 1028
rect 11588 972 11592 1028
rect 11528 968 11592 972
rect 11528 808 11592 872
rect 11528 648 11592 712
rect 11528 548 11592 552
rect 11528 492 11532 548
rect 11532 492 11588 548
rect 11588 492 11592 548
rect 11528 488 11592 492
rect 11528 388 11592 392
rect 11528 332 11532 388
rect 11532 332 11588 388
rect 11588 332 11592 388
rect 11528 328 11592 332
rect 11528 228 11592 232
rect 11528 172 11532 228
rect 11532 172 11588 228
rect 11588 172 11592 228
rect 11528 168 11592 172
rect 11528 68 11592 72
rect 11528 12 11532 68
rect 11532 12 11588 68
rect 11588 12 11592 68
rect 11528 8 11592 12
rect 11848 31428 11912 31432
rect 11848 31372 11852 31428
rect 11852 31372 11908 31428
rect 11908 31372 11912 31428
rect 11848 31368 11912 31372
rect 11848 31268 11912 31272
rect 11848 31212 11852 31268
rect 11852 31212 11908 31268
rect 11908 31212 11912 31268
rect 11848 31208 11912 31212
rect 11848 31108 11912 31112
rect 11848 31052 11852 31108
rect 11852 31052 11908 31108
rect 11908 31052 11912 31108
rect 11848 31048 11912 31052
rect 11848 30948 11912 30952
rect 11848 30892 11852 30948
rect 11852 30892 11908 30948
rect 11908 30892 11912 30948
rect 11848 30888 11912 30892
rect 11848 30788 11912 30792
rect 11848 30732 11852 30788
rect 11852 30732 11908 30788
rect 11908 30732 11912 30788
rect 11848 30728 11912 30732
rect 11848 30628 11912 30632
rect 11848 30572 11852 30628
rect 11852 30572 11908 30628
rect 11908 30572 11912 30628
rect 11848 30568 11912 30572
rect 11848 30468 11912 30472
rect 11848 30412 11852 30468
rect 11852 30412 11908 30468
rect 11908 30412 11912 30468
rect 11848 30408 11912 30412
rect 11848 30308 11912 30312
rect 11848 30252 11852 30308
rect 11852 30252 11908 30308
rect 11908 30252 11912 30308
rect 11848 30248 11912 30252
rect 11848 30088 11912 30152
rect 11848 29988 11912 29992
rect 11848 29932 11852 29988
rect 11852 29932 11908 29988
rect 11908 29932 11912 29988
rect 11848 29928 11912 29932
rect 11848 29828 11912 29832
rect 11848 29772 11852 29828
rect 11852 29772 11908 29828
rect 11908 29772 11912 29828
rect 11848 29768 11912 29772
rect 11848 29668 11912 29672
rect 11848 29612 11852 29668
rect 11852 29612 11908 29668
rect 11908 29612 11912 29668
rect 11848 29608 11912 29612
rect 11848 29508 11912 29512
rect 11848 29452 11852 29508
rect 11852 29452 11908 29508
rect 11908 29452 11912 29508
rect 11848 29448 11912 29452
rect 11848 29348 11912 29352
rect 11848 29292 11852 29348
rect 11852 29292 11908 29348
rect 11908 29292 11912 29348
rect 11848 29288 11912 29292
rect 11848 29188 11912 29192
rect 11848 29132 11852 29188
rect 11852 29132 11908 29188
rect 11908 29132 11912 29188
rect 11848 29128 11912 29132
rect 11848 29028 11912 29032
rect 11848 28972 11852 29028
rect 11852 28972 11908 29028
rect 11908 28972 11912 29028
rect 11848 28968 11912 28972
rect 11848 28868 11912 28872
rect 11848 28812 11852 28868
rect 11852 28812 11908 28868
rect 11908 28812 11912 28868
rect 11848 28808 11912 28812
rect 11848 28648 11912 28712
rect 11848 28488 11912 28552
rect 11848 28328 11912 28392
rect 11848 28168 11912 28232
rect 11848 28068 11912 28072
rect 11848 28012 11852 28068
rect 11852 28012 11908 28068
rect 11908 28012 11912 28068
rect 11848 28008 11912 28012
rect 11848 27908 11912 27912
rect 11848 27852 11852 27908
rect 11852 27852 11908 27908
rect 11908 27852 11912 27908
rect 11848 27848 11912 27852
rect 11848 27748 11912 27752
rect 11848 27692 11852 27748
rect 11852 27692 11908 27748
rect 11908 27692 11912 27748
rect 11848 27688 11912 27692
rect 11848 27588 11912 27592
rect 11848 27532 11852 27588
rect 11852 27532 11908 27588
rect 11908 27532 11912 27588
rect 11848 27528 11912 27532
rect 11848 27428 11912 27432
rect 11848 27372 11852 27428
rect 11852 27372 11908 27428
rect 11908 27372 11912 27428
rect 11848 27368 11912 27372
rect 11848 27268 11912 27272
rect 11848 27212 11852 27268
rect 11852 27212 11908 27268
rect 11908 27212 11912 27268
rect 11848 27208 11912 27212
rect 11848 27108 11912 27112
rect 11848 27052 11852 27108
rect 11852 27052 11908 27108
rect 11908 27052 11912 27108
rect 11848 27048 11912 27052
rect 11848 26948 11912 26952
rect 11848 26892 11852 26948
rect 11852 26892 11908 26948
rect 11908 26892 11912 26948
rect 11848 26888 11912 26892
rect 11848 26728 11912 26792
rect 11848 26568 11912 26632
rect 11848 26408 11912 26472
rect 11848 26248 11912 26312
rect 11848 26148 11912 26152
rect 11848 26092 11852 26148
rect 11852 26092 11908 26148
rect 11908 26092 11912 26148
rect 11848 26088 11912 26092
rect 11848 25988 11912 25992
rect 11848 25932 11852 25988
rect 11852 25932 11908 25988
rect 11908 25932 11912 25988
rect 11848 25928 11912 25932
rect 11848 25828 11912 25832
rect 11848 25772 11852 25828
rect 11852 25772 11908 25828
rect 11908 25772 11912 25828
rect 11848 25768 11912 25772
rect 11848 25668 11912 25672
rect 11848 25612 11852 25668
rect 11852 25612 11908 25668
rect 11908 25612 11912 25668
rect 11848 25608 11912 25612
rect 11848 25508 11912 25512
rect 11848 25452 11852 25508
rect 11852 25452 11908 25508
rect 11908 25452 11912 25508
rect 11848 25448 11912 25452
rect 11848 25348 11912 25352
rect 11848 25292 11852 25348
rect 11852 25292 11908 25348
rect 11908 25292 11912 25348
rect 11848 25288 11912 25292
rect 11848 25188 11912 25192
rect 11848 25132 11852 25188
rect 11852 25132 11908 25188
rect 11908 25132 11912 25188
rect 11848 25128 11912 25132
rect 11848 25028 11912 25032
rect 11848 24972 11852 25028
rect 11852 24972 11908 25028
rect 11908 24972 11912 25028
rect 11848 24968 11912 24972
rect 11848 24808 11912 24872
rect 11848 24708 11912 24712
rect 11848 24652 11852 24708
rect 11852 24652 11908 24708
rect 11908 24652 11912 24708
rect 11848 24648 11912 24652
rect 11848 24548 11912 24552
rect 11848 24492 11852 24548
rect 11852 24492 11908 24548
rect 11908 24492 11912 24548
rect 11848 24488 11912 24492
rect 11848 24388 11912 24392
rect 11848 24332 11852 24388
rect 11852 24332 11908 24388
rect 11908 24332 11912 24388
rect 11848 24328 11912 24332
rect 11848 24228 11912 24232
rect 11848 24172 11852 24228
rect 11852 24172 11908 24228
rect 11908 24172 11912 24228
rect 11848 24168 11912 24172
rect 11848 24068 11912 24072
rect 11848 24012 11852 24068
rect 11852 24012 11908 24068
rect 11908 24012 11912 24068
rect 11848 24008 11912 24012
rect 11848 23908 11912 23912
rect 11848 23852 11852 23908
rect 11852 23852 11908 23908
rect 11908 23852 11912 23908
rect 11848 23848 11912 23852
rect 11848 23748 11912 23752
rect 11848 23692 11852 23748
rect 11852 23692 11908 23748
rect 11908 23692 11912 23748
rect 11848 23688 11912 23692
rect 11848 23588 11912 23592
rect 11848 23532 11852 23588
rect 11852 23532 11908 23588
rect 11908 23532 11912 23588
rect 11848 23528 11912 23532
rect 11848 23428 11912 23432
rect 11848 23372 11852 23428
rect 11852 23372 11908 23428
rect 11908 23372 11912 23428
rect 11848 23368 11912 23372
rect 11848 23268 11912 23272
rect 11848 23212 11852 23268
rect 11852 23212 11908 23268
rect 11908 23212 11912 23268
rect 11848 23208 11912 23212
rect 11848 23108 11912 23112
rect 11848 23052 11852 23108
rect 11852 23052 11908 23108
rect 11908 23052 11912 23108
rect 11848 23048 11912 23052
rect 11848 22948 11912 22952
rect 11848 22892 11852 22948
rect 11852 22892 11908 22948
rect 11908 22892 11912 22948
rect 11848 22888 11912 22892
rect 11848 22788 11912 22792
rect 11848 22732 11852 22788
rect 11852 22732 11908 22788
rect 11908 22732 11912 22788
rect 11848 22728 11912 22732
rect 11848 22628 11912 22632
rect 11848 22572 11852 22628
rect 11852 22572 11908 22628
rect 11908 22572 11912 22628
rect 11848 22568 11912 22572
rect 11848 22468 11912 22472
rect 11848 22412 11852 22468
rect 11852 22412 11908 22468
rect 11908 22412 11912 22468
rect 11848 22408 11912 22412
rect 11848 22308 11912 22312
rect 11848 22252 11852 22308
rect 11852 22252 11908 22308
rect 11908 22252 11912 22308
rect 11848 22248 11912 22252
rect 11848 22148 11912 22152
rect 11848 22092 11852 22148
rect 11852 22092 11908 22148
rect 11908 22092 11912 22148
rect 11848 22088 11912 22092
rect 11848 21928 11912 21992
rect 11848 21828 11912 21832
rect 11848 21772 11852 21828
rect 11852 21772 11908 21828
rect 11908 21772 11912 21828
rect 11848 21768 11912 21772
rect 11848 21668 11912 21672
rect 11848 21612 11852 21668
rect 11852 21612 11908 21668
rect 11908 21612 11912 21668
rect 11848 21608 11912 21612
rect 11848 21508 11912 21512
rect 11848 21452 11852 21508
rect 11852 21452 11908 21508
rect 11908 21452 11912 21508
rect 11848 21448 11912 21452
rect 11848 21348 11912 21352
rect 11848 21292 11852 21348
rect 11852 21292 11908 21348
rect 11908 21292 11912 21348
rect 11848 21288 11912 21292
rect 11848 21188 11912 21192
rect 11848 21132 11852 21188
rect 11852 21132 11908 21188
rect 11908 21132 11912 21188
rect 11848 21128 11912 21132
rect 11848 21028 11912 21032
rect 11848 20972 11852 21028
rect 11852 20972 11908 21028
rect 11908 20972 11912 21028
rect 11848 20968 11912 20972
rect 11848 20868 11912 20872
rect 11848 20812 11852 20868
rect 11852 20812 11908 20868
rect 11908 20812 11912 20868
rect 11848 20808 11912 20812
rect 11848 20708 11912 20712
rect 11848 20652 11852 20708
rect 11852 20652 11908 20708
rect 11908 20652 11912 20708
rect 11848 20648 11912 20652
rect 11848 20488 11912 20552
rect 11848 20328 11912 20392
rect 11848 20168 11912 20232
rect 11848 20008 11912 20072
rect 11848 19908 11912 19912
rect 11848 19852 11852 19908
rect 11852 19852 11908 19908
rect 11908 19852 11912 19908
rect 11848 19848 11912 19852
rect 11848 19748 11912 19752
rect 11848 19692 11852 19748
rect 11852 19692 11908 19748
rect 11908 19692 11912 19748
rect 11848 19688 11912 19692
rect 11848 19588 11912 19592
rect 11848 19532 11852 19588
rect 11852 19532 11908 19588
rect 11908 19532 11912 19588
rect 11848 19528 11912 19532
rect 11848 19428 11912 19432
rect 11848 19372 11852 19428
rect 11852 19372 11908 19428
rect 11908 19372 11912 19428
rect 11848 19368 11912 19372
rect 11848 19268 11912 19272
rect 11848 19212 11852 19268
rect 11852 19212 11908 19268
rect 11908 19212 11912 19268
rect 11848 19208 11912 19212
rect 11848 19108 11912 19112
rect 11848 19052 11852 19108
rect 11852 19052 11908 19108
rect 11908 19052 11912 19108
rect 11848 19048 11912 19052
rect 11848 18948 11912 18952
rect 11848 18892 11852 18948
rect 11852 18892 11908 18948
rect 11908 18892 11912 18948
rect 11848 18888 11912 18892
rect 11848 18788 11912 18792
rect 11848 18732 11852 18788
rect 11852 18732 11908 18788
rect 11908 18732 11912 18788
rect 11848 18728 11912 18732
rect 11848 18568 11912 18632
rect 11848 18408 11912 18472
rect 11848 18248 11912 18312
rect 11848 18088 11912 18152
rect 11848 17988 11912 17992
rect 11848 17932 11852 17988
rect 11852 17932 11908 17988
rect 11908 17932 11912 17988
rect 11848 17928 11912 17932
rect 11848 17828 11912 17832
rect 11848 17772 11852 17828
rect 11852 17772 11908 17828
rect 11908 17772 11912 17828
rect 11848 17768 11912 17772
rect 11848 17668 11912 17672
rect 11848 17612 11852 17668
rect 11852 17612 11908 17668
rect 11908 17612 11912 17668
rect 11848 17608 11912 17612
rect 11848 17508 11912 17512
rect 11848 17452 11852 17508
rect 11852 17452 11908 17508
rect 11908 17452 11912 17508
rect 11848 17448 11912 17452
rect 11848 17348 11912 17352
rect 11848 17292 11852 17348
rect 11852 17292 11908 17348
rect 11908 17292 11912 17348
rect 11848 17288 11912 17292
rect 11848 17188 11912 17192
rect 11848 17132 11852 17188
rect 11852 17132 11908 17188
rect 11908 17132 11912 17188
rect 11848 17128 11912 17132
rect 11848 17028 11912 17032
rect 11848 16972 11852 17028
rect 11852 16972 11908 17028
rect 11908 16972 11912 17028
rect 11848 16968 11912 16972
rect 11848 16868 11912 16872
rect 11848 16812 11852 16868
rect 11852 16812 11908 16868
rect 11908 16812 11912 16868
rect 11848 16808 11912 16812
rect 11848 16648 11912 16712
rect 11848 16548 11912 16552
rect 11848 16492 11852 16548
rect 11852 16492 11908 16548
rect 11908 16492 11912 16548
rect 11848 16488 11912 16492
rect 11848 16388 11912 16392
rect 11848 16332 11852 16388
rect 11852 16332 11908 16388
rect 11908 16332 11912 16388
rect 11848 16328 11912 16332
rect 11848 16228 11912 16232
rect 11848 16172 11852 16228
rect 11852 16172 11908 16228
rect 11908 16172 11912 16228
rect 11848 16168 11912 16172
rect 11848 16068 11912 16072
rect 11848 16012 11852 16068
rect 11852 16012 11908 16068
rect 11908 16012 11912 16068
rect 11848 16008 11912 16012
rect 11848 15908 11912 15912
rect 11848 15852 11852 15908
rect 11852 15852 11908 15908
rect 11908 15852 11912 15908
rect 11848 15848 11912 15852
rect 11848 15748 11912 15752
rect 11848 15692 11852 15748
rect 11852 15692 11908 15748
rect 11908 15692 11912 15748
rect 11848 15688 11912 15692
rect 11848 15588 11912 15592
rect 11848 15532 11852 15588
rect 11852 15532 11908 15588
rect 11908 15532 11912 15588
rect 11848 15528 11912 15532
rect 11848 15428 11912 15432
rect 11848 15372 11852 15428
rect 11852 15372 11908 15428
rect 11908 15372 11912 15428
rect 11848 15368 11912 15372
rect 11848 15268 11912 15272
rect 11848 15212 11852 15268
rect 11852 15212 11908 15268
rect 11908 15212 11912 15268
rect 11848 15208 11912 15212
rect 11848 15108 11912 15112
rect 11848 15052 11852 15108
rect 11852 15052 11908 15108
rect 11908 15052 11912 15108
rect 11848 15048 11912 15052
rect 11848 14948 11912 14952
rect 11848 14892 11852 14948
rect 11852 14892 11908 14948
rect 11908 14892 11912 14948
rect 11848 14888 11912 14892
rect 11848 14788 11912 14792
rect 11848 14732 11852 14788
rect 11852 14732 11908 14788
rect 11908 14732 11912 14788
rect 11848 14728 11912 14732
rect 11848 14628 11912 14632
rect 11848 14572 11852 14628
rect 11852 14572 11908 14628
rect 11908 14572 11912 14628
rect 11848 14568 11912 14572
rect 11848 14468 11912 14472
rect 11848 14412 11852 14468
rect 11852 14412 11908 14468
rect 11908 14412 11912 14468
rect 11848 14408 11912 14412
rect 11848 14308 11912 14312
rect 11848 14252 11852 14308
rect 11852 14252 11908 14308
rect 11908 14252 11912 14308
rect 11848 14248 11912 14252
rect 11848 14148 11912 14152
rect 11848 14092 11852 14148
rect 11852 14092 11908 14148
rect 11908 14092 11912 14148
rect 11848 14088 11912 14092
rect 11848 13988 11912 13992
rect 11848 13932 11852 13988
rect 11852 13932 11908 13988
rect 11908 13932 11912 13988
rect 11848 13928 11912 13932
rect 11848 13768 11912 13832
rect 11848 13668 11912 13672
rect 11848 13612 11852 13668
rect 11852 13612 11908 13668
rect 11908 13612 11912 13668
rect 11848 13608 11912 13612
rect 11848 13508 11912 13512
rect 11848 13452 11852 13508
rect 11852 13452 11908 13508
rect 11908 13452 11912 13508
rect 11848 13448 11912 13452
rect 11848 13348 11912 13352
rect 11848 13292 11852 13348
rect 11852 13292 11908 13348
rect 11908 13292 11912 13348
rect 11848 13288 11912 13292
rect 11848 13188 11912 13192
rect 11848 13132 11852 13188
rect 11852 13132 11908 13188
rect 11908 13132 11912 13188
rect 11848 13128 11912 13132
rect 11848 13028 11912 13032
rect 11848 12972 11852 13028
rect 11852 12972 11908 13028
rect 11908 12972 11912 13028
rect 11848 12968 11912 12972
rect 11848 12868 11912 12872
rect 11848 12812 11852 12868
rect 11852 12812 11908 12868
rect 11908 12812 11912 12868
rect 11848 12808 11912 12812
rect 11848 12708 11912 12712
rect 11848 12652 11852 12708
rect 11852 12652 11908 12708
rect 11908 12652 11912 12708
rect 11848 12648 11912 12652
rect 11848 12548 11912 12552
rect 11848 12492 11852 12548
rect 11852 12492 11908 12548
rect 11908 12492 11912 12548
rect 11848 12488 11912 12492
rect 11848 12328 11912 12392
rect 11848 12168 11912 12232
rect 11848 12008 11912 12072
rect 11848 11848 11912 11912
rect 11848 11748 11912 11752
rect 11848 11692 11852 11748
rect 11852 11692 11908 11748
rect 11908 11692 11912 11748
rect 11848 11688 11912 11692
rect 11848 11588 11912 11592
rect 11848 11532 11852 11588
rect 11852 11532 11908 11588
rect 11908 11532 11912 11588
rect 11848 11528 11912 11532
rect 11848 11428 11912 11432
rect 11848 11372 11852 11428
rect 11852 11372 11908 11428
rect 11908 11372 11912 11428
rect 11848 11368 11912 11372
rect 11848 11268 11912 11272
rect 11848 11212 11852 11268
rect 11852 11212 11908 11268
rect 11908 11212 11912 11268
rect 11848 11208 11912 11212
rect 11848 11108 11912 11112
rect 11848 11052 11852 11108
rect 11852 11052 11908 11108
rect 11908 11052 11912 11108
rect 11848 11048 11912 11052
rect 11848 10948 11912 10952
rect 11848 10892 11852 10948
rect 11852 10892 11908 10948
rect 11908 10892 11912 10948
rect 11848 10888 11912 10892
rect 11848 10788 11912 10792
rect 11848 10732 11852 10788
rect 11852 10732 11908 10788
rect 11908 10732 11912 10788
rect 11848 10728 11912 10732
rect 11848 10628 11912 10632
rect 11848 10572 11852 10628
rect 11852 10572 11908 10628
rect 11908 10572 11912 10628
rect 11848 10568 11912 10572
rect 11848 10468 11912 10472
rect 11848 10412 11852 10468
rect 11852 10412 11908 10468
rect 11908 10412 11912 10468
rect 11848 10408 11912 10412
rect 11848 10308 11912 10312
rect 11848 10252 11852 10308
rect 11852 10252 11908 10308
rect 11908 10252 11912 10308
rect 11848 10248 11912 10252
rect 11848 10148 11912 10152
rect 11848 10092 11852 10148
rect 11852 10092 11908 10148
rect 11908 10092 11912 10148
rect 11848 10088 11912 10092
rect 11848 9988 11912 9992
rect 11848 9932 11852 9988
rect 11852 9932 11908 9988
rect 11908 9932 11912 9988
rect 11848 9928 11912 9932
rect 11848 9828 11912 9832
rect 11848 9772 11852 9828
rect 11852 9772 11908 9828
rect 11908 9772 11912 9828
rect 11848 9768 11912 9772
rect 11848 9608 11912 9672
rect 11848 9508 11912 9512
rect 11848 9452 11852 9508
rect 11852 9452 11908 9508
rect 11908 9452 11912 9508
rect 11848 9448 11912 9452
rect 11848 9348 11912 9352
rect 11848 9292 11852 9348
rect 11852 9292 11908 9348
rect 11908 9292 11912 9348
rect 11848 9288 11912 9292
rect 11848 9128 11912 9192
rect 11848 9028 11912 9032
rect 11848 8972 11852 9028
rect 11852 8972 11908 9028
rect 11908 8972 11912 9028
rect 11848 8968 11912 8972
rect 11848 8868 11912 8872
rect 11848 8812 11852 8868
rect 11852 8812 11908 8868
rect 11908 8812 11912 8868
rect 11848 8808 11912 8812
rect 11848 8708 11912 8712
rect 11848 8652 11852 8708
rect 11852 8652 11908 8708
rect 11908 8652 11912 8708
rect 11848 8648 11912 8652
rect 11848 8548 11912 8552
rect 11848 8492 11852 8548
rect 11852 8492 11908 8548
rect 11908 8492 11912 8548
rect 11848 8488 11912 8492
rect 11848 8388 11912 8392
rect 11848 8332 11852 8388
rect 11852 8332 11908 8388
rect 11908 8332 11912 8388
rect 11848 8328 11912 8332
rect 11848 8228 11912 8232
rect 11848 8172 11852 8228
rect 11852 8172 11908 8228
rect 11908 8172 11912 8228
rect 11848 8168 11912 8172
rect 11848 8068 11912 8072
rect 11848 8012 11852 8068
rect 11852 8012 11908 8068
rect 11908 8012 11912 8068
rect 11848 8008 11912 8012
rect 11848 7908 11912 7912
rect 11848 7852 11852 7908
rect 11852 7852 11908 7908
rect 11908 7852 11912 7908
rect 11848 7848 11912 7852
rect 11848 7748 11912 7752
rect 11848 7692 11852 7748
rect 11852 7692 11908 7748
rect 11908 7692 11912 7748
rect 11848 7688 11912 7692
rect 11848 7528 11912 7592
rect 11848 7428 11912 7432
rect 11848 7372 11852 7428
rect 11852 7372 11908 7428
rect 11908 7372 11912 7428
rect 11848 7368 11912 7372
rect 11848 7268 11912 7272
rect 11848 7212 11852 7268
rect 11852 7212 11908 7268
rect 11908 7212 11912 7268
rect 11848 7208 11912 7212
rect 11848 7048 11912 7112
rect 11848 6948 11912 6952
rect 11848 6892 11852 6948
rect 11852 6892 11908 6948
rect 11908 6892 11912 6948
rect 11848 6888 11912 6892
rect 11848 6788 11912 6792
rect 11848 6732 11852 6788
rect 11852 6732 11908 6788
rect 11908 6732 11912 6788
rect 11848 6728 11912 6732
rect 11848 6568 11912 6632
rect 11848 6468 11912 6472
rect 11848 6412 11852 6468
rect 11852 6412 11908 6468
rect 11908 6412 11912 6468
rect 11848 6408 11912 6412
rect 11848 6308 11912 6312
rect 11848 6252 11852 6308
rect 11852 6252 11908 6308
rect 11908 6252 11912 6308
rect 11848 6248 11912 6252
rect 11848 6148 11912 6152
rect 11848 6092 11852 6148
rect 11852 6092 11908 6148
rect 11908 6092 11912 6148
rect 11848 6088 11912 6092
rect 11848 5988 11912 5992
rect 11848 5932 11852 5988
rect 11852 5932 11908 5988
rect 11908 5932 11912 5988
rect 11848 5928 11912 5932
rect 11848 5828 11912 5832
rect 11848 5772 11852 5828
rect 11852 5772 11908 5828
rect 11908 5772 11912 5828
rect 11848 5768 11912 5772
rect 11848 5668 11912 5672
rect 11848 5612 11852 5668
rect 11852 5612 11908 5668
rect 11908 5612 11912 5668
rect 11848 5608 11912 5612
rect 11848 5508 11912 5512
rect 11848 5452 11852 5508
rect 11852 5452 11908 5508
rect 11908 5452 11912 5508
rect 11848 5448 11912 5452
rect 11848 5348 11912 5352
rect 11848 5292 11852 5348
rect 11852 5292 11908 5348
rect 11908 5292 11912 5348
rect 11848 5288 11912 5292
rect 11848 5188 11912 5192
rect 11848 5132 11852 5188
rect 11852 5132 11908 5188
rect 11908 5132 11912 5188
rect 11848 5128 11912 5132
rect 11848 5028 11912 5032
rect 11848 4972 11852 5028
rect 11852 4972 11908 5028
rect 11908 4972 11912 5028
rect 11848 4968 11912 4972
rect 11848 4868 11912 4872
rect 11848 4812 11852 4868
rect 11852 4812 11908 4868
rect 11908 4812 11912 4868
rect 11848 4808 11912 4812
rect 11848 4708 11912 4712
rect 11848 4652 11852 4708
rect 11852 4652 11908 4708
rect 11908 4652 11912 4708
rect 11848 4648 11912 4652
rect 11848 4548 11912 4552
rect 11848 4492 11852 4548
rect 11852 4492 11908 4548
rect 11908 4492 11912 4548
rect 11848 4488 11912 4492
rect 11848 4388 11912 4392
rect 11848 4332 11852 4388
rect 11852 4332 11908 4388
rect 11908 4332 11912 4388
rect 11848 4328 11912 4332
rect 11848 4228 11912 4232
rect 11848 4172 11852 4228
rect 11852 4172 11908 4228
rect 11908 4172 11912 4228
rect 11848 4168 11912 4172
rect 11848 4068 11912 4072
rect 11848 4012 11852 4068
rect 11852 4012 11908 4068
rect 11908 4012 11912 4068
rect 11848 4008 11912 4012
rect 11848 3908 11912 3912
rect 11848 3852 11852 3908
rect 11852 3852 11908 3908
rect 11908 3852 11912 3908
rect 11848 3848 11912 3852
rect 11848 3688 11912 3752
rect 11848 3528 11912 3592
rect 11848 3428 11912 3432
rect 11848 3372 11852 3428
rect 11852 3372 11908 3428
rect 11908 3372 11912 3428
rect 11848 3368 11912 3372
rect 11848 3268 11912 3272
rect 11848 3212 11852 3268
rect 11852 3212 11908 3268
rect 11908 3212 11912 3268
rect 11848 3208 11912 3212
rect 11848 3108 11912 3112
rect 11848 3052 11852 3108
rect 11852 3052 11908 3108
rect 11908 3052 11912 3108
rect 11848 3048 11912 3052
rect 11848 2948 11912 2952
rect 11848 2892 11852 2948
rect 11852 2892 11908 2948
rect 11908 2892 11912 2948
rect 11848 2888 11912 2892
rect 11848 2788 11912 2792
rect 11848 2732 11852 2788
rect 11852 2732 11908 2788
rect 11908 2732 11912 2788
rect 11848 2728 11912 2732
rect 11848 2628 11912 2632
rect 11848 2572 11852 2628
rect 11852 2572 11908 2628
rect 11908 2572 11912 2628
rect 11848 2568 11912 2572
rect 11848 2468 11912 2472
rect 11848 2412 11852 2468
rect 11852 2412 11908 2468
rect 11908 2412 11912 2468
rect 11848 2408 11912 2412
rect 11848 2308 11912 2312
rect 11848 2252 11852 2308
rect 11852 2252 11908 2308
rect 11908 2252 11912 2308
rect 11848 2248 11912 2252
rect 11848 2148 11912 2152
rect 11848 2092 11852 2148
rect 11852 2092 11908 2148
rect 11908 2092 11912 2148
rect 11848 2088 11912 2092
rect 11848 1988 11912 1992
rect 11848 1932 11852 1988
rect 11852 1932 11908 1988
rect 11908 1932 11912 1988
rect 11848 1928 11912 1932
rect 11848 1768 11912 1832
rect 11848 1668 11912 1672
rect 11848 1612 11852 1668
rect 11852 1612 11908 1668
rect 11908 1612 11912 1668
rect 11848 1608 11912 1612
rect 11848 1508 11912 1512
rect 11848 1452 11852 1508
rect 11852 1452 11908 1508
rect 11908 1452 11912 1508
rect 11848 1448 11912 1452
rect 11848 1348 11912 1352
rect 11848 1292 11852 1348
rect 11852 1292 11908 1348
rect 11908 1292 11912 1348
rect 11848 1288 11912 1292
rect 11848 1188 11912 1192
rect 11848 1132 11852 1188
rect 11852 1132 11908 1188
rect 11908 1132 11912 1188
rect 11848 1128 11912 1132
rect 11848 1028 11912 1032
rect 11848 972 11852 1028
rect 11852 972 11908 1028
rect 11908 972 11912 1028
rect 11848 968 11912 972
rect 11848 808 11912 872
rect 11848 648 11912 712
rect 11848 548 11912 552
rect 11848 492 11852 548
rect 11852 492 11908 548
rect 11908 492 11912 548
rect 11848 488 11912 492
rect 11848 388 11912 392
rect 11848 332 11852 388
rect 11852 332 11908 388
rect 11908 332 11912 388
rect 11848 328 11912 332
rect 11848 228 11912 232
rect 11848 172 11852 228
rect 11852 172 11908 228
rect 11908 172 11912 228
rect 11848 168 11912 172
rect 11848 68 11912 72
rect 11848 12 11852 68
rect 11852 12 11908 68
rect 11908 12 11912 68
rect 11848 8 11912 12
rect 11528 -152 11592 -88
rect 11528 -232 11592 -168
rect 11528 -312 11592 -248
rect 11528 -392 11592 -328
rect 11528 -472 11592 -408
rect 11848 -152 11912 -88
rect 11848 -232 11912 -168
rect 11848 -312 11912 -248
rect 11848 -392 11912 -328
rect 11848 -472 11912 -408
rect 12008 31428 12072 31432
rect 12008 31372 12012 31428
rect 12012 31372 12068 31428
rect 12068 31372 12072 31428
rect 12008 31368 12072 31372
rect 12008 31268 12072 31272
rect 12008 31212 12012 31268
rect 12012 31212 12068 31268
rect 12068 31212 12072 31268
rect 12008 31208 12072 31212
rect 12008 31108 12072 31112
rect 12008 31052 12012 31108
rect 12012 31052 12068 31108
rect 12068 31052 12072 31108
rect 12008 31048 12072 31052
rect 12008 30948 12072 30952
rect 12008 30892 12012 30948
rect 12012 30892 12068 30948
rect 12068 30892 12072 30948
rect 12008 30888 12072 30892
rect 12008 30788 12072 30792
rect 12008 30732 12012 30788
rect 12012 30732 12068 30788
rect 12068 30732 12072 30788
rect 12008 30728 12072 30732
rect 12008 30628 12072 30632
rect 12008 30572 12012 30628
rect 12012 30572 12068 30628
rect 12068 30572 12072 30628
rect 12008 30568 12072 30572
rect 12008 30468 12072 30472
rect 12008 30412 12012 30468
rect 12012 30412 12068 30468
rect 12068 30412 12072 30468
rect 12008 30408 12072 30412
rect 12008 30308 12072 30312
rect 12008 30252 12012 30308
rect 12012 30252 12068 30308
rect 12068 30252 12072 30308
rect 12008 30248 12072 30252
rect 12008 30088 12072 30152
rect 12008 29988 12072 29992
rect 12008 29932 12012 29988
rect 12012 29932 12068 29988
rect 12068 29932 12072 29988
rect 12008 29928 12072 29932
rect 12008 29828 12072 29832
rect 12008 29772 12012 29828
rect 12012 29772 12068 29828
rect 12068 29772 12072 29828
rect 12008 29768 12072 29772
rect 12008 29668 12072 29672
rect 12008 29612 12012 29668
rect 12012 29612 12068 29668
rect 12068 29612 12072 29668
rect 12008 29608 12072 29612
rect 12008 29508 12072 29512
rect 12008 29452 12012 29508
rect 12012 29452 12068 29508
rect 12068 29452 12072 29508
rect 12008 29448 12072 29452
rect 12008 29348 12072 29352
rect 12008 29292 12012 29348
rect 12012 29292 12068 29348
rect 12068 29292 12072 29348
rect 12008 29288 12072 29292
rect 12008 29188 12072 29192
rect 12008 29132 12012 29188
rect 12012 29132 12068 29188
rect 12068 29132 12072 29188
rect 12008 29128 12072 29132
rect 12008 29028 12072 29032
rect 12008 28972 12012 29028
rect 12012 28972 12068 29028
rect 12068 28972 12072 29028
rect 12008 28968 12072 28972
rect 12008 28868 12072 28872
rect 12008 28812 12012 28868
rect 12012 28812 12068 28868
rect 12068 28812 12072 28868
rect 12008 28808 12072 28812
rect 12008 28648 12072 28712
rect 12008 28488 12072 28552
rect 12008 28328 12072 28392
rect 12008 28168 12072 28232
rect 12008 28068 12072 28072
rect 12008 28012 12012 28068
rect 12012 28012 12068 28068
rect 12068 28012 12072 28068
rect 12008 28008 12072 28012
rect 12008 27908 12072 27912
rect 12008 27852 12012 27908
rect 12012 27852 12068 27908
rect 12068 27852 12072 27908
rect 12008 27848 12072 27852
rect 12008 27748 12072 27752
rect 12008 27692 12012 27748
rect 12012 27692 12068 27748
rect 12068 27692 12072 27748
rect 12008 27688 12072 27692
rect 12008 27588 12072 27592
rect 12008 27532 12012 27588
rect 12012 27532 12068 27588
rect 12068 27532 12072 27588
rect 12008 27528 12072 27532
rect 12008 27428 12072 27432
rect 12008 27372 12012 27428
rect 12012 27372 12068 27428
rect 12068 27372 12072 27428
rect 12008 27368 12072 27372
rect 12008 27268 12072 27272
rect 12008 27212 12012 27268
rect 12012 27212 12068 27268
rect 12068 27212 12072 27268
rect 12008 27208 12072 27212
rect 12008 27108 12072 27112
rect 12008 27052 12012 27108
rect 12012 27052 12068 27108
rect 12068 27052 12072 27108
rect 12008 27048 12072 27052
rect 12008 26948 12072 26952
rect 12008 26892 12012 26948
rect 12012 26892 12068 26948
rect 12068 26892 12072 26948
rect 12008 26888 12072 26892
rect 12008 26728 12072 26792
rect 12008 26568 12072 26632
rect 12008 26408 12072 26472
rect 12008 26248 12072 26312
rect 12008 26148 12072 26152
rect 12008 26092 12012 26148
rect 12012 26092 12068 26148
rect 12068 26092 12072 26148
rect 12008 26088 12072 26092
rect 12008 25988 12072 25992
rect 12008 25932 12012 25988
rect 12012 25932 12068 25988
rect 12068 25932 12072 25988
rect 12008 25928 12072 25932
rect 12008 25828 12072 25832
rect 12008 25772 12012 25828
rect 12012 25772 12068 25828
rect 12068 25772 12072 25828
rect 12008 25768 12072 25772
rect 12008 25668 12072 25672
rect 12008 25612 12012 25668
rect 12012 25612 12068 25668
rect 12068 25612 12072 25668
rect 12008 25608 12072 25612
rect 12008 25508 12072 25512
rect 12008 25452 12012 25508
rect 12012 25452 12068 25508
rect 12068 25452 12072 25508
rect 12008 25448 12072 25452
rect 12008 25348 12072 25352
rect 12008 25292 12012 25348
rect 12012 25292 12068 25348
rect 12068 25292 12072 25348
rect 12008 25288 12072 25292
rect 12008 25188 12072 25192
rect 12008 25132 12012 25188
rect 12012 25132 12068 25188
rect 12068 25132 12072 25188
rect 12008 25128 12072 25132
rect 12008 25028 12072 25032
rect 12008 24972 12012 25028
rect 12012 24972 12068 25028
rect 12068 24972 12072 25028
rect 12008 24968 12072 24972
rect 12008 24808 12072 24872
rect 12008 24708 12072 24712
rect 12008 24652 12012 24708
rect 12012 24652 12068 24708
rect 12068 24652 12072 24708
rect 12008 24648 12072 24652
rect 12008 24548 12072 24552
rect 12008 24492 12012 24548
rect 12012 24492 12068 24548
rect 12068 24492 12072 24548
rect 12008 24488 12072 24492
rect 12008 24388 12072 24392
rect 12008 24332 12012 24388
rect 12012 24332 12068 24388
rect 12068 24332 12072 24388
rect 12008 24328 12072 24332
rect 12008 24228 12072 24232
rect 12008 24172 12012 24228
rect 12012 24172 12068 24228
rect 12068 24172 12072 24228
rect 12008 24168 12072 24172
rect 12008 24068 12072 24072
rect 12008 24012 12012 24068
rect 12012 24012 12068 24068
rect 12068 24012 12072 24068
rect 12008 24008 12072 24012
rect 12008 23908 12072 23912
rect 12008 23852 12012 23908
rect 12012 23852 12068 23908
rect 12068 23852 12072 23908
rect 12008 23848 12072 23852
rect 12008 23748 12072 23752
rect 12008 23692 12012 23748
rect 12012 23692 12068 23748
rect 12068 23692 12072 23748
rect 12008 23688 12072 23692
rect 12008 23588 12072 23592
rect 12008 23532 12012 23588
rect 12012 23532 12068 23588
rect 12068 23532 12072 23588
rect 12008 23528 12072 23532
rect 12008 23428 12072 23432
rect 12008 23372 12012 23428
rect 12012 23372 12068 23428
rect 12068 23372 12072 23428
rect 12008 23368 12072 23372
rect 12008 23268 12072 23272
rect 12008 23212 12012 23268
rect 12012 23212 12068 23268
rect 12068 23212 12072 23268
rect 12008 23208 12072 23212
rect 12008 23108 12072 23112
rect 12008 23052 12012 23108
rect 12012 23052 12068 23108
rect 12068 23052 12072 23108
rect 12008 23048 12072 23052
rect 12008 22948 12072 22952
rect 12008 22892 12012 22948
rect 12012 22892 12068 22948
rect 12068 22892 12072 22948
rect 12008 22888 12072 22892
rect 12008 22788 12072 22792
rect 12008 22732 12012 22788
rect 12012 22732 12068 22788
rect 12068 22732 12072 22788
rect 12008 22728 12072 22732
rect 12008 22628 12072 22632
rect 12008 22572 12012 22628
rect 12012 22572 12068 22628
rect 12068 22572 12072 22628
rect 12008 22568 12072 22572
rect 12008 22468 12072 22472
rect 12008 22412 12012 22468
rect 12012 22412 12068 22468
rect 12068 22412 12072 22468
rect 12008 22408 12072 22412
rect 12008 22308 12072 22312
rect 12008 22252 12012 22308
rect 12012 22252 12068 22308
rect 12068 22252 12072 22308
rect 12008 22248 12072 22252
rect 12008 22148 12072 22152
rect 12008 22092 12012 22148
rect 12012 22092 12068 22148
rect 12068 22092 12072 22148
rect 12008 22088 12072 22092
rect 12008 21928 12072 21992
rect 12008 21828 12072 21832
rect 12008 21772 12012 21828
rect 12012 21772 12068 21828
rect 12068 21772 12072 21828
rect 12008 21768 12072 21772
rect 12008 21668 12072 21672
rect 12008 21612 12012 21668
rect 12012 21612 12068 21668
rect 12068 21612 12072 21668
rect 12008 21608 12072 21612
rect 12008 21508 12072 21512
rect 12008 21452 12012 21508
rect 12012 21452 12068 21508
rect 12068 21452 12072 21508
rect 12008 21448 12072 21452
rect 12008 21348 12072 21352
rect 12008 21292 12012 21348
rect 12012 21292 12068 21348
rect 12068 21292 12072 21348
rect 12008 21288 12072 21292
rect 12008 21188 12072 21192
rect 12008 21132 12012 21188
rect 12012 21132 12068 21188
rect 12068 21132 12072 21188
rect 12008 21128 12072 21132
rect 12008 21028 12072 21032
rect 12008 20972 12012 21028
rect 12012 20972 12068 21028
rect 12068 20972 12072 21028
rect 12008 20968 12072 20972
rect 12008 20868 12072 20872
rect 12008 20812 12012 20868
rect 12012 20812 12068 20868
rect 12068 20812 12072 20868
rect 12008 20808 12072 20812
rect 12008 20708 12072 20712
rect 12008 20652 12012 20708
rect 12012 20652 12068 20708
rect 12068 20652 12072 20708
rect 12008 20648 12072 20652
rect 12008 20488 12072 20552
rect 12008 20328 12072 20392
rect 12008 20168 12072 20232
rect 12008 20008 12072 20072
rect 12008 19908 12072 19912
rect 12008 19852 12012 19908
rect 12012 19852 12068 19908
rect 12068 19852 12072 19908
rect 12008 19848 12072 19852
rect 12008 19748 12072 19752
rect 12008 19692 12012 19748
rect 12012 19692 12068 19748
rect 12068 19692 12072 19748
rect 12008 19688 12072 19692
rect 12008 19588 12072 19592
rect 12008 19532 12012 19588
rect 12012 19532 12068 19588
rect 12068 19532 12072 19588
rect 12008 19528 12072 19532
rect 12008 19428 12072 19432
rect 12008 19372 12012 19428
rect 12012 19372 12068 19428
rect 12068 19372 12072 19428
rect 12008 19368 12072 19372
rect 12008 19268 12072 19272
rect 12008 19212 12012 19268
rect 12012 19212 12068 19268
rect 12068 19212 12072 19268
rect 12008 19208 12072 19212
rect 12008 19108 12072 19112
rect 12008 19052 12012 19108
rect 12012 19052 12068 19108
rect 12068 19052 12072 19108
rect 12008 19048 12072 19052
rect 12008 18948 12072 18952
rect 12008 18892 12012 18948
rect 12012 18892 12068 18948
rect 12068 18892 12072 18948
rect 12008 18888 12072 18892
rect 12008 18788 12072 18792
rect 12008 18732 12012 18788
rect 12012 18732 12068 18788
rect 12068 18732 12072 18788
rect 12008 18728 12072 18732
rect 12008 18568 12072 18632
rect 12008 18408 12072 18472
rect 12008 18248 12072 18312
rect 12008 18088 12072 18152
rect 12008 17988 12072 17992
rect 12008 17932 12012 17988
rect 12012 17932 12068 17988
rect 12068 17932 12072 17988
rect 12008 17928 12072 17932
rect 12008 17828 12072 17832
rect 12008 17772 12012 17828
rect 12012 17772 12068 17828
rect 12068 17772 12072 17828
rect 12008 17768 12072 17772
rect 12008 17668 12072 17672
rect 12008 17612 12012 17668
rect 12012 17612 12068 17668
rect 12068 17612 12072 17668
rect 12008 17608 12072 17612
rect 12008 17508 12072 17512
rect 12008 17452 12012 17508
rect 12012 17452 12068 17508
rect 12068 17452 12072 17508
rect 12008 17448 12072 17452
rect 12008 17348 12072 17352
rect 12008 17292 12012 17348
rect 12012 17292 12068 17348
rect 12068 17292 12072 17348
rect 12008 17288 12072 17292
rect 12008 17188 12072 17192
rect 12008 17132 12012 17188
rect 12012 17132 12068 17188
rect 12068 17132 12072 17188
rect 12008 17128 12072 17132
rect 12008 17028 12072 17032
rect 12008 16972 12012 17028
rect 12012 16972 12068 17028
rect 12068 16972 12072 17028
rect 12008 16968 12072 16972
rect 12008 16868 12072 16872
rect 12008 16812 12012 16868
rect 12012 16812 12068 16868
rect 12068 16812 12072 16868
rect 12008 16808 12072 16812
rect 12008 16648 12072 16712
rect 12008 16548 12072 16552
rect 12008 16492 12012 16548
rect 12012 16492 12068 16548
rect 12068 16492 12072 16548
rect 12008 16488 12072 16492
rect 12008 16388 12072 16392
rect 12008 16332 12012 16388
rect 12012 16332 12068 16388
rect 12068 16332 12072 16388
rect 12008 16328 12072 16332
rect 12008 16228 12072 16232
rect 12008 16172 12012 16228
rect 12012 16172 12068 16228
rect 12068 16172 12072 16228
rect 12008 16168 12072 16172
rect 12008 16068 12072 16072
rect 12008 16012 12012 16068
rect 12012 16012 12068 16068
rect 12068 16012 12072 16068
rect 12008 16008 12072 16012
rect 12008 15908 12072 15912
rect 12008 15852 12012 15908
rect 12012 15852 12068 15908
rect 12068 15852 12072 15908
rect 12008 15848 12072 15852
rect 12008 15748 12072 15752
rect 12008 15692 12012 15748
rect 12012 15692 12068 15748
rect 12068 15692 12072 15748
rect 12008 15688 12072 15692
rect 12008 15588 12072 15592
rect 12008 15532 12012 15588
rect 12012 15532 12068 15588
rect 12068 15532 12072 15588
rect 12008 15528 12072 15532
rect 12008 15428 12072 15432
rect 12008 15372 12012 15428
rect 12012 15372 12068 15428
rect 12068 15372 12072 15428
rect 12008 15368 12072 15372
rect 12008 15268 12072 15272
rect 12008 15212 12012 15268
rect 12012 15212 12068 15268
rect 12068 15212 12072 15268
rect 12008 15208 12072 15212
rect 12008 15108 12072 15112
rect 12008 15052 12012 15108
rect 12012 15052 12068 15108
rect 12068 15052 12072 15108
rect 12008 15048 12072 15052
rect 12008 14948 12072 14952
rect 12008 14892 12012 14948
rect 12012 14892 12068 14948
rect 12068 14892 12072 14948
rect 12008 14888 12072 14892
rect 12008 14788 12072 14792
rect 12008 14732 12012 14788
rect 12012 14732 12068 14788
rect 12068 14732 12072 14788
rect 12008 14728 12072 14732
rect 12008 14628 12072 14632
rect 12008 14572 12012 14628
rect 12012 14572 12068 14628
rect 12068 14572 12072 14628
rect 12008 14568 12072 14572
rect 12008 14468 12072 14472
rect 12008 14412 12012 14468
rect 12012 14412 12068 14468
rect 12068 14412 12072 14468
rect 12008 14408 12072 14412
rect 12008 14308 12072 14312
rect 12008 14252 12012 14308
rect 12012 14252 12068 14308
rect 12068 14252 12072 14308
rect 12008 14248 12072 14252
rect 12008 14148 12072 14152
rect 12008 14092 12012 14148
rect 12012 14092 12068 14148
rect 12068 14092 12072 14148
rect 12008 14088 12072 14092
rect 12008 13988 12072 13992
rect 12008 13932 12012 13988
rect 12012 13932 12068 13988
rect 12068 13932 12072 13988
rect 12008 13928 12072 13932
rect 12008 13768 12072 13832
rect 12008 13668 12072 13672
rect 12008 13612 12012 13668
rect 12012 13612 12068 13668
rect 12068 13612 12072 13668
rect 12008 13608 12072 13612
rect 12008 13508 12072 13512
rect 12008 13452 12012 13508
rect 12012 13452 12068 13508
rect 12068 13452 12072 13508
rect 12008 13448 12072 13452
rect 12008 13348 12072 13352
rect 12008 13292 12012 13348
rect 12012 13292 12068 13348
rect 12068 13292 12072 13348
rect 12008 13288 12072 13292
rect 12008 13188 12072 13192
rect 12008 13132 12012 13188
rect 12012 13132 12068 13188
rect 12068 13132 12072 13188
rect 12008 13128 12072 13132
rect 12008 13028 12072 13032
rect 12008 12972 12012 13028
rect 12012 12972 12068 13028
rect 12068 12972 12072 13028
rect 12008 12968 12072 12972
rect 12008 12868 12072 12872
rect 12008 12812 12012 12868
rect 12012 12812 12068 12868
rect 12068 12812 12072 12868
rect 12008 12808 12072 12812
rect 12008 12708 12072 12712
rect 12008 12652 12012 12708
rect 12012 12652 12068 12708
rect 12068 12652 12072 12708
rect 12008 12648 12072 12652
rect 12008 12548 12072 12552
rect 12008 12492 12012 12548
rect 12012 12492 12068 12548
rect 12068 12492 12072 12548
rect 12008 12488 12072 12492
rect 12008 12328 12072 12392
rect 12008 12168 12072 12232
rect 12008 12008 12072 12072
rect 12008 11848 12072 11912
rect 12008 11748 12072 11752
rect 12008 11692 12012 11748
rect 12012 11692 12068 11748
rect 12068 11692 12072 11748
rect 12008 11688 12072 11692
rect 12008 11588 12072 11592
rect 12008 11532 12012 11588
rect 12012 11532 12068 11588
rect 12068 11532 12072 11588
rect 12008 11528 12072 11532
rect 12008 11428 12072 11432
rect 12008 11372 12012 11428
rect 12012 11372 12068 11428
rect 12068 11372 12072 11428
rect 12008 11368 12072 11372
rect 12008 11268 12072 11272
rect 12008 11212 12012 11268
rect 12012 11212 12068 11268
rect 12068 11212 12072 11268
rect 12008 11208 12072 11212
rect 12008 11108 12072 11112
rect 12008 11052 12012 11108
rect 12012 11052 12068 11108
rect 12068 11052 12072 11108
rect 12008 11048 12072 11052
rect 12008 10948 12072 10952
rect 12008 10892 12012 10948
rect 12012 10892 12068 10948
rect 12068 10892 12072 10948
rect 12008 10888 12072 10892
rect 12008 10788 12072 10792
rect 12008 10732 12012 10788
rect 12012 10732 12068 10788
rect 12068 10732 12072 10788
rect 12008 10728 12072 10732
rect 12008 10628 12072 10632
rect 12008 10572 12012 10628
rect 12012 10572 12068 10628
rect 12068 10572 12072 10628
rect 12008 10568 12072 10572
rect 12008 10468 12072 10472
rect 12008 10412 12012 10468
rect 12012 10412 12068 10468
rect 12068 10412 12072 10468
rect 12008 10408 12072 10412
rect 12008 10308 12072 10312
rect 12008 10252 12012 10308
rect 12012 10252 12068 10308
rect 12068 10252 12072 10308
rect 12008 10248 12072 10252
rect 12008 10148 12072 10152
rect 12008 10092 12012 10148
rect 12012 10092 12068 10148
rect 12068 10092 12072 10148
rect 12008 10088 12072 10092
rect 12008 9988 12072 9992
rect 12008 9932 12012 9988
rect 12012 9932 12068 9988
rect 12068 9932 12072 9988
rect 12008 9928 12072 9932
rect 12008 9828 12072 9832
rect 12008 9772 12012 9828
rect 12012 9772 12068 9828
rect 12068 9772 12072 9828
rect 12008 9768 12072 9772
rect 12008 9608 12072 9672
rect 12008 9508 12072 9512
rect 12008 9452 12012 9508
rect 12012 9452 12068 9508
rect 12068 9452 12072 9508
rect 12008 9448 12072 9452
rect 12008 9348 12072 9352
rect 12008 9292 12012 9348
rect 12012 9292 12068 9348
rect 12068 9292 12072 9348
rect 12008 9288 12072 9292
rect 12008 9128 12072 9192
rect 12008 9028 12072 9032
rect 12008 8972 12012 9028
rect 12012 8972 12068 9028
rect 12068 8972 12072 9028
rect 12008 8968 12072 8972
rect 12008 8868 12072 8872
rect 12008 8812 12012 8868
rect 12012 8812 12068 8868
rect 12068 8812 12072 8868
rect 12008 8808 12072 8812
rect 12008 8708 12072 8712
rect 12008 8652 12012 8708
rect 12012 8652 12068 8708
rect 12068 8652 12072 8708
rect 12008 8648 12072 8652
rect 12008 8548 12072 8552
rect 12008 8492 12012 8548
rect 12012 8492 12068 8548
rect 12068 8492 12072 8548
rect 12008 8488 12072 8492
rect 12008 8388 12072 8392
rect 12008 8332 12012 8388
rect 12012 8332 12068 8388
rect 12068 8332 12072 8388
rect 12008 8328 12072 8332
rect 12008 8228 12072 8232
rect 12008 8172 12012 8228
rect 12012 8172 12068 8228
rect 12068 8172 12072 8228
rect 12008 8168 12072 8172
rect 12008 8068 12072 8072
rect 12008 8012 12012 8068
rect 12012 8012 12068 8068
rect 12068 8012 12072 8068
rect 12008 8008 12072 8012
rect 12008 7908 12072 7912
rect 12008 7852 12012 7908
rect 12012 7852 12068 7908
rect 12068 7852 12072 7908
rect 12008 7848 12072 7852
rect 12008 7748 12072 7752
rect 12008 7692 12012 7748
rect 12012 7692 12068 7748
rect 12068 7692 12072 7748
rect 12008 7688 12072 7692
rect 12008 7528 12072 7592
rect 12008 7428 12072 7432
rect 12008 7372 12012 7428
rect 12012 7372 12068 7428
rect 12068 7372 12072 7428
rect 12008 7368 12072 7372
rect 12008 7268 12072 7272
rect 12008 7212 12012 7268
rect 12012 7212 12068 7268
rect 12068 7212 12072 7268
rect 12008 7208 12072 7212
rect 12008 7048 12072 7112
rect 12008 6948 12072 6952
rect 12008 6892 12012 6948
rect 12012 6892 12068 6948
rect 12068 6892 12072 6948
rect 12008 6888 12072 6892
rect 12008 6788 12072 6792
rect 12008 6732 12012 6788
rect 12012 6732 12068 6788
rect 12068 6732 12072 6788
rect 12008 6728 12072 6732
rect 12008 6568 12072 6632
rect 12008 6468 12072 6472
rect 12008 6412 12012 6468
rect 12012 6412 12068 6468
rect 12068 6412 12072 6468
rect 12008 6408 12072 6412
rect 12008 6308 12072 6312
rect 12008 6252 12012 6308
rect 12012 6252 12068 6308
rect 12068 6252 12072 6308
rect 12008 6248 12072 6252
rect 12008 6148 12072 6152
rect 12008 6092 12012 6148
rect 12012 6092 12068 6148
rect 12068 6092 12072 6148
rect 12008 6088 12072 6092
rect 12008 5988 12072 5992
rect 12008 5932 12012 5988
rect 12012 5932 12068 5988
rect 12068 5932 12072 5988
rect 12008 5928 12072 5932
rect 12008 5828 12072 5832
rect 12008 5772 12012 5828
rect 12012 5772 12068 5828
rect 12068 5772 12072 5828
rect 12008 5768 12072 5772
rect 12008 5668 12072 5672
rect 12008 5612 12012 5668
rect 12012 5612 12068 5668
rect 12068 5612 12072 5668
rect 12008 5608 12072 5612
rect 12008 5508 12072 5512
rect 12008 5452 12012 5508
rect 12012 5452 12068 5508
rect 12068 5452 12072 5508
rect 12008 5448 12072 5452
rect 12008 5348 12072 5352
rect 12008 5292 12012 5348
rect 12012 5292 12068 5348
rect 12068 5292 12072 5348
rect 12008 5288 12072 5292
rect 12008 5188 12072 5192
rect 12008 5132 12012 5188
rect 12012 5132 12068 5188
rect 12068 5132 12072 5188
rect 12008 5128 12072 5132
rect 12008 5028 12072 5032
rect 12008 4972 12012 5028
rect 12012 4972 12068 5028
rect 12068 4972 12072 5028
rect 12008 4968 12072 4972
rect 12008 4868 12072 4872
rect 12008 4812 12012 4868
rect 12012 4812 12068 4868
rect 12068 4812 12072 4868
rect 12008 4808 12072 4812
rect 12008 4708 12072 4712
rect 12008 4652 12012 4708
rect 12012 4652 12068 4708
rect 12068 4652 12072 4708
rect 12008 4648 12072 4652
rect 12008 4548 12072 4552
rect 12008 4492 12012 4548
rect 12012 4492 12068 4548
rect 12068 4492 12072 4548
rect 12008 4488 12072 4492
rect 12008 4388 12072 4392
rect 12008 4332 12012 4388
rect 12012 4332 12068 4388
rect 12068 4332 12072 4388
rect 12008 4328 12072 4332
rect 12008 4228 12072 4232
rect 12008 4172 12012 4228
rect 12012 4172 12068 4228
rect 12068 4172 12072 4228
rect 12008 4168 12072 4172
rect 12008 4068 12072 4072
rect 12008 4012 12012 4068
rect 12012 4012 12068 4068
rect 12068 4012 12072 4068
rect 12008 4008 12072 4012
rect 12008 3908 12072 3912
rect 12008 3852 12012 3908
rect 12012 3852 12068 3908
rect 12068 3852 12072 3908
rect 12008 3848 12072 3852
rect 12008 3688 12072 3752
rect 12008 3528 12072 3592
rect 12008 3428 12072 3432
rect 12008 3372 12012 3428
rect 12012 3372 12068 3428
rect 12068 3372 12072 3428
rect 12008 3368 12072 3372
rect 12008 3268 12072 3272
rect 12008 3212 12012 3268
rect 12012 3212 12068 3268
rect 12068 3212 12072 3268
rect 12008 3208 12072 3212
rect 12008 3108 12072 3112
rect 12008 3052 12012 3108
rect 12012 3052 12068 3108
rect 12068 3052 12072 3108
rect 12008 3048 12072 3052
rect 12008 2948 12072 2952
rect 12008 2892 12012 2948
rect 12012 2892 12068 2948
rect 12068 2892 12072 2948
rect 12008 2888 12072 2892
rect 12008 2788 12072 2792
rect 12008 2732 12012 2788
rect 12012 2732 12068 2788
rect 12068 2732 12072 2788
rect 12008 2728 12072 2732
rect 12008 2628 12072 2632
rect 12008 2572 12012 2628
rect 12012 2572 12068 2628
rect 12068 2572 12072 2628
rect 12008 2568 12072 2572
rect 12008 2468 12072 2472
rect 12008 2412 12012 2468
rect 12012 2412 12068 2468
rect 12068 2412 12072 2468
rect 12008 2408 12072 2412
rect 12008 2308 12072 2312
rect 12008 2252 12012 2308
rect 12012 2252 12068 2308
rect 12068 2252 12072 2308
rect 12008 2248 12072 2252
rect 12008 2148 12072 2152
rect 12008 2092 12012 2148
rect 12012 2092 12068 2148
rect 12068 2092 12072 2148
rect 12008 2088 12072 2092
rect 12008 1988 12072 1992
rect 12008 1932 12012 1988
rect 12012 1932 12068 1988
rect 12068 1932 12072 1988
rect 12008 1928 12072 1932
rect 12008 1768 12072 1832
rect 12008 1668 12072 1672
rect 12008 1612 12012 1668
rect 12012 1612 12068 1668
rect 12068 1612 12072 1668
rect 12008 1608 12072 1612
rect 12008 1508 12072 1512
rect 12008 1452 12012 1508
rect 12012 1452 12068 1508
rect 12068 1452 12072 1508
rect 12008 1448 12072 1452
rect 12008 1348 12072 1352
rect 12008 1292 12012 1348
rect 12012 1292 12068 1348
rect 12068 1292 12072 1348
rect 12008 1288 12072 1292
rect 12008 1188 12072 1192
rect 12008 1132 12012 1188
rect 12012 1132 12068 1188
rect 12068 1132 12072 1188
rect 12008 1128 12072 1132
rect 12008 1028 12072 1032
rect 12008 972 12012 1028
rect 12012 972 12068 1028
rect 12068 972 12072 1028
rect 12008 968 12072 972
rect 12008 808 12072 872
rect 12008 648 12072 712
rect 12008 548 12072 552
rect 12008 492 12012 548
rect 12012 492 12068 548
rect 12068 492 12072 548
rect 12008 488 12072 492
rect 12008 388 12072 392
rect 12008 332 12012 388
rect 12012 332 12068 388
rect 12068 332 12072 388
rect 12008 328 12072 332
rect 12008 228 12072 232
rect 12008 172 12012 228
rect 12012 172 12068 228
rect 12068 172 12072 228
rect 12008 168 12072 172
rect 12008 68 12072 72
rect 12008 12 12012 68
rect 12012 12 12068 68
rect 12068 12 12072 68
rect 12008 8 12072 12
rect 12328 31428 12392 31432
rect 12328 31372 12332 31428
rect 12332 31372 12388 31428
rect 12388 31372 12392 31428
rect 12328 31368 12392 31372
rect 12328 31268 12392 31272
rect 12328 31212 12332 31268
rect 12332 31212 12388 31268
rect 12388 31212 12392 31268
rect 12328 31208 12392 31212
rect 12328 31108 12392 31112
rect 12328 31052 12332 31108
rect 12332 31052 12388 31108
rect 12388 31052 12392 31108
rect 12328 31048 12392 31052
rect 12328 30948 12392 30952
rect 12328 30892 12332 30948
rect 12332 30892 12388 30948
rect 12388 30892 12392 30948
rect 12328 30888 12392 30892
rect 12328 30788 12392 30792
rect 12328 30732 12332 30788
rect 12332 30732 12388 30788
rect 12388 30732 12392 30788
rect 12328 30728 12392 30732
rect 12328 30628 12392 30632
rect 12328 30572 12332 30628
rect 12332 30572 12388 30628
rect 12388 30572 12392 30628
rect 12328 30568 12392 30572
rect 12328 30468 12392 30472
rect 12328 30412 12332 30468
rect 12332 30412 12388 30468
rect 12388 30412 12392 30468
rect 12328 30408 12392 30412
rect 12328 30308 12392 30312
rect 12328 30252 12332 30308
rect 12332 30252 12388 30308
rect 12388 30252 12392 30308
rect 12328 30248 12392 30252
rect 12328 30088 12392 30152
rect 12328 29988 12392 29992
rect 12328 29932 12332 29988
rect 12332 29932 12388 29988
rect 12388 29932 12392 29988
rect 12328 29928 12392 29932
rect 12328 29828 12392 29832
rect 12328 29772 12332 29828
rect 12332 29772 12388 29828
rect 12388 29772 12392 29828
rect 12328 29768 12392 29772
rect 12328 29668 12392 29672
rect 12328 29612 12332 29668
rect 12332 29612 12388 29668
rect 12388 29612 12392 29668
rect 12328 29608 12392 29612
rect 12328 29508 12392 29512
rect 12328 29452 12332 29508
rect 12332 29452 12388 29508
rect 12388 29452 12392 29508
rect 12328 29448 12392 29452
rect 12328 29348 12392 29352
rect 12328 29292 12332 29348
rect 12332 29292 12388 29348
rect 12388 29292 12392 29348
rect 12328 29288 12392 29292
rect 12328 29188 12392 29192
rect 12328 29132 12332 29188
rect 12332 29132 12388 29188
rect 12388 29132 12392 29188
rect 12328 29128 12392 29132
rect 12328 29028 12392 29032
rect 12328 28972 12332 29028
rect 12332 28972 12388 29028
rect 12388 28972 12392 29028
rect 12328 28968 12392 28972
rect 12328 28868 12392 28872
rect 12328 28812 12332 28868
rect 12332 28812 12388 28868
rect 12388 28812 12392 28868
rect 12328 28808 12392 28812
rect 12328 28648 12392 28712
rect 12328 28488 12392 28552
rect 12328 28328 12392 28392
rect 12328 28168 12392 28232
rect 12328 28068 12392 28072
rect 12328 28012 12332 28068
rect 12332 28012 12388 28068
rect 12388 28012 12392 28068
rect 12328 28008 12392 28012
rect 12328 27908 12392 27912
rect 12328 27852 12332 27908
rect 12332 27852 12388 27908
rect 12388 27852 12392 27908
rect 12328 27848 12392 27852
rect 12328 27748 12392 27752
rect 12328 27692 12332 27748
rect 12332 27692 12388 27748
rect 12388 27692 12392 27748
rect 12328 27688 12392 27692
rect 12328 27588 12392 27592
rect 12328 27532 12332 27588
rect 12332 27532 12388 27588
rect 12388 27532 12392 27588
rect 12328 27528 12392 27532
rect 12328 27428 12392 27432
rect 12328 27372 12332 27428
rect 12332 27372 12388 27428
rect 12388 27372 12392 27428
rect 12328 27368 12392 27372
rect 12328 27268 12392 27272
rect 12328 27212 12332 27268
rect 12332 27212 12388 27268
rect 12388 27212 12392 27268
rect 12328 27208 12392 27212
rect 12328 27108 12392 27112
rect 12328 27052 12332 27108
rect 12332 27052 12388 27108
rect 12388 27052 12392 27108
rect 12328 27048 12392 27052
rect 12328 26948 12392 26952
rect 12328 26892 12332 26948
rect 12332 26892 12388 26948
rect 12388 26892 12392 26948
rect 12328 26888 12392 26892
rect 12328 26728 12392 26792
rect 12328 26568 12392 26632
rect 12328 26408 12392 26472
rect 12328 26248 12392 26312
rect 12328 26148 12392 26152
rect 12328 26092 12332 26148
rect 12332 26092 12388 26148
rect 12388 26092 12392 26148
rect 12328 26088 12392 26092
rect 12328 25988 12392 25992
rect 12328 25932 12332 25988
rect 12332 25932 12388 25988
rect 12388 25932 12392 25988
rect 12328 25928 12392 25932
rect 12328 25828 12392 25832
rect 12328 25772 12332 25828
rect 12332 25772 12388 25828
rect 12388 25772 12392 25828
rect 12328 25768 12392 25772
rect 12328 25668 12392 25672
rect 12328 25612 12332 25668
rect 12332 25612 12388 25668
rect 12388 25612 12392 25668
rect 12328 25608 12392 25612
rect 12328 25508 12392 25512
rect 12328 25452 12332 25508
rect 12332 25452 12388 25508
rect 12388 25452 12392 25508
rect 12328 25448 12392 25452
rect 12328 25348 12392 25352
rect 12328 25292 12332 25348
rect 12332 25292 12388 25348
rect 12388 25292 12392 25348
rect 12328 25288 12392 25292
rect 12328 25188 12392 25192
rect 12328 25132 12332 25188
rect 12332 25132 12388 25188
rect 12388 25132 12392 25188
rect 12328 25128 12392 25132
rect 12328 25028 12392 25032
rect 12328 24972 12332 25028
rect 12332 24972 12388 25028
rect 12388 24972 12392 25028
rect 12328 24968 12392 24972
rect 12328 24808 12392 24872
rect 12328 24708 12392 24712
rect 12328 24652 12332 24708
rect 12332 24652 12388 24708
rect 12388 24652 12392 24708
rect 12328 24648 12392 24652
rect 12328 24548 12392 24552
rect 12328 24492 12332 24548
rect 12332 24492 12388 24548
rect 12388 24492 12392 24548
rect 12328 24488 12392 24492
rect 12328 24388 12392 24392
rect 12328 24332 12332 24388
rect 12332 24332 12388 24388
rect 12388 24332 12392 24388
rect 12328 24328 12392 24332
rect 12328 24228 12392 24232
rect 12328 24172 12332 24228
rect 12332 24172 12388 24228
rect 12388 24172 12392 24228
rect 12328 24168 12392 24172
rect 12328 24068 12392 24072
rect 12328 24012 12332 24068
rect 12332 24012 12388 24068
rect 12388 24012 12392 24068
rect 12328 24008 12392 24012
rect 12328 23908 12392 23912
rect 12328 23852 12332 23908
rect 12332 23852 12388 23908
rect 12388 23852 12392 23908
rect 12328 23848 12392 23852
rect 12328 23748 12392 23752
rect 12328 23692 12332 23748
rect 12332 23692 12388 23748
rect 12388 23692 12392 23748
rect 12328 23688 12392 23692
rect 12328 23588 12392 23592
rect 12328 23532 12332 23588
rect 12332 23532 12388 23588
rect 12388 23532 12392 23588
rect 12328 23528 12392 23532
rect 12328 23428 12392 23432
rect 12328 23372 12332 23428
rect 12332 23372 12388 23428
rect 12388 23372 12392 23428
rect 12328 23368 12392 23372
rect 12328 23268 12392 23272
rect 12328 23212 12332 23268
rect 12332 23212 12388 23268
rect 12388 23212 12392 23268
rect 12328 23208 12392 23212
rect 12328 23108 12392 23112
rect 12328 23052 12332 23108
rect 12332 23052 12388 23108
rect 12388 23052 12392 23108
rect 12328 23048 12392 23052
rect 12328 22948 12392 22952
rect 12328 22892 12332 22948
rect 12332 22892 12388 22948
rect 12388 22892 12392 22948
rect 12328 22888 12392 22892
rect 12328 22788 12392 22792
rect 12328 22732 12332 22788
rect 12332 22732 12388 22788
rect 12388 22732 12392 22788
rect 12328 22728 12392 22732
rect 12328 22628 12392 22632
rect 12328 22572 12332 22628
rect 12332 22572 12388 22628
rect 12388 22572 12392 22628
rect 12328 22568 12392 22572
rect 12328 22468 12392 22472
rect 12328 22412 12332 22468
rect 12332 22412 12388 22468
rect 12388 22412 12392 22468
rect 12328 22408 12392 22412
rect 12328 22308 12392 22312
rect 12328 22252 12332 22308
rect 12332 22252 12388 22308
rect 12388 22252 12392 22308
rect 12328 22248 12392 22252
rect 12328 22148 12392 22152
rect 12328 22092 12332 22148
rect 12332 22092 12388 22148
rect 12388 22092 12392 22148
rect 12328 22088 12392 22092
rect 12328 21928 12392 21992
rect 12328 21828 12392 21832
rect 12328 21772 12332 21828
rect 12332 21772 12388 21828
rect 12388 21772 12392 21828
rect 12328 21768 12392 21772
rect 12328 21668 12392 21672
rect 12328 21612 12332 21668
rect 12332 21612 12388 21668
rect 12388 21612 12392 21668
rect 12328 21608 12392 21612
rect 12328 21508 12392 21512
rect 12328 21452 12332 21508
rect 12332 21452 12388 21508
rect 12388 21452 12392 21508
rect 12328 21448 12392 21452
rect 12328 21348 12392 21352
rect 12328 21292 12332 21348
rect 12332 21292 12388 21348
rect 12388 21292 12392 21348
rect 12328 21288 12392 21292
rect 12328 21188 12392 21192
rect 12328 21132 12332 21188
rect 12332 21132 12388 21188
rect 12388 21132 12392 21188
rect 12328 21128 12392 21132
rect 12328 21028 12392 21032
rect 12328 20972 12332 21028
rect 12332 20972 12388 21028
rect 12388 20972 12392 21028
rect 12328 20968 12392 20972
rect 12328 20868 12392 20872
rect 12328 20812 12332 20868
rect 12332 20812 12388 20868
rect 12388 20812 12392 20868
rect 12328 20808 12392 20812
rect 12328 20708 12392 20712
rect 12328 20652 12332 20708
rect 12332 20652 12388 20708
rect 12388 20652 12392 20708
rect 12328 20648 12392 20652
rect 12328 20488 12392 20552
rect 12328 20328 12392 20392
rect 12328 20168 12392 20232
rect 12328 20008 12392 20072
rect 12328 19908 12392 19912
rect 12328 19852 12332 19908
rect 12332 19852 12388 19908
rect 12388 19852 12392 19908
rect 12328 19848 12392 19852
rect 12328 19748 12392 19752
rect 12328 19692 12332 19748
rect 12332 19692 12388 19748
rect 12388 19692 12392 19748
rect 12328 19688 12392 19692
rect 12328 19588 12392 19592
rect 12328 19532 12332 19588
rect 12332 19532 12388 19588
rect 12388 19532 12392 19588
rect 12328 19528 12392 19532
rect 12328 19428 12392 19432
rect 12328 19372 12332 19428
rect 12332 19372 12388 19428
rect 12388 19372 12392 19428
rect 12328 19368 12392 19372
rect 12328 19268 12392 19272
rect 12328 19212 12332 19268
rect 12332 19212 12388 19268
rect 12388 19212 12392 19268
rect 12328 19208 12392 19212
rect 12328 19108 12392 19112
rect 12328 19052 12332 19108
rect 12332 19052 12388 19108
rect 12388 19052 12392 19108
rect 12328 19048 12392 19052
rect 12328 18948 12392 18952
rect 12328 18892 12332 18948
rect 12332 18892 12388 18948
rect 12388 18892 12392 18948
rect 12328 18888 12392 18892
rect 12328 18788 12392 18792
rect 12328 18732 12332 18788
rect 12332 18732 12388 18788
rect 12388 18732 12392 18788
rect 12328 18728 12392 18732
rect 12328 18568 12392 18632
rect 12328 18408 12392 18472
rect 12328 18248 12392 18312
rect 12328 18088 12392 18152
rect 12328 17988 12392 17992
rect 12328 17932 12332 17988
rect 12332 17932 12388 17988
rect 12388 17932 12392 17988
rect 12328 17928 12392 17932
rect 12328 17828 12392 17832
rect 12328 17772 12332 17828
rect 12332 17772 12388 17828
rect 12388 17772 12392 17828
rect 12328 17768 12392 17772
rect 12328 17668 12392 17672
rect 12328 17612 12332 17668
rect 12332 17612 12388 17668
rect 12388 17612 12392 17668
rect 12328 17608 12392 17612
rect 12328 17508 12392 17512
rect 12328 17452 12332 17508
rect 12332 17452 12388 17508
rect 12388 17452 12392 17508
rect 12328 17448 12392 17452
rect 12328 17348 12392 17352
rect 12328 17292 12332 17348
rect 12332 17292 12388 17348
rect 12388 17292 12392 17348
rect 12328 17288 12392 17292
rect 12328 17188 12392 17192
rect 12328 17132 12332 17188
rect 12332 17132 12388 17188
rect 12388 17132 12392 17188
rect 12328 17128 12392 17132
rect 12328 17028 12392 17032
rect 12328 16972 12332 17028
rect 12332 16972 12388 17028
rect 12388 16972 12392 17028
rect 12328 16968 12392 16972
rect 12328 16868 12392 16872
rect 12328 16812 12332 16868
rect 12332 16812 12388 16868
rect 12388 16812 12392 16868
rect 12328 16808 12392 16812
rect 12328 16648 12392 16712
rect 12328 16548 12392 16552
rect 12328 16492 12332 16548
rect 12332 16492 12388 16548
rect 12388 16492 12392 16548
rect 12328 16488 12392 16492
rect 12328 16388 12392 16392
rect 12328 16332 12332 16388
rect 12332 16332 12388 16388
rect 12388 16332 12392 16388
rect 12328 16328 12392 16332
rect 12328 16228 12392 16232
rect 12328 16172 12332 16228
rect 12332 16172 12388 16228
rect 12388 16172 12392 16228
rect 12328 16168 12392 16172
rect 12328 16068 12392 16072
rect 12328 16012 12332 16068
rect 12332 16012 12388 16068
rect 12388 16012 12392 16068
rect 12328 16008 12392 16012
rect 12328 15908 12392 15912
rect 12328 15852 12332 15908
rect 12332 15852 12388 15908
rect 12388 15852 12392 15908
rect 12328 15848 12392 15852
rect 12328 15748 12392 15752
rect 12328 15692 12332 15748
rect 12332 15692 12388 15748
rect 12388 15692 12392 15748
rect 12328 15688 12392 15692
rect 12328 15588 12392 15592
rect 12328 15532 12332 15588
rect 12332 15532 12388 15588
rect 12388 15532 12392 15588
rect 12328 15528 12392 15532
rect 12328 15428 12392 15432
rect 12328 15372 12332 15428
rect 12332 15372 12388 15428
rect 12388 15372 12392 15428
rect 12328 15368 12392 15372
rect 12328 15268 12392 15272
rect 12328 15212 12332 15268
rect 12332 15212 12388 15268
rect 12388 15212 12392 15268
rect 12328 15208 12392 15212
rect 12328 15108 12392 15112
rect 12328 15052 12332 15108
rect 12332 15052 12388 15108
rect 12388 15052 12392 15108
rect 12328 15048 12392 15052
rect 12328 14948 12392 14952
rect 12328 14892 12332 14948
rect 12332 14892 12388 14948
rect 12388 14892 12392 14948
rect 12328 14888 12392 14892
rect 12328 14788 12392 14792
rect 12328 14732 12332 14788
rect 12332 14732 12388 14788
rect 12388 14732 12392 14788
rect 12328 14728 12392 14732
rect 12328 14628 12392 14632
rect 12328 14572 12332 14628
rect 12332 14572 12388 14628
rect 12388 14572 12392 14628
rect 12328 14568 12392 14572
rect 12328 14468 12392 14472
rect 12328 14412 12332 14468
rect 12332 14412 12388 14468
rect 12388 14412 12392 14468
rect 12328 14408 12392 14412
rect 12328 14308 12392 14312
rect 12328 14252 12332 14308
rect 12332 14252 12388 14308
rect 12388 14252 12392 14308
rect 12328 14248 12392 14252
rect 12328 14148 12392 14152
rect 12328 14092 12332 14148
rect 12332 14092 12388 14148
rect 12388 14092 12392 14148
rect 12328 14088 12392 14092
rect 12328 13988 12392 13992
rect 12328 13932 12332 13988
rect 12332 13932 12388 13988
rect 12388 13932 12392 13988
rect 12328 13928 12392 13932
rect 12328 13768 12392 13832
rect 12328 13668 12392 13672
rect 12328 13612 12332 13668
rect 12332 13612 12388 13668
rect 12388 13612 12392 13668
rect 12328 13608 12392 13612
rect 12328 13508 12392 13512
rect 12328 13452 12332 13508
rect 12332 13452 12388 13508
rect 12388 13452 12392 13508
rect 12328 13448 12392 13452
rect 12328 13348 12392 13352
rect 12328 13292 12332 13348
rect 12332 13292 12388 13348
rect 12388 13292 12392 13348
rect 12328 13288 12392 13292
rect 12328 13188 12392 13192
rect 12328 13132 12332 13188
rect 12332 13132 12388 13188
rect 12388 13132 12392 13188
rect 12328 13128 12392 13132
rect 12328 13028 12392 13032
rect 12328 12972 12332 13028
rect 12332 12972 12388 13028
rect 12388 12972 12392 13028
rect 12328 12968 12392 12972
rect 12328 12868 12392 12872
rect 12328 12812 12332 12868
rect 12332 12812 12388 12868
rect 12388 12812 12392 12868
rect 12328 12808 12392 12812
rect 12328 12708 12392 12712
rect 12328 12652 12332 12708
rect 12332 12652 12388 12708
rect 12388 12652 12392 12708
rect 12328 12648 12392 12652
rect 12328 12548 12392 12552
rect 12328 12492 12332 12548
rect 12332 12492 12388 12548
rect 12388 12492 12392 12548
rect 12328 12488 12392 12492
rect 12328 12328 12392 12392
rect 12328 12168 12392 12232
rect 12328 12008 12392 12072
rect 12328 11848 12392 11912
rect 12328 11748 12392 11752
rect 12328 11692 12332 11748
rect 12332 11692 12388 11748
rect 12388 11692 12392 11748
rect 12328 11688 12392 11692
rect 12328 11588 12392 11592
rect 12328 11532 12332 11588
rect 12332 11532 12388 11588
rect 12388 11532 12392 11588
rect 12328 11528 12392 11532
rect 12328 11428 12392 11432
rect 12328 11372 12332 11428
rect 12332 11372 12388 11428
rect 12388 11372 12392 11428
rect 12328 11368 12392 11372
rect 12328 11268 12392 11272
rect 12328 11212 12332 11268
rect 12332 11212 12388 11268
rect 12388 11212 12392 11268
rect 12328 11208 12392 11212
rect 12328 11108 12392 11112
rect 12328 11052 12332 11108
rect 12332 11052 12388 11108
rect 12388 11052 12392 11108
rect 12328 11048 12392 11052
rect 12328 10948 12392 10952
rect 12328 10892 12332 10948
rect 12332 10892 12388 10948
rect 12388 10892 12392 10948
rect 12328 10888 12392 10892
rect 12328 10788 12392 10792
rect 12328 10732 12332 10788
rect 12332 10732 12388 10788
rect 12388 10732 12392 10788
rect 12328 10728 12392 10732
rect 12328 10628 12392 10632
rect 12328 10572 12332 10628
rect 12332 10572 12388 10628
rect 12388 10572 12392 10628
rect 12328 10568 12392 10572
rect 12328 10468 12392 10472
rect 12328 10412 12332 10468
rect 12332 10412 12388 10468
rect 12388 10412 12392 10468
rect 12328 10408 12392 10412
rect 12328 10308 12392 10312
rect 12328 10252 12332 10308
rect 12332 10252 12388 10308
rect 12388 10252 12392 10308
rect 12328 10248 12392 10252
rect 12328 10148 12392 10152
rect 12328 10092 12332 10148
rect 12332 10092 12388 10148
rect 12388 10092 12392 10148
rect 12328 10088 12392 10092
rect 12328 9988 12392 9992
rect 12328 9932 12332 9988
rect 12332 9932 12388 9988
rect 12388 9932 12392 9988
rect 12328 9928 12392 9932
rect 12328 9828 12392 9832
rect 12328 9772 12332 9828
rect 12332 9772 12388 9828
rect 12388 9772 12392 9828
rect 12328 9768 12392 9772
rect 12328 9608 12392 9672
rect 12328 9508 12392 9512
rect 12328 9452 12332 9508
rect 12332 9452 12388 9508
rect 12388 9452 12392 9508
rect 12328 9448 12392 9452
rect 12328 9348 12392 9352
rect 12328 9292 12332 9348
rect 12332 9292 12388 9348
rect 12388 9292 12392 9348
rect 12328 9288 12392 9292
rect 12328 9128 12392 9192
rect 12328 9028 12392 9032
rect 12328 8972 12332 9028
rect 12332 8972 12388 9028
rect 12388 8972 12392 9028
rect 12328 8968 12392 8972
rect 12328 8868 12392 8872
rect 12328 8812 12332 8868
rect 12332 8812 12388 8868
rect 12388 8812 12392 8868
rect 12328 8808 12392 8812
rect 12328 8708 12392 8712
rect 12328 8652 12332 8708
rect 12332 8652 12388 8708
rect 12388 8652 12392 8708
rect 12328 8648 12392 8652
rect 12328 8548 12392 8552
rect 12328 8492 12332 8548
rect 12332 8492 12388 8548
rect 12388 8492 12392 8548
rect 12328 8488 12392 8492
rect 12328 8388 12392 8392
rect 12328 8332 12332 8388
rect 12332 8332 12388 8388
rect 12388 8332 12392 8388
rect 12328 8328 12392 8332
rect 12328 8228 12392 8232
rect 12328 8172 12332 8228
rect 12332 8172 12388 8228
rect 12388 8172 12392 8228
rect 12328 8168 12392 8172
rect 12328 8068 12392 8072
rect 12328 8012 12332 8068
rect 12332 8012 12388 8068
rect 12388 8012 12392 8068
rect 12328 8008 12392 8012
rect 12328 7908 12392 7912
rect 12328 7852 12332 7908
rect 12332 7852 12388 7908
rect 12388 7852 12392 7908
rect 12328 7848 12392 7852
rect 12328 7748 12392 7752
rect 12328 7692 12332 7748
rect 12332 7692 12388 7748
rect 12388 7692 12392 7748
rect 12328 7688 12392 7692
rect 12328 7528 12392 7592
rect 12328 7428 12392 7432
rect 12328 7372 12332 7428
rect 12332 7372 12388 7428
rect 12388 7372 12392 7428
rect 12328 7368 12392 7372
rect 12328 7268 12392 7272
rect 12328 7212 12332 7268
rect 12332 7212 12388 7268
rect 12388 7212 12392 7268
rect 12328 7208 12392 7212
rect 12328 7048 12392 7112
rect 12328 6948 12392 6952
rect 12328 6892 12332 6948
rect 12332 6892 12388 6948
rect 12388 6892 12392 6948
rect 12328 6888 12392 6892
rect 12328 6788 12392 6792
rect 12328 6732 12332 6788
rect 12332 6732 12388 6788
rect 12388 6732 12392 6788
rect 12328 6728 12392 6732
rect 12328 6568 12392 6632
rect 12328 6468 12392 6472
rect 12328 6412 12332 6468
rect 12332 6412 12388 6468
rect 12388 6412 12392 6468
rect 12328 6408 12392 6412
rect 12328 6308 12392 6312
rect 12328 6252 12332 6308
rect 12332 6252 12388 6308
rect 12388 6252 12392 6308
rect 12328 6248 12392 6252
rect 12328 6148 12392 6152
rect 12328 6092 12332 6148
rect 12332 6092 12388 6148
rect 12388 6092 12392 6148
rect 12328 6088 12392 6092
rect 12328 5988 12392 5992
rect 12328 5932 12332 5988
rect 12332 5932 12388 5988
rect 12388 5932 12392 5988
rect 12328 5928 12392 5932
rect 12328 5828 12392 5832
rect 12328 5772 12332 5828
rect 12332 5772 12388 5828
rect 12388 5772 12392 5828
rect 12328 5768 12392 5772
rect 12328 5668 12392 5672
rect 12328 5612 12332 5668
rect 12332 5612 12388 5668
rect 12388 5612 12392 5668
rect 12328 5608 12392 5612
rect 12328 5508 12392 5512
rect 12328 5452 12332 5508
rect 12332 5452 12388 5508
rect 12388 5452 12392 5508
rect 12328 5448 12392 5452
rect 12328 5348 12392 5352
rect 12328 5292 12332 5348
rect 12332 5292 12388 5348
rect 12388 5292 12392 5348
rect 12328 5288 12392 5292
rect 12328 5188 12392 5192
rect 12328 5132 12332 5188
rect 12332 5132 12388 5188
rect 12388 5132 12392 5188
rect 12328 5128 12392 5132
rect 12328 5028 12392 5032
rect 12328 4972 12332 5028
rect 12332 4972 12388 5028
rect 12388 4972 12392 5028
rect 12328 4968 12392 4972
rect 12328 4868 12392 4872
rect 12328 4812 12332 4868
rect 12332 4812 12388 4868
rect 12388 4812 12392 4868
rect 12328 4808 12392 4812
rect 12328 4708 12392 4712
rect 12328 4652 12332 4708
rect 12332 4652 12388 4708
rect 12388 4652 12392 4708
rect 12328 4648 12392 4652
rect 12328 4548 12392 4552
rect 12328 4492 12332 4548
rect 12332 4492 12388 4548
rect 12388 4492 12392 4548
rect 12328 4488 12392 4492
rect 12328 4388 12392 4392
rect 12328 4332 12332 4388
rect 12332 4332 12388 4388
rect 12388 4332 12392 4388
rect 12328 4328 12392 4332
rect 12328 4228 12392 4232
rect 12328 4172 12332 4228
rect 12332 4172 12388 4228
rect 12388 4172 12392 4228
rect 12328 4168 12392 4172
rect 12328 4068 12392 4072
rect 12328 4012 12332 4068
rect 12332 4012 12388 4068
rect 12388 4012 12392 4068
rect 12328 4008 12392 4012
rect 12328 3908 12392 3912
rect 12328 3852 12332 3908
rect 12332 3852 12388 3908
rect 12388 3852 12392 3908
rect 12328 3848 12392 3852
rect 12328 3688 12392 3752
rect 12328 3528 12392 3592
rect 12328 3428 12392 3432
rect 12328 3372 12332 3428
rect 12332 3372 12388 3428
rect 12388 3372 12392 3428
rect 12328 3368 12392 3372
rect 12328 3268 12392 3272
rect 12328 3212 12332 3268
rect 12332 3212 12388 3268
rect 12388 3212 12392 3268
rect 12328 3208 12392 3212
rect 12328 3108 12392 3112
rect 12328 3052 12332 3108
rect 12332 3052 12388 3108
rect 12388 3052 12392 3108
rect 12328 3048 12392 3052
rect 12328 2948 12392 2952
rect 12328 2892 12332 2948
rect 12332 2892 12388 2948
rect 12388 2892 12392 2948
rect 12328 2888 12392 2892
rect 12328 2788 12392 2792
rect 12328 2732 12332 2788
rect 12332 2732 12388 2788
rect 12388 2732 12392 2788
rect 12328 2728 12392 2732
rect 12328 2628 12392 2632
rect 12328 2572 12332 2628
rect 12332 2572 12388 2628
rect 12388 2572 12392 2628
rect 12328 2568 12392 2572
rect 12328 2468 12392 2472
rect 12328 2412 12332 2468
rect 12332 2412 12388 2468
rect 12388 2412 12392 2468
rect 12328 2408 12392 2412
rect 12328 2308 12392 2312
rect 12328 2252 12332 2308
rect 12332 2252 12388 2308
rect 12388 2252 12392 2308
rect 12328 2248 12392 2252
rect 12328 2148 12392 2152
rect 12328 2092 12332 2148
rect 12332 2092 12388 2148
rect 12388 2092 12392 2148
rect 12328 2088 12392 2092
rect 12328 1988 12392 1992
rect 12328 1932 12332 1988
rect 12332 1932 12388 1988
rect 12388 1932 12392 1988
rect 12328 1928 12392 1932
rect 12328 1768 12392 1832
rect 12328 1668 12392 1672
rect 12328 1612 12332 1668
rect 12332 1612 12388 1668
rect 12388 1612 12392 1668
rect 12328 1608 12392 1612
rect 12328 1508 12392 1512
rect 12328 1452 12332 1508
rect 12332 1452 12388 1508
rect 12388 1452 12392 1508
rect 12328 1448 12392 1452
rect 12328 1348 12392 1352
rect 12328 1292 12332 1348
rect 12332 1292 12388 1348
rect 12388 1292 12392 1348
rect 12328 1288 12392 1292
rect 12328 1188 12392 1192
rect 12328 1132 12332 1188
rect 12332 1132 12388 1188
rect 12388 1132 12392 1188
rect 12328 1128 12392 1132
rect 12328 1028 12392 1032
rect 12328 972 12332 1028
rect 12332 972 12388 1028
rect 12388 972 12392 1028
rect 12328 968 12392 972
rect 12328 808 12392 872
rect 12328 648 12392 712
rect 12328 548 12392 552
rect 12328 492 12332 548
rect 12332 492 12388 548
rect 12388 492 12392 548
rect 12328 488 12392 492
rect 12328 388 12392 392
rect 12328 332 12332 388
rect 12332 332 12388 388
rect 12388 332 12392 388
rect 12328 328 12392 332
rect 12328 228 12392 232
rect 12328 172 12332 228
rect 12332 172 12388 228
rect 12388 172 12392 228
rect 12328 168 12392 172
rect 12328 68 12392 72
rect 12328 12 12332 68
rect 12332 12 12388 68
rect 12388 12 12392 68
rect 12328 8 12392 12
rect 12008 -1112 12072 -1048
rect 12008 -1192 12072 -1128
rect 12008 -1272 12072 -1208
rect 12008 -1352 12072 -1288
rect 12008 -1432 12072 -1368
rect 12328 -1112 12392 -1048
rect 12328 -1192 12392 -1128
rect 12328 -1272 12392 -1208
rect 12328 -1352 12392 -1288
rect 12328 -1432 12392 -1368
rect 9288 -2072 9352 -2008
rect 20568 -2072 20632 -2008
rect 408 -2232 472 -2168
rect 2488 -2232 2552 -2168
rect 2648 -2232 2712 -2168
rect 4728 -2232 4792 -2168
rect 4888 -2232 4952 -2168
rect 6968 -2232 7032 -2168
rect 7128 -2232 7192 -2168
rect 9208 -2232 9272 -2168
rect 9368 -2232 9432 -2168
rect 11448 -2232 11512 -2168
rect 11608 -2232 11672 -2168
rect 13688 -2232 13752 -2168
rect 13848 -2232 13912 -2168
rect 15928 -2232 15992 -2168
rect 16088 -2232 16152 -2168
rect 18168 -2232 18232 -2168
rect 18328 -2232 18392 -2168
rect 20408 -2232 20472 -2168
rect 248 -4632 312 -4568
rect 20568 -4632 20632 -4568
<< mimcap >>
rect 480 -2488 2480 -2400
rect 480 -4312 568 -2488
rect 2392 -4312 2480 -2488
rect 480 -4400 2480 -4312
rect 2720 -2488 4720 -2400
rect 2720 -4312 2808 -2488
rect 4632 -4312 4720 -2488
rect 2720 -4400 4720 -4312
rect 4960 -2488 6960 -2400
rect 4960 -4312 5048 -2488
rect 6872 -4312 6960 -2488
rect 4960 -4400 6960 -4312
rect 7200 -2488 9200 -2400
rect 7200 -4312 7288 -2488
rect 9112 -4312 9200 -2488
rect 7200 -4400 9200 -4312
rect 9440 -2488 11440 -2400
rect 9440 -4312 9528 -2488
rect 11352 -4312 11440 -2488
rect 9440 -4400 11440 -4312
rect 11680 -2488 13680 -2400
rect 11680 -4312 11768 -2488
rect 13592 -4312 13680 -2488
rect 11680 -4400 13680 -4312
rect 13920 -2488 15920 -2400
rect 13920 -4312 14008 -2488
rect 15832 -4312 15920 -2488
rect 13920 -4400 15920 -4312
rect 16160 -2488 18160 -2400
rect 16160 -4312 16248 -2488
rect 18072 -4312 18160 -2488
rect 16160 -4400 18160 -4312
rect 18400 -2488 20400 -2400
rect 18400 -4312 18488 -2488
rect 20312 -4312 20400 -2488
rect 18400 -4400 20400 -4312
<< mimcapcontact >>
rect 568 -4312 2392 -2488
rect 2808 -4312 4632 -2488
rect 5048 -4312 6872 -2488
rect 7288 -4312 9112 -2488
rect 9528 -4312 11352 -2488
rect 11768 -4312 13592 -2488
rect 14008 -4312 15832 -2488
rect 16248 -4312 18072 -2488
rect 18488 -4312 20312 -2488
<< metal4 >>
rect 8480 31432 8880 31440
rect 8480 31368 8488 31432
rect 8552 31368 8808 31432
rect 8872 31368 8880 31432
rect 8480 31360 8880 31368
rect 8960 31432 9360 31440
rect 8960 31368 8968 31432
rect 9032 31368 9288 31432
rect 9352 31368 9360 31432
rect 8960 31360 9360 31368
rect 9440 31432 11440 31440
rect 9440 31368 9448 31432
rect 9512 31368 9768 31432
rect 9832 31368 10088 31432
rect 10152 31368 10408 31432
rect 10472 31368 10728 31432
rect 10792 31368 11048 31432
rect 11112 31368 11368 31432
rect 11432 31368 11440 31432
rect 9440 31360 11440 31368
rect 11520 31432 11920 31440
rect 11520 31368 11528 31432
rect 11592 31368 11848 31432
rect 11912 31368 11920 31432
rect 11520 31360 11920 31368
rect 12000 31432 12400 31440
rect 12000 31368 12008 31432
rect 12072 31368 12328 31432
rect 12392 31368 12400 31432
rect 12000 31360 12400 31368
rect 8480 31272 8880 31280
rect 8480 31208 8488 31272
rect 8552 31208 8808 31272
rect 8872 31208 8880 31272
rect 8480 31200 8880 31208
rect 8960 31272 9360 31280
rect 8960 31208 8968 31272
rect 9032 31208 9288 31272
rect 9352 31208 9360 31272
rect 8960 31200 9360 31208
rect 9440 31272 11440 31280
rect 9440 31208 9448 31272
rect 9512 31208 9768 31272
rect 9832 31208 10088 31272
rect 10152 31208 10408 31272
rect 10472 31208 10728 31272
rect 10792 31208 11048 31272
rect 11112 31208 11368 31272
rect 11432 31208 11440 31272
rect 9440 31200 11440 31208
rect 11520 31272 11920 31280
rect 11520 31208 11528 31272
rect 11592 31208 11848 31272
rect 11912 31208 11920 31272
rect 11520 31200 11920 31208
rect 12000 31272 12400 31280
rect 12000 31208 12008 31272
rect 12072 31208 12328 31272
rect 12392 31208 12400 31272
rect 12000 31200 12400 31208
rect 8480 31112 8880 31120
rect 8480 31048 8488 31112
rect 8552 31048 8808 31112
rect 8872 31048 8880 31112
rect 8480 31040 8880 31048
rect 8960 31112 9360 31120
rect 8960 31048 8968 31112
rect 9032 31048 9288 31112
rect 9352 31048 9360 31112
rect 8960 31040 9360 31048
rect 9440 31112 11440 31120
rect 9440 31048 9448 31112
rect 9512 31048 9768 31112
rect 9832 31048 10088 31112
rect 10152 31048 10408 31112
rect 10472 31048 10728 31112
rect 10792 31048 11048 31112
rect 11112 31048 11368 31112
rect 11432 31048 11440 31112
rect 9440 31040 11440 31048
rect 11520 31112 11920 31120
rect 11520 31048 11528 31112
rect 11592 31048 11848 31112
rect 11912 31048 11920 31112
rect 11520 31040 11920 31048
rect 12000 31112 12400 31120
rect 12000 31048 12008 31112
rect 12072 31048 12328 31112
rect 12392 31048 12400 31112
rect 12000 31040 12400 31048
rect 8480 30952 8880 30960
rect 8480 30888 8488 30952
rect 8552 30888 8808 30952
rect 8872 30888 8880 30952
rect 8480 30880 8880 30888
rect 8960 30952 9360 30960
rect 8960 30888 8968 30952
rect 9032 30888 9288 30952
rect 9352 30888 9360 30952
rect 8960 30880 9360 30888
rect 9440 30952 11440 30960
rect 9440 30888 9448 30952
rect 9512 30888 9768 30952
rect 9832 30888 10088 30952
rect 10152 30888 10408 30952
rect 10472 30888 10728 30952
rect 10792 30888 11048 30952
rect 11112 30888 11368 30952
rect 11432 30888 11440 30952
rect 9440 30880 11440 30888
rect 11520 30952 11920 30960
rect 11520 30888 11528 30952
rect 11592 30888 11848 30952
rect 11912 30888 11920 30952
rect 11520 30880 11920 30888
rect 12000 30952 12400 30960
rect 12000 30888 12008 30952
rect 12072 30888 12328 30952
rect 12392 30888 12400 30952
rect 12000 30880 12400 30888
rect 8480 30792 8880 30800
rect 8480 30728 8488 30792
rect 8552 30728 8808 30792
rect 8872 30728 8880 30792
rect 8480 30720 8880 30728
rect 8960 30792 9360 30800
rect 8960 30728 8968 30792
rect 9032 30728 9288 30792
rect 9352 30728 9360 30792
rect 8960 30720 9360 30728
rect 9440 30792 11440 30800
rect 9440 30728 9448 30792
rect 9512 30728 9768 30792
rect 9832 30728 10088 30792
rect 10152 30728 10408 30792
rect 10472 30728 10728 30792
rect 10792 30728 11048 30792
rect 11112 30728 11368 30792
rect 11432 30728 11440 30792
rect 9440 30720 11440 30728
rect 11520 30792 11920 30800
rect 11520 30728 11528 30792
rect 11592 30728 11848 30792
rect 11912 30728 11920 30792
rect 11520 30720 11920 30728
rect 12000 30792 12400 30800
rect 12000 30728 12008 30792
rect 12072 30728 12328 30792
rect 12392 30728 12400 30792
rect 12000 30720 12400 30728
rect 8480 30632 8880 30640
rect 8480 30568 8488 30632
rect 8552 30568 8808 30632
rect 8872 30568 8880 30632
rect 8480 30560 8880 30568
rect 8960 30632 9360 30640
rect 8960 30568 8968 30632
rect 9032 30568 9288 30632
rect 9352 30568 9360 30632
rect 8960 30560 9360 30568
rect 9440 30632 11440 30640
rect 9440 30568 9448 30632
rect 9512 30568 9768 30632
rect 9832 30568 10088 30632
rect 10152 30568 10408 30632
rect 10472 30568 10728 30632
rect 10792 30568 11048 30632
rect 11112 30568 11368 30632
rect 11432 30568 11440 30632
rect 9440 30560 11440 30568
rect 11520 30632 11920 30640
rect 11520 30568 11528 30632
rect 11592 30568 11848 30632
rect 11912 30568 11920 30632
rect 11520 30560 11920 30568
rect 12000 30632 12400 30640
rect 12000 30568 12008 30632
rect 12072 30568 12328 30632
rect 12392 30568 12400 30632
rect 12000 30560 12400 30568
rect 8480 30472 8880 30480
rect 8480 30408 8488 30472
rect 8552 30408 8808 30472
rect 8872 30408 8880 30472
rect 8480 30400 8880 30408
rect 8960 30472 9360 30480
rect 8960 30408 8968 30472
rect 9032 30408 9288 30472
rect 9352 30408 9360 30472
rect 8960 30400 9360 30408
rect 9440 30472 11440 30480
rect 9440 30408 9448 30472
rect 9512 30408 9768 30472
rect 9832 30408 10088 30472
rect 10152 30408 10408 30472
rect 10472 30408 10728 30472
rect 10792 30408 11048 30472
rect 11112 30408 11368 30472
rect 11432 30408 11440 30472
rect 9440 30400 11440 30408
rect 11520 30472 11920 30480
rect 11520 30408 11528 30472
rect 11592 30408 11848 30472
rect 11912 30408 11920 30472
rect 11520 30400 11920 30408
rect 12000 30472 12400 30480
rect 12000 30408 12008 30472
rect 12072 30408 12328 30472
rect 12392 30408 12400 30472
rect 12000 30400 12400 30408
rect 8480 30312 8880 30320
rect 8480 30248 8488 30312
rect 8552 30248 8808 30312
rect 8872 30248 8880 30312
rect 8480 30240 8880 30248
rect 8960 30312 9360 30320
rect 8960 30248 8968 30312
rect 9032 30248 9288 30312
rect 9352 30248 9360 30312
rect 8960 30240 9360 30248
rect 9440 30312 11440 30320
rect 9440 30248 9448 30312
rect 9512 30248 9768 30312
rect 9832 30248 10088 30312
rect 10152 30248 10408 30312
rect 10472 30248 10728 30312
rect 10792 30248 11048 30312
rect 11112 30248 11368 30312
rect 11432 30248 11440 30312
rect 9440 30240 11440 30248
rect 11520 30312 11920 30320
rect 11520 30248 11528 30312
rect 11592 30248 11848 30312
rect 11912 30248 11920 30312
rect 11520 30240 11920 30248
rect 12000 30312 12400 30320
rect 12000 30248 12008 30312
rect 12072 30248 12328 30312
rect 12392 30248 12400 30312
rect 12000 30240 12400 30248
rect 8480 30152 8880 30160
rect 8480 30088 8488 30152
rect 8552 30088 8808 30152
rect 8872 30088 8880 30152
rect 8480 30080 8880 30088
rect 8960 30152 9360 30160
rect 8960 30088 8968 30152
rect 9032 30088 9288 30152
rect 9352 30088 9360 30152
rect 8960 30080 9360 30088
rect 9440 30152 11440 30160
rect 9440 30088 9448 30152
rect 9512 30088 9768 30152
rect 9832 30088 10088 30152
rect 10152 30088 10408 30152
rect 10472 30088 10728 30152
rect 10792 30088 11048 30152
rect 11112 30088 11368 30152
rect 11432 30088 11440 30152
rect 9440 30080 11440 30088
rect 11520 30152 11920 30160
rect 11520 30088 11528 30152
rect 11592 30088 11848 30152
rect 11912 30088 11920 30152
rect 11520 30080 11920 30088
rect 12000 30152 12400 30160
rect 12000 30088 12008 30152
rect 12072 30088 12328 30152
rect 12392 30088 12400 30152
rect 12000 30080 12400 30088
rect 8480 29992 8880 30000
rect 8480 29928 8488 29992
rect 8552 29928 8808 29992
rect 8872 29928 8880 29992
rect 8480 29920 8880 29928
rect 8960 29992 9360 30000
rect 8960 29928 8968 29992
rect 9032 29928 9288 29992
rect 9352 29928 9360 29992
rect 8960 29920 9360 29928
rect 9440 29992 11440 30000
rect 9440 29928 9448 29992
rect 9512 29928 9768 29992
rect 9832 29928 10088 29992
rect 10152 29928 10408 29992
rect 10472 29928 10728 29992
rect 10792 29928 11048 29992
rect 11112 29928 11368 29992
rect 11432 29928 11440 29992
rect 9440 29920 11440 29928
rect 11520 29992 11920 30000
rect 11520 29928 11528 29992
rect 11592 29928 11848 29992
rect 11912 29928 11920 29992
rect 11520 29920 11920 29928
rect 12000 29992 12400 30000
rect 12000 29928 12008 29992
rect 12072 29928 12328 29992
rect 12392 29928 12400 29992
rect 12000 29920 12400 29928
rect 8480 29832 8880 29840
rect 8480 29768 8488 29832
rect 8552 29768 8808 29832
rect 8872 29768 8880 29832
rect 8480 29760 8880 29768
rect 8960 29832 9360 29840
rect 8960 29768 8968 29832
rect 9032 29768 9288 29832
rect 9352 29768 9360 29832
rect 8960 29760 9360 29768
rect 9440 29832 11440 29840
rect 9440 29768 9448 29832
rect 9512 29768 9768 29832
rect 9832 29768 10088 29832
rect 10152 29768 10408 29832
rect 10472 29768 10728 29832
rect 10792 29768 11048 29832
rect 11112 29768 11368 29832
rect 11432 29768 11440 29832
rect 9440 29760 11440 29768
rect 11520 29832 11920 29840
rect 11520 29768 11528 29832
rect 11592 29768 11848 29832
rect 11912 29768 11920 29832
rect 11520 29760 11920 29768
rect 12000 29832 12400 29840
rect 12000 29768 12008 29832
rect 12072 29768 12328 29832
rect 12392 29768 12400 29832
rect 12000 29760 12400 29768
rect 8480 29672 8880 29680
rect 8480 29608 8488 29672
rect 8552 29608 8808 29672
rect 8872 29608 8880 29672
rect 8480 29600 8880 29608
rect 8960 29672 9360 29680
rect 8960 29608 8968 29672
rect 9032 29608 9288 29672
rect 9352 29608 9360 29672
rect 8960 29600 9360 29608
rect 9440 29672 11440 29680
rect 9440 29608 9448 29672
rect 9512 29608 9768 29672
rect 9832 29608 10088 29672
rect 10152 29608 10408 29672
rect 10472 29608 10728 29672
rect 10792 29608 11048 29672
rect 11112 29608 11368 29672
rect 11432 29608 11440 29672
rect 9440 29600 11440 29608
rect 11520 29672 11920 29680
rect 11520 29608 11528 29672
rect 11592 29608 11848 29672
rect 11912 29608 11920 29672
rect 11520 29600 11920 29608
rect 12000 29672 12400 29680
rect 12000 29608 12008 29672
rect 12072 29608 12328 29672
rect 12392 29608 12400 29672
rect 12000 29600 12400 29608
rect 8480 29512 8880 29520
rect 8480 29448 8488 29512
rect 8552 29448 8808 29512
rect 8872 29448 8880 29512
rect 8480 29440 8880 29448
rect 8960 29512 9360 29520
rect 8960 29448 8968 29512
rect 9032 29448 9288 29512
rect 9352 29448 9360 29512
rect 8960 29440 9360 29448
rect 9440 29512 11440 29520
rect 9440 29448 9448 29512
rect 9512 29448 9768 29512
rect 9832 29448 10088 29512
rect 10152 29448 10408 29512
rect 10472 29448 10728 29512
rect 10792 29448 11048 29512
rect 11112 29448 11368 29512
rect 11432 29448 11440 29512
rect 9440 29440 11440 29448
rect 11520 29512 11920 29520
rect 11520 29448 11528 29512
rect 11592 29448 11848 29512
rect 11912 29448 11920 29512
rect 11520 29440 11920 29448
rect 12000 29512 12400 29520
rect 12000 29448 12008 29512
rect 12072 29448 12328 29512
rect 12392 29448 12400 29512
rect 12000 29440 12400 29448
rect 8480 29352 8880 29360
rect 8480 29288 8488 29352
rect 8552 29288 8808 29352
rect 8872 29288 8880 29352
rect 8480 29280 8880 29288
rect 8960 29352 9360 29360
rect 8960 29288 8968 29352
rect 9032 29288 9288 29352
rect 9352 29288 9360 29352
rect 8960 29280 9360 29288
rect 9440 29352 11440 29360
rect 9440 29288 9448 29352
rect 9512 29288 9768 29352
rect 9832 29288 10088 29352
rect 10152 29288 10408 29352
rect 10472 29288 10728 29352
rect 10792 29288 11048 29352
rect 11112 29288 11368 29352
rect 11432 29288 11440 29352
rect 9440 29280 11440 29288
rect 11520 29352 11920 29360
rect 11520 29288 11528 29352
rect 11592 29288 11848 29352
rect 11912 29288 11920 29352
rect 11520 29280 11920 29288
rect 12000 29352 12400 29360
rect 12000 29288 12008 29352
rect 12072 29288 12328 29352
rect 12392 29288 12400 29352
rect 12000 29280 12400 29288
rect 8480 29192 8880 29200
rect 8480 29128 8488 29192
rect 8552 29128 8808 29192
rect 8872 29128 8880 29192
rect 8480 29120 8880 29128
rect 8960 29192 9360 29200
rect 8960 29128 8968 29192
rect 9032 29128 9288 29192
rect 9352 29128 9360 29192
rect 8960 29120 9360 29128
rect 9440 29192 11440 29200
rect 9440 29128 9448 29192
rect 9512 29128 9768 29192
rect 9832 29128 10088 29192
rect 10152 29128 10408 29192
rect 10472 29128 10728 29192
rect 10792 29128 11048 29192
rect 11112 29128 11368 29192
rect 11432 29128 11440 29192
rect 9440 29120 11440 29128
rect 11520 29192 11920 29200
rect 11520 29128 11528 29192
rect 11592 29128 11848 29192
rect 11912 29128 11920 29192
rect 11520 29120 11920 29128
rect 12000 29192 12400 29200
rect 12000 29128 12008 29192
rect 12072 29128 12328 29192
rect 12392 29128 12400 29192
rect 12000 29120 12400 29128
rect 8480 29032 8880 29040
rect 8480 28968 8488 29032
rect 8552 28968 8808 29032
rect 8872 28968 8880 29032
rect 8480 28960 8880 28968
rect 8960 29032 9360 29040
rect 8960 28968 8968 29032
rect 9032 28968 9288 29032
rect 9352 28968 9360 29032
rect 8960 28960 9360 28968
rect 9440 29032 11440 29040
rect 9440 28968 9448 29032
rect 9512 28968 9768 29032
rect 9832 28968 10088 29032
rect 10152 28968 10408 29032
rect 10472 28968 10728 29032
rect 10792 28968 11048 29032
rect 11112 28968 11368 29032
rect 11432 28968 11440 29032
rect 9440 28960 11440 28968
rect 11520 29032 11920 29040
rect 11520 28968 11528 29032
rect 11592 28968 11848 29032
rect 11912 28968 11920 29032
rect 11520 28960 11920 28968
rect 12000 29032 12400 29040
rect 12000 28968 12008 29032
rect 12072 28968 12328 29032
rect 12392 28968 12400 29032
rect 12000 28960 12400 28968
rect 8480 28872 8880 28880
rect 8480 28808 8488 28872
rect 8552 28808 8808 28872
rect 8872 28808 8880 28872
rect 8480 28800 8880 28808
rect 8960 28872 9360 28880
rect 8960 28808 8968 28872
rect 9032 28808 9288 28872
rect 9352 28808 9360 28872
rect 8960 28800 9360 28808
rect 9440 28872 11440 28880
rect 9440 28808 9448 28872
rect 9512 28808 9768 28872
rect 9832 28808 10088 28872
rect 10152 28808 10408 28872
rect 10472 28808 10728 28872
rect 10792 28808 11048 28872
rect 11112 28808 11368 28872
rect 11432 28808 11440 28872
rect 9440 28800 11440 28808
rect 11520 28872 11920 28880
rect 11520 28808 11528 28872
rect 11592 28808 11848 28872
rect 11912 28808 11920 28872
rect 11520 28800 11920 28808
rect 12000 28872 12400 28880
rect 12000 28808 12008 28872
rect 12072 28808 12328 28872
rect 12392 28808 12400 28872
rect 12000 28800 12400 28808
rect 8480 28712 8880 28720
rect 8480 28648 8488 28712
rect 8552 28648 8808 28712
rect 8872 28648 8880 28712
rect 8480 28640 8880 28648
rect 8960 28712 9360 28720
rect 8960 28648 8968 28712
rect 9032 28648 9288 28712
rect 9352 28648 9360 28712
rect 8960 28640 9360 28648
rect 9440 28712 11440 28720
rect 9440 28648 9448 28712
rect 9512 28648 9768 28712
rect 9832 28648 10088 28712
rect 10152 28648 10408 28712
rect 10472 28648 10728 28712
rect 10792 28648 11048 28712
rect 11112 28648 11368 28712
rect 11432 28648 11440 28712
rect 9440 28640 11440 28648
rect 11520 28712 11920 28720
rect 11520 28648 11528 28712
rect 11592 28648 11848 28712
rect 11912 28648 11920 28712
rect 11520 28640 11920 28648
rect 12000 28712 12400 28720
rect 12000 28648 12008 28712
rect 12072 28648 12328 28712
rect 12392 28648 12400 28712
rect 12000 28640 12400 28648
rect 8480 28552 8880 28560
rect 8480 28488 8488 28552
rect 8552 28488 8808 28552
rect 8872 28488 8880 28552
rect 8480 28480 8880 28488
rect 8960 28552 9360 28560
rect 8960 28488 8968 28552
rect 9032 28488 9288 28552
rect 9352 28488 9360 28552
rect 8960 28480 9360 28488
rect 9440 28552 11440 28560
rect 9440 28488 9448 28552
rect 9512 28488 9768 28552
rect 9832 28488 10088 28552
rect 10152 28488 10408 28552
rect 10472 28488 10728 28552
rect 10792 28488 11048 28552
rect 11112 28488 11368 28552
rect 11432 28488 11440 28552
rect 9440 28480 11440 28488
rect 11520 28552 11920 28560
rect 11520 28488 11528 28552
rect 11592 28488 11848 28552
rect 11912 28488 11920 28552
rect 11520 28480 11920 28488
rect 12000 28552 12400 28560
rect 12000 28488 12008 28552
rect 12072 28488 12328 28552
rect 12392 28488 12400 28552
rect 12000 28480 12400 28488
rect 8480 28392 8880 28400
rect 8480 28328 8488 28392
rect 8552 28328 8808 28392
rect 8872 28328 8880 28392
rect 8480 28320 8880 28328
rect 8960 28392 9360 28400
rect 8960 28328 8968 28392
rect 9032 28328 9288 28392
rect 9352 28328 9360 28392
rect 8960 28320 9360 28328
rect 9440 28392 11440 28400
rect 9440 28328 9448 28392
rect 9512 28328 9768 28392
rect 9832 28328 10088 28392
rect 10152 28328 10408 28392
rect 10472 28328 10728 28392
rect 10792 28328 11048 28392
rect 11112 28328 11368 28392
rect 11432 28328 11440 28392
rect 9440 28320 11440 28328
rect 11520 28392 11920 28400
rect 11520 28328 11528 28392
rect 11592 28328 11848 28392
rect 11912 28328 11920 28392
rect 11520 28320 11920 28328
rect 12000 28392 12400 28400
rect 12000 28328 12008 28392
rect 12072 28328 12328 28392
rect 12392 28328 12400 28392
rect 12000 28320 12400 28328
rect 8480 28232 8880 28240
rect 8480 28168 8488 28232
rect 8552 28168 8808 28232
rect 8872 28168 8880 28232
rect 8480 28160 8880 28168
rect 8960 28232 9360 28240
rect 8960 28168 8968 28232
rect 9032 28168 9288 28232
rect 9352 28168 9360 28232
rect 8960 28160 9360 28168
rect 9440 28232 11440 28240
rect 9440 28168 9448 28232
rect 9512 28168 9768 28232
rect 9832 28168 10088 28232
rect 10152 28168 10408 28232
rect 10472 28168 10728 28232
rect 10792 28168 11048 28232
rect 11112 28168 11368 28232
rect 11432 28168 11440 28232
rect 9440 28160 11440 28168
rect 11520 28232 11920 28240
rect 11520 28168 11528 28232
rect 11592 28168 11848 28232
rect 11912 28168 11920 28232
rect 11520 28160 11920 28168
rect 12000 28232 12400 28240
rect 12000 28168 12008 28232
rect 12072 28168 12328 28232
rect 12392 28168 12400 28232
rect 12000 28160 12400 28168
rect 8480 28072 8880 28080
rect 8480 28008 8488 28072
rect 8552 28008 8808 28072
rect 8872 28008 8880 28072
rect 8480 28000 8880 28008
rect 8960 28072 9360 28080
rect 8960 28008 8968 28072
rect 9032 28008 9288 28072
rect 9352 28008 9360 28072
rect 8960 28000 9360 28008
rect 9440 28072 11440 28080
rect 9440 28008 9448 28072
rect 9512 28008 9768 28072
rect 9832 28008 10088 28072
rect 10152 28008 10408 28072
rect 10472 28008 10728 28072
rect 10792 28008 11048 28072
rect 11112 28008 11368 28072
rect 11432 28008 11440 28072
rect 9440 28000 11440 28008
rect 11520 28072 11920 28080
rect 11520 28008 11528 28072
rect 11592 28008 11848 28072
rect 11912 28008 11920 28072
rect 11520 28000 11920 28008
rect 12000 28072 12400 28080
rect 12000 28008 12008 28072
rect 12072 28008 12328 28072
rect 12392 28008 12400 28072
rect 12000 28000 12400 28008
rect 8480 27912 8880 27920
rect 8480 27848 8488 27912
rect 8552 27848 8808 27912
rect 8872 27848 8880 27912
rect 8480 27840 8880 27848
rect 8960 27912 9360 27920
rect 8960 27848 8968 27912
rect 9032 27848 9288 27912
rect 9352 27848 9360 27912
rect 8960 27840 9360 27848
rect 9440 27912 11440 27920
rect 9440 27848 9448 27912
rect 9512 27848 9768 27912
rect 9832 27848 10088 27912
rect 10152 27848 10408 27912
rect 10472 27848 10728 27912
rect 10792 27848 11048 27912
rect 11112 27848 11368 27912
rect 11432 27848 11440 27912
rect 9440 27840 11440 27848
rect 11520 27912 11920 27920
rect 11520 27848 11528 27912
rect 11592 27848 11848 27912
rect 11912 27848 11920 27912
rect 11520 27840 11920 27848
rect 12000 27912 12400 27920
rect 12000 27848 12008 27912
rect 12072 27848 12328 27912
rect 12392 27848 12400 27912
rect 12000 27840 12400 27848
rect 8480 27752 8880 27760
rect 8480 27688 8488 27752
rect 8552 27688 8808 27752
rect 8872 27688 8880 27752
rect 8480 27680 8880 27688
rect 8960 27752 9360 27760
rect 8960 27688 8968 27752
rect 9032 27688 9288 27752
rect 9352 27688 9360 27752
rect 8960 27680 9360 27688
rect 9440 27752 11440 27760
rect 9440 27688 9448 27752
rect 9512 27688 9768 27752
rect 9832 27688 10088 27752
rect 10152 27688 10408 27752
rect 10472 27688 10728 27752
rect 10792 27688 11048 27752
rect 11112 27688 11368 27752
rect 11432 27688 11440 27752
rect 9440 27680 11440 27688
rect 11520 27752 11920 27760
rect 11520 27688 11528 27752
rect 11592 27688 11848 27752
rect 11912 27688 11920 27752
rect 11520 27680 11920 27688
rect 12000 27752 12400 27760
rect 12000 27688 12008 27752
rect 12072 27688 12328 27752
rect 12392 27688 12400 27752
rect 12000 27680 12400 27688
rect 8480 27592 8880 27600
rect 8480 27528 8488 27592
rect 8552 27528 8808 27592
rect 8872 27528 8880 27592
rect 8480 27520 8880 27528
rect 8960 27592 9360 27600
rect 8960 27528 8968 27592
rect 9032 27528 9288 27592
rect 9352 27528 9360 27592
rect 8960 27520 9360 27528
rect 9440 27592 11440 27600
rect 9440 27528 9448 27592
rect 9512 27528 9768 27592
rect 9832 27528 10088 27592
rect 10152 27528 10408 27592
rect 10472 27528 10728 27592
rect 10792 27528 11048 27592
rect 11112 27528 11368 27592
rect 11432 27528 11440 27592
rect 9440 27520 11440 27528
rect 11520 27592 11920 27600
rect 11520 27528 11528 27592
rect 11592 27528 11848 27592
rect 11912 27528 11920 27592
rect 11520 27520 11920 27528
rect 12000 27592 12400 27600
rect 12000 27528 12008 27592
rect 12072 27528 12328 27592
rect 12392 27528 12400 27592
rect 12000 27520 12400 27528
rect 8480 27432 8880 27440
rect 8480 27368 8488 27432
rect 8552 27368 8808 27432
rect 8872 27368 8880 27432
rect 8480 27360 8880 27368
rect 8960 27432 9360 27440
rect 8960 27368 8968 27432
rect 9032 27368 9288 27432
rect 9352 27368 9360 27432
rect 8960 27360 9360 27368
rect 9440 27432 11440 27440
rect 9440 27368 9448 27432
rect 9512 27368 9768 27432
rect 9832 27368 10088 27432
rect 10152 27368 10408 27432
rect 10472 27368 10728 27432
rect 10792 27368 11048 27432
rect 11112 27368 11368 27432
rect 11432 27368 11440 27432
rect 9440 27360 11440 27368
rect 11520 27432 11920 27440
rect 11520 27368 11528 27432
rect 11592 27368 11848 27432
rect 11912 27368 11920 27432
rect 11520 27360 11920 27368
rect 12000 27432 12400 27440
rect 12000 27368 12008 27432
rect 12072 27368 12328 27432
rect 12392 27368 12400 27432
rect 12000 27360 12400 27368
rect 8480 27272 8880 27280
rect 8480 27208 8488 27272
rect 8552 27208 8808 27272
rect 8872 27208 8880 27272
rect 8480 27200 8880 27208
rect 8960 27272 9360 27280
rect 8960 27208 8968 27272
rect 9032 27208 9288 27272
rect 9352 27208 9360 27272
rect 8960 27200 9360 27208
rect 9440 27272 11440 27280
rect 9440 27208 9448 27272
rect 9512 27208 9768 27272
rect 9832 27208 10088 27272
rect 10152 27208 10408 27272
rect 10472 27208 10728 27272
rect 10792 27208 11048 27272
rect 11112 27208 11368 27272
rect 11432 27208 11440 27272
rect 9440 27200 11440 27208
rect 11520 27272 11920 27280
rect 11520 27208 11528 27272
rect 11592 27208 11848 27272
rect 11912 27208 11920 27272
rect 11520 27200 11920 27208
rect 12000 27272 12400 27280
rect 12000 27208 12008 27272
rect 12072 27208 12328 27272
rect 12392 27208 12400 27272
rect 12000 27200 12400 27208
rect 8480 27112 8880 27120
rect 8480 27048 8488 27112
rect 8552 27048 8808 27112
rect 8872 27048 8880 27112
rect 8480 27040 8880 27048
rect 8960 27112 9360 27120
rect 8960 27048 8968 27112
rect 9032 27048 9288 27112
rect 9352 27048 9360 27112
rect 8960 27040 9360 27048
rect 9440 27112 11440 27120
rect 9440 27048 9448 27112
rect 9512 27048 9768 27112
rect 9832 27048 10088 27112
rect 10152 27048 10408 27112
rect 10472 27048 10728 27112
rect 10792 27048 11048 27112
rect 11112 27048 11368 27112
rect 11432 27048 11440 27112
rect 9440 27040 11440 27048
rect 11520 27112 11920 27120
rect 11520 27048 11528 27112
rect 11592 27048 11848 27112
rect 11912 27048 11920 27112
rect 11520 27040 11920 27048
rect 12000 27112 12400 27120
rect 12000 27048 12008 27112
rect 12072 27048 12328 27112
rect 12392 27048 12400 27112
rect 12000 27040 12400 27048
rect 8480 26952 8880 26960
rect 8480 26888 8488 26952
rect 8552 26888 8808 26952
rect 8872 26888 8880 26952
rect 8480 26880 8880 26888
rect 8960 26952 9360 26960
rect 8960 26888 8968 26952
rect 9032 26888 9288 26952
rect 9352 26888 9360 26952
rect 8960 26880 9360 26888
rect 9440 26952 11440 26960
rect 9440 26888 9448 26952
rect 9512 26888 9768 26952
rect 9832 26888 10088 26952
rect 10152 26888 10408 26952
rect 10472 26888 10728 26952
rect 10792 26888 11048 26952
rect 11112 26888 11368 26952
rect 11432 26888 11440 26952
rect 9440 26880 11440 26888
rect 11520 26952 11920 26960
rect 11520 26888 11528 26952
rect 11592 26888 11848 26952
rect 11912 26888 11920 26952
rect 11520 26880 11920 26888
rect 12000 26952 12400 26960
rect 12000 26888 12008 26952
rect 12072 26888 12328 26952
rect 12392 26888 12400 26952
rect 12000 26880 12400 26888
rect 8480 26792 8880 26800
rect 8480 26728 8488 26792
rect 8552 26728 8808 26792
rect 8872 26728 8880 26792
rect 8480 26720 8880 26728
rect 8960 26792 9360 26800
rect 8960 26728 8968 26792
rect 9032 26728 9288 26792
rect 9352 26728 9360 26792
rect 8960 26720 9360 26728
rect 9440 26792 11440 26800
rect 9440 26728 9448 26792
rect 9512 26728 9768 26792
rect 9832 26728 10088 26792
rect 10152 26728 10408 26792
rect 10472 26728 10728 26792
rect 10792 26728 11048 26792
rect 11112 26728 11368 26792
rect 11432 26728 11440 26792
rect 9440 26720 11440 26728
rect 11520 26792 11920 26800
rect 11520 26728 11528 26792
rect 11592 26728 11848 26792
rect 11912 26728 11920 26792
rect 11520 26720 11920 26728
rect 12000 26792 12400 26800
rect 12000 26728 12008 26792
rect 12072 26728 12328 26792
rect 12392 26728 12400 26792
rect 12000 26720 12400 26728
rect 8480 26632 8880 26640
rect 8480 26568 8488 26632
rect 8552 26568 8808 26632
rect 8872 26568 8880 26632
rect 8480 26560 8880 26568
rect 8960 26632 9360 26640
rect 8960 26568 8968 26632
rect 9032 26568 9288 26632
rect 9352 26568 9360 26632
rect 8960 26560 9360 26568
rect 9440 26632 11440 26640
rect 9440 26568 9448 26632
rect 9512 26568 9768 26632
rect 9832 26568 10088 26632
rect 10152 26568 10408 26632
rect 10472 26568 10728 26632
rect 10792 26568 11048 26632
rect 11112 26568 11368 26632
rect 11432 26568 11440 26632
rect 9440 26560 11440 26568
rect 11520 26632 11920 26640
rect 11520 26568 11528 26632
rect 11592 26568 11848 26632
rect 11912 26568 11920 26632
rect 11520 26560 11920 26568
rect 12000 26632 12400 26640
rect 12000 26568 12008 26632
rect 12072 26568 12328 26632
rect 12392 26568 12400 26632
rect 12000 26560 12400 26568
rect 8480 26472 8880 26480
rect 8480 26408 8488 26472
rect 8552 26408 8808 26472
rect 8872 26408 8880 26472
rect 8480 26400 8880 26408
rect 8960 26472 9360 26480
rect 8960 26408 8968 26472
rect 9032 26408 9288 26472
rect 9352 26408 9360 26472
rect 8960 26400 9360 26408
rect 9440 26472 11440 26480
rect 9440 26408 9448 26472
rect 9512 26408 9768 26472
rect 9832 26408 10088 26472
rect 10152 26408 10408 26472
rect 10472 26408 10728 26472
rect 10792 26408 11048 26472
rect 11112 26408 11368 26472
rect 11432 26408 11440 26472
rect 9440 26400 11440 26408
rect 11520 26472 11920 26480
rect 11520 26408 11528 26472
rect 11592 26408 11848 26472
rect 11912 26408 11920 26472
rect 11520 26400 11920 26408
rect 12000 26472 12400 26480
rect 12000 26408 12008 26472
rect 12072 26408 12328 26472
rect 12392 26408 12400 26472
rect 12000 26400 12400 26408
rect 8480 26312 8880 26320
rect 8480 26248 8488 26312
rect 8552 26248 8808 26312
rect 8872 26248 8880 26312
rect 8480 26240 8880 26248
rect 8960 26312 9360 26320
rect 8960 26248 8968 26312
rect 9032 26248 9288 26312
rect 9352 26248 9360 26312
rect 8960 26240 9360 26248
rect 9440 26312 11440 26320
rect 9440 26248 9448 26312
rect 9512 26248 9768 26312
rect 9832 26248 10088 26312
rect 10152 26248 10408 26312
rect 10472 26248 10728 26312
rect 10792 26248 11048 26312
rect 11112 26248 11368 26312
rect 11432 26248 11440 26312
rect 9440 26240 11440 26248
rect 11520 26312 11920 26320
rect 11520 26248 11528 26312
rect 11592 26248 11848 26312
rect 11912 26248 11920 26312
rect 11520 26240 11920 26248
rect 12000 26312 12400 26320
rect 12000 26248 12008 26312
rect 12072 26248 12328 26312
rect 12392 26248 12400 26312
rect 12000 26240 12400 26248
rect 8480 26152 8880 26160
rect 8480 26088 8488 26152
rect 8552 26088 8808 26152
rect 8872 26088 8880 26152
rect 8480 26080 8880 26088
rect 8960 26152 9360 26160
rect 8960 26088 8968 26152
rect 9032 26088 9288 26152
rect 9352 26088 9360 26152
rect 8960 26080 9360 26088
rect 9440 26152 11440 26160
rect 9440 26088 9448 26152
rect 9512 26088 9768 26152
rect 9832 26088 10088 26152
rect 10152 26088 10408 26152
rect 10472 26088 10728 26152
rect 10792 26088 11048 26152
rect 11112 26088 11368 26152
rect 11432 26088 11440 26152
rect 9440 26080 11440 26088
rect 11520 26152 11920 26160
rect 11520 26088 11528 26152
rect 11592 26088 11848 26152
rect 11912 26088 11920 26152
rect 11520 26080 11920 26088
rect 12000 26152 12400 26160
rect 12000 26088 12008 26152
rect 12072 26088 12328 26152
rect 12392 26088 12400 26152
rect 12000 26080 12400 26088
rect 8480 25992 8880 26000
rect 8480 25928 8488 25992
rect 8552 25928 8808 25992
rect 8872 25928 8880 25992
rect 8480 25920 8880 25928
rect 8960 25992 9360 26000
rect 8960 25928 8968 25992
rect 9032 25928 9288 25992
rect 9352 25928 9360 25992
rect 8960 25920 9360 25928
rect 9440 25992 11440 26000
rect 9440 25928 9448 25992
rect 9512 25928 9768 25992
rect 9832 25928 10088 25992
rect 10152 25928 10408 25992
rect 10472 25928 10728 25992
rect 10792 25928 11048 25992
rect 11112 25928 11368 25992
rect 11432 25928 11440 25992
rect 9440 25920 11440 25928
rect 11520 25992 11920 26000
rect 11520 25928 11528 25992
rect 11592 25928 11848 25992
rect 11912 25928 11920 25992
rect 11520 25920 11920 25928
rect 12000 25992 12400 26000
rect 12000 25928 12008 25992
rect 12072 25928 12328 25992
rect 12392 25928 12400 25992
rect 12000 25920 12400 25928
rect 8480 25832 8880 25840
rect 8480 25768 8488 25832
rect 8552 25768 8808 25832
rect 8872 25768 8880 25832
rect 8480 25760 8880 25768
rect 8960 25832 9360 25840
rect 8960 25768 8968 25832
rect 9032 25768 9288 25832
rect 9352 25768 9360 25832
rect 8960 25760 9360 25768
rect 9440 25832 11440 25840
rect 9440 25768 9448 25832
rect 9512 25768 9768 25832
rect 9832 25768 10088 25832
rect 10152 25768 10408 25832
rect 10472 25768 10728 25832
rect 10792 25768 11048 25832
rect 11112 25768 11368 25832
rect 11432 25768 11440 25832
rect 9440 25760 11440 25768
rect 11520 25832 11920 25840
rect 11520 25768 11528 25832
rect 11592 25768 11848 25832
rect 11912 25768 11920 25832
rect 11520 25760 11920 25768
rect 12000 25832 12400 25840
rect 12000 25768 12008 25832
rect 12072 25768 12328 25832
rect 12392 25768 12400 25832
rect 12000 25760 12400 25768
rect 8480 25672 8880 25680
rect 8480 25608 8488 25672
rect 8552 25608 8808 25672
rect 8872 25608 8880 25672
rect 8480 25600 8880 25608
rect 8960 25672 9360 25680
rect 8960 25608 8968 25672
rect 9032 25608 9288 25672
rect 9352 25608 9360 25672
rect 8960 25600 9360 25608
rect 9440 25672 11440 25680
rect 9440 25608 9448 25672
rect 9512 25608 9768 25672
rect 9832 25608 10088 25672
rect 10152 25608 10408 25672
rect 10472 25608 10728 25672
rect 10792 25608 11048 25672
rect 11112 25608 11368 25672
rect 11432 25608 11440 25672
rect 9440 25600 11440 25608
rect 11520 25672 11920 25680
rect 11520 25608 11528 25672
rect 11592 25608 11848 25672
rect 11912 25608 11920 25672
rect 11520 25600 11920 25608
rect 12000 25672 12400 25680
rect 12000 25608 12008 25672
rect 12072 25608 12328 25672
rect 12392 25608 12400 25672
rect 12000 25600 12400 25608
rect 8480 25512 8880 25520
rect 8480 25448 8488 25512
rect 8552 25448 8808 25512
rect 8872 25448 8880 25512
rect 8480 25440 8880 25448
rect 8960 25512 9360 25520
rect 8960 25448 8968 25512
rect 9032 25448 9288 25512
rect 9352 25448 9360 25512
rect 8960 25440 9360 25448
rect 9440 25512 11440 25520
rect 9440 25448 9448 25512
rect 9512 25448 9768 25512
rect 9832 25448 10088 25512
rect 10152 25448 10408 25512
rect 10472 25448 10728 25512
rect 10792 25448 11048 25512
rect 11112 25448 11368 25512
rect 11432 25448 11440 25512
rect 9440 25440 11440 25448
rect 11520 25512 11920 25520
rect 11520 25448 11528 25512
rect 11592 25448 11848 25512
rect 11912 25448 11920 25512
rect 11520 25440 11920 25448
rect 12000 25512 12400 25520
rect 12000 25448 12008 25512
rect 12072 25448 12328 25512
rect 12392 25448 12400 25512
rect 12000 25440 12400 25448
rect 8480 25352 8880 25360
rect 8480 25288 8488 25352
rect 8552 25288 8808 25352
rect 8872 25288 8880 25352
rect 8480 25280 8880 25288
rect 8960 25352 9360 25360
rect 8960 25288 8968 25352
rect 9032 25288 9288 25352
rect 9352 25288 9360 25352
rect 8960 25280 9360 25288
rect 9440 25352 11440 25360
rect 9440 25288 9448 25352
rect 9512 25288 9768 25352
rect 9832 25288 10088 25352
rect 10152 25288 10408 25352
rect 10472 25288 10728 25352
rect 10792 25288 11048 25352
rect 11112 25288 11368 25352
rect 11432 25288 11440 25352
rect 9440 25280 11440 25288
rect 11520 25352 11920 25360
rect 11520 25288 11528 25352
rect 11592 25288 11848 25352
rect 11912 25288 11920 25352
rect 11520 25280 11920 25288
rect 12000 25352 12400 25360
rect 12000 25288 12008 25352
rect 12072 25288 12328 25352
rect 12392 25288 12400 25352
rect 12000 25280 12400 25288
rect 8480 25192 8880 25200
rect 8480 25128 8488 25192
rect 8552 25128 8808 25192
rect 8872 25128 8880 25192
rect 8480 25120 8880 25128
rect 8960 25192 9360 25200
rect 8960 25128 8968 25192
rect 9032 25128 9288 25192
rect 9352 25128 9360 25192
rect 8960 25120 9360 25128
rect 9440 25192 11440 25200
rect 9440 25128 9448 25192
rect 9512 25128 9768 25192
rect 9832 25128 10088 25192
rect 10152 25128 10408 25192
rect 10472 25128 10728 25192
rect 10792 25128 11048 25192
rect 11112 25128 11368 25192
rect 11432 25128 11440 25192
rect 9440 25120 11440 25128
rect 11520 25192 11920 25200
rect 11520 25128 11528 25192
rect 11592 25128 11848 25192
rect 11912 25128 11920 25192
rect 11520 25120 11920 25128
rect 12000 25192 12400 25200
rect 12000 25128 12008 25192
rect 12072 25128 12328 25192
rect 12392 25128 12400 25192
rect 12000 25120 12400 25128
rect 8480 25032 8880 25040
rect 8480 24968 8488 25032
rect 8552 24968 8808 25032
rect 8872 24968 8880 25032
rect 8480 24960 8880 24968
rect 8960 25032 9360 25040
rect 8960 24968 8968 25032
rect 9032 24968 9288 25032
rect 9352 24968 9360 25032
rect 8960 24960 9360 24968
rect 9440 25032 11440 25040
rect 9440 24968 9448 25032
rect 9512 24968 9768 25032
rect 9832 24968 10088 25032
rect 10152 24968 10408 25032
rect 10472 24968 10728 25032
rect 10792 24968 11048 25032
rect 11112 24968 11368 25032
rect 11432 24968 11440 25032
rect 9440 24960 11440 24968
rect 11520 25032 11920 25040
rect 11520 24968 11528 25032
rect 11592 24968 11848 25032
rect 11912 24968 11920 25032
rect 11520 24960 11920 24968
rect 12000 25032 12400 25040
rect 12000 24968 12008 25032
rect 12072 24968 12328 25032
rect 12392 24968 12400 25032
rect 12000 24960 12400 24968
rect 8480 24872 8880 24880
rect 8480 24808 8488 24872
rect 8552 24808 8808 24872
rect 8872 24808 8880 24872
rect 8480 24800 8880 24808
rect 8960 24872 9360 24880
rect 8960 24808 8968 24872
rect 9032 24808 9288 24872
rect 9352 24808 9360 24872
rect 8960 24800 9360 24808
rect 9440 24872 11440 24880
rect 9440 24808 9448 24872
rect 9512 24808 9768 24872
rect 9832 24808 10088 24872
rect 10152 24808 10408 24872
rect 10472 24808 10728 24872
rect 10792 24808 11048 24872
rect 11112 24808 11368 24872
rect 11432 24808 11440 24872
rect 9440 24800 11440 24808
rect 11520 24872 11920 24880
rect 11520 24808 11528 24872
rect 11592 24808 11848 24872
rect 11912 24808 11920 24872
rect 11520 24800 11920 24808
rect 12000 24872 12400 24880
rect 12000 24808 12008 24872
rect 12072 24808 12328 24872
rect 12392 24808 12400 24872
rect 12000 24800 12400 24808
rect 8480 24712 8880 24720
rect 8480 24648 8488 24712
rect 8552 24648 8808 24712
rect 8872 24648 8880 24712
rect 8480 24640 8880 24648
rect 8960 24712 9360 24720
rect 8960 24648 8968 24712
rect 9032 24648 9288 24712
rect 9352 24648 9360 24712
rect 8960 24640 9360 24648
rect 9440 24712 11440 24720
rect 9440 24648 9448 24712
rect 9512 24648 9768 24712
rect 9832 24648 10088 24712
rect 10152 24648 10408 24712
rect 10472 24648 10728 24712
rect 10792 24648 11048 24712
rect 11112 24648 11368 24712
rect 11432 24648 11440 24712
rect 9440 24640 11440 24648
rect 11520 24712 11920 24720
rect 11520 24648 11528 24712
rect 11592 24648 11848 24712
rect 11912 24648 11920 24712
rect 11520 24640 11920 24648
rect 12000 24712 12400 24720
rect 12000 24648 12008 24712
rect 12072 24648 12328 24712
rect 12392 24648 12400 24712
rect 12000 24640 12400 24648
rect 8480 24552 8880 24560
rect 8480 24488 8488 24552
rect 8552 24488 8808 24552
rect 8872 24488 8880 24552
rect 8480 24480 8880 24488
rect 8960 24552 9360 24560
rect 8960 24488 8968 24552
rect 9032 24488 9288 24552
rect 9352 24488 9360 24552
rect 8960 24480 9360 24488
rect 9440 24552 11440 24560
rect 9440 24488 9448 24552
rect 9512 24488 9768 24552
rect 9832 24488 10088 24552
rect 10152 24488 10408 24552
rect 10472 24488 10728 24552
rect 10792 24488 11048 24552
rect 11112 24488 11368 24552
rect 11432 24488 11440 24552
rect 9440 24480 11440 24488
rect 11520 24552 11920 24560
rect 11520 24488 11528 24552
rect 11592 24488 11848 24552
rect 11912 24488 11920 24552
rect 11520 24480 11920 24488
rect 12000 24552 12400 24560
rect 12000 24488 12008 24552
rect 12072 24488 12328 24552
rect 12392 24488 12400 24552
rect 12000 24480 12400 24488
rect 8480 24392 8880 24400
rect 8480 24328 8488 24392
rect 8552 24328 8808 24392
rect 8872 24328 8880 24392
rect 8480 24320 8880 24328
rect 8960 24392 9360 24400
rect 8960 24328 8968 24392
rect 9032 24328 9288 24392
rect 9352 24328 9360 24392
rect 8960 24320 9360 24328
rect 9440 24392 11440 24400
rect 9440 24328 9448 24392
rect 9512 24328 9768 24392
rect 9832 24328 10088 24392
rect 10152 24328 10408 24392
rect 10472 24328 10728 24392
rect 10792 24328 11048 24392
rect 11112 24328 11368 24392
rect 11432 24328 11440 24392
rect 9440 24320 11440 24328
rect 11520 24392 11920 24400
rect 11520 24328 11528 24392
rect 11592 24328 11848 24392
rect 11912 24328 11920 24392
rect 11520 24320 11920 24328
rect 12000 24392 12400 24400
rect 12000 24328 12008 24392
rect 12072 24328 12328 24392
rect 12392 24328 12400 24392
rect 12000 24320 12400 24328
rect 8480 24232 8880 24240
rect 8480 24168 8488 24232
rect 8552 24168 8808 24232
rect 8872 24168 8880 24232
rect 8480 24160 8880 24168
rect 8960 24232 9360 24240
rect 8960 24168 8968 24232
rect 9032 24168 9288 24232
rect 9352 24168 9360 24232
rect 8960 24160 9360 24168
rect 9440 24232 11440 24240
rect 9440 24168 9448 24232
rect 9512 24168 9768 24232
rect 9832 24168 10088 24232
rect 10152 24168 10408 24232
rect 10472 24168 10728 24232
rect 10792 24168 11048 24232
rect 11112 24168 11368 24232
rect 11432 24168 11440 24232
rect 9440 24160 11440 24168
rect 11520 24232 11920 24240
rect 11520 24168 11528 24232
rect 11592 24168 11848 24232
rect 11912 24168 11920 24232
rect 11520 24160 11920 24168
rect 12000 24232 12400 24240
rect 12000 24168 12008 24232
rect 12072 24168 12328 24232
rect 12392 24168 12400 24232
rect 12000 24160 12400 24168
rect 8480 24072 8880 24080
rect 8480 24008 8488 24072
rect 8552 24008 8808 24072
rect 8872 24008 8880 24072
rect 8480 24000 8880 24008
rect 8960 24072 9360 24080
rect 8960 24008 8968 24072
rect 9032 24008 9288 24072
rect 9352 24008 9360 24072
rect 8960 24000 9360 24008
rect 9440 24072 11440 24080
rect 9440 24008 9448 24072
rect 9512 24008 9768 24072
rect 9832 24008 10088 24072
rect 10152 24008 10408 24072
rect 10472 24008 10728 24072
rect 10792 24008 11048 24072
rect 11112 24008 11368 24072
rect 11432 24008 11440 24072
rect 9440 24000 11440 24008
rect 11520 24072 11920 24080
rect 11520 24008 11528 24072
rect 11592 24008 11848 24072
rect 11912 24008 11920 24072
rect 11520 24000 11920 24008
rect 12000 24072 12400 24080
rect 12000 24008 12008 24072
rect 12072 24008 12328 24072
rect 12392 24008 12400 24072
rect 12000 24000 12400 24008
rect 8480 23912 8880 23920
rect 8480 23848 8488 23912
rect 8552 23848 8808 23912
rect 8872 23848 8880 23912
rect 8480 23840 8880 23848
rect 8960 23912 9360 23920
rect 8960 23848 8968 23912
rect 9032 23848 9288 23912
rect 9352 23848 9360 23912
rect 8960 23840 9360 23848
rect 9440 23912 11440 23920
rect 9440 23848 9448 23912
rect 9512 23848 9768 23912
rect 9832 23848 10088 23912
rect 10152 23848 10408 23912
rect 10472 23848 10728 23912
rect 10792 23848 11048 23912
rect 11112 23848 11368 23912
rect 11432 23848 11440 23912
rect 9440 23840 11440 23848
rect 11520 23912 11920 23920
rect 11520 23848 11528 23912
rect 11592 23848 11848 23912
rect 11912 23848 11920 23912
rect 11520 23840 11920 23848
rect 12000 23912 12400 23920
rect 12000 23848 12008 23912
rect 12072 23848 12328 23912
rect 12392 23848 12400 23912
rect 12000 23840 12400 23848
rect 8480 23752 8880 23760
rect 8480 23688 8488 23752
rect 8552 23688 8808 23752
rect 8872 23688 8880 23752
rect 8480 23680 8880 23688
rect 8960 23752 9360 23760
rect 8960 23688 8968 23752
rect 9032 23688 9288 23752
rect 9352 23688 9360 23752
rect 8960 23680 9360 23688
rect 9440 23752 11440 23760
rect 9440 23688 9448 23752
rect 9512 23688 9768 23752
rect 9832 23688 10088 23752
rect 10152 23688 10408 23752
rect 10472 23688 10728 23752
rect 10792 23688 11048 23752
rect 11112 23688 11368 23752
rect 11432 23688 11440 23752
rect 9440 23680 11440 23688
rect 11520 23752 11920 23760
rect 11520 23688 11528 23752
rect 11592 23688 11848 23752
rect 11912 23688 11920 23752
rect 11520 23680 11920 23688
rect 12000 23752 12400 23760
rect 12000 23688 12008 23752
rect 12072 23688 12328 23752
rect 12392 23688 12400 23752
rect 12000 23680 12400 23688
rect 8480 23592 8880 23600
rect 8480 23528 8488 23592
rect 8552 23528 8808 23592
rect 8872 23528 8880 23592
rect 8480 23520 8880 23528
rect 8960 23592 9360 23600
rect 8960 23528 8968 23592
rect 9032 23528 9288 23592
rect 9352 23528 9360 23592
rect 8960 23520 9360 23528
rect 9440 23592 11440 23600
rect 9440 23528 9448 23592
rect 9512 23528 9768 23592
rect 9832 23528 10088 23592
rect 10152 23528 10408 23592
rect 10472 23528 10728 23592
rect 10792 23528 11048 23592
rect 11112 23528 11368 23592
rect 11432 23528 11440 23592
rect 9440 23520 11440 23528
rect 11520 23592 11920 23600
rect 11520 23528 11528 23592
rect 11592 23528 11848 23592
rect 11912 23528 11920 23592
rect 11520 23520 11920 23528
rect 12000 23592 12400 23600
rect 12000 23528 12008 23592
rect 12072 23528 12328 23592
rect 12392 23528 12400 23592
rect 12000 23520 12400 23528
rect 8480 23432 8880 23440
rect 8480 23368 8488 23432
rect 8552 23368 8808 23432
rect 8872 23368 8880 23432
rect 8480 23360 8880 23368
rect 8960 23432 9360 23440
rect 8960 23368 8968 23432
rect 9032 23368 9288 23432
rect 9352 23368 9360 23432
rect 8960 23360 9360 23368
rect 9440 23432 11440 23440
rect 9440 23368 9448 23432
rect 9512 23368 9768 23432
rect 9832 23368 10088 23432
rect 10152 23368 10408 23432
rect 10472 23368 10728 23432
rect 10792 23368 11048 23432
rect 11112 23368 11368 23432
rect 11432 23368 11440 23432
rect 9440 23360 11440 23368
rect 11520 23432 11920 23440
rect 11520 23368 11528 23432
rect 11592 23368 11848 23432
rect 11912 23368 11920 23432
rect 11520 23360 11920 23368
rect 12000 23432 12400 23440
rect 12000 23368 12008 23432
rect 12072 23368 12328 23432
rect 12392 23368 12400 23432
rect 12000 23360 12400 23368
rect 8480 23272 8880 23280
rect 8480 23208 8488 23272
rect 8552 23208 8808 23272
rect 8872 23208 8880 23272
rect 8480 23200 8880 23208
rect 8960 23272 9360 23280
rect 8960 23208 8968 23272
rect 9032 23208 9288 23272
rect 9352 23208 9360 23272
rect 8960 23200 9360 23208
rect 9440 23272 11440 23280
rect 9440 23208 9448 23272
rect 9512 23208 9768 23272
rect 9832 23208 10088 23272
rect 10152 23208 10408 23272
rect 10472 23208 10728 23272
rect 10792 23208 11048 23272
rect 11112 23208 11368 23272
rect 11432 23208 11440 23272
rect 9440 23200 11440 23208
rect 11520 23272 11920 23280
rect 11520 23208 11528 23272
rect 11592 23208 11848 23272
rect 11912 23208 11920 23272
rect 11520 23200 11920 23208
rect 12000 23272 12400 23280
rect 12000 23208 12008 23272
rect 12072 23208 12328 23272
rect 12392 23208 12400 23272
rect 12000 23200 12400 23208
rect 8480 23112 8880 23120
rect 8480 23048 8488 23112
rect 8552 23048 8808 23112
rect 8872 23048 8880 23112
rect 8480 23040 8880 23048
rect 8960 23112 9360 23120
rect 8960 23048 8968 23112
rect 9032 23048 9288 23112
rect 9352 23048 9360 23112
rect 8960 23040 9360 23048
rect 9440 23112 11440 23120
rect 9440 23048 9448 23112
rect 9512 23048 9768 23112
rect 9832 23048 10088 23112
rect 10152 23048 10408 23112
rect 10472 23048 10728 23112
rect 10792 23048 11048 23112
rect 11112 23048 11368 23112
rect 11432 23048 11440 23112
rect 9440 23040 11440 23048
rect 11520 23112 11920 23120
rect 11520 23048 11528 23112
rect 11592 23048 11848 23112
rect 11912 23048 11920 23112
rect 11520 23040 11920 23048
rect 12000 23112 12400 23120
rect 12000 23048 12008 23112
rect 12072 23048 12328 23112
rect 12392 23048 12400 23112
rect 12000 23040 12400 23048
rect 8480 22952 8880 22960
rect 8480 22888 8488 22952
rect 8552 22888 8808 22952
rect 8872 22888 8880 22952
rect 8480 22880 8880 22888
rect 8960 22952 9360 22960
rect 8960 22888 8968 22952
rect 9032 22888 9288 22952
rect 9352 22888 9360 22952
rect 8960 22880 9360 22888
rect 9440 22952 11440 22960
rect 9440 22888 9448 22952
rect 9512 22888 9768 22952
rect 9832 22888 10088 22952
rect 10152 22888 10408 22952
rect 10472 22888 10728 22952
rect 10792 22888 11048 22952
rect 11112 22888 11368 22952
rect 11432 22888 11440 22952
rect 9440 22880 11440 22888
rect 11520 22952 11920 22960
rect 11520 22888 11528 22952
rect 11592 22888 11848 22952
rect 11912 22888 11920 22952
rect 11520 22880 11920 22888
rect 12000 22952 12400 22960
rect 12000 22888 12008 22952
rect 12072 22888 12328 22952
rect 12392 22888 12400 22952
rect 12000 22880 12400 22888
rect 8480 22792 8880 22800
rect 8480 22728 8488 22792
rect 8552 22728 8808 22792
rect 8872 22728 8880 22792
rect 8480 22720 8880 22728
rect 8960 22792 9360 22800
rect 8960 22728 8968 22792
rect 9032 22728 9288 22792
rect 9352 22728 9360 22792
rect 8960 22720 9360 22728
rect 9440 22792 11440 22800
rect 9440 22728 9448 22792
rect 9512 22728 9768 22792
rect 9832 22728 10088 22792
rect 10152 22728 10408 22792
rect 10472 22728 10728 22792
rect 10792 22728 11048 22792
rect 11112 22728 11368 22792
rect 11432 22728 11440 22792
rect 9440 22720 11440 22728
rect 11520 22792 11920 22800
rect 11520 22728 11528 22792
rect 11592 22728 11848 22792
rect 11912 22728 11920 22792
rect 11520 22720 11920 22728
rect 12000 22792 12400 22800
rect 12000 22728 12008 22792
rect 12072 22728 12328 22792
rect 12392 22728 12400 22792
rect 12000 22720 12400 22728
rect 8480 22632 8880 22640
rect 8480 22568 8488 22632
rect 8552 22568 8808 22632
rect 8872 22568 8880 22632
rect 8480 22560 8880 22568
rect 8960 22632 9360 22640
rect 8960 22568 8968 22632
rect 9032 22568 9288 22632
rect 9352 22568 9360 22632
rect 8960 22560 9360 22568
rect 9440 22632 11440 22640
rect 9440 22568 9448 22632
rect 9512 22568 9768 22632
rect 9832 22568 10088 22632
rect 10152 22568 10408 22632
rect 10472 22568 10728 22632
rect 10792 22568 11048 22632
rect 11112 22568 11368 22632
rect 11432 22568 11440 22632
rect 9440 22560 11440 22568
rect 11520 22632 11920 22640
rect 11520 22568 11528 22632
rect 11592 22568 11848 22632
rect 11912 22568 11920 22632
rect 11520 22560 11920 22568
rect 12000 22632 12400 22640
rect 12000 22568 12008 22632
rect 12072 22568 12328 22632
rect 12392 22568 12400 22632
rect 12000 22560 12400 22568
rect 8480 22472 8880 22480
rect 8480 22408 8488 22472
rect 8552 22408 8808 22472
rect 8872 22408 8880 22472
rect 8480 22400 8880 22408
rect 8960 22472 9360 22480
rect 8960 22408 8968 22472
rect 9032 22408 9288 22472
rect 9352 22408 9360 22472
rect 8960 22400 9360 22408
rect 9440 22472 11440 22480
rect 9440 22408 9448 22472
rect 9512 22408 9768 22472
rect 9832 22408 10088 22472
rect 10152 22408 10408 22472
rect 10472 22408 10728 22472
rect 10792 22408 11048 22472
rect 11112 22408 11368 22472
rect 11432 22408 11440 22472
rect 9440 22400 11440 22408
rect 11520 22472 11920 22480
rect 11520 22408 11528 22472
rect 11592 22408 11848 22472
rect 11912 22408 11920 22472
rect 11520 22400 11920 22408
rect 12000 22472 12400 22480
rect 12000 22408 12008 22472
rect 12072 22408 12328 22472
rect 12392 22408 12400 22472
rect 12000 22400 12400 22408
rect 8480 22312 8880 22320
rect 8480 22248 8488 22312
rect 8552 22248 8808 22312
rect 8872 22248 8880 22312
rect 8480 22240 8880 22248
rect 8960 22312 9360 22320
rect 8960 22248 8968 22312
rect 9032 22248 9288 22312
rect 9352 22248 9360 22312
rect 8960 22240 9360 22248
rect 9440 22312 11440 22320
rect 9440 22248 9448 22312
rect 9512 22248 9768 22312
rect 9832 22248 10088 22312
rect 10152 22248 10408 22312
rect 10472 22248 10728 22312
rect 10792 22248 11048 22312
rect 11112 22248 11368 22312
rect 11432 22248 11440 22312
rect 9440 22240 11440 22248
rect 11520 22312 11920 22320
rect 11520 22248 11528 22312
rect 11592 22248 11848 22312
rect 11912 22248 11920 22312
rect 11520 22240 11920 22248
rect 12000 22312 12400 22320
rect 12000 22248 12008 22312
rect 12072 22248 12328 22312
rect 12392 22248 12400 22312
rect 12000 22240 12400 22248
rect 8480 22152 8880 22160
rect 8480 22088 8488 22152
rect 8552 22088 8808 22152
rect 8872 22088 8880 22152
rect 8480 22080 8880 22088
rect 8960 22152 9360 22160
rect 8960 22088 8968 22152
rect 9032 22088 9288 22152
rect 9352 22088 9360 22152
rect 8960 22080 9360 22088
rect 9440 22152 11440 22160
rect 9440 22088 9448 22152
rect 9512 22088 9768 22152
rect 9832 22088 10088 22152
rect 10152 22088 10408 22152
rect 10472 22088 10728 22152
rect 10792 22088 11048 22152
rect 11112 22088 11368 22152
rect 11432 22088 11440 22152
rect 9440 22080 11440 22088
rect 11520 22152 11920 22160
rect 11520 22088 11528 22152
rect 11592 22088 11848 22152
rect 11912 22088 11920 22152
rect 11520 22080 11920 22088
rect 12000 22152 12400 22160
rect 12000 22088 12008 22152
rect 12072 22088 12328 22152
rect 12392 22088 12400 22152
rect 12000 22080 12400 22088
rect 8480 21992 8880 22000
rect 8480 21928 8488 21992
rect 8552 21928 8808 21992
rect 8872 21928 8880 21992
rect 8480 21920 8880 21928
rect 8960 21992 9360 22000
rect 8960 21928 8968 21992
rect 9032 21928 9288 21992
rect 9352 21928 9360 21992
rect 8960 21920 9360 21928
rect 9440 21992 11440 22000
rect 9440 21928 9448 21992
rect 9512 21928 9768 21992
rect 9832 21928 10088 21992
rect 10152 21928 10408 21992
rect 10472 21928 10728 21992
rect 10792 21928 11048 21992
rect 11112 21928 11368 21992
rect 11432 21928 11440 21992
rect 9440 21920 11440 21928
rect 11520 21992 11920 22000
rect 11520 21928 11528 21992
rect 11592 21928 11848 21992
rect 11912 21928 11920 21992
rect 11520 21920 11920 21928
rect 12000 21992 12400 22000
rect 12000 21928 12008 21992
rect 12072 21928 12328 21992
rect 12392 21928 12400 21992
rect 12000 21920 12400 21928
rect 8480 21832 8880 21840
rect 8480 21768 8488 21832
rect 8552 21768 8808 21832
rect 8872 21768 8880 21832
rect 8480 21760 8880 21768
rect 8960 21832 9360 21840
rect 8960 21768 8968 21832
rect 9032 21768 9288 21832
rect 9352 21768 9360 21832
rect 8960 21760 9360 21768
rect 9440 21832 11440 21840
rect 9440 21768 9448 21832
rect 9512 21768 9768 21832
rect 9832 21768 10088 21832
rect 10152 21768 10408 21832
rect 10472 21768 10728 21832
rect 10792 21768 11048 21832
rect 11112 21768 11368 21832
rect 11432 21768 11440 21832
rect 9440 21760 11440 21768
rect 11520 21832 11920 21840
rect 11520 21768 11528 21832
rect 11592 21768 11848 21832
rect 11912 21768 11920 21832
rect 11520 21760 11920 21768
rect 12000 21832 12400 21840
rect 12000 21768 12008 21832
rect 12072 21768 12328 21832
rect 12392 21768 12400 21832
rect 12000 21760 12400 21768
rect 8480 21672 8880 21680
rect 8480 21608 8488 21672
rect 8552 21608 8808 21672
rect 8872 21608 8880 21672
rect 8480 21600 8880 21608
rect 8960 21672 9360 21680
rect 8960 21608 8968 21672
rect 9032 21608 9288 21672
rect 9352 21608 9360 21672
rect 8960 21600 9360 21608
rect 9440 21672 11440 21680
rect 9440 21608 9448 21672
rect 9512 21608 9768 21672
rect 9832 21608 10088 21672
rect 10152 21608 10408 21672
rect 10472 21608 10728 21672
rect 10792 21608 11048 21672
rect 11112 21608 11368 21672
rect 11432 21608 11440 21672
rect 9440 21600 11440 21608
rect 11520 21672 11920 21680
rect 11520 21608 11528 21672
rect 11592 21608 11848 21672
rect 11912 21608 11920 21672
rect 11520 21600 11920 21608
rect 12000 21672 12400 21680
rect 12000 21608 12008 21672
rect 12072 21608 12328 21672
rect 12392 21608 12400 21672
rect 12000 21600 12400 21608
rect 8480 21512 8880 21520
rect 8480 21448 8488 21512
rect 8552 21448 8808 21512
rect 8872 21448 8880 21512
rect 8480 21440 8880 21448
rect 8960 21512 9360 21520
rect 8960 21448 8968 21512
rect 9032 21448 9288 21512
rect 9352 21448 9360 21512
rect 8960 21440 9360 21448
rect 9440 21512 11440 21520
rect 9440 21448 9448 21512
rect 9512 21448 9768 21512
rect 9832 21448 10088 21512
rect 10152 21448 10408 21512
rect 10472 21448 10728 21512
rect 10792 21448 11048 21512
rect 11112 21448 11368 21512
rect 11432 21448 11440 21512
rect 9440 21440 11440 21448
rect 11520 21512 11920 21520
rect 11520 21448 11528 21512
rect 11592 21448 11848 21512
rect 11912 21448 11920 21512
rect 11520 21440 11920 21448
rect 12000 21512 12400 21520
rect 12000 21448 12008 21512
rect 12072 21448 12328 21512
rect 12392 21448 12400 21512
rect 12000 21440 12400 21448
rect 8480 21352 8880 21360
rect 8480 21288 8488 21352
rect 8552 21288 8808 21352
rect 8872 21288 8880 21352
rect 8480 21280 8880 21288
rect 8960 21352 9360 21360
rect 8960 21288 8968 21352
rect 9032 21288 9288 21352
rect 9352 21288 9360 21352
rect 8960 21280 9360 21288
rect 9440 21352 11440 21360
rect 9440 21288 9448 21352
rect 9512 21288 9768 21352
rect 9832 21288 10088 21352
rect 10152 21288 10408 21352
rect 10472 21288 10728 21352
rect 10792 21288 11048 21352
rect 11112 21288 11368 21352
rect 11432 21288 11440 21352
rect 9440 21280 11440 21288
rect 11520 21352 11920 21360
rect 11520 21288 11528 21352
rect 11592 21288 11848 21352
rect 11912 21288 11920 21352
rect 11520 21280 11920 21288
rect 12000 21352 12400 21360
rect 12000 21288 12008 21352
rect 12072 21288 12328 21352
rect 12392 21288 12400 21352
rect 12000 21280 12400 21288
rect 8480 21192 8880 21200
rect 8480 21128 8488 21192
rect 8552 21128 8808 21192
rect 8872 21128 8880 21192
rect 8480 21120 8880 21128
rect 8960 21192 9360 21200
rect 8960 21128 8968 21192
rect 9032 21128 9288 21192
rect 9352 21128 9360 21192
rect 8960 21120 9360 21128
rect 9440 21192 11440 21200
rect 9440 21128 9448 21192
rect 9512 21128 9768 21192
rect 9832 21128 10088 21192
rect 10152 21128 10408 21192
rect 10472 21128 10728 21192
rect 10792 21128 11048 21192
rect 11112 21128 11368 21192
rect 11432 21128 11440 21192
rect 9440 21120 11440 21128
rect 11520 21192 11920 21200
rect 11520 21128 11528 21192
rect 11592 21128 11848 21192
rect 11912 21128 11920 21192
rect 11520 21120 11920 21128
rect 12000 21192 12400 21200
rect 12000 21128 12008 21192
rect 12072 21128 12328 21192
rect 12392 21128 12400 21192
rect 12000 21120 12400 21128
rect 8480 21032 8880 21040
rect 8480 20968 8488 21032
rect 8552 20968 8808 21032
rect 8872 20968 8880 21032
rect 8480 20960 8880 20968
rect 8960 21032 9360 21040
rect 8960 20968 8968 21032
rect 9032 20968 9288 21032
rect 9352 20968 9360 21032
rect 8960 20960 9360 20968
rect 9440 21032 11440 21040
rect 9440 20968 9448 21032
rect 9512 20968 9768 21032
rect 9832 20968 10088 21032
rect 10152 20968 10408 21032
rect 10472 20968 10728 21032
rect 10792 20968 11048 21032
rect 11112 20968 11368 21032
rect 11432 20968 11440 21032
rect 9440 20960 11440 20968
rect 11520 21032 11920 21040
rect 11520 20968 11528 21032
rect 11592 20968 11848 21032
rect 11912 20968 11920 21032
rect 11520 20960 11920 20968
rect 12000 21032 12400 21040
rect 12000 20968 12008 21032
rect 12072 20968 12328 21032
rect 12392 20968 12400 21032
rect 12000 20960 12400 20968
rect 8480 20872 8880 20880
rect 8480 20808 8488 20872
rect 8552 20808 8808 20872
rect 8872 20808 8880 20872
rect 8480 20800 8880 20808
rect 8960 20872 9360 20880
rect 8960 20808 8968 20872
rect 9032 20808 9288 20872
rect 9352 20808 9360 20872
rect 8960 20800 9360 20808
rect 9440 20872 11440 20880
rect 9440 20808 9448 20872
rect 9512 20808 9768 20872
rect 9832 20808 10088 20872
rect 10152 20808 10408 20872
rect 10472 20808 10728 20872
rect 10792 20808 11048 20872
rect 11112 20808 11368 20872
rect 11432 20808 11440 20872
rect 9440 20800 11440 20808
rect 11520 20872 11920 20880
rect 11520 20808 11528 20872
rect 11592 20808 11848 20872
rect 11912 20808 11920 20872
rect 11520 20800 11920 20808
rect 12000 20872 12400 20880
rect 12000 20808 12008 20872
rect 12072 20808 12328 20872
rect 12392 20808 12400 20872
rect 12000 20800 12400 20808
rect 8480 20712 8880 20720
rect 8480 20648 8488 20712
rect 8552 20648 8808 20712
rect 8872 20648 8880 20712
rect 8480 20640 8880 20648
rect 8960 20712 9360 20720
rect 8960 20648 8968 20712
rect 9032 20648 9288 20712
rect 9352 20648 9360 20712
rect 8960 20640 9360 20648
rect 9440 20712 11440 20720
rect 9440 20648 9448 20712
rect 9512 20648 9768 20712
rect 9832 20648 10088 20712
rect 10152 20648 10408 20712
rect 10472 20648 10728 20712
rect 10792 20648 11048 20712
rect 11112 20648 11368 20712
rect 11432 20648 11440 20712
rect 9440 20640 11440 20648
rect 11520 20712 11920 20720
rect 11520 20648 11528 20712
rect 11592 20648 11848 20712
rect 11912 20648 11920 20712
rect 11520 20640 11920 20648
rect 12000 20712 12400 20720
rect 12000 20648 12008 20712
rect 12072 20648 12328 20712
rect 12392 20648 12400 20712
rect 12000 20640 12400 20648
rect 8480 20552 8880 20560
rect 8480 20488 8488 20552
rect 8552 20488 8808 20552
rect 8872 20488 8880 20552
rect 8480 20480 8880 20488
rect 8960 20552 9360 20560
rect 8960 20488 8968 20552
rect 9032 20488 9288 20552
rect 9352 20488 9360 20552
rect 8960 20480 9360 20488
rect 9440 20552 11440 20560
rect 9440 20488 9448 20552
rect 9512 20488 9768 20552
rect 9832 20488 10088 20552
rect 10152 20488 10408 20552
rect 10472 20488 10728 20552
rect 10792 20488 11048 20552
rect 11112 20488 11368 20552
rect 11432 20488 11440 20552
rect 9440 20480 11440 20488
rect 11520 20552 11920 20560
rect 11520 20488 11528 20552
rect 11592 20488 11848 20552
rect 11912 20488 11920 20552
rect 11520 20480 11920 20488
rect 12000 20552 12400 20560
rect 12000 20488 12008 20552
rect 12072 20488 12328 20552
rect 12392 20488 12400 20552
rect 12000 20480 12400 20488
rect 8480 20392 8880 20400
rect 8480 20328 8488 20392
rect 8552 20328 8808 20392
rect 8872 20328 8880 20392
rect 8480 20320 8880 20328
rect 8960 20392 9360 20400
rect 8960 20328 8968 20392
rect 9032 20328 9288 20392
rect 9352 20328 9360 20392
rect 8960 20320 9360 20328
rect 9440 20392 11440 20400
rect 9440 20328 9448 20392
rect 9512 20328 9768 20392
rect 9832 20328 10088 20392
rect 10152 20328 10408 20392
rect 10472 20328 10728 20392
rect 10792 20328 11048 20392
rect 11112 20328 11368 20392
rect 11432 20328 11440 20392
rect 9440 20320 11440 20328
rect 11520 20392 11920 20400
rect 11520 20328 11528 20392
rect 11592 20328 11848 20392
rect 11912 20328 11920 20392
rect 11520 20320 11920 20328
rect 12000 20392 12400 20400
rect 12000 20328 12008 20392
rect 12072 20328 12328 20392
rect 12392 20328 12400 20392
rect 12000 20320 12400 20328
rect 8480 20232 8880 20240
rect 8480 20168 8488 20232
rect 8552 20168 8808 20232
rect 8872 20168 8880 20232
rect 8480 20160 8880 20168
rect 8960 20232 9360 20240
rect 8960 20168 8968 20232
rect 9032 20168 9288 20232
rect 9352 20168 9360 20232
rect 8960 20160 9360 20168
rect 9440 20232 11440 20240
rect 9440 20168 9448 20232
rect 9512 20168 9768 20232
rect 9832 20168 10088 20232
rect 10152 20168 10408 20232
rect 10472 20168 10728 20232
rect 10792 20168 11048 20232
rect 11112 20168 11368 20232
rect 11432 20168 11440 20232
rect 9440 20160 11440 20168
rect 11520 20232 11920 20240
rect 11520 20168 11528 20232
rect 11592 20168 11848 20232
rect 11912 20168 11920 20232
rect 11520 20160 11920 20168
rect 12000 20232 12400 20240
rect 12000 20168 12008 20232
rect 12072 20168 12328 20232
rect 12392 20168 12400 20232
rect 12000 20160 12400 20168
rect 8480 20072 8880 20080
rect 8480 20008 8488 20072
rect 8552 20008 8808 20072
rect 8872 20008 8880 20072
rect 8480 20000 8880 20008
rect 8960 20072 9360 20080
rect 8960 20008 8968 20072
rect 9032 20008 9288 20072
rect 9352 20008 9360 20072
rect 8960 20000 9360 20008
rect 9440 20072 11440 20080
rect 9440 20008 9448 20072
rect 9512 20008 9768 20072
rect 9832 20008 10088 20072
rect 10152 20008 10408 20072
rect 10472 20008 10728 20072
rect 10792 20008 11048 20072
rect 11112 20008 11368 20072
rect 11432 20008 11440 20072
rect 9440 20000 11440 20008
rect 11520 20072 11920 20080
rect 11520 20008 11528 20072
rect 11592 20008 11848 20072
rect 11912 20008 11920 20072
rect 11520 20000 11920 20008
rect 12000 20072 12400 20080
rect 12000 20008 12008 20072
rect 12072 20008 12328 20072
rect 12392 20008 12400 20072
rect 12000 20000 12400 20008
rect 8480 19912 8880 19920
rect 8480 19848 8488 19912
rect 8552 19848 8808 19912
rect 8872 19848 8880 19912
rect 8480 19840 8880 19848
rect 8960 19912 9360 19920
rect 8960 19848 8968 19912
rect 9032 19848 9288 19912
rect 9352 19848 9360 19912
rect 8960 19840 9360 19848
rect 9440 19912 11440 19920
rect 9440 19848 9448 19912
rect 9512 19848 9768 19912
rect 9832 19848 10088 19912
rect 10152 19848 10408 19912
rect 10472 19848 10728 19912
rect 10792 19848 11048 19912
rect 11112 19848 11368 19912
rect 11432 19848 11440 19912
rect 9440 19840 11440 19848
rect 11520 19912 11920 19920
rect 11520 19848 11528 19912
rect 11592 19848 11848 19912
rect 11912 19848 11920 19912
rect 11520 19840 11920 19848
rect 12000 19912 12400 19920
rect 12000 19848 12008 19912
rect 12072 19848 12328 19912
rect 12392 19848 12400 19912
rect 12000 19840 12400 19848
rect 8480 19752 8880 19760
rect 8480 19688 8488 19752
rect 8552 19688 8808 19752
rect 8872 19688 8880 19752
rect 8480 19680 8880 19688
rect 8960 19752 9360 19760
rect 8960 19688 8968 19752
rect 9032 19688 9288 19752
rect 9352 19688 9360 19752
rect 8960 19680 9360 19688
rect 9440 19752 11440 19760
rect 9440 19688 9448 19752
rect 9512 19688 9768 19752
rect 9832 19688 10088 19752
rect 10152 19688 10408 19752
rect 10472 19688 10728 19752
rect 10792 19688 11048 19752
rect 11112 19688 11368 19752
rect 11432 19688 11440 19752
rect 9440 19680 11440 19688
rect 11520 19752 11920 19760
rect 11520 19688 11528 19752
rect 11592 19688 11848 19752
rect 11912 19688 11920 19752
rect 11520 19680 11920 19688
rect 12000 19752 12400 19760
rect 12000 19688 12008 19752
rect 12072 19688 12328 19752
rect 12392 19688 12400 19752
rect 12000 19680 12400 19688
rect 8480 19592 8880 19600
rect 8480 19528 8488 19592
rect 8552 19528 8808 19592
rect 8872 19528 8880 19592
rect 8480 19520 8880 19528
rect 8960 19592 9360 19600
rect 8960 19528 8968 19592
rect 9032 19528 9288 19592
rect 9352 19528 9360 19592
rect 8960 19520 9360 19528
rect 9440 19592 11440 19600
rect 9440 19528 9448 19592
rect 9512 19528 9768 19592
rect 9832 19528 10088 19592
rect 10152 19528 10408 19592
rect 10472 19528 10728 19592
rect 10792 19528 11048 19592
rect 11112 19528 11368 19592
rect 11432 19528 11440 19592
rect 9440 19520 11440 19528
rect 11520 19592 11920 19600
rect 11520 19528 11528 19592
rect 11592 19528 11848 19592
rect 11912 19528 11920 19592
rect 11520 19520 11920 19528
rect 12000 19592 12400 19600
rect 12000 19528 12008 19592
rect 12072 19528 12328 19592
rect 12392 19528 12400 19592
rect 12000 19520 12400 19528
rect 8480 19432 8880 19440
rect 8480 19368 8488 19432
rect 8552 19368 8808 19432
rect 8872 19368 8880 19432
rect 8480 19360 8880 19368
rect 8960 19432 9360 19440
rect 8960 19368 8968 19432
rect 9032 19368 9288 19432
rect 9352 19368 9360 19432
rect 8960 19360 9360 19368
rect 9440 19432 11440 19440
rect 9440 19368 9448 19432
rect 9512 19368 9768 19432
rect 9832 19368 10088 19432
rect 10152 19368 10408 19432
rect 10472 19368 10728 19432
rect 10792 19368 11048 19432
rect 11112 19368 11368 19432
rect 11432 19368 11440 19432
rect 9440 19360 11440 19368
rect 11520 19432 11920 19440
rect 11520 19368 11528 19432
rect 11592 19368 11848 19432
rect 11912 19368 11920 19432
rect 11520 19360 11920 19368
rect 12000 19432 12400 19440
rect 12000 19368 12008 19432
rect 12072 19368 12328 19432
rect 12392 19368 12400 19432
rect 12000 19360 12400 19368
rect 8480 19272 8880 19280
rect 8480 19208 8488 19272
rect 8552 19208 8808 19272
rect 8872 19208 8880 19272
rect 8480 19200 8880 19208
rect 8960 19272 9360 19280
rect 8960 19208 8968 19272
rect 9032 19208 9288 19272
rect 9352 19208 9360 19272
rect 8960 19200 9360 19208
rect 9440 19272 11440 19280
rect 9440 19208 9448 19272
rect 9512 19208 9768 19272
rect 9832 19208 10088 19272
rect 10152 19208 10408 19272
rect 10472 19208 10728 19272
rect 10792 19208 11048 19272
rect 11112 19208 11368 19272
rect 11432 19208 11440 19272
rect 9440 19200 11440 19208
rect 11520 19272 11920 19280
rect 11520 19208 11528 19272
rect 11592 19208 11848 19272
rect 11912 19208 11920 19272
rect 11520 19200 11920 19208
rect 12000 19272 12400 19280
rect 12000 19208 12008 19272
rect 12072 19208 12328 19272
rect 12392 19208 12400 19272
rect 12000 19200 12400 19208
rect 8480 19112 8880 19120
rect 8480 19048 8488 19112
rect 8552 19048 8808 19112
rect 8872 19048 8880 19112
rect 8480 19040 8880 19048
rect 8960 19112 9360 19120
rect 8960 19048 8968 19112
rect 9032 19048 9288 19112
rect 9352 19048 9360 19112
rect 8960 19040 9360 19048
rect 9440 19112 11440 19120
rect 9440 19048 9448 19112
rect 9512 19048 9768 19112
rect 9832 19048 10088 19112
rect 10152 19048 10408 19112
rect 10472 19048 10728 19112
rect 10792 19048 11048 19112
rect 11112 19048 11368 19112
rect 11432 19048 11440 19112
rect 9440 19040 11440 19048
rect 11520 19112 11920 19120
rect 11520 19048 11528 19112
rect 11592 19048 11848 19112
rect 11912 19048 11920 19112
rect 11520 19040 11920 19048
rect 12000 19112 12400 19120
rect 12000 19048 12008 19112
rect 12072 19048 12328 19112
rect 12392 19048 12400 19112
rect 12000 19040 12400 19048
rect 8480 18952 8880 18960
rect 8480 18888 8488 18952
rect 8552 18888 8808 18952
rect 8872 18888 8880 18952
rect 8480 18880 8880 18888
rect 8960 18952 9360 18960
rect 8960 18888 8968 18952
rect 9032 18888 9288 18952
rect 9352 18888 9360 18952
rect 8960 18880 9360 18888
rect 9440 18952 11440 18960
rect 9440 18888 9448 18952
rect 9512 18888 9768 18952
rect 9832 18888 10088 18952
rect 10152 18888 10408 18952
rect 10472 18888 10728 18952
rect 10792 18888 11048 18952
rect 11112 18888 11368 18952
rect 11432 18888 11440 18952
rect 9440 18880 11440 18888
rect 11520 18952 11920 18960
rect 11520 18888 11528 18952
rect 11592 18888 11848 18952
rect 11912 18888 11920 18952
rect 11520 18880 11920 18888
rect 12000 18952 12400 18960
rect 12000 18888 12008 18952
rect 12072 18888 12328 18952
rect 12392 18888 12400 18952
rect 12000 18880 12400 18888
rect 8480 18792 8880 18800
rect 8480 18728 8488 18792
rect 8552 18728 8808 18792
rect 8872 18728 8880 18792
rect 8480 18720 8880 18728
rect 8960 18792 9360 18800
rect 8960 18728 8968 18792
rect 9032 18728 9288 18792
rect 9352 18728 9360 18792
rect 8960 18720 9360 18728
rect 9440 18792 11440 18800
rect 9440 18728 9448 18792
rect 9512 18728 9768 18792
rect 9832 18728 10088 18792
rect 10152 18728 10408 18792
rect 10472 18728 10728 18792
rect 10792 18728 11048 18792
rect 11112 18728 11368 18792
rect 11432 18728 11440 18792
rect 9440 18720 11440 18728
rect 11520 18792 11920 18800
rect 11520 18728 11528 18792
rect 11592 18728 11848 18792
rect 11912 18728 11920 18792
rect 11520 18720 11920 18728
rect 12000 18792 12400 18800
rect 12000 18728 12008 18792
rect 12072 18728 12328 18792
rect 12392 18728 12400 18792
rect 12000 18720 12400 18728
rect 8480 18632 8880 18640
rect 8480 18568 8488 18632
rect 8552 18568 8808 18632
rect 8872 18568 8880 18632
rect 8480 18560 8880 18568
rect 8960 18632 9360 18640
rect 8960 18568 8968 18632
rect 9032 18568 9288 18632
rect 9352 18568 9360 18632
rect 8960 18560 9360 18568
rect 9440 18632 11440 18640
rect 9440 18568 9448 18632
rect 9512 18568 9768 18632
rect 9832 18568 10088 18632
rect 10152 18568 10408 18632
rect 10472 18568 10728 18632
rect 10792 18568 11048 18632
rect 11112 18568 11368 18632
rect 11432 18568 11440 18632
rect 9440 18560 11440 18568
rect 11520 18632 11920 18640
rect 11520 18568 11528 18632
rect 11592 18568 11848 18632
rect 11912 18568 11920 18632
rect 11520 18560 11920 18568
rect 12000 18632 12400 18640
rect 12000 18568 12008 18632
rect 12072 18568 12328 18632
rect 12392 18568 12400 18632
rect 12000 18560 12400 18568
rect 8480 18472 8880 18480
rect 8480 18408 8488 18472
rect 8552 18408 8808 18472
rect 8872 18408 8880 18472
rect 8480 18400 8880 18408
rect 8960 18472 9360 18480
rect 8960 18408 8968 18472
rect 9032 18408 9288 18472
rect 9352 18408 9360 18472
rect 8960 18400 9360 18408
rect 9440 18472 11440 18480
rect 9440 18408 9448 18472
rect 9512 18408 9768 18472
rect 9832 18408 10088 18472
rect 10152 18408 10408 18472
rect 10472 18408 10728 18472
rect 10792 18408 11048 18472
rect 11112 18408 11368 18472
rect 11432 18408 11440 18472
rect 9440 18400 11440 18408
rect 11520 18472 11920 18480
rect 11520 18408 11528 18472
rect 11592 18408 11848 18472
rect 11912 18408 11920 18472
rect 11520 18400 11920 18408
rect 12000 18472 12400 18480
rect 12000 18408 12008 18472
rect 12072 18408 12328 18472
rect 12392 18408 12400 18472
rect 12000 18400 12400 18408
rect 8480 18312 8880 18320
rect 8480 18248 8488 18312
rect 8552 18248 8808 18312
rect 8872 18248 8880 18312
rect 8480 18240 8880 18248
rect 8960 18312 9360 18320
rect 8960 18248 8968 18312
rect 9032 18248 9288 18312
rect 9352 18248 9360 18312
rect 8960 18240 9360 18248
rect 9440 18312 11440 18320
rect 9440 18248 9448 18312
rect 9512 18248 9768 18312
rect 9832 18248 10088 18312
rect 10152 18248 10408 18312
rect 10472 18248 10728 18312
rect 10792 18248 11048 18312
rect 11112 18248 11368 18312
rect 11432 18248 11440 18312
rect 9440 18240 11440 18248
rect 11520 18312 11920 18320
rect 11520 18248 11528 18312
rect 11592 18248 11848 18312
rect 11912 18248 11920 18312
rect 11520 18240 11920 18248
rect 12000 18312 12400 18320
rect 12000 18248 12008 18312
rect 12072 18248 12328 18312
rect 12392 18248 12400 18312
rect 12000 18240 12400 18248
rect 8480 18152 8880 18160
rect 8480 18088 8488 18152
rect 8552 18088 8808 18152
rect 8872 18088 8880 18152
rect 8480 18080 8880 18088
rect 8960 18152 9360 18160
rect 8960 18088 8968 18152
rect 9032 18088 9288 18152
rect 9352 18088 9360 18152
rect 8960 18080 9360 18088
rect 9440 18152 11440 18160
rect 9440 18088 9448 18152
rect 9512 18088 9768 18152
rect 9832 18088 10088 18152
rect 10152 18088 10408 18152
rect 10472 18088 10728 18152
rect 10792 18088 11048 18152
rect 11112 18088 11368 18152
rect 11432 18088 11440 18152
rect 9440 18080 11440 18088
rect 11520 18152 11920 18160
rect 11520 18088 11528 18152
rect 11592 18088 11848 18152
rect 11912 18088 11920 18152
rect 11520 18080 11920 18088
rect 12000 18152 12400 18160
rect 12000 18088 12008 18152
rect 12072 18088 12328 18152
rect 12392 18088 12400 18152
rect 12000 18080 12400 18088
rect 8480 17992 8880 18000
rect 8480 17928 8488 17992
rect 8552 17928 8808 17992
rect 8872 17928 8880 17992
rect 8480 17920 8880 17928
rect 8960 17992 9360 18000
rect 8960 17928 8968 17992
rect 9032 17928 9288 17992
rect 9352 17928 9360 17992
rect 8960 17920 9360 17928
rect 9440 17992 11440 18000
rect 9440 17928 9448 17992
rect 9512 17928 9768 17992
rect 9832 17928 10088 17992
rect 10152 17928 10408 17992
rect 10472 17928 10728 17992
rect 10792 17928 11048 17992
rect 11112 17928 11368 17992
rect 11432 17928 11440 17992
rect 9440 17920 11440 17928
rect 11520 17992 11920 18000
rect 11520 17928 11528 17992
rect 11592 17928 11848 17992
rect 11912 17928 11920 17992
rect 11520 17920 11920 17928
rect 12000 17992 12400 18000
rect 12000 17928 12008 17992
rect 12072 17928 12328 17992
rect 12392 17928 12400 17992
rect 12000 17920 12400 17928
rect 8480 17832 8880 17840
rect 8480 17768 8488 17832
rect 8552 17768 8808 17832
rect 8872 17768 8880 17832
rect 8480 17760 8880 17768
rect 8960 17832 9360 17840
rect 8960 17768 8968 17832
rect 9032 17768 9288 17832
rect 9352 17768 9360 17832
rect 8960 17760 9360 17768
rect 9440 17832 11440 17840
rect 9440 17768 9448 17832
rect 9512 17768 9768 17832
rect 9832 17768 10088 17832
rect 10152 17768 10408 17832
rect 10472 17768 10728 17832
rect 10792 17768 11048 17832
rect 11112 17768 11368 17832
rect 11432 17768 11440 17832
rect 9440 17760 11440 17768
rect 11520 17832 11920 17840
rect 11520 17768 11528 17832
rect 11592 17768 11848 17832
rect 11912 17768 11920 17832
rect 11520 17760 11920 17768
rect 12000 17832 12400 17840
rect 12000 17768 12008 17832
rect 12072 17768 12328 17832
rect 12392 17768 12400 17832
rect 12000 17760 12400 17768
rect 8480 17672 8880 17680
rect 8480 17608 8488 17672
rect 8552 17608 8808 17672
rect 8872 17608 8880 17672
rect 8480 17600 8880 17608
rect 8960 17672 9360 17680
rect 8960 17608 8968 17672
rect 9032 17608 9288 17672
rect 9352 17608 9360 17672
rect 8960 17600 9360 17608
rect 9440 17672 11440 17680
rect 9440 17608 9448 17672
rect 9512 17608 9768 17672
rect 9832 17608 10088 17672
rect 10152 17608 10408 17672
rect 10472 17608 10728 17672
rect 10792 17608 11048 17672
rect 11112 17608 11368 17672
rect 11432 17608 11440 17672
rect 9440 17600 11440 17608
rect 11520 17672 11920 17680
rect 11520 17608 11528 17672
rect 11592 17608 11848 17672
rect 11912 17608 11920 17672
rect 11520 17600 11920 17608
rect 12000 17672 12400 17680
rect 12000 17608 12008 17672
rect 12072 17608 12328 17672
rect 12392 17608 12400 17672
rect 12000 17600 12400 17608
rect 8480 17512 8880 17520
rect 8480 17448 8488 17512
rect 8552 17448 8808 17512
rect 8872 17448 8880 17512
rect 8480 17440 8880 17448
rect 8960 17512 9360 17520
rect 8960 17448 8968 17512
rect 9032 17448 9288 17512
rect 9352 17448 9360 17512
rect 8960 17440 9360 17448
rect 9440 17512 11440 17520
rect 9440 17448 9448 17512
rect 9512 17448 9768 17512
rect 9832 17448 10088 17512
rect 10152 17448 10408 17512
rect 10472 17448 10728 17512
rect 10792 17448 11048 17512
rect 11112 17448 11368 17512
rect 11432 17448 11440 17512
rect 9440 17440 11440 17448
rect 11520 17512 11920 17520
rect 11520 17448 11528 17512
rect 11592 17448 11848 17512
rect 11912 17448 11920 17512
rect 11520 17440 11920 17448
rect 12000 17512 12400 17520
rect 12000 17448 12008 17512
rect 12072 17448 12328 17512
rect 12392 17448 12400 17512
rect 12000 17440 12400 17448
rect 8480 17352 8880 17360
rect 8480 17288 8488 17352
rect 8552 17288 8808 17352
rect 8872 17288 8880 17352
rect 8480 17280 8880 17288
rect 8960 17352 9360 17360
rect 8960 17288 8968 17352
rect 9032 17288 9288 17352
rect 9352 17288 9360 17352
rect 8960 17280 9360 17288
rect 9440 17352 11440 17360
rect 9440 17288 9448 17352
rect 9512 17288 9768 17352
rect 9832 17288 10088 17352
rect 10152 17288 10408 17352
rect 10472 17288 10728 17352
rect 10792 17288 11048 17352
rect 11112 17288 11368 17352
rect 11432 17288 11440 17352
rect 9440 17280 11440 17288
rect 11520 17352 11920 17360
rect 11520 17288 11528 17352
rect 11592 17288 11848 17352
rect 11912 17288 11920 17352
rect 11520 17280 11920 17288
rect 12000 17352 12400 17360
rect 12000 17288 12008 17352
rect 12072 17288 12328 17352
rect 12392 17288 12400 17352
rect 12000 17280 12400 17288
rect 8480 17192 8880 17200
rect 8480 17128 8488 17192
rect 8552 17128 8808 17192
rect 8872 17128 8880 17192
rect 8480 17120 8880 17128
rect 8960 17192 9360 17200
rect 8960 17128 8968 17192
rect 9032 17128 9288 17192
rect 9352 17128 9360 17192
rect 8960 17120 9360 17128
rect 9440 17192 11440 17200
rect 9440 17128 9448 17192
rect 9512 17128 9768 17192
rect 9832 17128 10088 17192
rect 10152 17128 10408 17192
rect 10472 17128 10728 17192
rect 10792 17128 11048 17192
rect 11112 17128 11368 17192
rect 11432 17128 11440 17192
rect 9440 17120 11440 17128
rect 11520 17192 11920 17200
rect 11520 17128 11528 17192
rect 11592 17128 11848 17192
rect 11912 17128 11920 17192
rect 11520 17120 11920 17128
rect 12000 17192 12400 17200
rect 12000 17128 12008 17192
rect 12072 17128 12328 17192
rect 12392 17128 12400 17192
rect 12000 17120 12400 17128
rect 8480 17032 8880 17040
rect 8480 16968 8488 17032
rect 8552 16968 8808 17032
rect 8872 16968 8880 17032
rect 8480 16960 8880 16968
rect 8960 17032 9360 17040
rect 8960 16968 8968 17032
rect 9032 16968 9288 17032
rect 9352 16968 9360 17032
rect 8960 16960 9360 16968
rect 9440 17032 11440 17040
rect 9440 16968 9448 17032
rect 9512 16968 9768 17032
rect 9832 16968 10088 17032
rect 10152 16968 10408 17032
rect 10472 16968 10728 17032
rect 10792 16968 11048 17032
rect 11112 16968 11368 17032
rect 11432 16968 11440 17032
rect 9440 16960 11440 16968
rect 11520 17032 11920 17040
rect 11520 16968 11528 17032
rect 11592 16968 11848 17032
rect 11912 16968 11920 17032
rect 11520 16960 11920 16968
rect 12000 17032 12400 17040
rect 12000 16968 12008 17032
rect 12072 16968 12328 17032
rect 12392 16968 12400 17032
rect 12000 16960 12400 16968
rect 8480 16872 8880 16880
rect 8480 16808 8488 16872
rect 8552 16808 8808 16872
rect 8872 16808 8880 16872
rect 8480 16800 8880 16808
rect 8960 16872 9360 16880
rect 8960 16808 8968 16872
rect 9032 16808 9288 16872
rect 9352 16808 9360 16872
rect 8960 16800 9360 16808
rect 9440 16872 11440 16880
rect 9440 16808 9448 16872
rect 9512 16808 9768 16872
rect 9832 16808 10088 16872
rect 10152 16808 10408 16872
rect 10472 16808 10728 16872
rect 10792 16808 11048 16872
rect 11112 16808 11368 16872
rect 11432 16808 11440 16872
rect 9440 16800 11440 16808
rect 11520 16872 11920 16880
rect 11520 16808 11528 16872
rect 11592 16808 11848 16872
rect 11912 16808 11920 16872
rect 11520 16800 11920 16808
rect 12000 16872 12400 16880
rect 12000 16808 12008 16872
rect 12072 16808 12328 16872
rect 12392 16808 12400 16872
rect 12000 16800 12400 16808
rect 8480 16712 8880 16720
rect 8480 16648 8488 16712
rect 8552 16648 8808 16712
rect 8872 16648 8880 16712
rect 8480 16640 8880 16648
rect 8960 16712 9360 16720
rect 8960 16648 8968 16712
rect 9032 16648 9288 16712
rect 9352 16648 9360 16712
rect 8960 16640 9360 16648
rect 9440 16712 11440 16720
rect 9440 16648 9448 16712
rect 9512 16648 9768 16712
rect 9832 16648 10088 16712
rect 10152 16648 10408 16712
rect 10472 16648 10728 16712
rect 10792 16648 11048 16712
rect 11112 16648 11368 16712
rect 11432 16648 11440 16712
rect 9440 16640 11440 16648
rect 11520 16712 11920 16720
rect 11520 16648 11528 16712
rect 11592 16648 11848 16712
rect 11912 16648 11920 16712
rect 11520 16640 11920 16648
rect 12000 16712 12400 16720
rect 12000 16648 12008 16712
rect 12072 16648 12328 16712
rect 12392 16648 12400 16712
rect 12000 16640 12400 16648
rect 8480 16552 8880 16560
rect 8480 16488 8488 16552
rect 8552 16488 8808 16552
rect 8872 16488 8880 16552
rect 8480 16480 8880 16488
rect 8960 16552 9360 16560
rect 8960 16488 8968 16552
rect 9032 16488 9288 16552
rect 9352 16488 9360 16552
rect 8960 16480 9360 16488
rect 9440 16552 11440 16560
rect 9440 16488 9448 16552
rect 9512 16488 9768 16552
rect 9832 16488 10088 16552
rect 10152 16488 10408 16552
rect 10472 16488 10728 16552
rect 10792 16488 11048 16552
rect 11112 16488 11368 16552
rect 11432 16488 11440 16552
rect 9440 16480 11440 16488
rect 11520 16552 11920 16560
rect 11520 16488 11528 16552
rect 11592 16488 11848 16552
rect 11912 16488 11920 16552
rect 11520 16480 11920 16488
rect 12000 16552 12400 16560
rect 12000 16488 12008 16552
rect 12072 16488 12328 16552
rect 12392 16488 12400 16552
rect 12000 16480 12400 16488
rect 8480 16392 8880 16400
rect 8480 16328 8488 16392
rect 8552 16328 8808 16392
rect 8872 16328 8880 16392
rect 8480 16320 8880 16328
rect 8960 16392 9360 16400
rect 8960 16328 8968 16392
rect 9032 16328 9288 16392
rect 9352 16328 9360 16392
rect 8960 16320 9360 16328
rect 9440 16392 11440 16400
rect 9440 16328 9448 16392
rect 9512 16328 9768 16392
rect 9832 16328 10088 16392
rect 10152 16328 10408 16392
rect 10472 16328 10728 16392
rect 10792 16328 11048 16392
rect 11112 16328 11368 16392
rect 11432 16328 11440 16392
rect 9440 16320 11440 16328
rect 11520 16392 11920 16400
rect 11520 16328 11528 16392
rect 11592 16328 11848 16392
rect 11912 16328 11920 16392
rect 11520 16320 11920 16328
rect 12000 16392 12400 16400
rect 12000 16328 12008 16392
rect 12072 16328 12328 16392
rect 12392 16328 12400 16392
rect 12000 16320 12400 16328
rect 8480 16232 8880 16240
rect 8480 16168 8488 16232
rect 8552 16168 8808 16232
rect 8872 16168 8880 16232
rect 8480 16160 8880 16168
rect 8960 16232 9360 16240
rect 8960 16168 8968 16232
rect 9032 16168 9288 16232
rect 9352 16168 9360 16232
rect 8960 16160 9360 16168
rect 9440 16232 11440 16240
rect 9440 16168 9448 16232
rect 9512 16168 9768 16232
rect 9832 16168 10088 16232
rect 10152 16168 10408 16232
rect 10472 16168 10728 16232
rect 10792 16168 11048 16232
rect 11112 16168 11368 16232
rect 11432 16168 11440 16232
rect 9440 16160 11440 16168
rect 11520 16232 11920 16240
rect 11520 16168 11528 16232
rect 11592 16168 11848 16232
rect 11912 16168 11920 16232
rect 11520 16160 11920 16168
rect 12000 16232 12400 16240
rect 12000 16168 12008 16232
rect 12072 16168 12328 16232
rect 12392 16168 12400 16232
rect 12000 16160 12400 16168
rect 8480 16072 8880 16080
rect 8480 16008 8488 16072
rect 8552 16008 8808 16072
rect 8872 16008 8880 16072
rect 8480 16000 8880 16008
rect 8960 16072 9360 16080
rect 8960 16008 8968 16072
rect 9032 16008 9288 16072
rect 9352 16008 9360 16072
rect 8960 16000 9360 16008
rect 9440 16072 11440 16080
rect 9440 16008 9448 16072
rect 9512 16008 9768 16072
rect 9832 16008 10088 16072
rect 10152 16008 10408 16072
rect 10472 16008 10728 16072
rect 10792 16008 11048 16072
rect 11112 16008 11368 16072
rect 11432 16008 11440 16072
rect 9440 16000 11440 16008
rect 11520 16072 11920 16080
rect 11520 16008 11528 16072
rect 11592 16008 11848 16072
rect 11912 16008 11920 16072
rect 11520 16000 11920 16008
rect 12000 16072 12400 16080
rect 12000 16008 12008 16072
rect 12072 16008 12328 16072
rect 12392 16008 12400 16072
rect 12000 16000 12400 16008
rect 8480 15912 8880 15920
rect 8480 15848 8488 15912
rect 8552 15848 8808 15912
rect 8872 15848 8880 15912
rect 8480 15840 8880 15848
rect 8960 15912 9360 15920
rect 8960 15848 8968 15912
rect 9032 15848 9288 15912
rect 9352 15848 9360 15912
rect 8960 15840 9360 15848
rect 9440 15912 11440 15920
rect 9440 15848 9448 15912
rect 9512 15848 9768 15912
rect 9832 15848 10088 15912
rect 10152 15848 10408 15912
rect 10472 15848 10728 15912
rect 10792 15848 11048 15912
rect 11112 15848 11368 15912
rect 11432 15848 11440 15912
rect 9440 15840 11440 15848
rect 11520 15912 11920 15920
rect 11520 15848 11528 15912
rect 11592 15848 11848 15912
rect 11912 15848 11920 15912
rect 11520 15840 11920 15848
rect 12000 15912 12400 15920
rect 12000 15848 12008 15912
rect 12072 15848 12328 15912
rect 12392 15848 12400 15912
rect 12000 15840 12400 15848
rect 8480 15752 8880 15760
rect 8480 15688 8488 15752
rect 8552 15688 8808 15752
rect 8872 15688 8880 15752
rect 8480 15680 8880 15688
rect 8960 15752 9360 15760
rect 8960 15688 8968 15752
rect 9032 15688 9288 15752
rect 9352 15688 9360 15752
rect 8960 15680 9360 15688
rect 9440 15752 11440 15760
rect 9440 15688 9448 15752
rect 9512 15688 9768 15752
rect 9832 15688 10088 15752
rect 10152 15688 10408 15752
rect 10472 15688 10728 15752
rect 10792 15688 11048 15752
rect 11112 15688 11368 15752
rect 11432 15688 11440 15752
rect 9440 15680 11440 15688
rect 11520 15752 11920 15760
rect 11520 15688 11528 15752
rect 11592 15688 11848 15752
rect 11912 15688 11920 15752
rect 11520 15680 11920 15688
rect 12000 15752 12400 15760
rect 12000 15688 12008 15752
rect 12072 15688 12328 15752
rect 12392 15688 12400 15752
rect 12000 15680 12400 15688
rect 8480 15592 8880 15600
rect 8480 15528 8488 15592
rect 8552 15528 8808 15592
rect 8872 15528 8880 15592
rect 8480 15520 8880 15528
rect 8960 15592 9360 15600
rect 8960 15528 8968 15592
rect 9032 15528 9288 15592
rect 9352 15528 9360 15592
rect 8960 15520 9360 15528
rect 9440 15592 11440 15600
rect 9440 15528 9448 15592
rect 9512 15528 9768 15592
rect 9832 15528 10088 15592
rect 10152 15528 10408 15592
rect 10472 15528 10728 15592
rect 10792 15528 11048 15592
rect 11112 15528 11368 15592
rect 11432 15528 11440 15592
rect 9440 15520 11440 15528
rect 11520 15592 11920 15600
rect 11520 15528 11528 15592
rect 11592 15528 11848 15592
rect 11912 15528 11920 15592
rect 11520 15520 11920 15528
rect 12000 15592 12400 15600
rect 12000 15528 12008 15592
rect 12072 15528 12328 15592
rect 12392 15528 12400 15592
rect 12000 15520 12400 15528
rect 8480 15432 8880 15440
rect 8480 15368 8488 15432
rect 8552 15368 8808 15432
rect 8872 15368 8880 15432
rect 8480 15360 8880 15368
rect 8960 15432 9360 15440
rect 8960 15368 8968 15432
rect 9032 15368 9288 15432
rect 9352 15368 9360 15432
rect 8960 15360 9360 15368
rect 9440 15432 11440 15440
rect 9440 15368 9448 15432
rect 9512 15368 9768 15432
rect 9832 15368 10088 15432
rect 10152 15368 10408 15432
rect 10472 15368 10728 15432
rect 10792 15368 11048 15432
rect 11112 15368 11368 15432
rect 11432 15368 11440 15432
rect 9440 15360 11440 15368
rect 11520 15432 11920 15440
rect 11520 15368 11528 15432
rect 11592 15368 11848 15432
rect 11912 15368 11920 15432
rect 11520 15360 11920 15368
rect 12000 15432 12400 15440
rect 12000 15368 12008 15432
rect 12072 15368 12328 15432
rect 12392 15368 12400 15432
rect 12000 15360 12400 15368
rect 8480 15272 8880 15280
rect 8480 15208 8488 15272
rect 8552 15208 8808 15272
rect 8872 15208 8880 15272
rect 8480 15200 8880 15208
rect 8960 15272 9360 15280
rect 8960 15208 8968 15272
rect 9032 15208 9288 15272
rect 9352 15208 9360 15272
rect 8960 15200 9360 15208
rect 9440 15272 11440 15280
rect 9440 15208 9448 15272
rect 9512 15208 9768 15272
rect 9832 15208 10088 15272
rect 10152 15208 10408 15272
rect 10472 15208 10728 15272
rect 10792 15208 11048 15272
rect 11112 15208 11368 15272
rect 11432 15208 11440 15272
rect 9440 15200 11440 15208
rect 11520 15272 11920 15280
rect 11520 15208 11528 15272
rect 11592 15208 11848 15272
rect 11912 15208 11920 15272
rect 11520 15200 11920 15208
rect 12000 15272 12400 15280
rect 12000 15208 12008 15272
rect 12072 15208 12328 15272
rect 12392 15208 12400 15272
rect 12000 15200 12400 15208
rect 8480 15112 8880 15120
rect 8480 15048 8488 15112
rect 8552 15048 8808 15112
rect 8872 15048 8880 15112
rect 8480 15040 8880 15048
rect 8960 15112 9360 15120
rect 8960 15048 8968 15112
rect 9032 15048 9288 15112
rect 9352 15048 9360 15112
rect 8960 15040 9360 15048
rect 9440 15112 11440 15120
rect 9440 15048 9448 15112
rect 9512 15048 9768 15112
rect 9832 15048 10088 15112
rect 10152 15048 10408 15112
rect 10472 15048 10728 15112
rect 10792 15048 11048 15112
rect 11112 15048 11368 15112
rect 11432 15048 11440 15112
rect 9440 15040 11440 15048
rect 11520 15112 11920 15120
rect 11520 15048 11528 15112
rect 11592 15048 11848 15112
rect 11912 15048 11920 15112
rect 11520 15040 11920 15048
rect 12000 15112 12400 15120
rect 12000 15048 12008 15112
rect 12072 15048 12328 15112
rect 12392 15048 12400 15112
rect 12000 15040 12400 15048
rect 8480 14952 8880 14960
rect 8480 14888 8488 14952
rect 8552 14888 8808 14952
rect 8872 14888 8880 14952
rect 8480 14880 8880 14888
rect 8960 14952 9360 14960
rect 8960 14888 8968 14952
rect 9032 14888 9288 14952
rect 9352 14888 9360 14952
rect 8960 14880 9360 14888
rect 9440 14952 11440 14960
rect 9440 14888 9448 14952
rect 9512 14888 9768 14952
rect 9832 14888 10088 14952
rect 10152 14888 10408 14952
rect 10472 14888 10728 14952
rect 10792 14888 11048 14952
rect 11112 14888 11368 14952
rect 11432 14888 11440 14952
rect 9440 14880 11440 14888
rect 11520 14952 11920 14960
rect 11520 14888 11528 14952
rect 11592 14888 11848 14952
rect 11912 14888 11920 14952
rect 11520 14880 11920 14888
rect 12000 14952 12400 14960
rect 12000 14888 12008 14952
rect 12072 14888 12328 14952
rect 12392 14888 12400 14952
rect 12000 14880 12400 14888
rect 8480 14792 8880 14800
rect 8480 14728 8488 14792
rect 8552 14728 8808 14792
rect 8872 14728 8880 14792
rect 8480 14720 8880 14728
rect 8960 14792 9360 14800
rect 8960 14728 8968 14792
rect 9032 14728 9288 14792
rect 9352 14728 9360 14792
rect 8960 14720 9360 14728
rect 9440 14792 11440 14800
rect 9440 14728 9448 14792
rect 9512 14728 9768 14792
rect 9832 14728 10088 14792
rect 10152 14728 10408 14792
rect 10472 14728 10728 14792
rect 10792 14728 11048 14792
rect 11112 14728 11368 14792
rect 11432 14728 11440 14792
rect 9440 14720 11440 14728
rect 11520 14792 11920 14800
rect 11520 14728 11528 14792
rect 11592 14728 11848 14792
rect 11912 14728 11920 14792
rect 11520 14720 11920 14728
rect 12000 14792 12400 14800
rect 12000 14728 12008 14792
rect 12072 14728 12328 14792
rect 12392 14728 12400 14792
rect 12000 14720 12400 14728
rect 8480 14632 8880 14640
rect 8480 14568 8488 14632
rect 8552 14568 8808 14632
rect 8872 14568 8880 14632
rect 8480 14560 8880 14568
rect 8960 14632 9360 14640
rect 8960 14568 8968 14632
rect 9032 14568 9288 14632
rect 9352 14568 9360 14632
rect 8960 14560 9360 14568
rect 9440 14632 11440 14640
rect 9440 14568 9448 14632
rect 9512 14568 9768 14632
rect 9832 14568 10088 14632
rect 10152 14568 10408 14632
rect 10472 14568 10728 14632
rect 10792 14568 11048 14632
rect 11112 14568 11368 14632
rect 11432 14568 11440 14632
rect 9440 14560 11440 14568
rect 11520 14632 11920 14640
rect 11520 14568 11528 14632
rect 11592 14568 11848 14632
rect 11912 14568 11920 14632
rect 11520 14560 11920 14568
rect 12000 14632 12400 14640
rect 12000 14568 12008 14632
rect 12072 14568 12328 14632
rect 12392 14568 12400 14632
rect 12000 14560 12400 14568
rect 8480 14472 8880 14480
rect 8480 14408 8488 14472
rect 8552 14408 8808 14472
rect 8872 14408 8880 14472
rect 8480 14400 8880 14408
rect 8960 14472 9360 14480
rect 8960 14408 8968 14472
rect 9032 14408 9288 14472
rect 9352 14408 9360 14472
rect 8960 14400 9360 14408
rect 9440 14472 11440 14480
rect 9440 14408 9448 14472
rect 9512 14408 9768 14472
rect 9832 14408 10088 14472
rect 10152 14408 10408 14472
rect 10472 14408 10728 14472
rect 10792 14408 11048 14472
rect 11112 14408 11368 14472
rect 11432 14408 11440 14472
rect 9440 14400 11440 14408
rect 11520 14472 11920 14480
rect 11520 14408 11528 14472
rect 11592 14408 11848 14472
rect 11912 14408 11920 14472
rect 11520 14400 11920 14408
rect 12000 14472 12400 14480
rect 12000 14408 12008 14472
rect 12072 14408 12328 14472
rect 12392 14408 12400 14472
rect 12000 14400 12400 14408
rect 8480 14312 8880 14320
rect 8480 14248 8488 14312
rect 8552 14248 8808 14312
rect 8872 14248 8880 14312
rect 8480 14240 8880 14248
rect 8960 14312 9360 14320
rect 8960 14248 8968 14312
rect 9032 14248 9288 14312
rect 9352 14248 9360 14312
rect 8960 14240 9360 14248
rect 9440 14312 11440 14320
rect 9440 14248 9448 14312
rect 9512 14248 9768 14312
rect 9832 14248 10088 14312
rect 10152 14248 10408 14312
rect 10472 14248 10728 14312
rect 10792 14248 11048 14312
rect 11112 14248 11368 14312
rect 11432 14248 11440 14312
rect 9440 14240 11440 14248
rect 11520 14312 11920 14320
rect 11520 14248 11528 14312
rect 11592 14248 11848 14312
rect 11912 14248 11920 14312
rect 11520 14240 11920 14248
rect 12000 14312 12400 14320
rect 12000 14248 12008 14312
rect 12072 14248 12328 14312
rect 12392 14248 12400 14312
rect 12000 14240 12400 14248
rect 8480 14152 8880 14160
rect 8480 14088 8488 14152
rect 8552 14088 8808 14152
rect 8872 14088 8880 14152
rect 8480 14080 8880 14088
rect 8960 14152 9360 14160
rect 8960 14088 8968 14152
rect 9032 14088 9288 14152
rect 9352 14088 9360 14152
rect 8960 14080 9360 14088
rect 9440 14152 11440 14160
rect 9440 14088 9448 14152
rect 9512 14088 9768 14152
rect 9832 14088 10088 14152
rect 10152 14088 10408 14152
rect 10472 14088 10728 14152
rect 10792 14088 11048 14152
rect 11112 14088 11368 14152
rect 11432 14088 11440 14152
rect 9440 14080 11440 14088
rect 11520 14152 11920 14160
rect 11520 14088 11528 14152
rect 11592 14088 11848 14152
rect 11912 14088 11920 14152
rect 11520 14080 11920 14088
rect 12000 14152 12400 14160
rect 12000 14088 12008 14152
rect 12072 14088 12328 14152
rect 12392 14088 12400 14152
rect 12000 14080 12400 14088
rect 8480 13992 8880 14000
rect 8480 13928 8488 13992
rect 8552 13928 8808 13992
rect 8872 13928 8880 13992
rect 8480 13920 8880 13928
rect 8960 13992 9360 14000
rect 8960 13928 8968 13992
rect 9032 13928 9288 13992
rect 9352 13928 9360 13992
rect 8960 13920 9360 13928
rect 9440 13992 11440 14000
rect 9440 13928 9448 13992
rect 9512 13928 9768 13992
rect 9832 13928 10088 13992
rect 10152 13928 10408 13992
rect 10472 13928 10728 13992
rect 10792 13928 11048 13992
rect 11112 13928 11368 13992
rect 11432 13928 11440 13992
rect 9440 13920 11440 13928
rect 11520 13992 11920 14000
rect 11520 13928 11528 13992
rect 11592 13928 11848 13992
rect 11912 13928 11920 13992
rect 11520 13920 11920 13928
rect 12000 13992 12400 14000
rect 12000 13928 12008 13992
rect 12072 13928 12328 13992
rect 12392 13928 12400 13992
rect 12000 13920 12400 13928
rect 8480 13832 8880 13840
rect 8480 13768 8488 13832
rect 8552 13768 8808 13832
rect 8872 13768 8880 13832
rect 8480 13760 8880 13768
rect 8960 13832 9360 13840
rect 8960 13768 8968 13832
rect 9032 13768 9288 13832
rect 9352 13768 9360 13832
rect 8960 13760 9360 13768
rect 9440 13832 11440 13840
rect 9440 13768 9448 13832
rect 9512 13768 9768 13832
rect 9832 13768 10088 13832
rect 10152 13768 10408 13832
rect 10472 13768 10728 13832
rect 10792 13768 11048 13832
rect 11112 13768 11368 13832
rect 11432 13768 11440 13832
rect 9440 13760 11440 13768
rect 11520 13832 11920 13840
rect 11520 13768 11528 13832
rect 11592 13768 11848 13832
rect 11912 13768 11920 13832
rect 11520 13760 11920 13768
rect 12000 13832 12400 13840
rect 12000 13768 12008 13832
rect 12072 13768 12328 13832
rect 12392 13768 12400 13832
rect 12000 13760 12400 13768
rect 8480 13672 8880 13680
rect 8480 13608 8488 13672
rect 8552 13608 8808 13672
rect 8872 13608 8880 13672
rect 8480 13600 8880 13608
rect 8960 13672 9360 13680
rect 8960 13608 8968 13672
rect 9032 13608 9288 13672
rect 9352 13608 9360 13672
rect 8960 13600 9360 13608
rect 9440 13672 11440 13680
rect 9440 13608 9448 13672
rect 9512 13608 9768 13672
rect 9832 13608 10088 13672
rect 10152 13608 10408 13672
rect 10472 13608 10728 13672
rect 10792 13608 11048 13672
rect 11112 13608 11368 13672
rect 11432 13608 11440 13672
rect 9440 13600 11440 13608
rect 11520 13672 11920 13680
rect 11520 13608 11528 13672
rect 11592 13608 11848 13672
rect 11912 13608 11920 13672
rect 11520 13600 11920 13608
rect 12000 13672 12400 13680
rect 12000 13608 12008 13672
rect 12072 13608 12328 13672
rect 12392 13608 12400 13672
rect 12000 13600 12400 13608
rect 8480 13512 8880 13520
rect 8480 13448 8488 13512
rect 8552 13448 8808 13512
rect 8872 13448 8880 13512
rect 8480 13440 8880 13448
rect 8960 13512 9360 13520
rect 8960 13448 8968 13512
rect 9032 13448 9288 13512
rect 9352 13448 9360 13512
rect 8960 13440 9360 13448
rect 9440 13512 11440 13520
rect 9440 13448 9448 13512
rect 9512 13448 9768 13512
rect 9832 13448 10088 13512
rect 10152 13448 10408 13512
rect 10472 13448 10728 13512
rect 10792 13448 11048 13512
rect 11112 13448 11368 13512
rect 11432 13448 11440 13512
rect 9440 13440 11440 13448
rect 11520 13512 11920 13520
rect 11520 13448 11528 13512
rect 11592 13448 11848 13512
rect 11912 13448 11920 13512
rect 11520 13440 11920 13448
rect 12000 13512 12400 13520
rect 12000 13448 12008 13512
rect 12072 13448 12328 13512
rect 12392 13448 12400 13512
rect 12000 13440 12400 13448
rect 8480 13352 8880 13360
rect 8480 13288 8488 13352
rect 8552 13288 8808 13352
rect 8872 13288 8880 13352
rect 8480 13280 8880 13288
rect 8960 13352 9360 13360
rect 8960 13288 8968 13352
rect 9032 13288 9288 13352
rect 9352 13288 9360 13352
rect 8960 13280 9360 13288
rect 9440 13352 11440 13360
rect 9440 13288 9448 13352
rect 9512 13288 9768 13352
rect 9832 13288 10088 13352
rect 10152 13288 10408 13352
rect 10472 13288 10728 13352
rect 10792 13288 11048 13352
rect 11112 13288 11368 13352
rect 11432 13288 11440 13352
rect 9440 13280 11440 13288
rect 11520 13352 11920 13360
rect 11520 13288 11528 13352
rect 11592 13288 11848 13352
rect 11912 13288 11920 13352
rect 11520 13280 11920 13288
rect 12000 13352 12400 13360
rect 12000 13288 12008 13352
rect 12072 13288 12328 13352
rect 12392 13288 12400 13352
rect 12000 13280 12400 13288
rect 8480 13192 8880 13200
rect 8480 13128 8488 13192
rect 8552 13128 8808 13192
rect 8872 13128 8880 13192
rect 8480 13120 8880 13128
rect 8960 13192 9360 13200
rect 8960 13128 8968 13192
rect 9032 13128 9288 13192
rect 9352 13128 9360 13192
rect 8960 13120 9360 13128
rect 9440 13192 11440 13200
rect 9440 13128 9448 13192
rect 9512 13128 9768 13192
rect 9832 13128 10088 13192
rect 10152 13128 10408 13192
rect 10472 13128 10728 13192
rect 10792 13128 11048 13192
rect 11112 13128 11368 13192
rect 11432 13128 11440 13192
rect 9440 13120 11440 13128
rect 11520 13192 11920 13200
rect 11520 13128 11528 13192
rect 11592 13128 11848 13192
rect 11912 13128 11920 13192
rect 11520 13120 11920 13128
rect 12000 13192 12400 13200
rect 12000 13128 12008 13192
rect 12072 13128 12328 13192
rect 12392 13128 12400 13192
rect 12000 13120 12400 13128
rect 8480 13032 8880 13040
rect 8480 12968 8488 13032
rect 8552 12968 8808 13032
rect 8872 12968 8880 13032
rect 8480 12960 8880 12968
rect 8960 13032 9360 13040
rect 8960 12968 8968 13032
rect 9032 12968 9288 13032
rect 9352 12968 9360 13032
rect 8960 12960 9360 12968
rect 9440 13032 11440 13040
rect 9440 12968 9448 13032
rect 9512 12968 9768 13032
rect 9832 12968 10088 13032
rect 10152 12968 10408 13032
rect 10472 12968 10728 13032
rect 10792 12968 11048 13032
rect 11112 12968 11368 13032
rect 11432 12968 11440 13032
rect 9440 12960 11440 12968
rect 11520 13032 11920 13040
rect 11520 12968 11528 13032
rect 11592 12968 11848 13032
rect 11912 12968 11920 13032
rect 11520 12960 11920 12968
rect 12000 13032 12400 13040
rect 12000 12968 12008 13032
rect 12072 12968 12328 13032
rect 12392 12968 12400 13032
rect 12000 12960 12400 12968
rect 8480 12872 8880 12880
rect 8480 12808 8488 12872
rect 8552 12808 8808 12872
rect 8872 12808 8880 12872
rect 8480 12800 8880 12808
rect 8960 12872 9360 12880
rect 8960 12808 8968 12872
rect 9032 12808 9288 12872
rect 9352 12808 9360 12872
rect 8960 12800 9360 12808
rect 9440 12872 11440 12880
rect 9440 12808 9448 12872
rect 9512 12808 9768 12872
rect 9832 12808 10088 12872
rect 10152 12808 10408 12872
rect 10472 12808 10728 12872
rect 10792 12808 11048 12872
rect 11112 12808 11368 12872
rect 11432 12808 11440 12872
rect 9440 12800 11440 12808
rect 11520 12872 11920 12880
rect 11520 12808 11528 12872
rect 11592 12808 11848 12872
rect 11912 12808 11920 12872
rect 11520 12800 11920 12808
rect 12000 12872 12400 12880
rect 12000 12808 12008 12872
rect 12072 12808 12328 12872
rect 12392 12808 12400 12872
rect 12000 12800 12400 12808
rect 8480 12712 8880 12720
rect 8480 12648 8488 12712
rect 8552 12648 8808 12712
rect 8872 12648 8880 12712
rect 8480 12640 8880 12648
rect 8960 12712 9360 12720
rect 8960 12648 8968 12712
rect 9032 12648 9288 12712
rect 9352 12648 9360 12712
rect 8960 12640 9360 12648
rect 9440 12712 11440 12720
rect 9440 12648 9448 12712
rect 9512 12648 9768 12712
rect 9832 12648 10088 12712
rect 10152 12648 10408 12712
rect 10472 12648 10728 12712
rect 10792 12648 11048 12712
rect 11112 12648 11368 12712
rect 11432 12648 11440 12712
rect 9440 12640 11440 12648
rect 11520 12712 11920 12720
rect 11520 12648 11528 12712
rect 11592 12648 11848 12712
rect 11912 12648 11920 12712
rect 11520 12640 11920 12648
rect 12000 12712 12400 12720
rect 12000 12648 12008 12712
rect 12072 12648 12328 12712
rect 12392 12648 12400 12712
rect 12000 12640 12400 12648
rect 8480 12552 8880 12560
rect 8480 12488 8488 12552
rect 8552 12488 8808 12552
rect 8872 12488 8880 12552
rect 8480 12480 8880 12488
rect 8960 12552 9360 12560
rect 8960 12488 8968 12552
rect 9032 12488 9288 12552
rect 9352 12488 9360 12552
rect 8960 12480 9360 12488
rect 9440 12552 11440 12560
rect 9440 12488 9448 12552
rect 9512 12488 9768 12552
rect 9832 12488 10088 12552
rect 10152 12488 10408 12552
rect 10472 12488 10728 12552
rect 10792 12488 11048 12552
rect 11112 12488 11368 12552
rect 11432 12488 11440 12552
rect 9440 12480 11440 12488
rect 11520 12552 11920 12560
rect 11520 12488 11528 12552
rect 11592 12488 11848 12552
rect 11912 12488 11920 12552
rect 11520 12480 11920 12488
rect 12000 12552 12400 12560
rect 12000 12488 12008 12552
rect 12072 12488 12328 12552
rect 12392 12488 12400 12552
rect 12000 12480 12400 12488
rect 8480 12392 8880 12400
rect 8480 12328 8488 12392
rect 8552 12328 8808 12392
rect 8872 12328 8880 12392
rect 8480 12320 8880 12328
rect 8960 12392 9360 12400
rect 8960 12328 8968 12392
rect 9032 12328 9288 12392
rect 9352 12328 9360 12392
rect 8960 12320 9360 12328
rect 9440 12392 11440 12400
rect 9440 12328 9448 12392
rect 9512 12328 9768 12392
rect 9832 12328 10088 12392
rect 10152 12328 10408 12392
rect 10472 12328 10728 12392
rect 10792 12328 11048 12392
rect 11112 12328 11368 12392
rect 11432 12328 11440 12392
rect 9440 12320 11440 12328
rect 11520 12392 11920 12400
rect 11520 12328 11528 12392
rect 11592 12328 11848 12392
rect 11912 12328 11920 12392
rect 11520 12320 11920 12328
rect 12000 12392 12400 12400
rect 12000 12328 12008 12392
rect 12072 12328 12328 12392
rect 12392 12328 12400 12392
rect 12000 12320 12400 12328
rect 8480 12232 8880 12240
rect 8480 12168 8488 12232
rect 8552 12168 8808 12232
rect 8872 12168 8880 12232
rect 8480 12160 8880 12168
rect 8960 12232 9360 12240
rect 8960 12168 8968 12232
rect 9032 12168 9288 12232
rect 9352 12168 9360 12232
rect 8960 12160 9360 12168
rect 9440 12232 11440 12240
rect 9440 12168 9448 12232
rect 9512 12168 9768 12232
rect 9832 12168 10088 12232
rect 10152 12168 10408 12232
rect 10472 12168 10728 12232
rect 10792 12168 11048 12232
rect 11112 12168 11368 12232
rect 11432 12168 11440 12232
rect 9440 12160 11440 12168
rect 11520 12232 11920 12240
rect 11520 12168 11528 12232
rect 11592 12168 11848 12232
rect 11912 12168 11920 12232
rect 11520 12160 11920 12168
rect 12000 12232 12400 12240
rect 12000 12168 12008 12232
rect 12072 12168 12328 12232
rect 12392 12168 12400 12232
rect 12000 12160 12400 12168
rect 8480 12072 8880 12080
rect 8480 12008 8488 12072
rect 8552 12008 8808 12072
rect 8872 12008 8880 12072
rect 8480 12000 8880 12008
rect 8960 12072 9360 12080
rect 8960 12008 8968 12072
rect 9032 12008 9288 12072
rect 9352 12008 9360 12072
rect 8960 12000 9360 12008
rect 9440 12072 11440 12080
rect 9440 12008 9448 12072
rect 9512 12008 9768 12072
rect 9832 12008 10088 12072
rect 10152 12008 10408 12072
rect 10472 12008 10728 12072
rect 10792 12008 11048 12072
rect 11112 12008 11368 12072
rect 11432 12008 11440 12072
rect 9440 12000 11440 12008
rect 11520 12072 11920 12080
rect 11520 12008 11528 12072
rect 11592 12008 11848 12072
rect 11912 12008 11920 12072
rect 11520 12000 11920 12008
rect 12000 12072 12400 12080
rect 12000 12008 12008 12072
rect 12072 12008 12328 12072
rect 12392 12008 12400 12072
rect 12000 12000 12400 12008
rect 8480 11912 8880 11920
rect 8480 11848 8488 11912
rect 8552 11848 8808 11912
rect 8872 11848 8880 11912
rect 8480 11840 8880 11848
rect 8960 11912 9360 11920
rect 8960 11848 8968 11912
rect 9032 11848 9288 11912
rect 9352 11848 9360 11912
rect 8960 11840 9360 11848
rect 9440 11912 11440 11920
rect 9440 11848 9448 11912
rect 9512 11848 9768 11912
rect 9832 11848 10088 11912
rect 10152 11848 10408 11912
rect 10472 11848 10728 11912
rect 10792 11848 11048 11912
rect 11112 11848 11368 11912
rect 11432 11848 11440 11912
rect 9440 11840 11440 11848
rect 11520 11912 11920 11920
rect 11520 11848 11528 11912
rect 11592 11848 11848 11912
rect 11912 11848 11920 11912
rect 11520 11840 11920 11848
rect 12000 11912 12400 11920
rect 12000 11848 12008 11912
rect 12072 11848 12328 11912
rect 12392 11848 12400 11912
rect 12000 11840 12400 11848
rect 8480 11752 8880 11760
rect 8480 11688 8488 11752
rect 8552 11688 8808 11752
rect 8872 11688 8880 11752
rect 8480 11680 8880 11688
rect 8960 11752 9360 11760
rect 8960 11688 8968 11752
rect 9032 11688 9288 11752
rect 9352 11688 9360 11752
rect 8960 11680 9360 11688
rect 9440 11752 11440 11760
rect 9440 11688 9448 11752
rect 9512 11688 9768 11752
rect 9832 11688 10088 11752
rect 10152 11688 10408 11752
rect 10472 11688 10728 11752
rect 10792 11688 11048 11752
rect 11112 11688 11368 11752
rect 11432 11688 11440 11752
rect 9440 11680 11440 11688
rect 11520 11752 11920 11760
rect 11520 11688 11528 11752
rect 11592 11688 11848 11752
rect 11912 11688 11920 11752
rect 11520 11680 11920 11688
rect 12000 11752 12400 11760
rect 12000 11688 12008 11752
rect 12072 11688 12328 11752
rect 12392 11688 12400 11752
rect 12000 11680 12400 11688
rect 8480 11592 8880 11600
rect 8480 11528 8488 11592
rect 8552 11528 8808 11592
rect 8872 11528 8880 11592
rect 8480 11520 8880 11528
rect 8960 11592 9360 11600
rect 8960 11528 8968 11592
rect 9032 11528 9288 11592
rect 9352 11528 9360 11592
rect 8960 11520 9360 11528
rect 9440 11592 11440 11600
rect 9440 11528 9448 11592
rect 9512 11528 9768 11592
rect 9832 11528 10088 11592
rect 10152 11528 10408 11592
rect 10472 11528 10728 11592
rect 10792 11528 11048 11592
rect 11112 11528 11368 11592
rect 11432 11528 11440 11592
rect 9440 11520 11440 11528
rect 11520 11592 11920 11600
rect 11520 11528 11528 11592
rect 11592 11528 11848 11592
rect 11912 11528 11920 11592
rect 11520 11520 11920 11528
rect 12000 11592 12400 11600
rect 12000 11528 12008 11592
rect 12072 11528 12328 11592
rect 12392 11528 12400 11592
rect 12000 11520 12400 11528
rect 8480 11432 8880 11440
rect 8480 11368 8488 11432
rect 8552 11368 8808 11432
rect 8872 11368 8880 11432
rect 8480 11360 8880 11368
rect 8960 11432 9360 11440
rect 8960 11368 8968 11432
rect 9032 11368 9288 11432
rect 9352 11368 9360 11432
rect 8960 11360 9360 11368
rect 9440 11432 11440 11440
rect 9440 11368 9448 11432
rect 9512 11368 9768 11432
rect 9832 11368 10088 11432
rect 10152 11368 10408 11432
rect 10472 11368 10728 11432
rect 10792 11368 11048 11432
rect 11112 11368 11368 11432
rect 11432 11368 11440 11432
rect 9440 11360 11440 11368
rect 11520 11432 11920 11440
rect 11520 11368 11528 11432
rect 11592 11368 11848 11432
rect 11912 11368 11920 11432
rect 11520 11360 11920 11368
rect 12000 11432 12400 11440
rect 12000 11368 12008 11432
rect 12072 11368 12328 11432
rect 12392 11368 12400 11432
rect 12000 11360 12400 11368
rect 8480 11272 8880 11280
rect 8480 11208 8488 11272
rect 8552 11208 8808 11272
rect 8872 11208 8880 11272
rect 8480 11200 8880 11208
rect 8960 11272 9360 11280
rect 8960 11208 8968 11272
rect 9032 11208 9288 11272
rect 9352 11208 9360 11272
rect 8960 11200 9360 11208
rect 9440 11272 11440 11280
rect 9440 11208 9448 11272
rect 9512 11208 9768 11272
rect 9832 11208 10088 11272
rect 10152 11208 10408 11272
rect 10472 11208 10728 11272
rect 10792 11208 11048 11272
rect 11112 11208 11368 11272
rect 11432 11208 11440 11272
rect 9440 11200 11440 11208
rect 11520 11272 11920 11280
rect 11520 11208 11528 11272
rect 11592 11208 11848 11272
rect 11912 11208 11920 11272
rect 11520 11200 11920 11208
rect 12000 11272 12400 11280
rect 12000 11208 12008 11272
rect 12072 11208 12328 11272
rect 12392 11208 12400 11272
rect 12000 11200 12400 11208
rect 8480 11112 8880 11120
rect 8480 11048 8488 11112
rect 8552 11048 8808 11112
rect 8872 11048 8880 11112
rect 8480 11040 8880 11048
rect 8960 11112 9360 11120
rect 8960 11048 8968 11112
rect 9032 11048 9288 11112
rect 9352 11048 9360 11112
rect 8960 11040 9360 11048
rect 9440 11112 11440 11120
rect 9440 11048 9448 11112
rect 9512 11048 9768 11112
rect 9832 11048 10088 11112
rect 10152 11048 10408 11112
rect 10472 11048 10728 11112
rect 10792 11048 11048 11112
rect 11112 11048 11368 11112
rect 11432 11048 11440 11112
rect 9440 11040 11440 11048
rect 11520 11112 11920 11120
rect 11520 11048 11528 11112
rect 11592 11048 11848 11112
rect 11912 11048 11920 11112
rect 11520 11040 11920 11048
rect 12000 11112 12400 11120
rect 12000 11048 12008 11112
rect 12072 11048 12328 11112
rect 12392 11048 12400 11112
rect 12000 11040 12400 11048
rect 8480 10952 8880 10960
rect 8480 10888 8488 10952
rect 8552 10888 8808 10952
rect 8872 10888 8880 10952
rect 8480 10880 8880 10888
rect 8960 10952 9360 10960
rect 8960 10888 8968 10952
rect 9032 10888 9288 10952
rect 9352 10888 9360 10952
rect 8960 10880 9360 10888
rect 9440 10952 11440 10960
rect 9440 10888 9448 10952
rect 9512 10888 9768 10952
rect 9832 10888 10088 10952
rect 10152 10888 10408 10952
rect 10472 10888 10728 10952
rect 10792 10888 11048 10952
rect 11112 10888 11368 10952
rect 11432 10888 11440 10952
rect 9440 10880 11440 10888
rect 11520 10952 11920 10960
rect 11520 10888 11528 10952
rect 11592 10888 11848 10952
rect 11912 10888 11920 10952
rect 11520 10880 11920 10888
rect 12000 10952 12400 10960
rect 12000 10888 12008 10952
rect 12072 10888 12328 10952
rect 12392 10888 12400 10952
rect 12000 10880 12400 10888
rect 8480 10792 8880 10800
rect 8480 10728 8488 10792
rect 8552 10728 8808 10792
rect 8872 10728 8880 10792
rect 8480 10720 8880 10728
rect 8960 10792 9360 10800
rect 8960 10728 8968 10792
rect 9032 10728 9288 10792
rect 9352 10728 9360 10792
rect 8960 10720 9360 10728
rect 9440 10792 11440 10800
rect 9440 10728 9448 10792
rect 9512 10728 9768 10792
rect 9832 10728 10088 10792
rect 10152 10728 10408 10792
rect 10472 10728 10728 10792
rect 10792 10728 11048 10792
rect 11112 10728 11368 10792
rect 11432 10728 11440 10792
rect 9440 10720 11440 10728
rect 11520 10792 11920 10800
rect 11520 10728 11528 10792
rect 11592 10728 11848 10792
rect 11912 10728 11920 10792
rect 11520 10720 11920 10728
rect 12000 10792 12400 10800
rect 12000 10728 12008 10792
rect 12072 10728 12328 10792
rect 12392 10728 12400 10792
rect 12000 10720 12400 10728
rect 8480 10632 8880 10640
rect 8480 10568 8488 10632
rect 8552 10568 8808 10632
rect 8872 10568 8880 10632
rect 8480 10560 8880 10568
rect 8960 10632 9360 10640
rect 8960 10568 8968 10632
rect 9032 10568 9288 10632
rect 9352 10568 9360 10632
rect 8960 10560 9360 10568
rect 9440 10632 11440 10640
rect 9440 10568 9448 10632
rect 9512 10568 9768 10632
rect 9832 10568 10088 10632
rect 10152 10568 10408 10632
rect 10472 10568 10728 10632
rect 10792 10568 11048 10632
rect 11112 10568 11368 10632
rect 11432 10568 11440 10632
rect 9440 10560 11440 10568
rect 11520 10632 11920 10640
rect 11520 10568 11528 10632
rect 11592 10568 11848 10632
rect 11912 10568 11920 10632
rect 11520 10560 11920 10568
rect 12000 10632 12400 10640
rect 12000 10568 12008 10632
rect 12072 10568 12328 10632
rect 12392 10568 12400 10632
rect 12000 10560 12400 10568
rect 8480 10472 8880 10480
rect 8480 10408 8488 10472
rect 8552 10408 8808 10472
rect 8872 10408 8880 10472
rect 8480 10400 8880 10408
rect 8960 10472 9360 10480
rect 8960 10408 8968 10472
rect 9032 10408 9288 10472
rect 9352 10408 9360 10472
rect 8960 10400 9360 10408
rect 9440 10472 11440 10480
rect 9440 10408 9448 10472
rect 9512 10408 9768 10472
rect 9832 10408 10088 10472
rect 10152 10408 10408 10472
rect 10472 10408 10728 10472
rect 10792 10408 11048 10472
rect 11112 10408 11368 10472
rect 11432 10408 11440 10472
rect 9440 10400 11440 10408
rect 11520 10472 11920 10480
rect 11520 10408 11528 10472
rect 11592 10408 11848 10472
rect 11912 10408 11920 10472
rect 11520 10400 11920 10408
rect 12000 10472 12400 10480
rect 12000 10408 12008 10472
rect 12072 10408 12328 10472
rect 12392 10408 12400 10472
rect 12000 10400 12400 10408
rect 8480 10312 8880 10320
rect 8480 10248 8488 10312
rect 8552 10248 8808 10312
rect 8872 10248 8880 10312
rect 8480 10240 8880 10248
rect 8960 10312 9360 10320
rect 8960 10248 8968 10312
rect 9032 10248 9288 10312
rect 9352 10248 9360 10312
rect 8960 10240 9360 10248
rect 9440 10312 11440 10320
rect 9440 10248 9448 10312
rect 9512 10248 9768 10312
rect 9832 10248 10088 10312
rect 10152 10248 10408 10312
rect 10472 10248 10728 10312
rect 10792 10248 11048 10312
rect 11112 10248 11368 10312
rect 11432 10248 11440 10312
rect 9440 10240 11440 10248
rect 11520 10312 11920 10320
rect 11520 10248 11528 10312
rect 11592 10248 11848 10312
rect 11912 10248 11920 10312
rect 11520 10240 11920 10248
rect 12000 10312 12400 10320
rect 12000 10248 12008 10312
rect 12072 10248 12328 10312
rect 12392 10248 12400 10312
rect 12000 10240 12400 10248
rect 8480 10152 8880 10160
rect 8480 10088 8488 10152
rect 8552 10088 8808 10152
rect 8872 10088 8880 10152
rect 8480 10080 8880 10088
rect 8960 10152 9360 10160
rect 8960 10088 8968 10152
rect 9032 10088 9288 10152
rect 9352 10088 9360 10152
rect 8960 10080 9360 10088
rect 9440 10152 11440 10160
rect 9440 10088 9448 10152
rect 9512 10088 9768 10152
rect 9832 10088 10088 10152
rect 10152 10088 10408 10152
rect 10472 10088 10728 10152
rect 10792 10088 11048 10152
rect 11112 10088 11368 10152
rect 11432 10088 11440 10152
rect 9440 10080 11440 10088
rect 11520 10152 11920 10160
rect 11520 10088 11528 10152
rect 11592 10088 11848 10152
rect 11912 10088 11920 10152
rect 11520 10080 11920 10088
rect 12000 10152 12400 10160
rect 12000 10088 12008 10152
rect 12072 10088 12328 10152
rect 12392 10088 12400 10152
rect 12000 10080 12400 10088
rect 8480 9992 8880 10000
rect 8480 9928 8488 9992
rect 8552 9928 8808 9992
rect 8872 9928 8880 9992
rect 8480 9920 8880 9928
rect 8960 9992 9360 10000
rect 8960 9928 8968 9992
rect 9032 9928 9288 9992
rect 9352 9928 9360 9992
rect 8960 9920 9360 9928
rect 9440 9992 11440 10000
rect 9440 9928 9448 9992
rect 9512 9928 9768 9992
rect 9832 9928 10088 9992
rect 10152 9928 10408 9992
rect 10472 9928 10728 9992
rect 10792 9928 11048 9992
rect 11112 9928 11368 9992
rect 11432 9928 11440 9992
rect 9440 9920 11440 9928
rect 11520 9992 11920 10000
rect 11520 9928 11528 9992
rect 11592 9928 11848 9992
rect 11912 9928 11920 9992
rect 11520 9920 11920 9928
rect 12000 9992 12400 10000
rect 12000 9928 12008 9992
rect 12072 9928 12328 9992
rect 12392 9928 12400 9992
rect 12000 9920 12400 9928
rect 8480 9832 8880 9840
rect 8480 9768 8488 9832
rect 8552 9768 8808 9832
rect 8872 9768 8880 9832
rect 8480 9760 8880 9768
rect 8960 9832 9360 9840
rect 8960 9768 8968 9832
rect 9032 9768 9288 9832
rect 9352 9768 9360 9832
rect 8960 9760 9360 9768
rect 9440 9832 11440 9840
rect 9440 9768 9448 9832
rect 9512 9768 9768 9832
rect 9832 9768 10088 9832
rect 10152 9768 10408 9832
rect 10472 9768 10728 9832
rect 10792 9768 11048 9832
rect 11112 9768 11368 9832
rect 11432 9768 11440 9832
rect 9440 9760 11440 9768
rect 11520 9832 11920 9840
rect 11520 9768 11528 9832
rect 11592 9768 11848 9832
rect 11912 9768 11920 9832
rect 11520 9760 11920 9768
rect 12000 9832 12400 9840
rect 12000 9768 12008 9832
rect 12072 9768 12328 9832
rect 12392 9768 12400 9832
rect 12000 9760 12400 9768
rect 8480 9672 8880 9680
rect 8480 9608 8488 9672
rect 8552 9608 8808 9672
rect 8872 9608 8880 9672
rect 8480 9600 8880 9608
rect 8960 9672 9360 9680
rect 8960 9608 8968 9672
rect 9032 9608 9288 9672
rect 9352 9608 9360 9672
rect 8960 9600 9360 9608
rect 9440 9672 11440 9680
rect 9440 9608 9448 9672
rect 9512 9608 9768 9672
rect 9832 9608 10088 9672
rect 10152 9608 10408 9672
rect 10472 9608 10728 9672
rect 10792 9608 11048 9672
rect 11112 9608 11368 9672
rect 11432 9608 11440 9672
rect 9440 9600 11440 9608
rect 11520 9672 11920 9680
rect 11520 9608 11528 9672
rect 11592 9608 11848 9672
rect 11912 9608 11920 9672
rect 11520 9600 11920 9608
rect 12000 9672 12400 9680
rect 12000 9608 12008 9672
rect 12072 9608 12328 9672
rect 12392 9608 12400 9672
rect 12000 9600 12400 9608
rect 8480 9512 8880 9520
rect 8480 9448 8488 9512
rect 8552 9448 8808 9512
rect 8872 9448 8880 9512
rect 8480 9440 8880 9448
rect 8960 9512 9360 9520
rect 8960 9448 8968 9512
rect 9032 9448 9288 9512
rect 9352 9448 9360 9512
rect 8960 9440 9360 9448
rect 9440 9512 11440 9520
rect 9440 9448 9448 9512
rect 9512 9448 9768 9512
rect 9832 9448 10088 9512
rect 10152 9448 10408 9512
rect 10472 9448 10728 9512
rect 10792 9448 11048 9512
rect 11112 9448 11368 9512
rect 11432 9448 11440 9512
rect 9440 9440 11440 9448
rect 11520 9512 11920 9520
rect 11520 9448 11528 9512
rect 11592 9448 11848 9512
rect 11912 9448 11920 9512
rect 11520 9440 11920 9448
rect 12000 9512 12400 9520
rect 12000 9448 12008 9512
rect 12072 9448 12328 9512
rect 12392 9448 12400 9512
rect 12000 9440 12400 9448
rect 8480 9352 8880 9360
rect 8480 9288 8488 9352
rect 8552 9288 8808 9352
rect 8872 9288 8880 9352
rect 8480 9280 8880 9288
rect 8960 9352 9360 9360
rect 8960 9288 8968 9352
rect 9032 9288 9288 9352
rect 9352 9288 9360 9352
rect 8960 9280 9360 9288
rect 9440 9352 11440 9360
rect 9440 9288 9448 9352
rect 9512 9288 9768 9352
rect 9832 9288 10088 9352
rect 10152 9288 10408 9352
rect 10472 9288 10728 9352
rect 10792 9288 11048 9352
rect 11112 9288 11368 9352
rect 11432 9288 11440 9352
rect 9440 9280 11440 9288
rect 11520 9352 11920 9360
rect 11520 9288 11528 9352
rect 11592 9288 11848 9352
rect 11912 9288 11920 9352
rect 11520 9280 11920 9288
rect 12000 9352 12400 9360
rect 12000 9288 12008 9352
rect 12072 9288 12328 9352
rect 12392 9288 12400 9352
rect 12000 9280 12400 9288
rect 8480 9192 8880 9200
rect 8480 9128 8488 9192
rect 8552 9128 8808 9192
rect 8872 9128 8880 9192
rect 8480 9120 8880 9128
rect 8960 9192 9360 9200
rect 8960 9128 8968 9192
rect 9032 9128 9288 9192
rect 9352 9128 9360 9192
rect 8960 9120 9360 9128
rect 9440 9192 11440 9200
rect 9440 9128 9448 9192
rect 9512 9128 9768 9192
rect 9832 9128 10088 9192
rect 10152 9128 10408 9192
rect 10472 9128 10728 9192
rect 10792 9128 11048 9192
rect 11112 9128 11368 9192
rect 11432 9128 11440 9192
rect 9440 9120 11440 9128
rect 11520 9192 11920 9200
rect 11520 9128 11528 9192
rect 11592 9128 11848 9192
rect 11912 9128 11920 9192
rect 11520 9120 11920 9128
rect 12000 9192 12400 9200
rect 12000 9128 12008 9192
rect 12072 9128 12328 9192
rect 12392 9128 12400 9192
rect 12000 9120 12400 9128
rect 8480 9032 8880 9040
rect 8480 8968 8488 9032
rect 8552 8968 8808 9032
rect 8872 8968 8880 9032
rect 8480 8960 8880 8968
rect 8960 9032 9360 9040
rect 8960 8968 8968 9032
rect 9032 8968 9288 9032
rect 9352 8968 9360 9032
rect 8960 8960 9360 8968
rect 9440 9032 11440 9040
rect 9440 8968 9448 9032
rect 9512 8968 9768 9032
rect 9832 8968 10088 9032
rect 10152 8968 10408 9032
rect 10472 8968 10728 9032
rect 10792 8968 11048 9032
rect 11112 8968 11368 9032
rect 11432 8968 11440 9032
rect 9440 8960 11440 8968
rect 11520 9032 11920 9040
rect 11520 8968 11528 9032
rect 11592 8968 11848 9032
rect 11912 8968 11920 9032
rect 11520 8960 11920 8968
rect 12000 9032 12400 9040
rect 12000 8968 12008 9032
rect 12072 8968 12328 9032
rect 12392 8968 12400 9032
rect 12000 8960 12400 8968
rect 8480 8872 8880 8880
rect 8480 8808 8488 8872
rect 8552 8808 8808 8872
rect 8872 8808 8880 8872
rect 8480 8800 8880 8808
rect 8960 8872 9360 8880
rect 8960 8808 8968 8872
rect 9032 8808 9288 8872
rect 9352 8808 9360 8872
rect 8960 8800 9360 8808
rect 9440 8872 11440 8880
rect 9440 8808 9448 8872
rect 9512 8808 9768 8872
rect 9832 8808 10088 8872
rect 10152 8808 10408 8872
rect 10472 8808 10728 8872
rect 10792 8808 11048 8872
rect 11112 8808 11368 8872
rect 11432 8808 11440 8872
rect 9440 8800 11440 8808
rect 11520 8872 11920 8880
rect 11520 8808 11528 8872
rect 11592 8808 11848 8872
rect 11912 8808 11920 8872
rect 11520 8800 11920 8808
rect 12000 8872 12400 8880
rect 12000 8808 12008 8872
rect 12072 8808 12328 8872
rect 12392 8808 12400 8872
rect 12000 8800 12400 8808
rect 8480 8712 8880 8720
rect 8480 8648 8488 8712
rect 8552 8648 8808 8712
rect 8872 8648 8880 8712
rect 8480 8640 8880 8648
rect 8960 8712 9360 8720
rect 8960 8648 8968 8712
rect 9032 8648 9288 8712
rect 9352 8648 9360 8712
rect 8960 8640 9360 8648
rect 9440 8712 11440 8720
rect 9440 8648 9448 8712
rect 9512 8648 9768 8712
rect 9832 8648 10088 8712
rect 10152 8648 10408 8712
rect 10472 8648 10728 8712
rect 10792 8648 11048 8712
rect 11112 8648 11368 8712
rect 11432 8648 11440 8712
rect 9440 8640 11440 8648
rect 11520 8712 11920 8720
rect 11520 8648 11528 8712
rect 11592 8648 11848 8712
rect 11912 8648 11920 8712
rect 11520 8640 11920 8648
rect 12000 8712 12400 8720
rect 12000 8648 12008 8712
rect 12072 8648 12328 8712
rect 12392 8648 12400 8712
rect 12000 8640 12400 8648
rect 8480 8552 8880 8560
rect 8480 8488 8488 8552
rect 8552 8488 8808 8552
rect 8872 8488 8880 8552
rect 8480 8480 8880 8488
rect 8960 8552 9360 8560
rect 8960 8488 8968 8552
rect 9032 8488 9288 8552
rect 9352 8488 9360 8552
rect 8960 8480 9360 8488
rect 9440 8552 11440 8560
rect 9440 8488 9448 8552
rect 9512 8488 9768 8552
rect 9832 8488 10088 8552
rect 10152 8488 10408 8552
rect 10472 8488 10728 8552
rect 10792 8488 11048 8552
rect 11112 8488 11368 8552
rect 11432 8488 11440 8552
rect 9440 8480 11440 8488
rect 11520 8552 11920 8560
rect 11520 8488 11528 8552
rect 11592 8488 11848 8552
rect 11912 8488 11920 8552
rect 11520 8480 11920 8488
rect 12000 8552 12400 8560
rect 12000 8488 12008 8552
rect 12072 8488 12328 8552
rect 12392 8488 12400 8552
rect 12000 8480 12400 8488
rect 8480 8392 8880 8400
rect 8480 8328 8488 8392
rect 8552 8328 8808 8392
rect 8872 8328 8880 8392
rect 8480 8320 8880 8328
rect 8960 8392 9360 8400
rect 8960 8328 8968 8392
rect 9032 8328 9288 8392
rect 9352 8328 9360 8392
rect 8960 8320 9360 8328
rect 9440 8392 11440 8400
rect 9440 8328 9448 8392
rect 9512 8328 9768 8392
rect 9832 8328 10088 8392
rect 10152 8328 10408 8392
rect 10472 8328 10728 8392
rect 10792 8328 11048 8392
rect 11112 8328 11368 8392
rect 11432 8328 11440 8392
rect 9440 8320 11440 8328
rect 11520 8392 11920 8400
rect 11520 8328 11528 8392
rect 11592 8328 11848 8392
rect 11912 8328 11920 8392
rect 11520 8320 11920 8328
rect 12000 8392 12400 8400
rect 12000 8328 12008 8392
rect 12072 8328 12328 8392
rect 12392 8328 12400 8392
rect 12000 8320 12400 8328
rect 8480 8232 8880 8240
rect 8480 8168 8488 8232
rect 8552 8168 8808 8232
rect 8872 8168 8880 8232
rect 8480 8160 8880 8168
rect 8960 8232 9360 8240
rect 8960 8168 8968 8232
rect 9032 8168 9288 8232
rect 9352 8168 9360 8232
rect 8960 8160 9360 8168
rect 9440 8232 11440 8240
rect 9440 8168 9448 8232
rect 9512 8168 9768 8232
rect 9832 8168 10088 8232
rect 10152 8168 10408 8232
rect 10472 8168 10728 8232
rect 10792 8168 11048 8232
rect 11112 8168 11368 8232
rect 11432 8168 11440 8232
rect 9440 8160 11440 8168
rect 11520 8232 11920 8240
rect 11520 8168 11528 8232
rect 11592 8168 11848 8232
rect 11912 8168 11920 8232
rect 11520 8160 11920 8168
rect 12000 8232 12400 8240
rect 12000 8168 12008 8232
rect 12072 8168 12328 8232
rect 12392 8168 12400 8232
rect 12000 8160 12400 8168
rect 8480 8072 8880 8080
rect 8480 8008 8488 8072
rect 8552 8008 8808 8072
rect 8872 8008 8880 8072
rect 8480 8000 8880 8008
rect 8960 8072 9360 8080
rect 8960 8008 8968 8072
rect 9032 8008 9288 8072
rect 9352 8008 9360 8072
rect 8960 8000 9360 8008
rect 9440 8072 11440 8080
rect 9440 8008 9448 8072
rect 9512 8008 9768 8072
rect 9832 8008 10088 8072
rect 10152 8008 10408 8072
rect 10472 8008 10728 8072
rect 10792 8008 11048 8072
rect 11112 8008 11368 8072
rect 11432 8008 11440 8072
rect 9440 8000 11440 8008
rect 11520 8072 11920 8080
rect 11520 8008 11528 8072
rect 11592 8008 11848 8072
rect 11912 8008 11920 8072
rect 11520 8000 11920 8008
rect 12000 8072 12400 8080
rect 12000 8008 12008 8072
rect 12072 8008 12328 8072
rect 12392 8008 12400 8072
rect 12000 8000 12400 8008
rect 8480 7912 8880 7920
rect 8480 7848 8488 7912
rect 8552 7848 8808 7912
rect 8872 7848 8880 7912
rect 8480 7840 8880 7848
rect 8960 7912 9360 7920
rect 8960 7848 8968 7912
rect 9032 7848 9288 7912
rect 9352 7848 9360 7912
rect 8960 7840 9360 7848
rect 9440 7912 11440 7920
rect 9440 7848 9448 7912
rect 9512 7848 9768 7912
rect 9832 7848 10088 7912
rect 10152 7848 10408 7912
rect 10472 7848 10728 7912
rect 10792 7848 11048 7912
rect 11112 7848 11368 7912
rect 11432 7848 11440 7912
rect 9440 7840 11440 7848
rect 11520 7912 11920 7920
rect 11520 7848 11528 7912
rect 11592 7848 11848 7912
rect 11912 7848 11920 7912
rect 11520 7840 11920 7848
rect 12000 7912 12400 7920
rect 12000 7848 12008 7912
rect 12072 7848 12328 7912
rect 12392 7848 12400 7912
rect 12000 7840 12400 7848
rect 8480 7752 8880 7760
rect 8480 7688 8488 7752
rect 8552 7688 8808 7752
rect 8872 7688 8880 7752
rect 8480 7680 8880 7688
rect 8960 7752 9360 7760
rect 8960 7688 8968 7752
rect 9032 7688 9288 7752
rect 9352 7688 9360 7752
rect 8960 7680 9360 7688
rect 9440 7752 11440 7760
rect 9440 7688 9448 7752
rect 9512 7688 9768 7752
rect 9832 7688 10088 7752
rect 10152 7688 10408 7752
rect 10472 7688 10728 7752
rect 10792 7688 11048 7752
rect 11112 7688 11368 7752
rect 11432 7688 11440 7752
rect 9440 7680 11440 7688
rect 11520 7752 11920 7760
rect 11520 7688 11528 7752
rect 11592 7688 11848 7752
rect 11912 7688 11920 7752
rect 11520 7680 11920 7688
rect 12000 7752 12400 7760
rect 12000 7688 12008 7752
rect 12072 7688 12328 7752
rect 12392 7688 12400 7752
rect 12000 7680 12400 7688
rect 8480 7592 8880 7600
rect 8480 7528 8488 7592
rect 8552 7528 8808 7592
rect 8872 7528 8880 7592
rect 8480 7520 8880 7528
rect 8960 7592 9360 7600
rect 8960 7528 8968 7592
rect 9032 7528 9288 7592
rect 9352 7528 9360 7592
rect 8960 7520 9360 7528
rect 9440 7592 11440 7600
rect 9440 7528 9448 7592
rect 9512 7528 9768 7592
rect 9832 7528 10088 7592
rect 10152 7528 10408 7592
rect 10472 7528 10728 7592
rect 10792 7528 11048 7592
rect 11112 7528 11368 7592
rect 11432 7528 11440 7592
rect 9440 7520 11440 7528
rect 11520 7592 11920 7600
rect 11520 7528 11528 7592
rect 11592 7528 11848 7592
rect 11912 7528 11920 7592
rect 11520 7520 11920 7528
rect 12000 7592 12400 7600
rect 12000 7528 12008 7592
rect 12072 7528 12328 7592
rect 12392 7528 12400 7592
rect 12000 7520 12400 7528
rect 8480 7432 8880 7440
rect 8480 7368 8488 7432
rect 8552 7368 8808 7432
rect 8872 7368 8880 7432
rect 8480 7360 8880 7368
rect 8960 7432 9360 7440
rect 8960 7368 8968 7432
rect 9032 7368 9288 7432
rect 9352 7368 9360 7432
rect 8960 7360 9360 7368
rect 9440 7432 11440 7440
rect 9440 7368 9448 7432
rect 9512 7368 9768 7432
rect 9832 7368 10088 7432
rect 10152 7368 10408 7432
rect 10472 7368 10728 7432
rect 10792 7368 11048 7432
rect 11112 7368 11368 7432
rect 11432 7368 11440 7432
rect 9440 7360 11440 7368
rect 11520 7432 11920 7440
rect 11520 7368 11528 7432
rect 11592 7368 11848 7432
rect 11912 7368 11920 7432
rect 11520 7360 11920 7368
rect 12000 7432 12400 7440
rect 12000 7368 12008 7432
rect 12072 7368 12328 7432
rect 12392 7368 12400 7432
rect 12000 7360 12400 7368
rect 8480 7272 8880 7280
rect 8480 7208 8488 7272
rect 8552 7208 8808 7272
rect 8872 7208 8880 7272
rect 8480 7200 8880 7208
rect 8960 7272 9360 7280
rect 8960 7208 8968 7272
rect 9032 7208 9288 7272
rect 9352 7208 9360 7272
rect 8960 7200 9360 7208
rect 9440 7272 11440 7280
rect 9440 7208 9448 7272
rect 9512 7208 9768 7272
rect 9832 7208 10088 7272
rect 10152 7208 10408 7272
rect 10472 7208 10728 7272
rect 10792 7208 11048 7272
rect 11112 7208 11368 7272
rect 11432 7208 11440 7272
rect 9440 7200 11440 7208
rect 11520 7272 11920 7280
rect 11520 7208 11528 7272
rect 11592 7208 11848 7272
rect 11912 7208 11920 7272
rect 11520 7200 11920 7208
rect 12000 7272 12400 7280
rect 12000 7208 12008 7272
rect 12072 7208 12328 7272
rect 12392 7208 12400 7272
rect 12000 7200 12400 7208
rect 8480 7112 8880 7120
rect 8480 7048 8488 7112
rect 8552 7048 8808 7112
rect 8872 7048 8880 7112
rect 8480 7040 8880 7048
rect 8960 7112 9360 7120
rect 8960 7048 8968 7112
rect 9032 7048 9288 7112
rect 9352 7048 9360 7112
rect 8960 7040 9360 7048
rect 9440 7112 11440 7120
rect 9440 7048 9448 7112
rect 9512 7048 9768 7112
rect 9832 7048 10088 7112
rect 10152 7048 10408 7112
rect 10472 7048 10728 7112
rect 10792 7048 11048 7112
rect 11112 7048 11368 7112
rect 11432 7048 11440 7112
rect 9440 7040 11440 7048
rect 11520 7112 11920 7120
rect 11520 7048 11528 7112
rect 11592 7048 11848 7112
rect 11912 7048 11920 7112
rect 11520 7040 11920 7048
rect 12000 7112 12400 7120
rect 12000 7048 12008 7112
rect 12072 7048 12328 7112
rect 12392 7048 12400 7112
rect 12000 7040 12400 7048
rect 8480 6952 8880 6960
rect 8480 6888 8488 6952
rect 8552 6888 8808 6952
rect 8872 6888 8880 6952
rect 8480 6880 8880 6888
rect 8960 6952 9360 6960
rect 8960 6888 8968 6952
rect 9032 6888 9288 6952
rect 9352 6888 9360 6952
rect 8960 6880 9360 6888
rect 9440 6952 11440 6960
rect 9440 6888 9448 6952
rect 9512 6888 9768 6952
rect 9832 6888 10088 6952
rect 10152 6888 10408 6952
rect 10472 6888 10728 6952
rect 10792 6888 11048 6952
rect 11112 6888 11368 6952
rect 11432 6888 11440 6952
rect 9440 6880 11440 6888
rect 11520 6952 11920 6960
rect 11520 6888 11528 6952
rect 11592 6888 11848 6952
rect 11912 6888 11920 6952
rect 11520 6880 11920 6888
rect 12000 6952 12400 6960
rect 12000 6888 12008 6952
rect 12072 6888 12328 6952
rect 12392 6888 12400 6952
rect 12000 6880 12400 6888
rect 8480 6792 8880 6800
rect 8480 6728 8488 6792
rect 8552 6728 8808 6792
rect 8872 6728 8880 6792
rect 8480 6720 8880 6728
rect 8960 6792 9360 6800
rect 8960 6728 8968 6792
rect 9032 6728 9288 6792
rect 9352 6728 9360 6792
rect 8960 6720 9360 6728
rect 9440 6792 11440 6800
rect 9440 6728 9448 6792
rect 9512 6728 9768 6792
rect 9832 6728 10088 6792
rect 10152 6728 10408 6792
rect 10472 6728 10728 6792
rect 10792 6728 11048 6792
rect 11112 6728 11368 6792
rect 11432 6728 11440 6792
rect 9440 6720 11440 6728
rect 11520 6792 11920 6800
rect 11520 6728 11528 6792
rect 11592 6728 11848 6792
rect 11912 6728 11920 6792
rect 11520 6720 11920 6728
rect 12000 6792 12400 6800
rect 12000 6728 12008 6792
rect 12072 6728 12328 6792
rect 12392 6728 12400 6792
rect 12000 6720 12400 6728
rect 8480 6632 8880 6640
rect 8480 6568 8488 6632
rect 8552 6568 8808 6632
rect 8872 6568 8880 6632
rect 8480 6560 8880 6568
rect 8960 6632 9360 6640
rect 8960 6568 8968 6632
rect 9032 6568 9288 6632
rect 9352 6568 9360 6632
rect 8960 6560 9360 6568
rect 9440 6632 11440 6640
rect 9440 6568 9448 6632
rect 9512 6568 9768 6632
rect 9832 6568 10088 6632
rect 10152 6568 10408 6632
rect 10472 6568 10728 6632
rect 10792 6568 11048 6632
rect 11112 6568 11368 6632
rect 11432 6568 11440 6632
rect 9440 6560 11440 6568
rect 11520 6632 11920 6640
rect 11520 6568 11528 6632
rect 11592 6568 11848 6632
rect 11912 6568 11920 6632
rect 11520 6560 11920 6568
rect 12000 6632 12400 6640
rect 12000 6568 12008 6632
rect 12072 6568 12328 6632
rect 12392 6568 12400 6632
rect 12000 6560 12400 6568
rect 8480 6472 8880 6480
rect 8480 6408 8488 6472
rect 8552 6408 8808 6472
rect 8872 6408 8880 6472
rect 8480 6400 8880 6408
rect 8960 6472 9360 6480
rect 8960 6408 8968 6472
rect 9032 6408 9288 6472
rect 9352 6408 9360 6472
rect 8960 6400 9360 6408
rect 9440 6472 11440 6480
rect 9440 6408 9448 6472
rect 9512 6408 9768 6472
rect 9832 6408 10088 6472
rect 10152 6408 10408 6472
rect 10472 6408 10728 6472
rect 10792 6408 11048 6472
rect 11112 6408 11368 6472
rect 11432 6408 11440 6472
rect 9440 6400 11440 6408
rect 11520 6472 11920 6480
rect 11520 6408 11528 6472
rect 11592 6408 11848 6472
rect 11912 6408 11920 6472
rect 11520 6400 11920 6408
rect 12000 6472 12400 6480
rect 12000 6408 12008 6472
rect 12072 6408 12328 6472
rect 12392 6408 12400 6472
rect 12000 6400 12400 6408
rect 8480 6312 8880 6320
rect 8480 6248 8488 6312
rect 8552 6248 8808 6312
rect 8872 6248 8880 6312
rect 8480 6240 8880 6248
rect 8960 6312 9360 6320
rect 8960 6248 8968 6312
rect 9032 6248 9288 6312
rect 9352 6248 9360 6312
rect 8960 6240 9360 6248
rect 9440 6312 11440 6320
rect 9440 6248 9448 6312
rect 9512 6248 9768 6312
rect 9832 6248 10088 6312
rect 10152 6248 10408 6312
rect 10472 6248 10728 6312
rect 10792 6248 11048 6312
rect 11112 6248 11368 6312
rect 11432 6248 11440 6312
rect 9440 6240 11440 6248
rect 11520 6312 11920 6320
rect 11520 6248 11528 6312
rect 11592 6248 11848 6312
rect 11912 6248 11920 6312
rect 11520 6240 11920 6248
rect 12000 6312 12400 6320
rect 12000 6248 12008 6312
rect 12072 6248 12328 6312
rect 12392 6248 12400 6312
rect 12000 6240 12400 6248
rect 8480 6152 8880 6160
rect 8480 6088 8488 6152
rect 8552 6088 8808 6152
rect 8872 6088 8880 6152
rect 8480 6080 8880 6088
rect 8960 6152 9360 6160
rect 8960 6088 8968 6152
rect 9032 6088 9288 6152
rect 9352 6088 9360 6152
rect 8960 6080 9360 6088
rect 9440 6152 11440 6160
rect 9440 6088 9448 6152
rect 9512 6088 9768 6152
rect 9832 6088 10088 6152
rect 10152 6088 10408 6152
rect 10472 6088 10728 6152
rect 10792 6088 11048 6152
rect 11112 6088 11368 6152
rect 11432 6088 11440 6152
rect 9440 6080 11440 6088
rect 11520 6152 11920 6160
rect 11520 6088 11528 6152
rect 11592 6088 11848 6152
rect 11912 6088 11920 6152
rect 11520 6080 11920 6088
rect 12000 6152 12400 6160
rect 12000 6088 12008 6152
rect 12072 6088 12328 6152
rect 12392 6088 12400 6152
rect 12000 6080 12400 6088
rect 8480 5992 8880 6000
rect 8480 5928 8488 5992
rect 8552 5928 8808 5992
rect 8872 5928 8880 5992
rect 8480 5920 8880 5928
rect 8960 5992 9360 6000
rect 8960 5928 8968 5992
rect 9032 5928 9288 5992
rect 9352 5928 9360 5992
rect 8960 5920 9360 5928
rect 9440 5992 11440 6000
rect 9440 5928 9448 5992
rect 9512 5928 9768 5992
rect 9832 5928 10088 5992
rect 10152 5928 10408 5992
rect 10472 5928 10728 5992
rect 10792 5928 11048 5992
rect 11112 5928 11368 5992
rect 11432 5928 11440 5992
rect 9440 5920 11440 5928
rect 11520 5992 11920 6000
rect 11520 5928 11528 5992
rect 11592 5928 11848 5992
rect 11912 5928 11920 5992
rect 11520 5920 11920 5928
rect 12000 5992 12400 6000
rect 12000 5928 12008 5992
rect 12072 5928 12328 5992
rect 12392 5928 12400 5992
rect 12000 5920 12400 5928
rect 8480 5832 8880 5840
rect 8480 5768 8488 5832
rect 8552 5768 8808 5832
rect 8872 5768 8880 5832
rect 8480 5760 8880 5768
rect 8960 5832 9360 5840
rect 8960 5768 8968 5832
rect 9032 5768 9288 5832
rect 9352 5768 9360 5832
rect 8960 5760 9360 5768
rect 9440 5832 11440 5840
rect 9440 5768 9448 5832
rect 9512 5768 9768 5832
rect 9832 5768 10088 5832
rect 10152 5768 10408 5832
rect 10472 5768 10728 5832
rect 10792 5768 11048 5832
rect 11112 5768 11368 5832
rect 11432 5768 11440 5832
rect 9440 5760 11440 5768
rect 11520 5832 11920 5840
rect 11520 5768 11528 5832
rect 11592 5768 11848 5832
rect 11912 5768 11920 5832
rect 11520 5760 11920 5768
rect 12000 5832 12400 5840
rect 12000 5768 12008 5832
rect 12072 5768 12328 5832
rect 12392 5768 12400 5832
rect 12000 5760 12400 5768
rect 8480 5672 8880 5680
rect 8480 5608 8488 5672
rect 8552 5608 8808 5672
rect 8872 5608 8880 5672
rect 8480 5600 8880 5608
rect 8960 5672 9360 5680
rect 8960 5608 8968 5672
rect 9032 5608 9288 5672
rect 9352 5608 9360 5672
rect 8960 5600 9360 5608
rect 9440 5672 11440 5680
rect 9440 5608 9448 5672
rect 9512 5608 9768 5672
rect 9832 5608 10088 5672
rect 10152 5608 10408 5672
rect 10472 5608 10728 5672
rect 10792 5608 11048 5672
rect 11112 5608 11368 5672
rect 11432 5608 11440 5672
rect 9440 5600 11440 5608
rect 11520 5672 11920 5680
rect 11520 5608 11528 5672
rect 11592 5608 11848 5672
rect 11912 5608 11920 5672
rect 11520 5600 11920 5608
rect 12000 5672 12400 5680
rect 12000 5608 12008 5672
rect 12072 5608 12328 5672
rect 12392 5608 12400 5672
rect 12000 5600 12400 5608
rect 8480 5512 8880 5520
rect 8480 5448 8488 5512
rect 8552 5448 8808 5512
rect 8872 5448 8880 5512
rect 8480 5440 8880 5448
rect 8960 5512 9360 5520
rect 8960 5448 8968 5512
rect 9032 5448 9288 5512
rect 9352 5448 9360 5512
rect 8960 5440 9360 5448
rect 9440 5512 11440 5520
rect 9440 5448 9448 5512
rect 9512 5448 9768 5512
rect 9832 5448 10088 5512
rect 10152 5448 10408 5512
rect 10472 5448 10728 5512
rect 10792 5448 11048 5512
rect 11112 5448 11368 5512
rect 11432 5448 11440 5512
rect 9440 5440 11440 5448
rect 11520 5512 11920 5520
rect 11520 5448 11528 5512
rect 11592 5448 11848 5512
rect 11912 5448 11920 5512
rect 11520 5440 11920 5448
rect 12000 5512 12400 5520
rect 12000 5448 12008 5512
rect 12072 5448 12328 5512
rect 12392 5448 12400 5512
rect 12000 5440 12400 5448
rect 8480 5352 8880 5360
rect 8480 5288 8488 5352
rect 8552 5288 8808 5352
rect 8872 5288 8880 5352
rect 8480 5280 8880 5288
rect 8960 5352 9360 5360
rect 8960 5288 8968 5352
rect 9032 5288 9288 5352
rect 9352 5288 9360 5352
rect 8960 5280 9360 5288
rect 9440 5352 11440 5360
rect 9440 5288 9448 5352
rect 9512 5288 9768 5352
rect 9832 5288 10088 5352
rect 10152 5288 10408 5352
rect 10472 5288 10728 5352
rect 10792 5288 11048 5352
rect 11112 5288 11368 5352
rect 11432 5288 11440 5352
rect 9440 5280 11440 5288
rect 11520 5352 11920 5360
rect 11520 5288 11528 5352
rect 11592 5288 11848 5352
rect 11912 5288 11920 5352
rect 11520 5280 11920 5288
rect 12000 5352 12400 5360
rect 12000 5288 12008 5352
rect 12072 5288 12328 5352
rect 12392 5288 12400 5352
rect 12000 5280 12400 5288
rect 8480 5192 8880 5200
rect 8480 5128 8488 5192
rect 8552 5128 8808 5192
rect 8872 5128 8880 5192
rect 8480 5120 8880 5128
rect 8960 5192 9360 5200
rect 8960 5128 8968 5192
rect 9032 5128 9288 5192
rect 9352 5128 9360 5192
rect 8960 5120 9360 5128
rect 9440 5192 11440 5200
rect 9440 5128 9448 5192
rect 9512 5128 9768 5192
rect 9832 5128 10088 5192
rect 10152 5128 10408 5192
rect 10472 5128 10728 5192
rect 10792 5128 11048 5192
rect 11112 5128 11368 5192
rect 11432 5128 11440 5192
rect 9440 5120 11440 5128
rect 11520 5192 11920 5200
rect 11520 5128 11528 5192
rect 11592 5128 11848 5192
rect 11912 5128 11920 5192
rect 11520 5120 11920 5128
rect 12000 5192 12400 5200
rect 12000 5128 12008 5192
rect 12072 5128 12328 5192
rect 12392 5128 12400 5192
rect 12000 5120 12400 5128
rect 8480 5032 8880 5040
rect 8480 4968 8488 5032
rect 8552 4968 8808 5032
rect 8872 4968 8880 5032
rect 8480 4960 8880 4968
rect 8960 5032 9360 5040
rect 8960 4968 8968 5032
rect 9032 4968 9288 5032
rect 9352 4968 9360 5032
rect 8960 4960 9360 4968
rect 9440 5032 11440 5040
rect 9440 4968 9448 5032
rect 9512 4968 9768 5032
rect 9832 4968 10088 5032
rect 10152 4968 10408 5032
rect 10472 4968 10728 5032
rect 10792 4968 11048 5032
rect 11112 4968 11368 5032
rect 11432 4968 11440 5032
rect 9440 4960 11440 4968
rect 11520 5032 11920 5040
rect 11520 4968 11528 5032
rect 11592 4968 11848 5032
rect 11912 4968 11920 5032
rect 11520 4960 11920 4968
rect 12000 5032 12400 5040
rect 12000 4968 12008 5032
rect 12072 4968 12328 5032
rect 12392 4968 12400 5032
rect 12000 4960 12400 4968
rect 8480 4872 8880 4880
rect 8480 4808 8488 4872
rect 8552 4808 8808 4872
rect 8872 4808 8880 4872
rect 8480 4800 8880 4808
rect 8960 4872 9360 4880
rect 8960 4808 8968 4872
rect 9032 4808 9288 4872
rect 9352 4808 9360 4872
rect 8960 4800 9360 4808
rect 9440 4872 11440 4880
rect 9440 4808 9448 4872
rect 9512 4808 9768 4872
rect 9832 4808 10088 4872
rect 10152 4808 10408 4872
rect 10472 4808 10728 4872
rect 10792 4808 11048 4872
rect 11112 4808 11368 4872
rect 11432 4808 11440 4872
rect 9440 4800 11440 4808
rect 11520 4872 11920 4880
rect 11520 4808 11528 4872
rect 11592 4808 11848 4872
rect 11912 4808 11920 4872
rect 11520 4800 11920 4808
rect 12000 4872 12400 4880
rect 12000 4808 12008 4872
rect 12072 4808 12328 4872
rect 12392 4808 12400 4872
rect 12000 4800 12400 4808
rect 8480 4712 8880 4720
rect 8480 4648 8488 4712
rect 8552 4648 8808 4712
rect 8872 4648 8880 4712
rect 8480 4640 8880 4648
rect 8960 4712 9360 4720
rect 8960 4648 8968 4712
rect 9032 4648 9288 4712
rect 9352 4648 9360 4712
rect 8960 4640 9360 4648
rect 9440 4712 11440 4720
rect 9440 4648 9448 4712
rect 9512 4648 9768 4712
rect 9832 4648 10088 4712
rect 10152 4648 10408 4712
rect 10472 4648 10728 4712
rect 10792 4648 11048 4712
rect 11112 4648 11368 4712
rect 11432 4648 11440 4712
rect 9440 4640 11440 4648
rect 11520 4712 11920 4720
rect 11520 4648 11528 4712
rect 11592 4648 11848 4712
rect 11912 4648 11920 4712
rect 11520 4640 11920 4648
rect 12000 4712 12400 4720
rect 12000 4648 12008 4712
rect 12072 4648 12328 4712
rect 12392 4648 12400 4712
rect 12000 4640 12400 4648
rect 8480 4552 8880 4560
rect 8480 4488 8488 4552
rect 8552 4488 8808 4552
rect 8872 4488 8880 4552
rect 8480 4480 8880 4488
rect 8960 4552 9360 4560
rect 8960 4488 8968 4552
rect 9032 4488 9288 4552
rect 9352 4488 9360 4552
rect 8960 4480 9360 4488
rect 9440 4552 11440 4560
rect 9440 4488 9448 4552
rect 9512 4488 9768 4552
rect 9832 4488 10088 4552
rect 10152 4488 10408 4552
rect 10472 4488 10728 4552
rect 10792 4488 11048 4552
rect 11112 4488 11368 4552
rect 11432 4488 11440 4552
rect 9440 4480 11440 4488
rect 11520 4552 11920 4560
rect 11520 4488 11528 4552
rect 11592 4488 11848 4552
rect 11912 4488 11920 4552
rect 11520 4480 11920 4488
rect 12000 4552 12400 4560
rect 12000 4488 12008 4552
rect 12072 4488 12328 4552
rect 12392 4488 12400 4552
rect 12000 4480 12400 4488
rect 8480 4392 8880 4400
rect 8480 4328 8488 4392
rect 8552 4328 8808 4392
rect 8872 4328 8880 4392
rect 8480 4320 8880 4328
rect 8960 4392 9360 4400
rect 8960 4328 8968 4392
rect 9032 4328 9288 4392
rect 9352 4328 9360 4392
rect 8960 4320 9360 4328
rect 9440 4392 11440 4400
rect 9440 4328 9448 4392
rect 9512 4328 9768 4392
rect 9832 4328 10088 4392
rect 10152 4328 10408 4392
rect 10472 4328 10728 4392
rect 10792 4328 11048 4392
rect 11112 4328 11368 4392
rect 11432 4328 11440 4392
rect 9440 4320 11440 4328
rect 11520 4392 11920 4400
rect 11520 4328 11528 4392
rect 11592 4328 11848 4392
rect 11912 4328 11920 4392
rect 11520 4320 11920 4328
rect 12000 4392 12400 4400
rect 12000 4328 12008 4392
rect 12072 4328 12328 4392
rect 12392 4328 12400 4392
rect 12000 4320 12400 4328
rect 8480 4232 8880 4240
rect 8480 4168 8488 4232
rect 8552 4168 8808 4232
rect 8872 4168 8880 4232
rect 8480 4160 8880 4168
rect 8960 4232 9360 4240
rect 8960 4168 8968 4232
rect 9032 4168 9288 4232
rect 9352 4168 9360 4232
rect 8960 4160 9360 4168
rect 9440 4232 11440 4240
rect 9440 4168 9448 4232
rect 9512 4168 9768 4232
rect 9832 4168 10088 4232
rect 10152 4168 10408 4232
rect 10472 4168 10728 4232
rect 10792 4168 11048 4232
rect 11112 4168 11368 4232
rect 11432 4168 11440 4232
rect 9440 4160 11440 4168
rect 11520 4232 11920 4240
rect 11520 4168 11528 4232
rect 11592 4168 11848 4232
rect 11912 4168 11920 4232
rect 11520 4160 11920 4168
rect 12000 4232 12400 4240
rect 12000 4168 12008 4232
rect 12072 4168 12328 4232
rect 12392 4168 12400 4232
rect 12000 4160 12400 4168
rect 8480 4072 8880 4080
rect 8480 4008 8488 4072
rect 8552 4008 8808 4072
rect 8872 4008 8880 4072
rect 8480 4000 8880 4008
rect 8960 4072 9360 4080
rect 8960 4008 8968 4072
rect 9032 4008 9288 4072
rect 9352 4008 9360 4072
rect 8960 4000 9360 4008
rect 9440 4072 11440 4080
rect 9440 4008 9448 4072
rect 9512 4008 9768 4072
rect 9832 4008 10088 4072
rect 10152 4008 10408 4072
rect 10472 4008 10728 4072
rect 10792 4008 11048 4072
rect 11112 4008 11368 4072
rect 11432 4008 11440 4072
rect 9440 4000 11440 4008
rect 11520 4072 11920 4080
rect 11520 4008 11528 4072
rect 11592 4008 11848 4072
rect 11912 4008 11920 4072
rect 11520 4000 11920 4008
rect 12000 4072 12400 4080
rect 12000 4008 12008 4072
rect 12072 4008 12328 4072
rect 12392 4008 12400 4072
rect 12000 4000 12400 4008
rect 8480 3912 8880 3920
rect 8480 3848 8488 3912
rect 8552 3848 8808 3912
rect 8872 3848 8880 3912
rect 8480 3840 8880 3848
rect 8960 3912 9360 3920
rect 8960 3848 8968 3912
rect 9032 3848 9288 3912
rect 9352 3848 9360 3912
rect 8960 3840 9360 3848
rect 9440 3912 11440 3920
rect 9440 3848 9448 3912
rect 9512 3848 9768 3912
rect 9832 3848 10088 3912
rect 10152 3848 10408 3912
rect 10472 3848 10728 3912
rect 10792 3848 11048 3912
rect 11112 3848 11368 3912
rect 11432 3848 11440 3912
rect 9440 3840 11440 3848
rect 11520 3912 11920 3920
rect 11520 3848 11528 3912
rect 11592 3848 11848 3912
rect 11912 3848 11920 3912
rect 11520 3840 11920 3848
rect 12000 3912 12400 3920
rect 12000 3848 12008 3912
rect 12072 3848 12328 3912
rect 12392 3848 12400 3912
rect 12000 3840 12400 3848
rect 8480 3752 8880 3760
rect 8480 3688 8488 3752
rect 8552 3688 8808 3752
rect 8872 3688 8880 3752
rect 8480 3680 8880 3688
rect 8960 3752 9360 3760
rect 8960 3688 8968 3752
rect 9032 3688 9288 3752
rect 9352 3688 9360 3752
rect 8960 3680 9360 3688
rect 9440 3752 11440 3760
rect 9440 3688 9448 3752
rect 9512 3688 9768 3752
rect 9832 3688 10088 3752
rect 10152 3688 10408 3752
rect 10472 3688 10728 3752
rect 10792 3688 11048 3752
rect 11112 3688 11368 3752
rect 11432 3688 11440 3752
rect 9440 3680 11440 3688
rect 11520 3752 11920 3760
rect 11520 3688 11528 3752
rect 11592 3688 11848 3752
rect 11912 3688 11920 3752
rect 11520 3680 11920 3688
rect 12000 3752 12400 3760
rect 12000 3688 12008 3752
rect 12072 3688 12328 3752
rect 12392 3688 12400 3752
rect 12000 3680 12400 3688
rect 8480 3592 8880 3600
rect 8480 3528 8488 3592
rect 8552 3528 8808 3592
rect 8872 3528 8880 3592
rect 8480 3520 8880 3528
rect 8960 3592 9360 3600
rect 8960 3528 8968 3592
rect 9032 3528 9288 3592
rect 9352 3528 9360 3592
rect 8960 3520 9360 3528
rect 9440 3592 11440 3600
rect 9440 3528 9448 3592
rect 9512 3528 9768 3592
rect 9832 3528 10088 3592
rect 10152 3528 10408 3592
rect 10472 3528 10728 3592
rect 10792 3528 11048 3592
rect 11112 3528 11368 3592
rect 11432 3528 11440 3592
rect 9440 3520 11440 3528
rect 11520 3592 11920 3600
rect 11520 3528 11528 3592
rect 11592 3528 11848 3592
rect 11912 3528 11920 3592
rect 11520 3520 11920 3528
rect 12000 3592 12400 3600
rect 12000 3528 12008 3592
rect 12072 3528 12328 3592
rect 12392 3528 12400 3592
rect 12000 3520 12400 3528
rect 8480 3432 8880 3440
rect 8480 3368 8488 3432
rect 8552 3368 8808 3432
rect 8872 3368 8880 3432
rect 8480 3360 8880 3368
rect 8960 3432 9360 3440
rect 8960 3368 8968 3432
rect 9032 3368 9288 3432
rect 9352 3368 9360 3432
rect 8960 3360 9360 3368
rect 9440 3432 11440 3440
rect 9440 3368 9448 3432
rect 9512 3368 9768 3432
rect 9832 3368 10088 3432
rect 10152 3368 10408 3432
rect 10472 3368 10728 3432
rect 10792 3368 11048 3432
rect 11112 3368 11368 3432
rect 11432 3368 11440 3432
rect 9440 3360 11440 3368
rect 11520 3432 11920 3440
rect 11520 3368 11528 3432
rect 11592 3368 11848 3432
rect 11912 3368 11920 3432
rect 11520 3360 11920 3368
rect 12000 3432 12400 3440
rect 12000 3368 12008 3432
rect 12072 3368 12328 3432
rect 12392 3368 12400 3432
rect 12000 3360 12400 3368
rect 8480 3272 8880 3280
rect 8480 3208 8488 3272
rect 8552 3208 8808 3272
rect 8872 3208 8880 3272
rect 8480 3200 8880 3208
rect 8960 3272 9360 3280
rect 8960 3208 8968 3272
rect 9032 3208 9288 3272
rect 9352 3208 9360 3272
rect 8960 3200 9360 3208
rect 9440 3272 11440 3280
rect 9440 3208 9448 3272
rect 9512 3208 9768 3272
rect 9832 3208 10088 3272
rect 10152 3208 10408 3272
rect 10472 3208 10728 3272
rect 10792 3208 11048 3272
rect 11112 3208 11368 3272
rect 11432 3208 11440 3272
rect 9440 3200 11440 3208
rect 11520 3272 11920 3280
rect 11520 3208 11528 3272
rect 11592 3208 11848 3272
rect 11912 3208 11920 3272
rect 11520 3200 11920 3208
rect 12000 3272 12400 3280
rect 12000 3208 12008 3272
rect 12072 3208 12328 3272
rect 12392 3208 12400 3272
rect 12000 3200 12400 3208
rect 8480 3112 8880 3120
rect 8480 3048 8488 3112
rect 8552 3048 8808 3112
rect 8872 3048 8880 3112
rect 8480 3040 8880 3048
rect 8960 3112 9360 3120
rect 8960 3048 8968 3112
rect 9032 3048 9288 3112
rect 9352 3048 9360 3112
rect 8960 3040 9360 3048
rect 9440 3112 11440 3120
rect 9440 3048 9448 3112
rect 9512 3048 9768 3112
rect 9832 3048 10088 3112
rect 10152 3048 10408 3112
rect 10472 3048 10728 3112
rect 10792 3048 11048 3112
rect 11112 3048 11368 3112
rect 11432 3048 11440 3112
rect 9440 3040 11440 3048
rect 11520 3112 11920 3120
rect 11520 3048 11528 3112
rect 11592 3048 11848 3112
rect 11912 3048 11920 3112
rect 11520 3040 11920 3048
rect 12000 3112 12400 3120
rect 12000 3048 12008 3112
rect 12072 3048 12328 3112
rect 12392 3048 12400 3112
rect 12000 3040 12400 3048
rect 8480 2952 8880 2960
rect 8480 2888 8488 2952
rect 8552 2888 8808 2952
rect 8872 2888 8880 2952
rect 8480 2880 8880 2888
rect 8960 2952 9360 2960
rect 8960 2888 8968 2952
rect 9032 2888 9288 2952
rect 9352 2888 9360 2952
rect 8960 2880 9360 2888
rect 9440 2952 11440 2960
rect 9440 2888 9448 2952
rect 9512 2888 9768 2952
rect 9832 2888 10088 2952
rect 10152 2888 10408 2952
rect 10472 2888 10728 2952
rect 10792 2888 11048 2952
rect 11112 2888 11368 2952
rect 11432 2888 11440 2952
rect 9440 2880 11440 2888
rect 11520 2952 11920 2960
rect 11520 2888 11528 2952
rect 11592 2888 11848 2952
rect 11912 2888 11920 2952
rect 11520 2880 11920 2888
rect 12000 2952 12400 2960
rect 12000 2888 12008 2952
rect 12072 2888 12328 2952
rect 12392 2888 12400 2952
rect 12000 2880 12400 2888
rect 8480 2792 8880 2800
rect 8480 2728 8488 2792
rect 8552 2728 8808 2792
rect 8872 2728 8880 2792
rect 8480 2720 8880 2728
rect 8960 2792 9360 2800
rect 8960 2728 8968 2792
rect 9032 2728 9288 2792
rect 9352 2728 9360 2792
rect 8960 2720 9360 2728
rect 9440 2792 11440 2800
rect 9440 2728 9448 2792
rect 9512 2728 9768 2792
rect 9832 2728 10088 2792
rect 10152 2728 10408 2792
rect 10472 2728 10728 2792
rect 10792 2728 11048 2792
rect 11112 2728 11368 2792
rect 11432 2728 11440 2792
rect 9440 2720 11440 2728
rect 11520 2792 11920 2800
rect 11520 2728 11528 2792
rect 11592 2728 11848 2792
rect 11912 2728 11920 2792
rect 11520 2720 11920 2728
rect 12000 2792 12400 2800
rect 12000 2728 12008 2792
rect 12072 2728 12328 2792
rect 12392 2728 12400 2792
rect 12000 2720 12400 2728
rect 8480 2632 8880 2640
rect 8480 2568 8488 2632
rect 8552 2568 8808 2632
rect 8872 2568 8880 2632
rect 8480 2560 8880 2568
rect 8960 2632 9360 2640
rect 8960 2568 8968 2632
rect 9032 2568 9288 2632
rect 9352 2568 9360 2632
rect 8960 2560 9360 2568
rect 9440 2632 11440 2640
rect 9440 2568 9448 2632
rect 9512 2568 9768 2632
rect 9832 2568 10088 2632
rect 10152 2568 10408 2632
rect 10472 2568 10728 2632
rect 10792 2568 11048 2632
rect 11112 2568 11368 2632
rect 11432 2568 11440 2632
rect 9440 2560 11440 2568
rect 11520 2632 11920 2640
rect 11520 2568 11528 2632
rect 11592 2568 11848 2632
rect 11912 2568 11920 2632
rect 11520 2560 11920 2568
rect 12000 2632 12400 2640
rect 12000 2568 12008 2632
rect 12072 2568 12328 2632
rect 12392 2568 12400 2632
rect 12000 2560 12400 2568
rect 8480 2472 8880 2480
rect 8480 2408 8488 2472
rect 8552 2408 8808 2472
rect 8872 2408 8880 2472
rect 8480 2400 8880 2408
rect 8960 2472 9360 2480
rect 8960 2408 8968 2472
rect 9032 2408 9288 2472
rect 9352 2408 9360 2472
rect 8960 2400 9360 2408
rect 9440 2472 11440 2480
rect 9440 2408 9448 2472
rect 9512 2408 9768 2472
rect 9832 2408 10088 2472
rect 10152 2408 10408 2472
rect 10472 2408 10728 2472
rect 10792 2408 11048 2472
rect 11112 2408 11368 2472
rect 11432 2408 11440 2472
rect 9440 2400 11440 2408
rect 11520 2472 11920 2480
rect 11520 2408 11528 2472
rect 11592 2408 11848 2472
rect 11912 2408 11920 2472
rect 11520 2400 11920 2408
rect 12000 2472 12400 2480
rect 12000 2408 12008 2472
rect 12072 2408 12328 2472
rect 12392 2408 12400 2472
rect 12000 2400 12400 2408
rect 8480 2312 8880 2320
rect 8480 2248 8488 2312
rect 8552 2248 8808 2312
rect 8872 2248 8880 2312
rect 8480 2240 8880 2248
rect 8960 2312 9360 2320
rect 8960 2248 8968 2312
rect 9032 2248 9288 2312
rect 9352 2248 9360 2312
rect 8960 2240 9360 2248
rect 9440 2312 11440 2320
rect 9440 2248 9448 2312
rect 9512 2248 9768 2312
rect 9832 2248 10088 2312
rect 10152 2248 10408 2312
rect 10472 2248 10728 2312
rect 10792 2248 11048 2312
rect 11112 2248 11368 2312
rect 11432 2248 11440 2312
rect 9440 2240 11440 2248
rect 11520 2312 11920 2320
rect 11520 2248 11528 2312
rect 11592 2248 11848 2312
rect 11912 2248 11920 2312
rect 11520 2240 11920 2248
rect 12000 2312 12400 2320
rect 12000 2248 12008 2312
rect 12072 2248 12328 2312
rect 12392 2248 12400 2312
rect 12000 2240 12400 2248
rect 8480 2152 8880 2160
rect 8480 2088 8488 2152
rect 8552 2088 8808 2152
rect 8872 2088 8880 2152
rect 8480 2080 8880 2088
rect 8960 2152 9360 2160
rect 8960 2088 8968 2152
rect 9032 2088 9288 2152
rect 9352 2088 9360 2152
rect 8960 2080 9360 2088
rect 9440 2152 11440 2160
rect 9440 2088 9448 2152
rect 9512 2088 9768 2152
rect 9832 2088 10088 2152
rect 10152 2088 10408 2152
rect 10472 2088 10728 2152
rect 10792 2088 11048 2152
rect 11112 2088 11368 2152
rect 11432 2088 11440 2152
rect 9440 2080 11440 2088
rect 11520 2152 11920 2160
rect 11520 2088 11528 2152
rect 11592 2088 11848 2152
rect 11912 2088 11920 2152
rect 11520 2080 11920 2088
rect 12000 2152 12400 2160
rect 12000 2088 12008 2152
rect 12072 2088 12328 2152
rect 12392 2088 12400 2152
rect 12000 2080 12400 2088
rect 8480 1992 8880 2000
rect 8480 1928 8488 1992
rect 8552 1928 8808 1992
rect 8872 1928 8880 1992
rect 8480 1920 8880 1928
rect 8960 1992 9360 2000
rect 8960 1928 8968 1992
rect 9032 1928 9288 1992
rect 9352 1928 9360 1992
rect 8960 1920 9360 1928
rect 9440 1992 11440 2000
rect 9440 1928 9448 1992
rect 9512 1928 9768 1992
rect 9832 1928 10088 1992
rect 10152 1928 10408 1992
rect 10472 1928 10728 1992
rect 10792 1928 11048 1992
rect 11112 1928 11368 1992
rect 11432 1928 11440 1992
rect 9440 1920 11440 1928
rect 11520 1992 11920 2000
rect 11520 1928 11528 1992
rect 11592 1928 11848 1992
rect 11912 1928 11920 1992
rect 11520 1920 11920 1928
rect 12000 1992 12400 2000
rect 12000 1928 12008 1992
rect 12072 1928 12328 1992
rect 12392 1928 12400 1992
rect 12000 1920 12400 1928
rect 8480 1832 8880 1840
rect 8480 1768 8488 1832
rect 8552 1768 8808 1832
rect 8872 1768 8880 1832
rect 8480 1760 8880 1768
rect 8960 1832 9360 1840
rect 8960 1768 8968 1832
rect 9032 1768 9288 1832
rect 9352 1768 9360 1832
rect 8960 1760 9360 1768
rect 9440 1832 11440 1840
rect 9440 1768 9448 1832
rect 9512 1768 9768 1832
rect 9832 1768 10088 1832
rect 10152 1768 10408 1832
rect 10472 1768 10728 1832
rect 10792 1768 11048 1832
rect 11112 1768 11368 1832
rect 11432 1768 11440 1832
rect 9440 1760 11440 1768
rect 11520 1832 11920 1840
rect 11520 1768 11528 1832
rect 11592 1768 11848 1832
rect 11912 1768 11920 1832
rect 11520 1760 11920 1768
rect 12000 1832 12400 1840
rect 12000 1768 12008 1832
rect 12072 1768 12328 1832
rect 12392 1768 12400 1832
rect 12000 1760 12400 1768
rect 8480 1672 8880 1680
rect 8480 1608 8488 1672
rect 8552 1608 8808 1672
rect 8872 1608 8880 1672
rect 8480 1600 8880 1608
rect 8960 1672 9360 1680
rect 8960 1608 8968 1672
rect 9032 1608 9288 1672
rect 9352 1608 9360 1672
rect 8960 1600 9360 1608
rect 9440 1672 11440 1680
rect 9440 1608 9448 1672
rect 9512 1608 9768 1672
rect 9832 1608 10088 1672
rect 10152 1608 10408 1672
rect 10472 1608 10728 1672
rect 10792 1608 11048 1672
rect 11112 1608 11368 1672
rect 11432 1608 11440 1672
rect 9440 1600 11440 1608
rect 11520 1672 11920 1680
rect 11520 1608 11528 1672
rect 11592 1608 11848 1672
rect 11912 1608 11920 1672
rect 11520 1600 11920 1608
rect 12000 1672 12400 1680
rect 12000 1608 12008 1672
rect 12072 1608 12328 1672
rect 12392 1608 12400 1672
rect 12000 1600 12400 1608
rect 8480 1512 8880 1520
rect 8480 1448 8488 1512
rect 8552 1448 8808 1512
rect 8872 1448 8880 1512
rect 8480 1440 8880 1448
rect 8960 1512 9360 1520
rect 8960 1448 8968 1512
rect 9032 1448 9288 1512
rect 9352 1448 9360 1512
rect 8960 1440 9360 1448
rect 9440 1512 11440 1520
rect 9440 1448 9448 1512
rect 9512 1448 9768 1512
rect 9832 1448 10088 1512
rect 10152 1448 10408 1512
rect 10472 1448 10728 1512
rect 10792 1448 11048 1512
rect 11112 1448 11368 1512
rect 11432 1448 11440 1512
rect 9440 1440 11440 1448
rect 11520 1512 11920 1520
rect 11520 1448 11528 1512
rect 11592 1448 11848 1512
rect 11912 1448 11920 1512
rect 11520 1440 11920 1448
rect 12000 1512 12400 1520
rect 12000 1448 12008 1512
rect 12072 1448 12328 1512
rect 12392 1448 12400 1512
rect 12000 1440 12400 1448
rect 8480 1352 8880 1360
rect 8480 1288 8488 1352
rect 8552 1288 8808 1352
rect 8872 1288 8880 1352
rect 8480 1280 8880 1288
rect 8960 1352 9360 1360
rect 8960 1288 8968 1352
rect 9032 1288 9288 1352
rect 9352 1288 9360 1352
rect 8960 1280 9360 1288
rect 9440 1352 11440 1360
rect 9440 1288 9448 1352
rect 9512 1288 9768 1352
rect 9832 1288 10088 1352
rect 10152 1288 10408 1352
rect 10472 1288 10728 1352
rect 10792 1288 11048 1352
rect 11112 1288 11368 1352
rect 11432 1288 11440 1352
rect 9440 1280 11440 1288
rect 11520 1352 11920 1360
rect 11520 1288 11528 1352
rect 11592 1288 11848 1352
rect 11912 1288 11920 1352
rect 11520 1280 11920 1288
rect 12000 1352 12400 1360
rect 12000 1288 12008 1352
rect 12072 1288 12328 1352
rect 12392 1288 12400 1352
rect 12000 1280 12400 1288
rect 8480 1192 8880 1200
rect 8480 1128 8488 1192
rect 8552 1128 8808 1192
rect 8872 1128 8880 1192
rect 8480 1120 8880 1128
rect 8960 1192 9360 1200
rect 8960 1128 8968 1192
rect 9032 1128 9288 1192
rect 9352 1128 9360 1192
rect 8960 1120 9360 1128
rect 9440 1192 11440 1200
rect 9440 1128 9448 1192
rect 9512 1128 9768 1192
rect 9832 1128 10088 1192
rect 10152 1128 10408 1192
rect 10472 1128 10728 1192
rect 10792 1128 11048 1192
rect 11112 1128 11368 1192
rect 11432 1128 11440 1192
rect 9440 1120 11440 1128
rect 11520 1192 11920 1200
rect 11520 1128 11528 1192
rect 11592 1128 11848 1192
rect 11912 1128 11920 1192
rect 11520 1120 11920 1128
rect 12000 1192 12400 1200
rect 12000 1128 12008 1192
rect 12072 1128 12328 1192
rect 12392 1128 12400 1192
rect 12000 1120 12400 1128
rect 8480 1032 8880 1040
rect 8480 968 8488 1032
rect 8552 968 8808 1032
rect 8872 968 8880 1032
rect 8480 960 8880 968
rect 8960 1032 9360 1040
rect 8960 968 8968 1032
rect 9032 968 9288 1032
rect 9352 968 9360 1032
rect 8960 960 9360 968
rect 9440 1032 11440 1040
rect 9440 968 9448 1032
rect 9512 968 9768 1032
rect 9832 968 10088 1032
rect 10152 968 10408 1032
rect 10472 968 10728 1032
rect 10792 968 11048 1032
rect 11112 968 11368 1032
rect 11432 968 11440 1032
rect 9440 960 11440 968
rect 11520 1032 11920 1040
rect 11520 968 11528 1032
rect 11592 968 11848 1032
rect 11912 968 11920 1032
rect 11520 960 11920 968
rect 12000 1032 12400 1040
rect 12000 968 12008 1032
rect 12072 968 12328 1032
rect 12392 968 12400 1032
rect 12000 960 12400 968
rect 8480 872 8880 880
rect 8480 808 8488 872
rect 8552 808 8808 872
rect 8872 808 8880 872
rect 8480 800 8880 808
rect 8960 872 9360 880
rect 8960 808 8968 872
rect 9032 808 9288 872
rect 9352 808 9360 872
rect 8960 800 9360 808
rect 9440 872 11440 880
rect 9440 808 9448 872
rect 9512 808 9768 872
rect 9832 808 10088 872
rect 10152 808 10408 872
rect 10472 808 10728 872
rect 10792 808 11048 872
rect 11112 808 11368 872
rect 11432 808 11440 872
rect 9440 800 11440 808
rect 11520 872 11920 880
rect 11520 808 11528 872
rect 11592 808 11848 872
rect 11912 808 11920 872
rect 11520 800 11920 808
rect 12000 872 12400 880
rect 12000 808 12008 872
rect 12072 808 12328 872
rect 12392 808 12400 872
rect 12000 800 12400 808
rect 8480 712 8880 720
rect 8480 648 8488 712
rect 8552 648 8808 712
rect 8872 648 8880 712
rect 8480 640 8880 648
rect 8960 712 9360 720
rect 8960 648 8968 712
rect 9032 648 9288 712
rect 9352 648 9360 712
rect 8960 640 9360 648
rect 9440 712 11440 720
rect 9440 648 9448 712
rect 9512 648 9768 712
rect 9832 648 10088 712
rect 10152 648 10408 712
rect 10472 648 10728 712
rect 10792 648 11048 712
rect 11112 648 11368 712
rect 11432 648 11440 712
rect 9440 640 11440 648
rect 11520 712 11920 720
rect 11520 648 11528 712
rect 11592 648 11848 712
rect 11912 648 11920 712
rect 11520 640 11920 648
rect 12000 712 12400 720
rect 12000 648 12008 712
rect 12072 648 12328 712
rect 12392 648 12400 712
rect 12000 640 12400 648
rect 8480 552 8880 560
rect 8480 488 8488 552
rect 8552 488 8808 552
rect 8872 488 8880 552
rect 8480 480 8880 488
rect 8960 552 9360 560
rect 8960 488 8968 552
rect 9032 488 9288 552
rect 9352 488 9360 552
rect 8960 480 9360 488
rect 9440 552 11440 560
rect 9440 488 9448 552
rect 9512 488 9768 552
rect 9832 488 10088 552
rect 10152 488 10408 552
rect 10472 488 10728 552
rect 10792 488 11048 552
rect 11112 488 11368 552
rect 11432 488 11440 552
rect 9440 480 11440 488
rect 11520 552 11920 560
rect 11520 488 11528 552
rect 11592 488 11848 552
rect 11912 488 11920 552
rect 11520 480 11920 488
rect 12000 552 12400 560
rect 12000 488 12008 552
rect 12072 488 12328 552
rect 12392 488 12400 552
rect 12000 480 12400 488
rect 8480 392 8880 400
rect 8480 328 8488 392
rect 8552 328 8808 392
rect 8872 328 8880 392
rect 8480 320 8880 328
rect 8960 392 9360 400
rect 8960 328 8968 392
rect 9032 328 9288 392
rect 9352 328 9360 392
rect 8960 320 9360 328
rect 9440 392 11440 400
rect 9440 328 9448 392
rect 9512 328 9768 392
rect 9832 328 10088 392
rect 10152 328 10408 392
rect 10472 328 10728 392
rect 10792 328 11048 392
rect 11112 328 11368 392
rect 11432 328 11440 392
rect 9440 320 11440 328
rect 11520 392 11920 400
rect 11520 328 11528 392
rect 11592 328 11848 392
rect 11912 328 11920 392
rect 11520 320 11920 328
rect 12000 392 12400 400
rect 12000 328 12008 392
rect 12072 328 12328 392
rect 12392 328 12400 392
rect 12000 320 12400 328
rect 8480 232 8880 240
rect 8480 168 8488 232
rect 8552 168 8808 232
rect 8872 168 8880 232
rect 8480 160 8880 168
rect 8960 232 9360 240
rect 8960 168 8968 232
rect 9032 168 9288 232
rect 9352 168 9360 232
rect 8960 160 9360 168
rect 9440 232 11440 240
rect 9440 168 9448 232
rect 9512 168 9768 232
rect 9832 168 10088 232
rect 10152 168 10408 232
rect 10472 168 10728 232
rect 10792 168 11048 232
rect 11112 168 11368 232
rect 11432 168 11440 232
rect 9440 160 11440 168
rect 11520 232 11920 240
rect 11520 168 11528 232
rect 11592 168 11848 232
rect 11912 168 11920 232
rect 11520 160 11920 168
rect 12000 232 12400 240
rect 12000 168 12008 232
rect 12072 168 12328 232
rect 12392 168 12400 232
rect 12000 160 12400 168
rect 8480 72 8880 80
rect 8480 8 8488 72
rect 8552 8 8808 72
rect 8872 8 8880 72
rect 8480 0 8880 8
rect 8960 72 9360 80
rect 8960 8 8968 72
rect 9032 8 9288 72
rect 9352 8 9360 72
rect 8960 0 9360 8
rect 9440 72 11440 80
rect 9440 8 9448 72
rect 9512 8 9768 72
rect 9832 8 10088 72
rect 10152 8 10408 72
rect 10472 8 10728 72
rect 10792 8 11048 72
rect 11112 8 11368 72
rect 11432 8 11440 72
rect 9440 0 11440 8
rect 11520 72 11920 80
rect 11520 8 11528 72
rect 11592 8 11848 72
rect 11912 8 11920 72
rect 11520 0 11920 8
rect 12000 72 12400 80
rect 12000 8 12008 72
rect 12072 8 12328 72
rect 12392 8 12400 72
rect 12000 0 12400 8
rect 0 -88 20880 -80
rect 0 -152 11528 -88
rect 11592 -152 11848 -88
rect 11912 -152 20880 -88
rect 0 -162 20880 -152
rect 0 -398 242 -162
rect 478 -398 7922 -162
rect 8158 -168 12722 -162
rect 8158 -232 11528 -168
rect 11592 -232 11848 -168
rect 11912 -232 12722 -168
rect 8158 -248 12722 -232
rect 8158 -312 11528 -248
rect 11592 -312 11848 -248
rect 11912 -312 12722 -248
rect 8158 -328 12722 -312
rect 8158 -392 11528 -328
rect 11592 -392 11848 -328
rect 11912 -392 12722 -328
rect 8158 -398 12722 -392
rect 12958 -398 20402 -162
rect 20638 -398 20880 -162
rect 0 -408 20880 -398
rect 0 -472 11528 -408
rect 11592 -472 11848 -408
rect 11912 -472 20880 -408
rect 0 -480 20880 -472
rect 0 -568 20880 -560
rect 0 -632 8968 -568
rect 9032 -632 9288 -568
rect 9352 -632 20880 -568
rect 0 -642 20880 -632
rect 0 -878 1202 -642
rect 1438 -878 6962 -642
rect 7198 -648 13682 -642
rect 7198 -712 8968 -648
rect 9032 -712 9288 -648
rect 9352 -712 13682 -648
rect 7198 -728 13682 -712
rect 7198 -792 8968 -728
rect 9032 -792 9288 -728
rect 9352 -792 13682 -728
rect 7198 -808 13682 -792
rect 7198 -872 8968 -808
rect 9032 -872 9288 -808
rect 9352 -872 13682 -808
rect 7198 -878 13682 -872
rect 13918 -878 19442 -642
rect 19678 -878 20880 -642
rect 0 -888 20880 -878
rect 0 -952 8968 -888
rect 9032 -952 9288 -888
rect 9352 -952 20880 -888
rect 0 -960 20880 -952
rect 0 -1048 20880 -1040
rect 0 -1112 9448 -1048
rect 9512 -1112 9768 -1048
rect 9832 -1112 10088 -1048
rect 10152 -1112 10408 -1048
rect 10472 -1112 10728 -1048
rect 10792 -1112 11048 -1048
rect 11112 -1112 11368 -1048
rect 11432 -1112 12008 -1048
rect 12072 -1112 12328 -1048
rect 12392 -1112 20880 -1048
rect 0 -1122 20880 -1112
rect 0 -1358 2162 -1122
rect 2398 -1358 4082 -1122
rect 4318 -1358 6002 -1122
rect 6238 -1128 14642 -1122
rect 6238 -1192 9448 -1128
rect 9512 -1192 9768 -1128
rect 9832 -1192 10088 -1128
rect 10152 -1192 10408 -1128
rect 10472 -1192 10728 -1128
rect 10792 -1192 11048 -1128
rect 11112 -1192 11368 -1128
rect 11432 -1192 12008 -1128
rect 12072 -1192 12328 -1128
rect 12392 -1192 14642 -1128
rect 6238 -1208 14642 -1192
rect 6238 -1272 9448 -1208
rect 9512 -1272 9768 -1208
rect 9832 -1272 10088 -1208
rect 10152 -1272 10408 -1208
rect 10472 -1272 10728 -1208
rect 10792 -1272 11048 -1208
rect 11112 -1272 11368 -1208
rect 11432 -1272 12008 -1208
rect 12072 -1272 12328 -1208
rect 12392 -1272 14642 -1208
rect 6238 -1288 14642 -1272
rect 6238 -1352 9448 -1288
rect 9512 -1352 9768 -1288
rect 9832 -1352 10088 -1288
rect 10152 -1352 10408 -1288
rect 10472 -1352 10728 -1288
rect 10792 -1352 11048 -1288
rect 11112 -1352 11368 -1288
rect 11432 -1352 12008 -1288
rect 12072 -1352 12328 -1288
rect 12392 -1352 14642 -1288
rect 6238 -1358 14642 -1352
rect 14878 -1358 16562 -1122
rect 16798 -1358 18482 -1122
rect 18718 -1358 20880 -1122
rect 0 -1368 20880 -1358
rect 0 -1432 9448 -1368
rect 9512 -1432 9768 -1368
rect 9832 -1432 10088 -1368
rect 10152 -1432 10408 -1368
rect 10472 -1432 10728 -1368
rect 10792 -1432 11048 -1368
rect 11112 -1432 11368 -1368
rect 11432 -1432 12008 -1368
rect 12072 -1432 12328 -1368
rect 12392 -1432 20880 -1368
rect 0 -1440 20880 -1432
rect 0 -1528 20880 -1520
rect 0 -1592 8488 -1528
rect 8552 -1592 8808 -1528
rect 8872 -1592 20880 -1528
rect 0 -1602 20880 -1592
rect 0 -1838 3122 -1602
rect 3358 -1838 5042 -1602
rect 5278 -1608 15602 -1602
rect 5278 -1672 8488 -1608
rect 8552 -1672 8808 -1608
rect 8872 -1672 15602 -1608
rect 5278 -1688 15602 -1672
rect 5278 -1752 8488 -1688
rect 8552 -1752 8808 -1688
rect 8872 -1752 15602 -1688
rect 5278 -1768 15602 -1752
rect 5278 -1832 8488 -1768
rect 8552 -1832 8808 -1768
rect 8872 -1832 15602 -1768
rect 5278 -1838 15602 -1832
rect 15838 -1838 17522 -1602
rect 17758 -1838 20880 -1602
rect 0 -1848 20880 -1838
rect 0 -1912 8488 -1848
rect 8552 -1912 8808 -1848
rect 8872 -1912 20880 -1848
rect 0 -1920 20880 -1912
rect 240 -2008 20640 -2000
rect 240 -2072 248 -2008
rect 312 -2072 8968 -2008
rect 9032 -2072 9288 -2008
rect 9352 -2072 20568 -2008
rect 20632 -2072 20640 -2008
rect 240 -2080 20640 -2072
rect 400 -2168 20560 -2160
rect 400 -2232 408 -2168
rect 472 -2232 2488 -2168
rect 2552 -2232 2648 -2168
rect 2712 -2232 4728 -2168
rect 4792 -2232 4888 -2168
rect 4952 -2232 6968 -2168
rect 7032 -2232 7128 -2168
rect 7192 -2232 9208 -2168
rect 9272 -2232 9368 -2168
rect 9432 -2232 11448 -2168
rect 11512 -2232 11608 -2168
rect 11672 -2232 13688 -2168
rect 13752 -2232 13848 -2168
rect 13912 -2232 15928 -2168
rect 15992 -2232 16088 -2168
rect 16152 -2232 18168 -2168
rect 18232 -2232 18328 -2168
rect 18392 -2232 20408 -2168
rect 20472 -2232 20560 -2168
rect 400 -2240 20560 -2232
rect 400 -2488 2560 -2320
rect 400 -4312 568 -2488
rect 2392 -4312 2560 -2488
rect 400 -4480 2560 -4312
rect 400 -4560 480 -4480
rect 2480 -4560 2560 -4480
rect 2640 -2488 4800 -2320
rect 2640 -4312 2808 -2488
rect 4632 -4312 4800 -2488
rect 2640 -4480 4800 -4312
rect 2640 -4560 2720 -4480
rect 4720 -4560 4800 -4480
rect 4880 -2488 7040 -2320
rect 4880 -4312 5048 -2488
rect 6872 -4312 7040 -2488
rect 4880 -4480 7040 -4312
rect 4880 -4560 4960 -4480
rect 6960 -4560 7040 -4480
rect 7120 -2488 9280 -2320
rect 7120 -4312 7288 -2488
rect 9112 -4312 9280 -2488
rect 7120 -4480 9280 -4312
rect 7120 -4560 7200 -4480
rect 9200 -4560 9280 -4480
rect 9360 -2488 11520 -2320
rect 9360 -4312 9528 -2488
rect 11352 -4312 11520 -2488
rect 9360 -4480 11520 -4312
rect 9360 -4560 9440 -4480
rect 11440 -4560 11520 -4480
rect 11600 -2488 13760 -2320
rect 11600 -4312 11768 -2488
rect 13592 -4312 13760 -2488
rect 11600 -4480 13760 -4312
rect 11600 -4560 11680 -4480
rect 13680 -4560 13760 -4480
rect 13840 -2488 16000 -2320
rect 13840 -4312 14008 -2488
rect 15832 -4312 16000 -2488
rect 13840 -4480 16000 -4312
rect 13840 -4560 13920 -4480
rect 15920 -4560 16000 -4480
rect 16080 -2488 18240 -2320
rect 16080 -4312 16248 -2488
rect 18072 -4312 18240 -2488
rect 16080 -4480 18240 -4312
rect 16080 -4560 16160 -4480
rect 18160 -4560 18240 -4480
rect 18320 -2488 20480 -2320
rect 18320 -4312 18488 -2488
rect 20312 -4312 20480 -2488
rect 18320 -4480 20480 -4312
rect 18320 -4560 18400 -4480
rect 20400 -4560 20480 -4480
rect 240 -4568 20640 -4560
rect 240 -4632 248 -4568
rect 312 -4632 20568 -4568
rect 20632 -4632 20640 -4568
rect 240 -4640 20640 -4632
<< via4 >>
rect 242 -398 478 -162
rect 7922 -398 8158 -162
rect 12722 -398 12958 -162
rect 20402 -398 20638 -162
rect 1202 -878 1438 -642
rect 6962 -878 7198 -642
rect 13682 -878 13918 -642
rect 19442 -878 19678 -642
rect 2162 -1358 2398 -1122
rect 4082 -1358 4318 -1122
rect 6002 -1358 6238 -1122
rect 14642 -1358 14878 -1122
rect 16562 -1358 16798 -1122
rect 18482 -1358 18718 -1122
rect 3122 -1838 3358 -1602
rect 5042 -1838 5278 -1602
rect 15602 -1838 15838 -1602
rect 17522 -1838 17758 -1602
<< metal5 >>
rect 160 -162 560 31600
rect 160 -398 242 -162
rect 478 -398 560 -162
rect 160 -1920 560 -398
rect 1120 -642 1520 31600
rect 1120 -878 1202 -642
rect 1438 -878 1520 -642
rect 1120 -1920 1520 -878
rect 2080 -1122 2480 31600
rect 2080 -1358 2162 -1122
rect 2398 -1358 2480 -1122
rect 2080 -1920 2480 -1358
rect 3040 -1602 3440 31600
rect 3040 -1838 3122 -1602
rect 3358 -1838 3440 -1602
rect 3040 -1920 3440 -1838
rect 4000 -1122 4400 31600
rect 4000 -1358 4082 -1122
rect 4318 -1358 4400 -1122
rect 4000 -1920 4400 -1358
rect 4960 -1602 5360 31600
rect 4960 -1838 5042 -1602
rect 5278 -1838 5360 -1602
rect 4960 -1920 5360 -1838
rect 5920 -1122 6320 31600
rect 5920 -1358 6002 -1122
rect 6238 -1358 6320 -1122
rect 5920 -1920 6320 -1358
rect 6880 -642 7280 31600
rect 6880 -878 6962 -642
rect 7198 -878 7280 -642
rect 6880 -1920 7280 -878
rect 7840 -162 8240 31600
rect 7840 -398 7922 -162
rect 8158 -398 8240 -162
rect 7840 -1920 8240 -398
rect 12640 -162 13040 31600
rect 12640 -398 12722 -162
rect 12958 -398 13040 -162
rect 12640 -1920 13040 -398
rect 13600 -642 14000 31600
rect 13600 -878 13682 -642
rect 13918 -878 14000 -642
rect 13600 -1920 14000 -878
rect 14560 -1122 14960 31600
rect 14560 -1358 14642 -1122
rect 14878 -1358 14960 -1122
rect 14560 -1920 14960 -1358
rect 15520 -1602 15920 31600
rect 15520 -1838 15602 -1602
rect 15838 -1838 15920 -1602
rect 15520 -1920 15920 -1838
rect 16480 -1122 16880 31600
rect 16480 -1358 16562 -1122
rect 16798 -1358 16880 -1122
rect 16480 -1920 16880 -1358
rect 17440 -1602 17840 31600
rect 17440 -1838 17522 -1602
rect 17758 -1838 17840 -1602
rect 17440 -1920 17840 -1838
rect 18400 -1122 18800 31600
rect 18400 -1358 18482 -1122
rect 18718 -1358 18800 -1122
rect 18400 -1920 18800 -1358
rect 19360 -642 19760 31600
rect 19360 -878 19442 -642
rect 19678 -878 19760 -642
rect 19360 -1920 19760 -878
rect 20320 -162 20720 31600
rect 20320 -398 20402 -162
rect 20638 -398 20720 -162
rect 20320 -1920 20720 -398
use inv_bias  biasp
timestamp 1638148091
transform 1 0 0 0 1 1040
box -26 -1066 8426 10106
use inv_bias  biasm
timestamp 1638148091
transform -1 0 20880 0 1 1040
box -26 -1066 8426 10106
use inv_2_2  ap
timestamp 1638148091
transform 1 0 0 0 1 11200
box -26 -26 8426 4026
use inv_1_4  bp
timestamp 1638148091
transform 1 0 0 0 -1 19280
box -26 -26 8426 4026
use inv_1_4  cp
timestamp 1638148091
transform 1 0 0 0 1 19360
box -26 -26 8426 4026
use inv_2_2  am
timestamp 1638148091
transform -1 0 20880 0 1 11200
box -26 -26 8426 4026
use inv_1_4  bm
timestamp 1638148091
transform -1 0 20880 0 -1 19280
box -26 -26 8426 4026
use inv_1_4  cm
timestamp 1638148091
transform -1 0 20880 0 1 19360
box -26 -26 8426 4026
use inv_2_2  fp
timestamp 1638148091
transform 1 0 0 0 1 27520
box -26 -26 8426 4026
use inv_1_4  d
timestamp 1638148091
transform 1 0 0 0 -1 27440
box -26 -26 8426 4026
use inv_2_2  fm
timestamp 1638148091
transform -1 0 20880 0 1 27520
box -26 -26 8426 4026
use inv_1_4  e
timestamp 1638148091
transform -1 0 20880 0 -1 27440
box -26 -26 8426 4026
<< labels >>
rlabel metal3 s 11200 0 11280 31520 4 im
port 1 nsew
rlabel metal3 s 9600 0 9680 31520 4 ip
port 2 nsew
rlabel metal3 s 10880 0 10960 31520 4 op
port 3 nsew
rlabel metal3 s 9920 0 10000 31520 4 om
port 4 nsew
rlabel metal3 s 10240 0 10320 31520 4 x
port 5 nsew
rlabel metal3 s 10560 0 10640 31520 4 y
port 6 nsew
rlabel metal3 s 8640 0 8720 31520 4 ib
port 7 nsew
rlabel metal3 s 12160 0 12240 31520 4 q
port 8 nsew
rlabel metal3 s 11680 0 11760 31520 4 z
port 9 nsew
rlabel metal3 s 9120 0 9200 31520 4 bp
port 10 nsew
rlabel metal5 s 160 -1920 560 31520 4 vdda
port 11 nsew
rlabel metal5 s 1120 -1920 1520 31520 4 vddx
port 12 nsew
rlabel metal5 s 2080 -1920 2480 31520 4 gnda
port 13 nsew
rlabel metal5 s 3040 -1920 3440 31520 4 vssa
port 14 nsew
<< end >>
