magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< locali >>
rect -960 41897 -880 41920
rect -960 41863 -937 41897
rect -903 41863 -880 41897
rect -960 41577 -880 41863
rect -960 41543 -937 41577
rect -903 41543 -880 41577
rect -960 41520 -880 41543
rect -800 41897 -720 41920
rect -800 41863 -777 41897
rect -743 41863 -720 41897
rect -800 41577 -720 41863
rect -800 41543 -777 41577
rect -743 41543 -720 41577
rect -800 41520 -720 41543
rect -640 41897 -560 41920
rect -640 41863 -617 41897
rect -583 41863 -560 41897
rect -640 41577 -560 41863
rect -640 41543 -617 41577
rect -583 41543 -560 41577
rect -640 41520 -560 41543
rect -480 41897 -400 41920
rect -480 41863 -457 41897
rect -423 41863 -400 41897
rect -480 41577 -400 41863
rect -480 41543 -457 41577
rect -423 41543 -400 41577
rect -480 41520 -400 41543
rect -320 41897 -240 41920
rect -320 41863 -297 41897
rect -263 41863 -240 41897
rect -320 41577 -240 41863
rect -320 41543 -297 41577
rect -263 41543 -240 41577
rect -320 41520 -240 41543
rect -160 41897 -80 41920
rect -160 41863 -137 41897
rect -103 41863 -80 41897
rect -160 41577 -80 41863
rect -160 41543 -137 41577
rect -103 41543 -80 41577
rect -160 41520 -80 41543
rect 0 41897 80 41920
rect 0 41863 23 41897
rect 57 41863 80 41897
rect 0 41577 80 41863
rect 0 41543 23 41577
rect 57 41543 80 41577
rect 0 41520 80 41543
rect 76720 40617 76800 40640
rect 76720 40583 76743 40617
rect 76777 40583 76800 40617
rect 76720 40297 76800 40583
rect 76720 40263 76743 40297
rect 76777 40263 76800 40297
rect 76720 40240 76800 40263
rect 76880 40617 76960 40640
rect 76880 40583 76903 40617
rect 76937 40583 76960 40617
rect 76880 40297 76960 40583
rect 76880 40263 76903 40297
rect 76937 40263 76960 40297
rect 76880 40240 76960 40263
rect -7040 38297 -6960 38320
rect -7040 38263 -7017 38297
rect -6983 38263 -6960 38297
rect -7040 37977 -6960 38263
rect -7040 37943 -7017 37977
rect -6983 37943 -6960 37977
rect -7040 37657 -6960 37943
rect -7040 37623 -7017 37657
rect -6983 37623 -6960 37657
rect -7040 37600 -6960 37623
rect -6880 38297 -6800 38320
rect -6880 38263 -6857 38297
rect -6823 38263 -6800 38297
rect -6880 37977 -6800 38263
rect -6880 37943 -6857 37977
rect -6823 37943 -6800 37977
rect -6880 37657 -6800 37943
rect -6880 37623 -6857 37657
rect -6823 37623 -6800 37657
rect -6880 37600 -6800 37623
rect -6720 38297 -6640 38320
rect -6720 38263 -6697 38297
rect -6663 38263 -6640 38297
rect -6720 37977 -6640 38263
rect -6720 37943 -6697 37977
rect -6663 37943 -6640 37977
rect -6720 37657 -6640 37943
rect -6720 37623 -6697 37657
rect -6663 37623 -6640 37657
rect -6720 37600 -6640 37623
rect -6560 38297 -6480 38320
rect -6560 38263 -6537 38297
rect -6503 38263 -6480 38297
rect -6560 37977 -6480 38263
rect -6560 37943 -6537 37977
rect -6503 37943 -6480 37977
rect -6560 37657 -6480 37943
rect -6560 37623 -6537 37657
rect -6503 37623 -6480 37657
rect -6560 37600 -6480 37623
rect -6400 38297 -6320 38320
rect -6400 38263 -6377 38297
rect -6343 38263 -6320 38297
rect -6400 37977 -6320 38263
rect -6400 37943 -6377 37977
rect -6343 37943 -6320 37977
rect -6400 37657 -6320 37943
rect -6400 37623 -6377 37657
rect -6343 37623 -6320 37657
rect -6400 37600 -6320 37623
rect -6240 38297 -6160 38320
rect -6240 38263 -6217 38297
rect -6183 38263 -6160 38297
rect -6240 37977 -6160 38263
rect -6240 37943 -6217 37977
rect -6183 37943 -6160 37977
rect -6240 37657 -6160 37943
rect -6240 37623 -6217 37657
rect -6183 37623 -6160 37657
rect -6240 37600 -6160 37623
rect -6080 38297 -6000 38320
rect -6080 38263 -6057 38297
rect -6023 38263 -6000 38297
rect -6080 37977 -6000 38263
rect -6080 37943 -6057 37977
rect -6023 37943 -6000 37977
rect -6080 37657 -6000 37943
rect -6080 37623 -6057 37657
rect -6023 37623 -6000 37657
rect -6080 37600 -6000 37623
rect -5920 38297 -5840 38320
rect -5920 38263 -5897 38297
rect -5863 38263 -5840 38297
rect -5920 37977 -5840 38263
rect -5920 37943 -5897 37977
rect -5863 37943 -5840 37977
rect -5920 37657 -5840 37943
rect -5920 37623 -5897 37657
rect -5863 37623 -5840 37657
rect -5920 37600 -5840 37623
rect -5760 38297 -5680 38320
rect -5760 38263 -5737 38297
rect -5703 38263 -5680 38297
rect -5760 37977 -5680 38263
rect -5760 37943 -5737 37977
rect -5703 37943 -5680 37977
rect -5760 37657 -5680 37943
rect -5760 37623 -5737 37657
rect -5703 37623 -5680 37657
rect -5760 37600 -5680 37623
rect -5600 38297 -5520 38320
rect -5600 38263 -5577 38297
rect -5543 38263 -5520 38297
rect -5600 37977 -5520 38263
rect -5600 37943 -5577 37977
rect -5543 37943 -5520 37977
rect -5600 37657 -5520 37943
rect -5600 37623 -5577 37657
rect -5543 37623 -5520 37657
rect -5600 37600 -5520 37623
rect -5440 38297 -5360 38320
rect -5440 38263 -5417 38297
rect -5383 38263 -5360 38297
rect -5440 37977 -5360 38263
rect -5440 37943 -5417 37977
rect -5383 37943 -5360 37977
rect -5440 37657 -5360 37943
rect -5440 37623 -5417 37657
rect -5383 37623 -5360 37657
rect -5440 37600 -5360 37623
rect -5280 38297 -5200 38320
rect -5280 38263 -5257 38297
rect -5223 38263 -5200 38297
rect -5280 37977 -5200 38263
rect -5280 37943 -5257 37977
rect -5223 37943 -5200 37977
rect -5280 37657 -5200 37943
rect -5280 37623 -5257 37657
rect -5223 37623 -5200 37657
rect -5280 37600 -5200 37623
rect -5120 38297 -5040 38320
rect -5120 38263 -5097 38297
rect -5063 38263 -5040 38297
rect -5120 37977 -5040 38263
rect -5120 37943 -5097 37977
rect -5063 37943 -5040 37977
rect -5120 37657 -5040 37943
rect -5120 37623 -5097 37657
rect -5063 37623 -5040 37657
rect -5120 37600 -5040 37623
rect -4960 38297 -4880 38320
rect -4960 38263 -4937 38297
rect -4903 38263 -4880 38297
rect -4960 37977 -4880 38263
rect -4960 37943 -4937 37977
rect -4903 37943 -4880 37977
rect -4960 37657 -4880 37943
rect -4960 37623 -4937 37657
rect -4903 37623 -4880 37657
rect -4960 37600 -4880 37623
rect -4800 38297 -4720 38320
rect -4800 38263 -4777 38297
rect -4743 38263 -4720 38297
rect -4800 37977 -4720 38263
rect -4800 37943 -4777 37977
rect -4743 37943 -4720 37977
rect -4800 37657 -4720 37943
rect -4800 37623 -4777 37657
rect -4743 37623 -4720 37657
rect -4800 37600 -4720 37623
rect -4640 38297 -4560 38320
rect -4640 38263 -4617 38297
rect -4583 38263 -4560 38297
rect -4640 37977 -4560 38263
rect -4640 37943 -4617 37977
rect -4583 37943 -4560 37977
rect -4640 37657 -4560 37943
rect -4640 37623 -4617 37657
rect -4583 37623 -4560 37657
rect -4640 37600 -4560 37623
rect -4480 38297 -4400 38320
rect -4480 38263 -4457 38297
rect -4423 38263 -4400 38297
rect -4480 37977 -4400 38263
rect -4480 37943 -4457 37977
rect -4423 37943 -4400 37977
rect -4480 37657 -4400 37943
rect -4480 37623 -4457 37657
rect -4423 37623 -4400 37657
rect -4480 37600 -4400 37623
rect -4320 38297 -4240 38320
rect -4320 38263 -4297 38297
rect -4263 38263 -4240 38297
rect -4320 37977 -4240 38263
rect -4320 37943 -4297 37977
rect -4263 37943 -4240 37977
rect -4320 37657 -4240 37943
rect -4320 37623 -4297 37657
rect -4263 37623 -4240 37657
rect -4320 37600 -4240 37623
rect -4160 38297 -4080 38320
rect -4160 38263 -4137 38297
rect -4103 38263 -4080 38297
rect -4160 37977 -4080 38263
rect -4160 37943 -4137 37977
rect -4103 37943 -4080 37977
rect -4160 37657 -4080 37943
rect -4160 37623 -4137 37657
rect -4103 37623 -4080 37657
rect -4160 37600 -4080 37623
rect -4000 38297 -3920 38320
rect -4000 38263 -3977 38297
rect -3943 38263 -3920 38297
rect -4000 37977 -3920 38263
rect -4000 37943 -3977 37977
rect -3943 37943 -3920 37977
rect -4000 37657 -3920 37943
rect -4000 37623 -3977 37657
rect -3943 37623 -3920 37657
rect -4000 37600 -3920 37623
rect -3840 38297 -3760 38320
rect -3840 38263 -3817 38297
rect -3783 38263 -3760 38297
rect -3840 37977 -3760 38263
rect -3840 37943 -3817 37977
rect -3783 37943 -3760 37977
rect -3840 37657 -3760 37943
rect -3840 37623 -3817 37657
rect -3783 37623 -3760 37657
rect -3840 37600 -3760 37623
rect -3680 38297 -3600 38320
rect -3680 38263 -3657 38297
rect -3623 38263 -3600 38297
rect -3680 37977 -3600 38263
rect -3680 37943 -3657 37977
rect -3623 37943 -3600 37977
rect -3680 37657 -3600 37943
rect -3680 37623 -3657 37657
rect -3623 37623 -3600 37657
rect -3680 37600 -3600 37623
rect -3520 38297 -3440 38320
rect -3520 38263 -3497 38297
rect -3463 38263 -3440 38297
rect -3520 37977 -3440 38263
rect -3520 37943 -3497 37977
rect -3463 37943 -3440 37977
rect -3520 37657 -3440 37943
rect -3520 37623 -3497 37657
rect -3463 37623 -3440 37657
rect -3520 37600 -3440 37623
rect -3360 38297 -3280 38320
rect -3360 38263 -3337 38297
rect -3303 38263 -3280 38297
rect -3360 37977 -3280 38263
rect -3360 37943 -3337 37977
rect -3303 37943 -3280 37977
rect -3360 37657 -3280 37943
rect -3360 37623 -3337 37657
rect -3303 37623 -3280 37657
rect -3360 37600 -3280 37623
rect -3200 38297 -3120 38320
rect -3200 38263 -3177 38297
rect -3143 38263 -3120 38297
rect -3200 37977 -3120 38263
rect -3200 37943 -3177 37977
rect -3143 37943 -3120 37977
rect -3200 37657 -3120 37943
rect -3200 37623 -3177 37657
rect -3143 37623 -3120 37657
rect -3200 37600 -3120 37623
rect -3040 38297 -2960 38320
rect -3040 38263 -3017 38297
rect -2983 38263 -2960 38297
rect -3040 37977 -2960 38263
rect -3040 37943 -3017 37977
rect -2983 37943 -2960 37977
rect -3040 37657 -2960 37943
rect -3040 37623 -3017 37657
rect -2983 37623 -2960 37657
rect -3040 37600 -2960 37623
rect -2880 38297 -2800 38320
rect -2880 38263 -2857 38297
rect -2823 38263 -2800 38297
rect -2880 37977 -2800 38263
rect -2880 37943 -2857 37977
rect -2823 37943 -2800 37977
rect -2880 37657 -2800 37943
rect -2880 37623 -2857 37657
rect -2823 37623 -2800 37657
rect -2880 37600 -2800 37623
rect -2720 38297 -2640 38320
rect -2720 38263 -2697 38297
rect -2663 38263 -2640 38297
rect -2720 37977 -2640 38263
rect -2720 37943 -2697 37977
rect -2663 37943 -2640 37977
rect -2720 37657 -2640 37943
rect -2720 37623 -2697 37657
rect -2663 37623 -2640 37657
rect -2720 37600 -2640 37623
rect -2560 38297 -2480 38320
rect -2560 38263 -2537 38297
rect -2503 38263 -2480 38297
rect -2560 37977 -2480 38263
rect -2560 37943 -2537 37977
rect -2503 37943 -2480 37977
rect -2560 37657 -2480 37943
rect -2560 37623 -2537 37657
rect -2503 37623 -2480 37657
rect -2560 37600 -2480 37623
rect -2400 38297 -2320 38320
rect -2400 38263 -2377 38297
rect -2343 38263 -2320 38297
rect -2400 37977 -2320 38263
rect -2400 37943 -2377 37977
rect -2343 37943 -2320 37977
rect -2400 37657 -2320 37943
rect -2400 37623 -2377 37657
rect -2343 37623 -2320 37657
rect -2400 37600 -2320 37623
rect -2240 38297 -2160 38320
rect -2240 38263 -2217 38297
rect -2183 38263 -2160 38297
rect -2240 37977 -2160 38263
rect -2240 37943 -2217 37977
rect -2183 37943 -2160 37977
rect -2240 37657 -2160 37943
rect -2240 37623 -2217 37657
rect -2183 37623 -2160 37657
rect -2240 37600 -2160 37623
rect -2080 38297 -2000 38320
rect -2080 38263 -2057 38297
rect -2023 38263 -2000 38297
rect -2080 37977 -2000 38263
rect -2080 37943 -2057 37977
rect -2023 37943 -2000 37977
rect -2080 37657 -2000 37943
rect -2080 37623 -2057 37657
rect -2023 37623 -2000 37657
rect -2080 37600 -2000 37623
rect -1920 38297 -1840 38320
rect -1920 38263 -1897 38297
rect -1863 38263 -1840 38297
rect -1920 37977 -1840 38263
rect -1920 37943 -1897 37977
rect -1863 37943 -1840 37977
rect -1920 37657 -1840 37943
rect -1920 37623 -1897 37657
rect -1863 37623 -1840 37657
rect -1920 37600 -1840 37623
rect -1760 38297 -1680 38320
rect -1760 38263 -1737 38297
rect -1703 38263 -1680 38297
rect -1760 37977 -1680 38263
rect -1760 37943 -1737 37977
rect -1703 37943 -1680 37977
rect -1760 37657 -1680 37943
rect -1760 37623 -1737 37657
rect -1703 37623 -1680 37657
rect -1760 37600 -1680 37623
rect -1600 38297 -1520 38320
rect -1600 38263 -1577 38297
rect -1543 38263 -1520 38297
rect -1600 37977 -1520 38263
rect -1600 37943 -1577 37977
rect -1543 37943 -1520 37977
rect -1600 37657 -1520 37943
rect -1600 37623 -1577 37657
rect -1543 37623 -1520 37657
rect -1600 37600 -1520 37623
rect -1440 38297 -1360 38320
rect -1440 38263 -1417 38297
rect -1383 38263 -1360 38297
rect -1440 37977 -1360 38263
rect -1440 37943 -1417 37977
rect -1383 37943 -1360 37977
rect -1440 37657 -1360 37943
rect -1440 37623 -1417 37657
rect -1383 37623 -1360 37657
rect -1440 37600 -1360 37623
rect -1280 38297 -1200 38320
rect -1280 38263 -1257 38297
rect -1223 38263 -1200 38297
rect -1280 37977 -1200 38263
rect -1280 37943 -1257 37977
rect -1223 37943 -1200 37977
rect -1280 37657 -1200 37943
rect -1280 37623 -1257 37657
rect -1223 37623 -1200 37657
rect -1280 37600 -1200 37623
rect -1120 38297 -1040 38320
rect -1120 38263 -1097 38297
rect -1063 38263 -1040 38297
rect -1120 37977 -1040 38263
rect -1120 37943 -1097 37977
rect -1063 37943 -1040 37977
rect -1120 37657 -1040 37943
rect -1120 37623 -1097 37657
rect -1063 37623 -1040 37657
rect -1120 37600 -1040 37623
rect -960 38297 -880 38320
rect -960 38263 -937 38297
rect -903 38263 -880 38297
rect -960 37977 -880 38263
rect -960 37943 -937 37977
rect -903 37943 -880 37977
rect -960 37657 -880 37943
rect -960 37623 -937 37657
rect -903 37623 -880 37657
rect -960 37600 -880 37623
rect -800 38297 -720 38320
rect -800 38263 -777 38297
rect -743 38263 -720 38297
rect -800 37977 -720 38263
rect -800 37943 -777 37977
rect -743 37943 -720 37977
rect -800 37657 -720 37943
rect -800 37623 -777 37657
rect -743 37623 -720 37657
rect -800 37600 -720 37623
rect -640 38297 -560 38320
rect -640 38263 -617 38297
rect -583 38263 -560 38297
rect -640 37977 -560 38263
rect -640 37943 -617 37977
rect -583 37943 -560 37977
rect -640 37657 -560 37943
rect -640 37623 -617 37657
rect -583 37623 -560 37657
rect -640 37600 -560 37623
rect -480 38297 -400 38320
rect -480 38263 -457 38297
rect -423 38263 -400 38297
rect -480 37977 -400 38263
rect -480 37943 -457 37977
rect -423 37943 -400 37977
rect -480 37657 -400 37943
rect -480 37623 -457 37657
rect -423 37623 -400 37657
rect -480 37600 -400 37623
rect -320 38297 -240 38320
rect -320 38263 -297 38297
rect -263 38263 -240 38297
rect -320 37977 -240 38263
rect -320 37943 -297 37977
rect -263 37943 -240 37977
rect -320 37657 -240 37943
rect -320 37623 -297 37657
rect -263 37623 -240 37657
rect -320 37600 -240 37623
rect -160 38297 -80 38320
rect -160 38263 -137 38297
rect -103 38263 -80 38297
rect -160 37977 -80 38263
rect -160 37943 -137 37977
rect -103 37943 -80 37977
rect -160 37657 -80 37943
rect -160 37623 -137 37657
rect -103 37623 -80 37657
rect -160 37600 -80 37623
rect 0 38297 80 38320
rect 0 38263 23 38297
rect 57 38263 80 38297
rect 0 37977 80 38263
rect 0 37943 23 37977
rect 57 37943 80 37977
rect 0 37657 80 37943
rect 0 37623 23 37657
rect 57 37623 80 37657
rect 0 37600 80 37623
rect 76720 36617 76800 36640
rect 76720 36583 76743 36617
rect 76777 36583 76800 36617
rect 76720 36297 76800 36583
rect 76720 36263 76743 36297
rect 76777 36263 76800 36297
rect 76720 36240 76800 36263
rect 76880 36617 76960 36640
rect 76880 36583 76903 36617
rect 76937 36583 76960 36617
rect 76880 36297 76960 36583
rect 76880 36263 76903 36297
rect 76937 36263 76960 36297
rect 76880 36240 76960 36263
rect -2560 35257 -2480 35280
rect -2560 35223 -2537 35257
rect -2503 35223 -2480 35257
rect -2560 34937 -2480 35223
rect -2560 34903 -2537 34937
rect -2503 34903 -2480 34937
rect -2560 34880 -2480 34903
rect -2400 35257 -2320 35280
rect -2400 35223 -2377 35257
rect -2343 35223 -2320 35257
rect -2400 34937 -2320 35223
rect -2400 34903 -2377 34937
rect -2343 34903 -2320 34937
rect -2400 34880 -2320 34903
rect -2240 35257 -2160 35280
rect -2240 35223 -2217 35257
rect -2183 35223 -2160 35257
rect -2240 34937 -2160 35223
rect -2240 34903 -2217 34937
rect -2183 34903 -2160 34937
rect -2240 34880 -2160 34903
rect -2080 35257 -2000 35280
rect -2080 35223 -2057 35257
rect -2023 35223 -2000 35257
rect -2080 34937 -2000 35223
rect -2080 34903 -2057 34937
rect -2023 34903 -2000 34937
rect -2080 34880 -2000 34903
rect -1920 35257 -1840 35280
rect -1920 35223 -1897 35257
rect -1863 35223 -1840 35257
rect -1920 34937 -1840 35223
rect -1920 34903 -1897 34937
rect -1863 34903 -1840 34937
rect -1920 34880 -1840 34903
rect -1760 35257 -1680 35280
rect -1760 35223 -1737 35257
rect -1703 35223 -1680 35257
rect -1760 34937 -1680 35223
rect -1760 34903 -1737 34937
rect -1703 34903 -1680 34937
rect -1760 34880 -1680 34903
rect -1600 35257 -1520 35280
rect -1600 35223 -1577 35257
rect -1543 35223 -1520 35257
rect -1600 34937 -1520 35223
rect -1600 34903 -1577 34937
rect -1543 34903 -1520 34937
rect -1600 34880 -1520 34903
rect -1440 35257 -1360 35280
rect -1440 35223 -1417 35257
rect -1383 35223 -1360 35257
rect -1440 34937 -1360 35223
rect -1440 34903 -1417 34937
rect -1383 34903 -1360 34937
rect -1440 34880 -1360 34903
rect -1280 35257 -1200 35280
rect -1280 35223 -1257 35257
rect -1223 35223 -1200 35257
rect -1280 34937 -1200 35223
rect -1280 34903 -1257 34937
rect -1223 34903 -1200 34937
rect -1280 34880 -1200 34903
rect -1120 35257 -1040 35280
rect -1120 35223 -1097 35257
rect -1063 35223 -1040 35257
rect -1120 34937 -1040 35223
rect -1120 34903 -1097 34937
rect -1063 34903 -1040 34937
rect -1120 34880 -1040 34903
rect -960 35257 -880 35280
rect -960 35223 -937 35257
rect -903 35223 -880 35257
rect -960 34937 -880 35223
rect -960 34903 -937 34937
rect -903 34903 -880 34937
rect -960 34880 -880 34903
rect -800 35257 -720 35280
rect -800 35223 -777 35257
rect -743 35223 -720 35257
rect -800 34937 -720 35223
rect -800 34903 -777 34937
rect -743 34903 -720 34937
rect -800 34880 -720 34903
rect -640 35257 -560 35280
rect -640 35223 -617 35257
rect -583 35223 -560 35257
rect -640 34937 -560 35223
rect -640 34903 -617 34937
rect -583 34903 -560 34937
rect -640 34880 -560 34903
rect -480 35257 -400 35280
rect -480 35223 -457 35257
rect -423 35223 -400 35257
rect -480 34937 -400 35223
rect -480 34903 -457 34937
rect -423 34903 -400 34937
rect -480 34880 -400 34903
rect -320 35257 -240 35280
rect -320 35223 -297 35257
rect -263 35223 -240 35257
rect -320 34937 -240 35223
rect -320 34903 -297 34937
rect -263 34903 -240 34937
rect -320 34880 -240 34903
rect -160 35257 -80 35280
rect -160 35223 -137 35257
rect -103 35223 -80 35257
rect -160 34937 -80 35223
rect -160 34903 -137 34937
rect -103 34903 -80 34937
rect -160 34880 -80 34903
rect 0 35257 80 35280
rect 0 35223 23 35257
rect 57 35223 80 35257
rect 0 34937 80 35223
rect 0 34903 23 34937
rect 57 34903 80 34937
rect 0 34880 80 34903
<< viali >>
rect -937 41863 -903 41897
rect -937 41543 -903 41577
rect -777 41863 -743 41897
rect -777 41543 -743 41577
rect -617 41863 -583 41897
rect -617 41543 -583 41577
rect -457 41863 -423 41897
rect -457 41543 -423 41577
rect -297 41863 -263 41897
rect -297 41543 -263 41577
rect -137 41863 -103 41897
rect -137 41543 -103 41577
rect 23 41863 57 41897
rect 23 41543 57 41577
rect 76743 40583 76777 40617
rect 76743 40263 76777 40297
rect 76903 40583 76937 40617
rect 76903 40263 76937 40297
rect -7017 38263 -6983 38297
rect -7017 37943 -6983 37977
rect -7017 37623 -6983 37657
rect -6857 38263 -6823 38297
rect -6857 37943 -6823 37977
rect -6857 37623 -6823 37657
rect -6697 38263 -6663 38297
rect -6697 37943 -6663 37977
rect -6697 37623 -6663 37657
rect -6537 38263 -6503 38297
rect -6537 37943 -6503 37977
rect -6537 37623 -6503 37657
rect -6377 38263 -6343 38297
rect -6377 37943 -6343 37977
rect -6377 37623 -6343 37657
rect -6217 38263 -6183 38297
rect -6217 37943 -6183 37977
rect -6217 37623 -6183 37657
rect -6057 38263 -6023 38297
rect -6057 37943 -6023 37977
rect -6057 37623 -6023 37657
rect -5897 38263 -5863 38297
rect -5897 37943 -5863 37977
rect -5897 37623 -5863 37657
rect -5737 38263 -5703 38297
rect -5737 37943 -5703 37977
rect -5737 37623 -5703 37657
rect -5577 38263 -5543 38297
rect -5577 37943 -5543 37977
rect -5577 37623 -5543 37657
rect -5417 38263 -5383 38297
rect -5417 37943 -5383 37977
rect -5417 37623 -5383 37657
rect -5257 38263 -5223 38297
rect -5257 37943 -5223 37977
rect -5257 37623 -5223 37657
rect -5097 38263 -5063 38297
rect -5097 37943 -5063 37977
rect -5097 37623 -5063 37657
rect -4937 38263 -4903 38297
rect -4937 37943 -4903 37977
rect -4937 37623 -4903 37657
rect -4777 38263 -4743 38297
rect -4777 37943 -4743 37977
rect -4777 37623 -4743 37657
rect -4617 38263 -4583 38297
rect -4617 37943 -4583 37977
rect -4617 37623 -4583 37657
rect -4457 38263 -4423 38297
rect -4457 37943 -4423 37977
rect -4457 37623 -4423 37657
rect -4297 38263 -4263 38297
rect -4297 37943 -4263 37977
rect -4297 37623 -4263 37657
rect -4137 38263 -4103 38297
rect -4137 37943 -4103 37977
rect -4137 37623 -4103 37657
rect -3977 38263 -3943 38297
rect -3977 37943 -3943 37977
rect -3977 37623 -3943 37657
rect -3817 38263 -3783 38297
rect -3817 37943 -3783 37977
rect -3817 37623 -3783 37657
rect -3657 38263 -3623 38297
rect -3657 37943 -3623 37977
rect -3657 37623 -3623 37657
rect -3497 38263 -3463 38297
rect -3497 37943 -3463 37977
rect -3497 37623 -3463 37657
rect -3337 38263 -3303 38297
rect -3337 37943 -3303 37977
rect -3337 37623 -3303 37657
rect -3177 38263 -3143 38297
rect -3177 37943 -3143 37977
rect -3177 37623 -3143 37657
rect -3017 38263 -2983 38297
rect -3017 37943 -2983 37977
rect -3017 37623 -2983 37657
rect -2857 38263 -2823 38297
rect -2857 37943 -2823 37977
rect -2857 37623 -2823 37657
rect -2697 38263 -2663 38297
rect -2697 37943 -2663 37977
rect -2697 37623 -2663 37657
rect -2537 38263 -2503 38297
rect -2537 37943 -2503 37977
rect -2537 37623 -2503 37657
rect -2377 38263 -2343 38297
rect -2377 37943 -2343 37977
rect -2377 37623 -2343 37657
rect -2217 38263 -2183 38297
rect -2217 37943 -2183 37977
rect -2217 37623 -2183 37657
rect -2057 38263 -2023 38297
rect -2057 37943 -2023 37977
rect -2057 37623 -2023 37657
rect -1897 38263 -1863 38297
rect -1897 37943 -1863 37977
rect -1897 37623 -1863 37657
rect -1737 38263 -1703 38297
rect -1737 37943 -1703 37977
rect -1737 37623 -1703 37657
rect -1577 38263 -1543 38297
rect -1577 37943 -1543 37977
rect -1577 37623 -1543 37657
rect -1417 38263 -1383 38297
rect -1417 37943 -1383 37977
rect -1417 37623 -1383 37657
rect -1257 38263 -1223 38297
rect -1257 37943 -1223 37977
rect -1257 37623 -1223 37657
rect -1097 38263 -1063 38297
rect -1097 37943 -1063 37977
rect -1097 37623 -1063 37657
rect -937 38263 -903 38297
rect -937 37943 -903 37977
rect -937 37623 -903 37657
rect -777 38263 -743 38297
rect -777 37943 -743 37977
rect -777 37623 -743 37657
rect -617 38263 -583 38297
rect -617 37943 -583 37977
rect -617 37623 -583 37657
rect -457 38263 -423 38297
rect -457 37943 -423 37977
rect -457 37623 -423 37657
rect -297 38263 -263 38297
rect -297 37943 -263 37977
rect -297 37623 -263 37657
rect -137 38263 -103 38297
rect -137 37943 -103 37977
rect -137 37623 -103 37657
rect 23 38263 57 38297
rect 23 37943 57 37977
rect 23 37623 57 37657
rect 76743 36583 76777 36617
rect 76743 36263 76777 36297
rect 76903 36583 76937 36617
rect 76903 36263 76937 36297
rect -2537 35223 -2503 35257
rect -2537 34903 -2503 34937
rect -2377 35223 -2343 35257
rect -2377 34903 -2343 34937
rect -2217 35223 -2183 35257
rect -2217 34903 -2183 34937
rect -2057 35223 -2023 35257
rect -2057 34903 -2023 34937
rect -1897 35223 -1863 35257
rect -1897 34903 -1863 34937
rect -1737 35223 -1703 35257
rect -1737 34903 -1703 34937
rect -1577 35223 -1543 35257
rect -1577 34903 -1543 34937
rect -1417 35223 -1383 35257
rect -1417 34903 -1383 34937
rect -1257 35223 -1223 35257
rect -1257 34903 -1223 34937
rect -1097 35223 -1063 35257
rect -1097 34903 -1063 34937
rect -937 35223 -903 35257
rect -937 34903 -903 34937
rect -777 35223 -743 35257
rect -777 34903 -743 34937
rect -617 35223 -583 35257
rect -617 34903 -583 34937
rect -457 35223 -423 35257
rect -457 34903 -423 34937
rect -297 35223 -263 35257
rect -297 34903 -263 34937
rect -137 35223 -103 35257
rect -137 34903 -103 34937
rect 23 35223 57 35257
rect 23 34903 57 34937
<< metal1 >>
rect -960 41906 -880 41920
rect -960 41854 -946 41906
rect -894 41854 -880 41906
rect -960 41840 -880 41854
rect -800 41906 -720 41920
rect -800 41854 -786 41906
rect -734 41854 -720 41906
rect -800 41840 -720 41854
rect -640 41906 -560 41920
rect -640 41854 -626 41906
rect -574 41854 -560 41906
rect -640 41840 -560 41854
rect -480 41906 -400 41920
rect -480 41854 -466 41906
rect -414 41854 -400 41906
rect -480 41840 -400 41854
rect -320 41906 -240 41920
rect -320 41854 -306 41906
rect -254 41854 -240 41906
rect -320 41840 -240 41854
rect -160 41906 -80 41920
rect -160 41854 -146 41906
rect -94 41854 -80 41906
rect -160 41840 -80 41854
rect 0 41906 80 41920
rect 0 41854 14 41906
rect 66 41854 80 41906
rect 0 41840 80 41854
rect -960 41586 -880 41600
rect -960 41534 -946 41586
rect -894 41534 -880 41586
rect -960 41520 -880 41534
rect -800 41586 -720 41600
rect -800 41534 -786 41586
rect -734 41534 -720 41586
rect -800 41520 -720 41534
rect -640 41586 -560 41600
rect -640 41534 -626 41586
rect -574 41534 -560 41586
rect -640 41520 -560 41534
rect -480 41586 -400 41600
rect -480 41534 -466 41586
rect -414 41534 -400 41586
rect -480 41520 -400 41534
rect -320 41586 -240 41600
rect -320 41534 -306 41586
rect -254 41534 -240 41586
rect -320 41520 -240 41534
rect -160 41586 -80 41600
rect -160 41534 -146 41586
rect -94 41534 -80 41586
rect -160 41520 -80 41534
rect 0 41586 80 41600
rect 0 41534 14 41586
rect 66 41534 80 41586
rect 0 41520 80 41534
rect 76720 40626 76800 40640
rect 76720 40574 76734 40626
rect 76786 40574 76800 40626
rect 76720 40560 76800 40574
rect 76880 40626 76960 40640
rect 76880 40574 76894 40626
rect 76946 40574 76960 40626
rect 76880 40560 76960 40574
rect 76720 40306 76800 40320
rect 76720 40254 76734 40306
rect 76786 40254 76800 40306
rect 76720 40240 76800 40254
rect 76880 40306 76960 40320
rect 76880 40254 76894 40306
rect 76946 40254 76960 40306
rect 76880 40240 76960 40254
rect -7040 38306 -6960 38320
rect -7040 38254 -7026 38306
rect -6974 38254 -6960 38306
rect -7040 38240 -6960 38254
rect -6880 38306 -6800 38320
rect -6880 38254 -6866 38306
rect -6814 38254 -6800 38306
rect -6880 38240 -6800 38254
rect -6720 38306 -6640 38320
rect -6720 38254 -6706 38306
rect -6654 38254 -6640 38306
rect -6720 38240 -6640 38254
rect -6560 38306 -6480 38320
rect -6560 38254 -6546 38306
rect -6494 38254 -6480 38306
rect -6560 38240 -6480 38254
rect -6400 38306 -6320 38320
rect -6400 38254 -6386 38306
rect -6334 38254 -6320 38306
rect -6400 38240 -6320 38254
rect -6240 38306 -6160 38320
rect -6240 38254 -6226 38306
rect -6174 38254 -6160 38306
rect -6240 38240 -6160 38254
rect -6080 38306 -6000 38320
rect -6080 38254 -6066 38306
rect -6014 38254 -6000 38306
rect -6080 38240 -6000 38254
rect -5920 38306 -5840 38320
rect -5920 38254 -5906 38306
rect -5854 38254 -5840 38306
rect -5920 38240 -5840 38254
rect -5760 38306 -5680 38320
rect -5760 38254 -5746 38306
rect -5694 38254 -5680 38306
rect -5760 38240 -5680 38254
rect -5600 38306 -5520 38320
rect -5600 38254 -5586 38306
rect -5534 38254 -5520 38306
rect -5600 38240 -5520 38254
rect -5440 38306 -5360 38320
rect -5440 38254 -5426 38306
rect -5374 38254 -5360 38306
rect -5440 38240 -5360 38254
rect -5280 38306 -5200 38320
rect -5280 38254 -5266 38306
rect -5214 38254 -5200 38306
rect -5280 38240 -5200 38254
rect -5120 38306 -5040 38320
rect -5120 38254 -5106 38306
rect -5054 38254 -5040 38306
rect -5120 38240 -5040 38254
rect -4960 38306 -4880 38320
rect -4960 38254 -4946 38306
rect -4894 38254 -4880 38306
rect -4960 38240 -4880 38254
rect -4800 38306 -4720 38320
rect -4800 38254 -4786 38306
rect -4734 38254 -4720 38306
rect -4800 38240 -4720 38254
rect -4640 38306 -4560 38320
rect -4640 38254 -4626 38306
rect -4574 38254 -4560 38306
rect -4640 38240 -4560 38254
rect -4480 38306 -4400 38320
rect -4480 38254 -4466 38306
rect -4414 38254 -4400 38306
rect -4480 38240 -4400 38254
rect -4320 38306 -4240 38320
rect -4320 38254 -4306 38306
rect -4254 38254 -4240 38306
rect -4320 38240 -4240 38254
rect -4160 38306 -4080 38320
rect -4160 38254 -4146 38306
rect -4094 38254 -4080 38306
rect -4160 38240 -4080 38254
rect -4000 38306 -3920 38320
rect -4000 38254 -3986 38306
rect -3934 38254 -3920 38306
rect -4000 38240 -3920 38254
rect -3840 38306 -3760 38320
rect -3840 38254 -3826 38306
rect -3774 38254 -3760 38306
rect -3840 38240 -3760 38254
rect -3680 38306 -3600 38320
rect -3680 38254 -3666 38306
rect -3614 38254 -3600 38306
rect -3680 38240 -3600 38254
rect -3520 38306 -3440 38320
rect -3520 38254 -3506 38306
rect -3454 38254 -3440 38306
rect -3520 38240 -3440 38254
rect -3360 38306 -3280 38320
rect -3360 38254 -3346 38306
rect -3294 38254 -3280 38306
rect -3360 38240 -3280 38254
rect -3200 38306 -3120 38320
rect -3200 38254 -3186 38306
rect -3134 38254 -3120 38306
rect -3200 38240 -3120 38254
rect -3040 38306 -2960 38320
rect -3040 38254 -3026 38306
rect -2974 38254 -2960 38306
rect -3040 38240 -2960 38254
rect -2880 38306 -2800 38320
rect -2880 38254 -2866 38306
rect -2814 38254 -2800 38306
rect -2880 38240 -2800 38254
rect -2720 38306 -2640 38320
rect -2720 38254 -2706 38306
rect -2654 38254 -2640 38306
rect -2720 38240 -2640 38254
rect -2560 38306 -2480 38320
rect -2560 38254 -2546 38306
rect -2494 38254 -2480 38306
rect -2560 38240 -2480 38254
rect -2400 38306 -2320 38320
rect -2400 38254 -2386 38306
rect -2334 38254 -2320 38306
rect -2400 38240 -2320 38254
rect -2240 38306 -2160 38320
rect -2240 38254 -2226 38306
rect -2174 38254 -2160 38306
rect -2240 38240 -2160 38254
rect -2080 38306 -2000 38320
rect -2080 38254 -2066 38306
rect -2014 38254 -2000 38306
rect -2080 38240 -2000 38254
rect -1920 38306 -1840 38320
rect -1920 38254 -1906 38306
rect -1854 38254 -1840 38306
rect -1920 38240 -1840 38254
rect -1760 38306 -1680 38320
rect -1760 38254 -1746 38306
rect -1694 38254 -1680 38306
rect -1760 38240 -1680 38254
rect -1600 38306 -1520 38320
rect -1600 38254 -1586 38306
rect -1534 38254 -1520 38306
rect -1600 38240 -1520 38254
rect -1440 38306 -1360 38320
rect -1440 38254 -1426 38306
rect -1374 38254 -1360 38306
rect -1440 38240 -1360 38254
rect -1280 38306 -1200 38320
rect -1280 38254 -1266 38306
rect -1214 38254 -1200 38306
rect -1280 38240 -1200 38254
rect -1120 38306 -1040 38320
rect -1120 38254 -1106 38306
rect -1054 38254 -1040 38306
rect -1120 38240 -1040 38254
rect -960 38306 -880 38320
rect -960 38254 -946 38306
rect -894 38254 -880 38306
rect -960 38240 -880 38254
rect -800 38306 -720 38320
rect -800 38254 -786 38306
rect -734 38254 -720 38306
rect -800 38240 -720 38254
rect -640 38306 -560 38320
rect -640 38254 -626 38306
rect -574 38254 -560 38306
rect -640 38240 -560 38254
rect -480 38306 -400 38320
rect -480 38254 -466 38306
rect -414 38254 -400 38306
rect -480 38240 -400 38254
rect -320 38306 -240 38320
rect -320 38254 -306 38306
rect -254 38254 -240 38306
rect -320 38240 -240 38254
rect -160 38306 -80 38320
rect -160 38254 -146 38306
rect -94 38254 -80 38306
rect -160 38240 -80 38254
rect 0 38306 80 38320
rect 0 38254 14 38306
rect 66 38254 80 38306
rect 0 38240 80 38254
rect -7040 37986 -6960 38000
rect -7040 37934 -7026 37986
rect -6974 37934 -6960 37986
rect -7040 37920 -6960 37934
rect -6880 37986 -6800 38000
rect -6880 37934 -6866 37986
rect -6814 37934 -6800 37986
rect -6880 37920 -6800 37934
rect -6720 37986 -6640 38000
rect -6720 37934 -6706 37986
rect -6654 37934 -6640 37986
rect -6720 37920 -6640 37934
rect -6560 37986 -6480 38000
rect -6560 37934 -6546 37986
rect -6494 37934 -6480 37986
rect -6560 37920 -6480 37934
rect -6400 37986 -6320 38000
rect -6400 37934 -6386 37986
rect -6334 37934 -6320 37986
rect -6400 37920 -6320 37934
rect -6240 37986 -6160 38000
rect -6240 37934 -6226 37986
rect -6174 37934 -6160 37986
rect -6240 37920 -6160 37934
rect -6080 37986 -6000 38000
rect -6080 37934 -6066 37986
rect -6014 37934 -6000 37986
rect -6080 37920 -6000 37934
rect -5920 37986 -5840 38000
rect -5920 37934 -5906 37986
rect -5854 37934 -5840 37986
rect -5920 37920 -5840 37934
rect -5760 37986 -5680 38000
rect -5760 37934 -5746 37986
rect -5694 37934 -5680 37986
rect -5760 37920 -5680 37934
rect -5600 37986 -5520 38000
rect -5600 37934 -5586 37986
rect -5534 37934 -5520 37986
rect -5600 37920 -5520 37934
rect -5440 37986 -5360 38000
rect -5440 37934 -5426 37986
rect -5374 37934 -5360 37986
rect -5440 37920 -5360 37934
rect -5280 37986 -5200 38000
rect -5280 37934 -5266 37986
rect -5214 37934 -5200 37986
rect -5280 37920 -5200 37934
rect -5120 37986 -5040 38000
rect -5120 37934 -5106 37986
rect -5054 37934 -5040 37986
rect -5120 37920 -5040 37934
rect -4960 37986 -4880 38000
rect -4960 37934 -4946 37986
rect -4894 37934 -4880 37986
rect -4960 37920 -4880 37934
rect -4800 37986 -4720 38000
rect -4800 37934 -4786 37986
rect -4734 37934 -4720 37986
rect -4800 37920 -4720 37934
rect -4640 37986 -4560 38000
rect -4640 37934 -4626 37986
rect -4574 37934 -4560 37986
rect -4640 37920 -4560 37934
rect -4480 37986 -4400 38000
rect -4480 37934 -4466 37986
rect -4414 37934 -4400 37986
rect -4480 37920 -4400 37934
rect -4320 37986 -4240 38000
rect -4320 37934 -4306 37986
rect -4254 37934 -4240 37986
rect -4320 37920 -4240 37934
rect -4160 37986 -4080 38000
rect -4160 37934 -4146 37986
rect -4094 37934 -4080 37986
rect -4160 37920 -4080 37934
rect -4000 37986 -3920 38000
rect -4000 37934 -3986 37986
rect -3934 37934 -3920 37986
rect -4000 37920 -3920 37934
rect -3840 37986 -3760 38000
rect -3840 37934 -3826 37986
rect -3774 37934 -3760 37986
rect -3840 37920 -3760 37934
rect -3680 37986 -3600 38000
rect -3680 37934 -3666 37986
rect -3614 37934 -3600 37986
rect -3680 37920 -3600 37934
rect -3520 37986 -3440 38000
rect -3520 37934 -3506 37986
rect -3454 37934 -3440 37986
rect -3520 37920 -3440 37934
rect -3360 37986 -3280 38000
rect -3360 37934 -3346 37986
rect -3294 37934 -3280 37986
rect -3360 37920 -3280 37934
rect -3200 37986 -3120 38000
rect -3200 37934 -3186 37986
rect -3134 37934 -3120 37986
rect -3200 37920 -3120 37934
rect -3040 37986 -2960 38000
rect -3040 37934 -3026 37986
rect -2974 37934 -2960 37986
rect -3040 37920 -2960 37934
rect -2880 37986 -2800 38000
rect -2880 37934 -2866 37986
rect -2814 37934 -2800 37986
rect -2880 37920 -2800 37934
rect -2720 37986 -2640 38000
rect -2720 37934 -2706 37986
rect -2654 37934 -2640 37986
rect -2720 37920 -2640 37934
rect -2560 37986 -2480 38000
rect -2560 37934 -2546 37986
rect -2494 37934 -2480 37986
rect -2560 37920 -2480 37934
rect -2400 37986 -2320 38000
rect -2400 37934 -2386 37986
rect -2334 37934 -2320 37986
rect -2400 37920 -2320 37934
rect -2240 37986 -2160 38000
rect -2240 37934 -2226 37986
rect -2174 37934 -2160 37986
rect -2240 37920 -2160 37934
rect -2080 37986 -2000 38000
rect -2080 37934 -2066 37986
rect -2014 37934 -2000 37986
rect -2080 37920 -2000 37934
rect -1920 37986 -1840 38000
rect -1920 37934 -1906 37986
rect -1854 37934 -1840 37986
rect -1920 37920 -1840 37934
rect -1760 37986 -1680 38000
rect -1760 37934 -1746 37986
rect -1694 37934 -1680 37986
rect -1760 37920 -1680 37934
rect -1600 37986 -1520 38000
rect -1600 37934 -1586 37986
rect -1534 37934 -1520 37986
rect -1600 37920 -1520 37934
rect -1440 37986 -1360 38000
rect -1440 37934 -1426 37986
rect -1374 37934 -1360 37986
rect -1440 37920 -1360 37934
rect -1280 37986 -1200 38000
rect -1280 37934 -1266 37986
rect -1214 37934 -1200 37986
rect -1280 37920 -1200 37934
rect -1120 37986 -1040 38000
rect -1120 37934 -1106 37986
rect -1054 37934 -1040 37986
rect -1120 37920 -1040 37934
rect -960 37986 -880 38000
rect -960 37934 -946 37986
rect -894 37934 -880 37986
rect -960 37920 -880 37934
rect -800 37986 -720 38000
rect -800 37934 -786 37986
rect -734 37934 -720 37986
rect -800 37920 -720 37934
rect -640 37986 -560 38000
rect -640 37934 -626 37986
rect -574 37934 -560 37986
rect -640 37920 -560 37934
rect -480 37986 -400 38000
rect -480 37934 -466 37986
rect -414 37934 -400 37986
rect -480 37920 -400 37934
rect -320 37986 -240 38000
rect -320 37934 -306 37986
rect -254 37934 -240 37986
rect -320 37920 -240 37934
rect -160 37986 -80 38000
rect -160 37934 -146 37986
rect -94 37934 -80 37986
rect -160 37920 -80 37934
rect 0 37986 80 38000
rect 0 37934 14 37986
rect 66 37934 80 37986
rect 0 37920 80 37934
rect -7040 37666 -6960 37680
rect -7040 37614 -7026 37666
rect -6974 37614 -6960 37666
rect -7040 37600 -6960 37614
rect -6880 37666 -6800 37680
rect -6880 37614 -6866 37666
rect -6814 37614 -6800 37666
rect -6880 37600 -6800 37614
rect -6720 37666 -6640 37680
rect -6720 37614 -6706 37666
rect -6654 37614 -6640 37666
rect -6720 37600 -6640 37614
rect -6560 37666 -6480 37680
rect -6560 37614 -6546 37666
rect -6494 37614 -6480 37666
rect -6560 37600 -6480 37614
rect -6400 37666 -6320 37680
rect -6400 37614 -6386 37666
rect -6334 37614 -6320 37666
rect -6400 37600 -6320 37614
rect -6240 37666 -6160 37680
rect -6240 37614 -6226 37666
rect -6174 37614 -6160 37666
rect -6240 37600 -6160 37614
rect -6080 37666 -6000 37680
rect -6080 37614 -6066 37666
rect -6014 37614 -6000 37666
rect -6080 37600 -6000 37614
rect -5920 37666 -5840 37680
rect -5920 37614 -5906 37666
rect -5854 37614 -5840 37666
rect -5920 37600 -5840 37614
rect -5760 37666 -5680 37680
rect -5760 37614 -5746 37666
rect -5694 37614 -5680 37666
rect -5760 37600 -5680 37614
rect -5600 37666 -5520 37680
rect -5600 37614 -5586 37666
rect -5534 37614 -5520 37666
rect -5600 37600 -5520 37614
rect -5440 37666 -5360 37680
rect -5440 37614 -5426 37666
rect -5374 37614 -5360 37666
rect -5440 37600 -5360 37614
rect -5280 37666 -5200 37680
rect -5280 37614 -5266 37666
rect -5214 37614 -5200 37666
rect -5280 37600 -5200 37614
rect -5120 37666 -5040 37680
rect -5120 37614 -5106 37666
rect -5054 37614 -5040 37666
rect -5120 37600 -5040 37614
rect -4960 37666 -4880 37680
rect -4960 37614 -4946 37666
rect -4894 37614 -4880 37666
rect -4960 37600 -4880 37614
rect -4800 37666 -4720 37680
rect -4800 37614 -4786 37666
rect -4734 37614 -4720 37666
rect -4800 37600 -4720 37614
rect -4640 37666 -4560 37680
rect -4640 37614 -4626 37666
rect -4574 37614 -4560 37666
rect -4640 37600 -4560 37614
rect -4480 37666 -4400 37680
rect -4480 37614 -4466 37666
rect -4414 37614 -4400 37666
rect -4480 37600 -4400 37614
rect -4320 37666 -4240 37680
rect -4320 37614 -4306 37666
rect -4254 37614 -4240 37666
rect -4320 37600 -4240 37614
rect -4160 37666 -4080 37680
rect -4160 37614 -4146 37666
rect -4094 37614 -4080 37666
rect -4160 37600 -4080 37614
rect -4000 37666 -3920 37680
rect -4000 37614 -3986 37666
rect -3934 37614 -3920 37666
rect -4000 37600 -3920 37614
rect -3840 37666 -3760 37680
rect -3840 37614 -3826 37666
rect -3774 37614 -3760 37666
rect -3840 37600 -3760 37614
rect -3680 37666 -3600 37680
rect -3680 37614 -3666 37666
rect -3614 37614 -3600 37666
rect -3680 37600 -3600 37614
rect -3520 37666 -3440 37680
rect -3520 37614 -3506 37666
rect -3454 37614 -3440 37666
rect -3520 37600 -3440 37614
rect -3360 37666 -3280 37680
rect -3360 37614 -3346 37666
rect -3294 37614 -3280 37666
rect -3360 37600 -3280 37614
rect -3200 37666 -3120 37680
rect -3200 37614 -3186 37666
rect -3134 37614 -3120 37666
rect -3200 37600 -3120 37614
rect -3040 37666 -2960 37680
rect -3040 37614 -3026 37666
rect -2974 37614 -2960 37666
rect -3040 37600 -2960 37614
rect -2880 37666 -2800 37680
rect -2880 37614 -2866 37666
rect -2814 37614 -2800 37666
rect -2880 37600 -2800 37614
rect -2720 37666 -2640 37680
rect -2720 37614 -2706 37666
rect -2654 37614 -2640 37666
rect -2720 37600 -2640 37614
rect -2560 37666 -2480 37680
rect -2560 37614 -2546 37666
rect -2494 37614 -2480 37666
rect -2560 37600 -2480 37614
rect -2400 37666 -2320 37680
rect -2400 37614 -2386 37666
rect -2334 37614 -2320 37666
rect -2400 37600 -2320 37614
rect -2240 37666 -2160 37680
rect -2240 37614 -2226 37666
rect -2174 37614 -2160 37666
rect -2240 37600 -2160 37614
rect -2080 37666 -2000 37680
rect -2080 37614 -2066 37666
rect -2014 37614 -2000 37666
rect -2080 37600 -2000 37614
rect -1920 37666 -1840 37680
rect -1920 37614 -1906 37666
rect -1854 37614 -1840 37666
rect -1920 37600 -1840 37614
rect -1760 37666 -1680 37680
rect -1760 37614 -1746 37666
rect -1694 37614 -1680 37666
rect -1760 37600 -1680 37614
rect -1600 37666 -1520 37680
rect -1600 37614 -1586 37666
rect -1534 37614 -1520 37666
rect -1600 37600 -1520 37614
rect -1440 37666 -1360 37680
rect -1440 37614 -1426 37666
rect -1374 37614 -1360 37666
rect -1440 37600 -1360 37614
rect -1280 37666 -1200 37680
rect -1280 37614 -1266 37666
rect -1214 37614 -1200 37666
rect -1280 37600 -1200 37614
rect -1120 37666 -1040 37680
rect -1120 37614 -1106 37666
rect -1054 37614 -1040 37666
rect -1120 37600 -1040 37614
rect -960 37666 -880 37680
rect -960 37614 -946 37666
rect -894 37614 -880 37666
rect -960 37600 -880 37614
rect -800 37666 -720 37680
rect -800 37614 -786 37666
rect -734 37614 -720 37666
rect -800 37600 -720 37614
rect -640 37666 -560 37680
rect -640 37614 -626 37666
rect -574 37614 -560 37666
rect -640 37600 -560 37614
rect -480 37666 -400 37680
rect -480 37614 -466 37666
rect -414 37614 -400 37666
rect -480 37600 -400 37614
rect -320 37666 -240 37680
rect -320 37614 -306 37666
rect -254 37614 -240 37666
rect -320 37600 -240 37614
rect -160 37666 -80 37680
rect -160 37614 -146 37666
rect -94 37614 -80 37666
rect -160 37600 -80 37614
rect 0 37666 80 37680
rect 0 37614 14 37666
rect 66 37614 80 37666
rect 0 37600 80 37614
rect 76720 36626 76800 36640
rect 76720 36574 76734 36626
rect 76786 36574 76800 36626
rect 76720 36560 76800 36574
rect 76880 36626 76960 36640
rect 76880 36574 76894 36626
rect 76946 36574 76960 36626
rect 76880 36560 76960 36574
rect 76720 36306 76800 36320
rect 76720 36254 76734 36306
rect 76786 36254 76800 36306
rect 76720 36240 76800 36254
rect 76880 36306 76960 36320
rect 76880 36254 76894 36306
rect 76946 36254 76960 36306
rect 76880 36240 76960 36254
rect -2560 35266 -2480 35280
rect -2560 35214 -2546 35266
rect -2494 35214 -2480 35266
rect -2560 35200 -2480 35214
rect -2400 35266 -2320 35280
rect -2400 35214 -2386 35266
rect -2334 35214 -2320 35266
rect -2400 35200 -2320 35214
rect -2240 35266 -2160 35280
rect -2240 35214 -2226 35266
rect -2174 35214 -2160 35266
rect -2240 35200 -2160 35214
rect -2080 35266 -2000 35280
rect -2080 35214 -2066 35266
rect -2014 35214 -2000 35266
rect -2080 35200 -2000 35214
rect -1920 35266 -1840 35280
rect -1920 35214 -1906 35266
rect -1854 35214 -1840 35266
rect -1920 35200 -1840 35214
rect -1760 35266 -1680 35280
rect -1760 35214 -1746 35266
rect -1694 35214 -1680 35266
rect -1760 35200 -1680 35214
rect -1600 35266 -1520 35280
rect -1600 35214 -1586 35266
rect -1534 35214 -1520 35266
rect -1600 35200 -1520 35214
rect -1440 35266 -1360 35280
rect -1440 35214 -1426 35266
rect -1374 35214 -1360 35266
rect -1440 35200 -1360 35214
rect -1280 35266 -1200 35280
rect -1280 35214 -1266 35266
rect -1214 35214 -1200 35266
rect -1280 35200 -1200 35214
rect -1120 35266 -1040 35280
rect -1120 35214 -1106 35266
rect -1054 35214 -1040 35266
rect -1120 35200 -1040 35214
rect -960 35266 -880 35280
rect -960 35214 -946 35266
rect -894 35214 -880 35266
rect -960 35200 -880 35214
rect -800 35266 -720 35280
rect -800 35214 -786 35266
rect -734 35214 -720 35266
rect -800 35200 -720 35214
rect -640 35266 -560 35280
rect -640 35214 -626 35266
rect -574 35214 -560 35266
rect -640 35200 -560 35214
rect -480 35266 -400 35280
rect -480 35214 -466 35266
rect -414 35214 -400 35266
rect -480 35200 -400 35214
rect -320 35266 -240 35280
rect -320 35214 -306 35266
rect -254 35214 -240 35266
rect -320 35200 -240 35214
rect -160 35266 -80 35280
rect -160 35214 -146 35266
rect -94 35214 -80 35266
rect -160 35200 -80 35214
rect 0 35266 80 35280
rect 0 35214 14 35266
rect 66 35214 80 35266
rect 0 35200 80 35214
rect -2560 34946 -2480 34960
rect -2560 34894 -2546 34946
rect -2494 34894 -2480 34946
rect -2560 34880 -2480 34894
rect -2400 34946 -2320 34960
rect -2400 34894 -2386 34946
rect -2334 34894 -2320 34946
rect -2400 34880 -2320 34894
rect -2240 34946 -2160 34960
rect -2240 34894 -2226 34946
rect -2174 34894 -2160 34946
rect -2240 34880 -2160 34894
rect -2080 34946 -2000 34960
rect -2080 34894 -2066 34946
rect -2014 34894 -2000 34946
rect -2080 34880 -2000 34894
rect -1920 34946 -1840 34960
rect -1920 34894 -1906 34946
rect -1854 34894 -1840 34946
rect -1920 34880 -1840 34894
rect -1760 34946 -1680 34960
rect -1760 34894 -1746 34946
rect -1694 34894 -1680 34946
rect -1760 34880 -1680 34894
rect -1600 34946 -1520 34960
rect -1600 34894 -1586 34946
rect -1534 34894 -1520 34946
rect -1600 34880 -1520 34894
rect -1440 34946 -1360 34960
rect -1440 34894 -1426 34946
rect -1374 34894 -1360 34946
rect -1440 34880 -1360 34894
rect -1280 34946 -1200 34960
rect -1280 34894 -1266 34946
rect -1214 34894 -1200 34946
rect -1280 34880 -1200 34894
rect -1120 34946 -1040 34960
rect -1120 34894 -1106 34946
rect -1054 34894 -1040 34946
rect -1120 34880 -1040 34894
rect -960 34946 -880 34960
rect -960 34894 -946 34946
rect -894 34894 -880 34946
rect -960 34880 -880 34894
rect -800 34946 -720 34960
rect -800 34894 -786 34946
rect -734 34894 -720 34946
rect -800 34880 -720 34894
rect -640 34946 -560 34960
rect -640 34894 -626 34946
rect -574 34894 -560 34946
rect -640 34880 -560 34894
rect -480 34946 -400 34960
rect -480 34894 -466 34946
rect -414 34894 -400 34946
rect -480 34880 -400 34894
rect -320 34946 -240 34960
rect -320 34894 -306 34946
rect -254 34894 -240 34946
rect -320 34880 -240 34894
rect -160 34946 -80 34960
rect -160 34894 -146 34946
rect -94 34894 -80 34946
rect -160 34880 -80 34894
rect 0 34946 80 34960
rect 0 34894 14 34946
rect 66 34894 80 34946
rect 0 34880 80 34894
<< via1 >>
rect -946 41897 -894 41906
rect -946 41863 -937 41897
rect -937 41863 -903 41897
rect -903 41863 -894 41897
rect -946 41854 -894 41863
rect -786 41897 -734 41906
rect -786 41863 -777 41897
rect -777 41863 -743 41897
rect -743 41863 -734 41897
rect -786 41854 -734 41863
rect -626 41897 -574 41906
rect -626 41863 -617 41897
rect -617 41863 -583 41897
rect -583 41863 -574 41897
rect -626 41854 -574 41863
rect -466 41897 -414 41906
rect -466 41863 -457 41897
rect -457 41863 -423 41897
rect -423 41863 -414 41897
rect -466 41854 -414 41863
rect -306 41897 -254 41906
rect -306 41863 -297 41897
rect -297 41863 -263 41897
rect -263 41863 -254 41897
rect -306 41854 -254 41863
rect -146 41897 -94 41906
rect -146 41863 -137 41897
rect -137 41863 -103 41897
rect -103 41863 -94 41897
rect -146 41854 -94 41863
rect 14 41897 66 41906
rect 14 41863 23 41897
rect 23 41863 57 41897
rect 57 41863 66 41897
rect 14 41854 66 41863
rect -946 41577 -894 41586
rect -946 41543 -937 41577
rect -937 41543 -903 41577
rect -903 41543 -894 41577
rect -946 41534 -894 41543
rect -786 41577 -734 41586
rect -786 41543 -777 41577
rect -777 41543 -743 41577
rect -743 41543 -734 41577
rect -786 41534 -734 41543
rect -626 41577 -574 41586
rect -626 41543 -617 41577
rect -617 41543 -583 41577
rect -583 41543 -574 41577
rect -626 41534 -574 41543
rect -466 41577 -414 41586
rect -466 41543 -457 41577
rect -457 41543 -423 41577
rect -423 41543 -414 41577
rect -466 41534 -414 41543
rect -306 41577 -254 41586
rect -306 41543 -297 41577
rect -297 41543 -263 41577
rect -263 41543 -254 41577
rect -306 41534 -254 41543
rect -146 41577 -94 41586
rect -146 41543 -137 41577
rect -137 41543 -103 41577
rect -103 41543 -94 41577
rect -146 41534 -94 41543
rect 14 41577 66 41586
rect 14 41543 23 41577
rect 23 41543 57 41577
rect 57 41543 66 41577
rect 14 41534 66 41543
rect 76734 40617 76786 40626
rect 76734 40583 76743 40617
rect 76743 40583 76777 40617
rect 76777 40583 76786 40617
rect 76734 40574 76786 40583
rect 76894 40617 76946 40626
rect 76894 40583 76903 40617
rect 76903 40583 76937 40617
rect 76937 40583 76946 40617
rect 76894 40574 76946 40583
rect 76734 40297 76786 40306
rect 76734 40263 76743 40297
rect 76743 40263 76777 40297
rect 76777 40263 76786 40297
rect 76734 40254 76786 40263
rect 76894 40297 76946 40306
rect 76894 40263 76903 40297
rect 76903 40263 76937 40297
rect 76937 40263 76946 40297
rect 76894 40254 76946 40263
rect -7026 38297 -6974 38306
rect -7026 38263 -7017 38297
rect -7017 38263 -6983 38297
rect -6983 38263 -6974 38297
rect -7026 38254 -6974 38263
rect -6866 38297 -6814 38306
rect -6866 38263 -6857 38297
rect -6857 38263 -6823 38297
rect -6823 38263 -6814 38297
rect -6866 38254 -6814 38263
rect -6706 38297 -6654 38306
rect -6706 38263 -6697 38297
rect -6697 38263 -6663 38297
rect -6663 38263 -6654 38297
rect -6706 38254 -6654 38263
rect -6546 38297 -6494 38306
rect -6546 38263 -6537 38297
rect -6537 38263 -6503 38297
rect -6503 38263 -6494 38297
rect -6546 38254 -6494 38263
rect -6386 38297 -6334 38306
rect -6386 38263 -6377 38297
rect -6377 38263 -6343 38297
rect -6343 38263 -6334 38297
rect -6386 38254 -6334 38263
rect -6226 38297 -6174 38306
rect -6226 38263 -6217 38297
rect -6217 38263 -6183 38297
rect -6183 38263 -6174 38297
rect -6226 38254 -6174 38263
rect -6066 38297 -6014 38306
rect -6066 38263 -6057 38297
rect -6057 38263 -6023 38297
rect -6023 38263 -6014 38297
rect -6066 38254 -6014 38263
rect -5906 38297 -5854 38306
rect -5906 38263 -5897 38297
rect -5897 38263 -5863 38297
rect -5863 38263 -5854 38297
rect -5906 38254 -5854 38263
rect -5746 38297 -5694 38306
rect -5746 38263 -5737 38297
rect -5737 38263 -5703 38297
rect -5703 38263 -5694 38297
rect -5746 38254 -5694 38263
rect -5586 38297 -5534 38306
rect -5586 38263 -5577 38297
rect -5577 38263 -5543 38297
rect -5543 38263 -5534 38297
rect -5586 38254 -5534 38263
rect -5426 38297 -5374 38306
rect -5426 38263 -5417 38297
rect -5417 38263 -5383 38297
rect -5383 38263 -5374 38297
rect -5426 38254 -5374 38263
rect -5266 38297 -5214 38306
rect -5266 38263 -5257 38297
rect -5257 38263 -5223 38297
rect -5223 38263 -5214 38297
rect -5266 38254 -5214 38263
rect -5106 38297 -5054 38306
rect -5106 38263 -5097 38297
rect -5097 38263 -5063 38297
rect -5063 38263 -5054 38297
rect -5106 38254 -5054 38263
rect -4946 38297 -4894 38306
rect -4946 38263 -4937 38297
rect -4937 38263 -4903 38297
rect -4903 38263 -4894 38297
rect -4946 38254 -4894 38263
rect -4786 38297 -4734 38306
rect -4786 38263 -4777 38297
rect -4777 38263 -4743 38297
rect -4743 38263 -4734 38297
rect -4786 38254 -4734 38263
rect -4626 38297 -4574 38306
rect -4626 38263 -4617 38297
rect -4617 38263 -4583 38297
rect -4583 38263 -4574 38297
rect -4626 38254 -4574 38263
rect -4466 38297 -4414 38306
rect -4466 38263 -4457 38297
rect -4457 38263 -4423 38297
rect -4423 38263 -4414 38297
rect -4466 38254 -4414 38263
rect -4306 38297 -4254 38306
rect -4306 38263 -4297 38297
rect -4297 38263 -4263 38297
rect -4263 38263 -4254 38297
rect -4306 38254 -4254 38263
rect -4146 38297 -4094 38306
rect -4146 38263 -4137 38297
rect -4137 38263 -4103 38297
rect -4103 38263 -4094 38297
rect -4146 38254 -4094 38263
rect -3986 38297 -3934 38306
rect -3986 38263 -3977 38297
rect -3977 38263 -3943 38297
rect -3943 38263 -3934 38297
rect -3986 38254 -3934 38263
rect -3826 38297 -3774 38306
rect -3826 38263 -3817 38297
rect -3817 38263 -3783 38297
rect -3783 38263 -3774 38297
rect -3826 38254 -3774 38263
rect -3666 38297 -3614 38306
rect -3666 38263 -3657 38297
rect -3657 38263 -3623 38297
rect -3623 38263 -3614 38297
rect -3666 38254 -3614 38263
rect -3506 38297 -3454 38306
rect -3506 38263 -3497 38297
rect -3497 38263 -3463 38297
rect -3463 38263 -3454 38297
rect -3506 38254 -3454 38263
rect -3346 38297 -3294 38306
rect -3346 38263 -3337 38297
rect -3337 38263 -3303 38297
rect -3303 38263 -3294 38297
rect -3346 38254 -3294 38263
rect -3186 38297 -3134 38306
rect -3186 38263 -3177 38297
rect -3177 38263 -3143 38297
rect -3143 38263 -3134 38297
rect -3186 38254 -3134 38263
rect -3026 38297 -2974 38306
rect -3026 38263 -3017 38297
rect -3017 38263 -2983 38297
rect -2983 38263 -2974 38297
rect -3026 38254 -2974 38263
rect -2866 38297 -2814 38306
rect -2866 38263 -2857 38297
rect -2857 38263 -2823 38297
rect -2823 38263 -2814 38297
rect -2866 38254 -2814 38263
rect -2706 38297 -2654 38306
rect -2706 38263 -2697 38297
rect -2697 38263 -2663 38297
rect -2663 38263 -2654 38297
rect -2706 38254 -2654 38263
rect -2546 38297 -2494 38306
rect -2546 38263 -2537 38297
rect -2537 38263 -2503 38297
rect -2503 38263 -2494 38297
rect -2546 38254 -2494 38263
rect -2386 38297 -2334 38306
rect -2386 38263 -2377 38297
rect -2377 38263 -2343 38297
rect -2343 38263 -2334 38297
rect -2386 38254 -2334 38263
rect -2226 38297 -2174 38306
rect -2226 38263 -2217 38297
rect -2217 38263 -2183 38297
rect -2183 38263 -2174 38297
rect -2226 38254 -2174 38263
rect -2066 38297 -2014 38306
rect -2066 38263 -2057 38297
rect -2057 38263 -2023 38297
rect -2023 38263 -2014 38297
rect -2066 38254 -2014 38263
rect -1906 38297 -1854 38306
rect -1906 38263 -1897 38297
rect -1897 38263 -1863 38297
rect -1863 38263 -1854 38297
rect -1906 38254 -1854 38263
rect -1746 38297 -1694 38306
rect -1746 38263 -1737 38297
rect -1737 38263 -1703 38297
rect -1703 38263 -1694 38297
rect -1746 38254 -1694 38263
rect -1586 38297 -1534 38306
rect -1586 38263 -1577 38297
rect -1577 38263 -1543 38297
rect -1543 38263 -1534 38297
rect -1586 38254 -1534 38263
rect -1426 38297 -1374 38306
rect -1426 38263 -1417 38297
rect -1417 38263 -1383 38297
rect -1383 38263 -1374 38297
rect -1426 38254 -1374 38263
rect -1266 38297 -1214 38306
rect -1266 38263 -1257 38297
rect -1257 38263 -1223 38297
rect -1223 38263 -1214 38297
rect -1266 38254 -1214 38263
rect -1106 38297 -1054 38306
rect -1106 38263 -1097 38297
rect -1097 38263 -1063 38297
rect -1063 38263 -1054 38297
rect -1106 38254 -1054 38263
rect -946 38297 -894 38306
rect -946 38263 -937 38297
rect -937 38263 -903 38297
rect -903 38263 -894 38297
rect -946 38254 -894 38263
rect -786 38297 -734 38306
rect -786 38263 -777 38297
rect -777 38263 -743 38297
rect -743 38263 -734 38297
rect -786 38254 -734 38263
rect -626 38297 -574 38306
rect -626 38263 -617 38297
rect -617 38263 -583 38297
rect -583 38263 -574 38297
rect -626 38254 -574 38263
rect -466 38297 -414 38306
rect -466 38263 -457 38297
rect -457 38263 -423 38297
rect -423 38263 -414 38297
rect -466 38254 -414 38263
rect -306 38297 -254 38306
rect -306 38263 -297 38297
rect -297 38263 -263 38297
rect -263 38263 -254 38297
rect -306 38254 -254 38263
rect -146 38297 -94 38306
rect -146 38263 -137 38297
rect -137 38263 -103 38297
rect -103 38263 -94 38297
rect -146 38254 -94 38263
rect 14 38297 66 38306
rect 14 38263 23 38297
rect 23 38263 57 38297
rect 57 38263 66 38297
rect 14 38254 66 38263
rect -7026 37977 -6974 37986
rect -7026 37943 -7017 37977
rect -7017 37943 -6983 37977
rect -6983 37943 -6974 37977
rect -7026 37934 -6974 37943
rect -6866 37977 -6814 37986
rect -6866 37943 -6857 37977
rect -6857 37943 -6823 37977
rect -6823 37943 -6814 37977
rect -6866 37934 -6814 37943
rect -6706 37977 -6654 37986
rect -6706 37943 -6697 37977
rect -6697 37943 -6663 37977
rect -6663 37943 -6654 37977
rect -6706 37934 -6654 37943
rect -6546 37977 -6494 37986
rect -6546 37943 -6537 37977
rect -6537 37943 -6503 37977
rect -6503 37943 -6494 37977
rect -6546 37934 -6494 37943
rect -6386 37977 -6334 37986
rect -6386 37943 -6377 37977
rect -6377 37943 -6343 37977
rect -6343 37943 -6334 37977
rect -6386 37934 -6334 37943
rect -6226 37977 -6174 37986
rect -6226 37943 -6217 37977
rect -6217 37943 -6183 37977
rect -6183 37943 -6174 37977
rect -6226 37934 -6174 37943
rect -6066 37977 -6014 37986
rect -6066 37943 -6057 37977
rect -6057 37943 -6023 37977
rect -6023 37943 -6014 37977
rect -6066 37934 -6014 37943
rect -5906 37977 -5854 37986
rect -5906 37943 -5897 37977
rect -5897 37943 -5863 37977
rect -5863 37943 -5854 37977
rect -5906 37934 -5854 37943
rect -5746 37977 -5694 37986
rect -5746 37943 -5737 37977
rect -5737 37943 -5703 37977
rect -5703 37943 -5694 37977
rect -5746 37934 -5694 37943
rect -5586 37977 -5534 37986
rect -5586 37943 -5577 37977
rect -5577 37943 -5543 37977
rect -5543 37943 -5534 37977
rect -5586 37934 -5534 37943
rect -5426 37977 -5374 37986
rect -5426 37943 -5417 37977
rect -5417 37943 -5383 37977
rect -5383 37943 -5374 37977
rect -5426 37934 -5374 37943
rect -5266 37977 -5214 37986
rect -5266 37943 -5257 37977
rect -5257 37943 -5223 37977
rect -5223 37943 -5214 37977
rect -5266 37934 -5214 37943
rect -5106 37977 -5054 37986
rect -5106 37943 -5097 37977
rect -5097 37943 -5063 37977
rect -5063 37943 -5054 37977
rect -5106 37934 -5054 37943
rect -4946 37977 -4894 37986
rect -4946 37943 -4937 37977
rect -4937 37943 -4903 37977
rect -4903 37943 -4894 37977
rect -4946 37934 -4894 37943
rect -4786 37977 -4734 37986
rect -4786 37943 -4777 37977
rect -4777 37943 -4743 37977
rect -4743 37943 -4734 37977
rect -4786 37934 -4734 37943
rect -4626 37977 -4574 37986
rect -4626 37943 -4617 37977
rect -4617 37943 -4583 37977
rect -4583 37943 -4574 37977
rect -4626 37934 -4574 37943
rect -4466 37977 -4414 37986
rect -4466 37943 -4457 37977
rect -4457 37943 -4423 37977
rect -4423 37943 -4414 37977
rect -4466 37934 -4414 37943
rect -4306 37977 -4254 37986
rect -4306 37943 -4297 37977
rect -4297 37943 -4263 37977
rect -4263 37943 -4254 37977
rect -4306 37934 -4254 37943
rect -4146 37977 -4094 37986
rect -4146 37943 -4137 37977
rect -4137 37943 -4103 37977
rect -4103 37943 -4094 37977
rect -4146 37934 -4094 37943
rect -3986 37977 -3934 37986
rect -3986 37943 -3977 37977
rect -3977 37943 -3943 37977
rect -3943 37943 -3934 37977
rect -3986 37934 -3934 37943
rect -3826 37977 -3774 37986
rect -3826 37943 -3817 37977
rect -3817 37943 -3783 37977
rect -3783 37943 -3774 37977
rect -3826 37934 -3774 37943
rect -3666 37977 -3614 37986
rect -3666 37943 -3657 37977
rect -3657 37943 -3623 37977
rect -3623 37943 -3614 37977
rect -3666 37934 -3614 37943
rect -3506 37977 -3454 37986
rect -3506 37943 -3497 37977
rect -3497 37943 -3463 37977
rect -3463 37943 -3454 37977
rect -3506 37934 -3454 37943
rect -3346 37977 -3294 37986
rect -3346 37943 -3337 37977
rect -3337 37943 -3303 37977
rect -3303 37943 -3294 37977
rect -3346 37934 -3294 37943
rect -3186 37977 -3134 37986
rect -3186 37943 -3177 37977
rect -3177 37943 -3143 37977
rect -3143 37943 -3134 37977
rect -3186 37934 -3134 37943
rect -3026 37977 -2974 37986
rect -3026 37943 -3017 37977
rect -3017 37943 -2983 37977
rect -2983 37943 -2974 37977
rect -3026 37934 -2974 37943
rect -2866 37977 -2814 37986
rect -2866 37943 -2857 37977
rect -2857 37943 -2823 37977
rect -2823 37943 -2814 37977
rect -2866 37934 -2814 37943
rect -2706 37977 -2654 37986
rect -2706 37943 -2697 37977
rect -2697 37943 -2663 37977
rect -2663 37943 -2654 37977
rect -2706 37934 -2654 37943
rect -2546 37977 -2494 37986
rect -2546 37943 -2537 37977
rect -2537 37943 -2503 37977
rect -2503 37943 -2494 37977
rect -2546 37934 -2494 37943
rect -2386 37977 -2334 37986
rect -2386 37943 -2377 37977
rect -2377 37943 -2343 37977
rect -2343 37943 -2334 37977
rect -2386 37934 -2334 37943
rect -2226 37977 -2174 37986
rect -2226 37943 -2217 37977
rect -2217 37943 -2183 37977
rect -2183 37943 -2174 37977
rect -2226 37934 -2174 37943
rect -2066 37977 -2014 37986
rect -2066 37943 -2057 37977
rect -2057 37943 -2023 37977
rect -2023 37943 -2014 37977
rect -2066 37934 -2014 37943
rect -1906 37977 -1854 37986
rect -1906 37943 -1897 37977
rect -1897 37943 -1863 37977
rect -1863 37943 -1854 37977
rect -1906 37934 -1854 37943
rect -1746 37977 -1694 37986
rect -1746 37943 -1737 37977
rect -1737 37943 -1703 37977
rect -1703 37943 -1694 37977
rect -1746 37934 -1694 37943
rect -1586 37977 -1534 37986
rect -1586 37943 -1577 37977
rect -1577 37943 -1543 37977
rect -1543 37943 -1534 37977
rect -1586 37934 -1534 37943
rect -1426 37977 -1374 37986
rect -1426 37943 -1417 37977
rect -1417 37943 -1383 37977
rect -1383 37943 -1374 37977
rect -1426 37934 -1374 37943
rect -1266 37977 -1214 37986
rect -1266 37943 -1257 37977
rect -1257 37943 -1223 37977
rect -1223 37943 -1214 37977
rect -1266 37934 -1214 37943
rect -1106 37977 -1054 37986
rect -1106 37943 -1097 37977
rect -1097 37943 -1063 37977
rect -1063 37943 -1054 37977
rect -1106 37934 -1054 37943
rect -946 37977 -894 37986
rect -946 37943 -937 37977
rect -937 37943 -903 37977
rect -903 37943 -894 37977
rect -946 37934 -894 37943
rect -786 37977 -734 37986
rect -786 37943 -777 37977
rect -777 37943 -743 37977
rect -743 37943 -734 37977
rect -786 37934 -734 37943
rect -626 37977 -574 37986
rect -626 37943 -617 37977
rect -617 37943 -583 37977
rect -583 37943 -574 37977
rect -626 37934 -574 37943
rect -466 37977 -414 37986
rect -466 37943 -457 37977
rect -457 37943 -423 37977
rect -423 37943 -414 37977
rect -466 37934 -414 37943
rect -306 37977 -254 37986
rect -306 37943 -297 37977
rect -297 37943 -263 37977
rect -263 37943 -254 37977
rect -306 37934 -254 37943
rect -146 37977 -94 37986
rect -146 37943 -137 37977
rect -137 37943 -103 37977
rect -103 37943 -94 37977
rect -146 37934 -94 37943
rect 14 37977 66 37986
rect 14 37943 23 37977
rect 23 37943 57 37977
rect 57 37943 66 37977
rect 14 37934 66 37943
rect -7026 37657 -6974 37666
rect -7026 37623 -7017 37657
rect -7017 37623 -6983 37657
rect -6983 37623 -6974 37657
rect -7026 37614 -6974 37623
rect -6866 37657 -6814 37666
rect -6866 37623 -6857 37657
rect -6857 37623 -6823 37657
rect -6823 37623 -6814 37657
rect -6866 37614 -6814 37623
rect -6706 37657 -6654 37666
rect -6706 37623 -6697 37657
rect -6697 37623 -6663 37657
rect -6663 37623 -6654 37657
rect -6706 37614 -6654 37623
rect -6546 37657 -6494 37666
rect -6546 37623 -6537 37657
rect -6537 37623 -6503 37657
rect -6503 37623 -6494 37657
rect -6546 37614 -6494 37623
rect -6386 37657 -6334 37666
rect -6386 37623 -6377 37657
rect -6377 37623 -6343 37657
rect -6343 37623 -6334 37657
rect -6386 37614 -6334 37623
rect -6226 37657 -6174 37666
rect -6226 37623 -6217 37657
rect -6217 37623 -6183 37657
rect -6183 37623 -6174 37657
rect -6226 37614 -6174 37623
rect -6066 37657 -6014 37666
rect -6066 37623 -6057 37657
rect -6057 37623 -6023 37657
rect -6023 37623 -6014 37657
rect -6066 37614 -6014 37623
rect -5906 37657 -5854 37666
rect -5906 37623 -5897 37657
rect -5897 37623 -5863 37657
rect -5863 37623 -5854 37657
rect -5906 37614 -5854 37623
rect -5746 37657 -5694 37666
rect -5746 37623 -5737 37657
rect -5737 37623 -5703 37657
rect -5703 37623 -5694 37657
rect -5746 37614 -5694 37623
rect -5586 37657 -5534 37666
rect -5586 37623 -5577 37657
rect -5577 37623 -5543 37657
rect -5543 37623 -5534 37657
rect -5586 37614 -5534 37623
rect -5426 37657 -5374 37666
rect -5426 37623 -5417 37657
rect -5417 37623 -5383 37657
rect -5383 37623 -5374 37657
rect -5426 37614 -5374 37623
rect -5266 37657 -5214 37666
rect -5266 37623 -5257 37657
rect -5257 37623 -5223 37657
rect -5223 37623 -5214 37657
rect -5266 37614 -5214 37623
rect -5106 37657 -5054 37666
rect -5106 37623 -5097 37657
rect -5097 37623 -5063 37657
rect -5063 37623 -5054 37657
rect -5106 37614 -5054 37623
rect -4946 37657 -4894 37666
rect -4946 37623 -4937 37657
rect -4937 37623 -4903 37657
rect -4903 37623 -4894 37657
rect -4946 37614 -4894 37623
rect -4786 37657 -4734 37666
rect -4786 37623 -4777 37657
rect -4777 37623 -4743 37657
rect -4743 37623 -4734 37657
rect -4786 37614 -4734 37623
rect -4626 37657 -4574 37666
rect -4626 37623 -4617 37657
rect -4617 37623 -4583 37657
rect -4583 37623 -4574 37657
rect -4626 37614 -4574 37623
rect -4466 37657 -4414 37666
rect -4466 37623 -4457 37657
rect -4457 37623 -4423 37657
rect -4423 37623 -4414 37657
rect -4466 37614 -4414 37623
rect -4306 37657 -4254 37666
rect -4306 37623 -4297 37657
rect -4297 37623 -4263 37657
rect -4263 37623 -4254 37657
rect -4306 37614 -4254 37623
rect -4146 37657 -4094 37666
rect -4146 37623 -4137 37657
rect -4137 37623 -4103 37657
rect -4103 37623 -4094 37657
rect -4146 37614 -4094 37623
rect -3986 37657 -3934 37666
rect -3986 37623 -3977 37657
rect -3977 37623 -3943 37657
rect -3943 37623 -3934 37657
rect -3986 37614 -3934 37623
rect -3826 37657 -3774 37666
rect -3826 37623 -3817 37657
rect -3817 37623 -3783 37657
rect -3783 37623 -3774 37657
rect -3826 37614 -3774 37623
rect -3666 37657 -3614 37666
rect -3666 37623 -3657 37657
rect -3657 37623 -3623 37657
rect -3623 37623 -3614 37657
rect -3666 37614 -3614 37623
rect -3506 37657 -3454 37666
rect -3506 37623 -3497 37657
rect -3497 37623 -3463 37657
rect -3463 37623 -3454 37657
rect -3506 37614 -3454 37623
rect -3346 37657 -3294 37666
rect -3346 37623 -3337 37657
rect -3337 37623 -3303 37657
rect -3303 37623 -3294 37657
rect -3346 37614 -3294 37623
rect -3186 37657 -3134 37666
rect -3186 37623 -3177 37657
rect -3177 37623 -3143 37657
rect -3143 37623 -3134 37657
rect -3186 37614 -3134 37623
rect -3026 37657 -2974 37666
rect -3026 37623 -3017 37657
rect -3017 37623 -2983 37657
rect -2983 37623 -2974 37657
rect -3026 37614 -2974 37623
rect -2866 37657 -2814 37666
rect -2866 37623 -2857 37657
rect -2857 37623 -2823 37657
rect -2823 37623 -2814 37657
rect -2866 37614 -2814 37623
rect -2706 37657 -2654 37666
rect -2706 37623 -2697 37657
rect -2697 37623 -2663 37657
rect -2663 37623 -2654 37657
rect -2706 37614 -2654 37623
rect -2546 37657 -2494 37666
rect -2546 37623 -2537 37657
rect -2537 37623 -2503 37657
rect -2503 37623 -2494 37657
rect -2546 37614 -2494 37623
rect -2386 37657 -2334 37666
rect -2386 37623 -2377 37657
rect -2377 37623 -2343 37657
rect -2343 37623 -2334 37657
rect -2386 37614 -2334 37623
rect -2226 37657 -2174 37666
rect -2226 37623 -2217 37657
rect -2217 37623 -2183 37657
rect -2183 37623 -2174 37657
rect -2226 37614 -2174 37623
rect -2066 37657 -2014 37666
rect -2066 37623 -2057 37657
rect -2057 37623 -2023 37657
rect -2023 37623 -2014 37657
rect -2066 37614 -2014 37623
rect -1906 37657 -1854 37666
rect -1906 37623 -1897 37657
rect -1897 37623 -1863 37657
rect -1863 37623 -1854 37657
rect -1906 37614 -1854 37623
rect -1746 37657 -1694 37666
rect -1746 37623 -1737 37657
rect -1737 37623 -1703 37657
rect -1703 37623 -1694 37657
rect -1746 37614 -1694 37623
rect -1586 37657 -1534 37666
rect -1586 37623 -1577 37657
rect -1577 37623 -1543 37657
rect -1543 37623 -1534 37657
rect -1586 37614 -1534 37623
rect -1426 37657 -1374 37666
rect -1426 37623 -1417 37657
rect -1417 37623 -1383 37657
rect -1383 37623 -1374 37657
rect -1426 37614 -1374 37623
rect -1266 37657 -1214 37666
rect -1266 37623 -1257 37657
rect -1257 37623 -1223 37657
rect -1223 37623 -1214 37657
rect -1266 37614 -1214 37623
rect -1106 37657 -1054 37666
rect -1106 37623 -1097 37657
rect -1097 37623 -1063 37657
rect -1063 37623 -1054 37657
rect -1106 37614 -1054 37623
rect -946 37657 -894 37666
rect -946 37623 -937 37657
rect -937 37623 -903 37657
rect -903 37623 -894 37657
rect -946 37614 -894 37623
rect -786 37657 -734 37666
rect -786 37623 -777 37657
rect -777 37623 -743 37657
rect -743 37623 -734 37657
rect -786 37614 -734 37623
rect -626 37657 -574 37666
rect -626 37623 -617 37657
rect -617 37623 -583 37657
rect -583 37623 -574 37657
rect -626 37614 -574 37623
rect -466 37657 -414 37666
rect -466 37623 -457 37657
rect -457 37623 -423 37657
rect -423 37623 -414 37657
rect -466 37614 -414 37623
rect -306 37657 -254 37666
rect -306 37623 -297 37657
rect -297 37623 -263 37657
rect -263 37623 -254 37657
rect -306 37614 -254 37623
rect -146 37657 -94 37666
rect -146 37623 -137 37657
rect -137 37623 -103 37657
rect -103 37623 -94 37657
rect -146 37614 -94 37623
rect 14 37657 66 37666
rect 14 37623 23 37657
rect 23 37623 57 37657
rect 57 37623 66 37657
rect 14 37614 66 37623
rect 76734 36617 76786 36626
rect 76734 36583 76743 36617
rect 76743 36583 76777 36617
rect 76777 36583 76786 36617
rect 76734 36574 76786 36583
rect 76894 36617 76946 36626
rect 76894 36583 76903 36617
rect 76903 36583 76937 36617
rect 76937 36583 76946 36617
rect 76894 36574 76946 36583
rect 76734 36297 76786 36306
rect 76734 36263 76743 36297
rect 76743 36263 76777 36297
rect 76777 36263 76786 36297
rect 76734 36254 76786 36263
rect 76894 36297 76946 36306
rect 76894 36263 76903 36297
rect 76903 36263 76937 36297
rect 76937 36263 76946 36297
rect 76894 36254 76946 36263
rect -2546 35257 -2494 35266
rect -2546 35223 -2537 35257
rect -2537 35223 -2503 35257
rect -2503 35223 -2494 35257
rect -2546 35214 -2494 35223
rect -2386 35257 -2334 35266
rect -2386 35223 -2377 35257
rect -2377 35223 -2343 35257
rect -2343 35223 -2334 35257
rect -2386 35214 -2334 35223
rect -2226 35257 -2174 35266
rect -2226 35223 -2217 35257
rect -2217 35223 -2183 35257
rect -2183 35223 -2174 35257
rect -2226 35214 -2174 35223
rect -2066 35257 -2014 35266
rect -2066 35223 -2057 35257
rect -2057 35223 -2023 35257
rect -2023 35223 -2014 35257
rect -2066 35214 -2014 35223
rect -1906 35257 -1854 35266
rect -1906 35223 -1897 35257
rect -1897 35223 -1863 35257
rect -1863 35223 -1854 35257
rect -1906 35214 -1854 35223
rect -1746 35257 -1694 35266
rect -1746 35223 -1737 35257
rect -1737 35223 -1703 35257
rect -1703 35223 -1694 35257
rect -1746 35214 -1694 35223
rect -1586 35257 -1534 35266
rect -1586 35223 -1577 35257
rect -1577 35223 -1543 35257
rect -1543 35223 -1534 35257
rect -1586 35214 -1534 35223
rect -1426 35257 -1374 35266
rect -1426 35223 -1417 35257
rect -1417 35223 -1383 35257
rect -1383 35223 -1374 35257
rect -1426 35214 -1374 35223
rect -1266 35257 -1214 35266
rect -1266 35223 -1257 35257
rect -1257 35223 -1223 35257
rect -1223 35223 -1214 35257
rect -1266 35214 -1214 35223
rect -1106 35257 -1054 35266
rect -1106 35223 -1097 35257
rect -1097 35223 -1063 35257
rect -1063 35223 -1054 35257
rect -1106 35214 -1054 35223
rect -946 35257 -894 35266
rect -946 35223 -937 35257
rect -937 35223 -903 35257
rect -903 35223 -894 35257
rect -946 35214 -894 35223
rect -786 35257 -734 35266
rect -786 35223 -777 35257
rect -777 35223 -743 35257
rect -743 35223 -734 35257
rect -786 35214 -734 35223
rect -626 35257 -574 35266
rect -626 35223 -617 35257
rect -617 35223 -583 35257
rect -583 35223 -574 35257
rect -626 35214 -574 35223
rect -466 35257 -414 35266
rect -466 35223 -457 35257
rect -457 35223 -423 35257
rect -423 35223 -414 35257
rect -466 35214 -414 35223
rect -306 35257 -254 35266
rect -306 35223 -297 35257
rect -297 35223 -263 35257
rect -263 35223 -254 35257
rect -306 35214 -254 35223
rect -146 35257 -94 35266
rect -146 35223 -137 35257
rect -137 35223 -103 35257
rect -103 35223 -94 35257
rect -146 35214 -94 35223
rect 14 35257 66 35266
rect 14 35223 23 35257
rect 23 35223 57 35257
rect 57 35223 66 35257
rect 14 35214 66 35223
rect -2546 34937 -2494 34946
rect -2546 34903 -2537 34937
rect -2537 34903 -2503 34937
rect -2503 34903 -2494 34937
rect -2546 34894 -2494 34903
rect -2386 34937 -2334 34946
rect -2386 34903 -2377 34937
rect -2377 34903 -2343 34937
rect -2343 34903 -2334 34937
rect -2386 34894 -2334 34903
rect -2226 34937 -2174 34946
rect -2226 34903 -2217 34937
rect -2217 34903 -2183 34937
rect -2183 34903 -2174 34937
rect -2226 34894 -2174 34903
rect -2066 34937 -2014 34946
rect -2066 34903 -2057 34937
rect -2057 34903 -2023 34937
rect -2023 34903 -2014 34937
rect -2066 34894 -2014 34903
rect -1906 34937 -1854 34946
rect -1906 34903 -1897 34937
rect -1897 34903 -1863 34937
rect -1863 34903 -1854 34937
rect -1906 34894 -1854 34903
rect -1746 34937 -1694 34946
rect -1746 34903 -1737 34937
rect -1737 34903 -1703 34937
rect -1703 34903 -1694 34937
rect -1746 34894 -1694 34903
rect -1586 34937 -1534 34946
rect -1586 34903 -1577 34937
rect -1577 34903 -1543 34937
rect -1543 34903 -1534 34937
rect -1586 34894 -1534 34903
rect -1426 34937 -1374 34946
rect -1426 34903 -1417 34937
rect -1417 34903 -1383 34937
rect -1383 34903 -1374 34937
rect -1426 34894 -1374 34903
rect -1266 34937 -1214 34946
rect -1266 34903 -1257 34937
rect -1257 34903 -1223 34937
rect -1223 34903 -1214 34937
rect -1266 34894 -1214 34903
rect -1106 34937 -1054 34946
rect -1106 34903 -1097 34937
rect -1097 34903 -1063 34937
rect -1063 34903 -1054 34937
rect -1106 34894 -1054 34903
rect -946 34937 -894 34946
rect -946 34903 -937 34937
rect -937 34903 -903 34937
rect -903 34903 -894 34937
rect -946 34894 -894 34903
rect -786 34937 -734 34946
rect -786 34903 -777 34937
rect -777 34903 -743 34937
rect -743 34903 -734 34937
rect -786 34894 -734 34903
rect -626 34937 -574 34946
rect -626 34903 -617 34937
rect -617 34903 -583 34937
rect -583 34903 -574 34937
rect -626 34894 -574 34903
rect -466 34937 -414 34946
rect -466 34903 -457 34937
rect -457 34903 -423 34937
rect -423 34903 -414 34937
rect -466 34894 -414 34903
rect -306 34937 -254 34946
rect -306 34903 -297 34937
rect -297 34903 -263 34937
rect -263 34903 -254 34937
rect -306 34894 -254 34903
rect -146 34937 -94 34946
rect -146 34903 -137 34937
rect -137 34903 -103 34937
rect -103 34903 -94 34937
rect -146 34894 -94 34903
rect 14 34937 66 34946
rect 14 34903 23 34937
rect 23 34903 57 34937
rect 57 34903 66 34937
rect 14 34894 66 34903
<< metal2 >>
rect 76880 44468 77440 44480
rect 76880 44412 76892 44468
rect 76948 44412 77440 44468
rect 76880 44400 77440 44412
rect 77040 43668 77440 43680
rect 77040 43612 77052 43668
rect 77108 43612 77372 43668
rect 77428 43612 77440 43668
rect 77040 43600 77440 43612
rect 77200 43508 77440 43520
rect 77200 43452 77212 43508
rect 77268 43452 77440 43508
rect 77200 43440 77440 43452
rect 77040 43348 77440 43360
rect 77040 43292 77052 43348
rect 77108 43292 77372 43348
rect 77428 43292 77440 43348
rect 77040 43280 77440 43292
rect 77040 43188 77440 43200
rect 77040 43132 77052 43188
rect 77108 43132 77372 43188
rect 77428 43132 77440 43188
rect 77040 43120 77440 43132
rect 77040 43028 77440 43040
rect 77040 42972 77052 43028
rect 77108 42972 77372 43028
rect 77428 42972 77440 43028
rect 77040 42960 77440 42972
rect 77040 42868 77440 42880
rect 77040 42812 77052 42868
rect 77108 42812 77372 42868
rect 77428 42812 77440 42868
rect 77040 42800 77440 42812
rect 77040 42708 77440 42720
rect 77040 42652 77052 42708
rect 77108 42652 77372 42708
rect 77428 42652 77440 42708
rect 77040 42640 77440 42652
rect 126640 42628 127040 42720
rect 77200 42548 77440 42560
rect 77200 42492 77212 42548
rect 77268 42492 77440 42548
rect 77200 42480 77440 42492
rect 126640 42412 126732 42628
rect 126948 42412 127040 42628
rect 77040 42388 77440 42400
rect 77040 42332 77052 42388
rect 77108 42332 77372 42388
rect 77428 42332 77440 42388
rect 77040 42320 77440 42332
rect 126640 42320 127040 42412
rect -1440 41828 -1040 41920
rect -960 41908 160 41920
rect -960 41852 -948 41908
rect -892 41852 -788 41908
rect -732 41852 -628 41908
rect -572 41852 -468 41908
rect -412 41852 -308 41908
rect -252 41852 -148 41908
rect -92 41852 12 41908
rect 68 41852 160 41908
rect -960 41840 160 41852
rect -1440 41612 -1348 41828
rect -1132 41760 -1040 41828
rect -1132 41680 80 41760
rect 76640 41748 76960 41760
rect 76640 41692 76892 41748
rect 76948 41692 76960 41748
rect 76640 41680 76960 41692
rect 77040 41748 77440 41760
rect 77040 41692 77052 41748
rect 77108 41692 77372 41748
rect 77428 41692 77440 41748
rect 77040 41680 77440 41692
rect -1132 41612 -1040 41680
rect -1440 41520 -1040 41612
rect -960 41588 160 41600
rect -960 41532 -948 41588
rect -892 41532 -788 41588
rect -732 41532 -628 41588
rect -572 41532 -468 41588
rect -412 41532 -308 41588
rect -252 41532 -148 41588
rect -92 41532 12 41588
rect 68 41532 160 41588
rect -960 41520 160 41532
rect 77200 41588 77440 41600
rect 77200 41532 77212 41588
rect 77268 41532 77440 41588
rect 77200 41520 77440 41532
rect 77040 41428 77440 41440
rect 77040 41372 77052 41428
rect 77108 41372 77372 41428
rect 77428 41372 77440 41428
rect 77040 41360 77440 41372
rect 77040 41268 77440 41280
rect 77040 41212 77052 41268
rect 77108 41212 77372 41268
rect 77428 41212 77440 41268
rect 77040 41200 77440 41212
rect 77040 41108 77440 41120
rect 77040 41052 77052 41108
rect 77108 41052 77372 41108
rect 77428 41052 77440 41108
rect 77040 41040 77440 41052
rect 77040 40948 77440 40960
rect 77040 40892 77052 40948
rect 77108 40892 77372 40948
rect 77428 40892 77440 40948
rect 77040 40880 77440 40892
rect 77040 40788 77440 40800
rect 77040 40732 77052 40788
rect 77108 40732 77372 40788
rect 77428 40732 77440 40788
rect 77040 40720 77440 40732
rect 76480 40628 77440 40640
rect 76480 40572 76732 40628
rect 76788 40572 76892 40628
rect 76948 40572 77052 40628
rect 77108 40572 77372 40628
rect 77428 40572 77440 40628
rect 76480 40560 77440 40572
rect 76640 40468 77440 40480
rect 76640 40412 77212 40468
rect 77268 40412 77440 40468
rect 76640 40400 77440 40412
rect 76480 40308 77440 40320
rect 76480 40252 76732 40308
rect 76788 40252 76892 40308
rect 76948 40252 77052 40308
rect 77108 40252 77372 40308
rect 77428 40252 77440 40308
rect 76480 40240 77440 40252
rect -7040 38308 160 38320
rect -7040 38252 -7028 38308
rect -6972 38252 -6868 38308
rect -6812 38252 -6708 38308
rect -6652 38252 -6548 38308
rect -6492 38252 -6388 38308
rect -6332 38306 -5748 38308
rect -6332 38254 -6226 38306
rect -6174 38254 -6066 38306
rect -6014 38254 -5906 38306
rect -5854 38254 -5748 38306
rect -6332 38252 -5748 38254
rect -5692 38252 -5588 38308
rect -5532 38252 -5428 38308
rect -5372 38252 -5268 38308
rect -5212 38252 -5108 38308
rect -5052 38252 -4948 38308
rect -4892 38252 -4788 38308
rect -4732 38306 -4148 38308
rect -4732 38254 -4626 38306
rect -4574 38254 -4466 38306
rect -4414 38254 -4306 38306
rect -4254 38254 -4148 38306
rect -4732 38252 -4148 38254
rect -4092 38252 -3988 38308
rect -3932 38252 -3828 38308
rect -3772 38252 -3668 38308
rect -3612 38252 -3508 38308
rect -3452 38252 -3348 38308
rect -3292 38252 -3188 38308
rect -3132 38252 -3028 38308
rect -2972 38252 -2868 38308
rect -2812 38252 -2708 38308
rect -2652 38252 -2548 38308
rect -2492 38252 -2388 38308
rect -2332 38252 -2228 38308
rect -2172 38252 -2068 38308
rect -2012 38252 -1908 38308
rect -1852 38252 -1748 38308
rect -1692 38252 -1588 38308
rect -1532 38252 -1428 38308
rect -1372 38252 -1268 38308
rect -1212 38252 -1108 38308
rect -1052 38252 -948 38308
rect -892 38252 -788 38308
rect -732 38252 -628 38308
rect -572 38252 -468 38308
rect -412 38252 -308 38308
rect -252 38252 -148 38308
rect -92 38252 12 38308
rect 68 38252 160 38308
rect -7040 38240 160 38252
rect -7040 38148 80 38160
rect -7040 38092 -6068 38148
rect -6012 38092 80 38148
rect -7040 38080 80 38092
rect -7040 37988 160 38000
rect -7040 37932 -7028 37988
rect -6972 37932 -6868 37988
rect -6812 37932 -6708 37988
rect -6652 37932 -6548 37988
rect -6492 37932 -6388 37988
rect -6332 37986 -5748 37988
rect -6332 37934 -6226 37986
rect -6174 37934 -6066 37986
rect -6014 37934 -5906 37986
rect -5854 37934 -5748 37986
rect -6332 37932 -5748 37934
rect -5692 37932 -5588 37988
rect -5532 37932 -5428 37988
rect -5372 37932 -5268 37988
rect -5212 37932 -5108 37988
rect -5052 37932 -4948 37988
rect -4892 37932 -4788 37988
rect -4732 37986 -4148 37988
rect -4732 37934 -4626 37986
rect -4574 37934 -4466 37986
rect -4414 37934 -4306 37986
rect -4254 37934 -4148 37986
rect -4732 37932 -4148 37934
rect -4092 37932 -3988 37988
rect -3932 37932 -3828 37988
rect -3772 37932 -3668 37988
rect -3612 37932 -3508 37988
rect -3452 37932 -3348 37988
rect -3292 37932 -3188 37988
rect -3132 37932 -3028 37988
rect -2972 37932 -2868 37988
rect -2812 37932 -2708 37988
rect -2652 37932 -2548 37988
rect -2492 37932 -2388 37988
rect -2332 37932 -2228 37988
rect -2172 37932 -2068 37988
rect -2012 37932 -1908 37988
rect -1852 37932 -1748 37988
rect -1692 37932 -1588 37988
rect -1532 37932 -1428 37988
rect -1372 37932 -1268 37988
rect -1212 37932 -1108 37988
rect -1052 37932 -948 37988
rect -892 37932 -788 37988
rect -732 37932 -628 37988
rect -572 37932 -468 37988
rect -412 37932 -308 37988
rect -252 37932 -148 37988
rect -92 37932 12 37988
rect 68 37932 160 37988
rect -7040 37920 160 37932
rect -7040 37828 80 37840
rect -7040 37772 -4468 37828
rect -4412 37772 80 37828
rect -7040 37760 80 37772
rect -7040 37668 160 37680
rect -7040 37612 -7028 37668
rect -6972 37612 -6868 37668
rect -6812 37612 -6708 37668
rect -6652 37612 -6548 37668
rect -6492 37612 -6388 37668
rect -6332 37666 -5748 37668
rect -6332 37614 -6226 37666
rect -6174 37614 -6066 37666
rect -6014 37614 -5906 37666
rect -5854 37614 -5748 37666
rect -6332 37612 -5748 37614
rect -5692 37612 -5588 37668
rect -5532 37612 -5428 37668
rect -5372 37612 -5268 37668
rect -5212 37612 -5108 37668
rect -5052 37612 -4948 37668
rect -4892 37612 -4788 37668
rect -4732 37666 -4148 37668
rect -4732 37614 -4626 37666
rect -4574 37614 -4466 37666
rect -4414 37614 -4306 37666
rect -4254 37614 -4148 37666
rect -4732 37612 -4148 37614
rect -4092 37612 -3988 37668
rect -3932 37612 -3828 37668
rect -3772 37612 -3668 37668
rect -3612 37612 -3508 37668
rect -3452 37612 -3348 37668
rect -3292 37612 -3188 37668
rect -3132 37612 -3028 37668
rect -2972 37612 -2868 37668
rect -2812 37612 -2708 37668
rect -2652 37612 -2548 37668
rect -2492 37612 -2388 37668
rect -2332 37612 -2228 37668
rect -2172 37612 -2068 37668
rect -2012 37612 -1908 37668
rect -1852 37612 -1748 37668
rect -1692 37612 -1588 37668
rect -1532 37612 -1428 37668
rect -1372 37612 -1268 37668
rect -1212 37612 -1108 37668
rect -1052 37612 -948 37668
rect -892 37612 -788 37668
rect -732 37612 -628 37668
rect -572 37612 -468 37668
rect -412 37612 -308 37668
rect -252 37612 -148 37668
rect -92 37612 12 37668
rect 68 37612 160 37668
rect -7040 37600 160 37612
rect 77040 36948 77440 36960
rect 77040 36892 77052 36948
rect 77108 36892 77372 36948
rect 77428 36892 77440 36948
rect 77040 36880 77440 36892
rect 77200 36788 77440 36800
rect 77200 36732 77212 36788
rect 77268 36732 77440 36788
rect 77200 36720 77440 36732
rect 76480 36628 77440 36640
rect 76480 36572 76732 36628
rect 76788 36572 76892 36628
rect 76948 36572 77052 36628
rect 77108 36572 77372 36628
rect 77428 36572 77440 36628
rect 76480 36560 77440 36572
rect 76640 36468 77280 36480
rect 76640 36412 77212 36468
rect 77268 36412 77280 36468
rect 76640 36400 77280 36412
rect 76480 36308 77440 36320
rect 76480 36252 76732 36308
rect 76788 36252 76892 36308
rect 76948 36252 77052 36308
rect 77108 36252 77372 36308
rect 77428 36252 77440 36308
rect 76480 36240 77440 36252
rect 77040 35988 77440 36000
rect 77040 35932 77052 35988
rect 77108 35932 77372 35988
rect 77428 35932 77440 35988
rect 77040 35920 77440 35932
rect 126640 35908 127040 36000
rect 77200 35828 77440 35840
rect 77200 35772 77212 35828
rect 77268 35772 77440 35828
rect 77200 35760 77440 35772
rect 126640 35692 126732 35908
rect 126948 35692 127040 35908
rect 77040 35668 77440 35680
rect 77040 35612 77052 35668
rect 77108 35612 77372 35668
rect 77428 35612 77440 35668
rect 77040 35600 77440 35612
rect 126640 35600 127040 35692
rect 77040 35508 77440 35520
rect 77040 35452 77052 35508
rect 77108 35452 77372 35508
rect 77428 35452 77440 35508
rect 77040 35440 77440 35452
rect 77040 35348 77440 35360
rect 77040 35292 77052 35348
rect 77108 35292 77372 35348
rect 77428 35292 77440 35348
rect 77040 35280 77440 35292
rect -3040 35188 -2640 35280
rect -2560 35268 160 35280
rect -2560 35212 -2548 35268
rect -2492 35212 -2388 35268
rect -2332 35212 -2228 35268
rect -2172 35212 -2068 35268
rect -2012 35212 -1908 35268
rect -1852 35212 -1748 35268
rect -1692 35212 -1588 35268
rect -1532 35212 -1428 35268
rect -1372 35212 -1268 35268
rect -1212 35212 -1108 35268
rect -1052 35212 -948 35268
rect -892 35212 -788 35268
rect -732 35212 -628 35268
rect -572 35212 -468 35268
rect -412 35212 -308 35268
rect -252 35212 -148 35268
rect -92 35212 12 35268
rect 68 35212 160 35268
rect -2560 35200 160 35212
rect -3040 34972 -2948 35188
rect -2732 35120 -2640 35188
rect 77040 35188 77440 35200
rect 77040 35132 77052 35188
rect 77108 35132 77372 35188
rect 77428 35132 77440 35188
rect 77040 35120 77440 35132
rect -2732 35040 80 35120
rect -2732 34972 -2640 35040
rect -3040 34880 -2640 34972
rect 77040 35028 77440 35040
rect 77040 34972 77052 35028
rect 77108 34972 77372 35028
rect 77428 34972 77440 35028
rect 77040 34960 77440 34972
rect -2560 34948 160 34960
rect -2560 34892 -2548 34948
rect -2492 34892 -2388 34948
rect -2332 34892 -2228 34948
rect -2172 34892 -2068 34948
rect -2012 34892 -1908 34948
rect -1852 34892 -1748 34948
rect -1692 34892 -1588 34948
rect -1532 34892 -1428 34948
rect -1372 34892 -1268 34948
rect -1212 34892 -1108 34948
rect -1052 34892 -948 34948
rect -892 34892 -788 34948
rect -732 34892 -628 34948
rect -572 34892 -468 34948
rect -412 34892 -308 34948
rect -252 34892 -148 34948
rect -92 34892 12 34948
rect 68 34892 160 34948
rect -2560 34880 160 34892
rect 77200 34868 77440 34880
rect 77200 34812 77212 34868
rect 77268 34812 77440 34868
rect 77200 34800 77440 34812
rect 77040 34708 77440 34720
rect 77040 34652 77052 34708
rect 77108 34652 77372 34708
rect 77428 34652 77440 34708
rect 77040 34640 77440 34652
<< via2 >>
rect 76892 44412 76948 44468
rect 77052 43612 77108 43668
rect 77372 43612 77428 43668
rect 77212 43452 77268 43508
rect 77052 43292 77108 43348
rect 77372 43292 77428 43348
rect 77052 43132 77108 43188
rect 77372 43132 77428 43188
rect 77052 42972 77108 43028
rect 77372 42972 77428 43028
rect 77052 42812 77108 42868
rect 77372 42812 77428 42868
rect 77052 42652 77108 42708
rect 77372 42652 77428 42708
rect 77212 42492 77268 42548
rect 126732 42412 126948 42628
rect 77052 42332 77108 42388
rect 77372 42332 77428 42388
rect -948 41906 -892 41908
rect -948 41854 -946 41906
rect -946 41854 -894 41906
rect -894 41854 -892 41906
rect -948 41852 -892 41854
rect -788 41906 -732 41908
rect -788 41854 -786 41906
rect -786 41854 -734 41906
rect -734 41854 -732 41906
rect -788 41852 -732 41854
rect -628 41906 -572 41908
rect -628 41854 -626 41906
rect -626 41854 -574 41906
rect -574 41854 -572 41906
rect -628 41852 -572 41854
rect -468 41906 -412 41908
rect -468 41854 -466 41906
rect -466 41854 -414 41906
rect -414 41854 -412 41906
rect -468 41852 -412 41854
rect -308 41906 -252 41908
rect -308 41854 -306 41906
rect -306 41854 -254 41906
rect -254 41854 -252 41906
rect -308 41852 -252 41854
rect -148 41906 -92 41908
rect -148 41854 -146 41906
rect -146 41854 -94 41906
rect -94 41854 -92 41906
rect -148 41852 -92 41854
rect 12 41906 68 41908
rect 12 41854 14 41906
rect 14 41854 66 41906
rect 66 41854 68 41906
rect 12 41852 68 41854
rect -1348 41612 -1132 41828
rect 76892 41692 76948 41748
rect 77052 41692 77108 41748
rect 77372 41692 77428 41748
rect -948 41586 -892 41588
rect -948 41534 -946 41586
rect -946 41534 -894 41586
rect -894 41534 -892 41586
rect -948 41532 -892 41534
rect -788 41586 -732 41588
rect -788 41534 -786 41586
rect -786 41534 -734 41586
rect -734 41534 -732 41586
rect -788 41532 -732 41534
rect -628 41586 -572 41588
rect -628 41534 -626 41586
rect -626 41534 -574 41586
rect -574 41534 -572 41586
rect -628 41532 -572 41534
rect -468 41586 -412 41588
rect -468 41534 -466 41586
rect -466 41534 -414 41586
rect -414 41534 -412 41586
rect -468 41532 -412 41534
rect -308 41586 -252 41588
rect -308 41534 -306 41586
rect -306 41534 -254 41586
rect -254 41534 -252 41586
rect -308 41532 -252 41534
rect -148 41586 -92 41588
rect -148 41534 -146 41586
rect -146 41534 -94 41586
rect -94 41534 -92 41586
rect -148 41532 -92 41534
rect 12 41586 68 41588
rect 12 41534 14 41586
rect 14 41534 66 41586
rect 66 41534 68 41586
rect 12 41532 68 41534
rect 77212 41532 77268 41588
rect 77052 41372 77108 41428
rect 77372 41372 77428 41428
rect 77052 41212 77108 41268
rect 77372 41212 77428 41268
rect 77052 41052 77108 41108
rect 77372 41052 77428 41108
rect 77052 40892 77108 40948
rect 77372 40892 77428 40948
rect 77052 40732 77108 40788
rect 77372 40732 77428 40788
rect 76732 40626 76788 40628
rect 76732 40574 76734 40626
rect 76734 40574 76786 40626
rect 76786 40574 76788 40626
rect 76732 40572 76788 40574
rect 76892 40626 76948 40628
rect 76892 40574 76894 40626
rect 76894 40574 76946 40626
rect 76946 40574 76948 40626
rect 76892 40572 76948 40574
rect 77052 40572 77108 40628
rect 77372 40572 77428 40628
rect 77212 40412 77268 40468
rect 76732 40306 76788 40308
rect 76732 40254 76734 40306
rect 76734 40254 76786 40306
rect 76786 40254 76788 40306
rect 76732 40252 76788 40254
rect 76892 40306 76948 40308
rect 76892 40254 76894 40306
rect 76894 40254 76946 40306
rect 76946 40254 76948 40306
rect 76892 40252 76948 40254
rect 77052 40252 77108 40308
rect 77372 40252 77428 40308
rect -7028 38306 -6972 38308
rect -7028 38254 -7026 38306
rect -7026 38254 -6974 38306
rect -6974 38254 -6972 38306
rect -7028 38252 -6972 38254
rect -6868 38306 -6812 38308
rect -6868 38254 -6866 38306
rect -6866 38254 -6814 38306
rect -6814 38254 -6812 38306
rect -6868 38252 -6812 38254
rect -6708 38306 -6652 38308
rect -6708 38254 -6706 38306
rect -6706 38254 -6654 38306
rect -6654 38254 -6652 38306
rect -6708 38252 -6652 38254
rect -6548 38306 -6492 38308
rect -6548 38254 -6546 38306
rect -6546 38254 -6494 38306
rect -6494 38254 -6492 38306
rect -6548 38252 -6492 38254
rect -6388 38306 -6332 38308
rect -5748 38306 -5692 38308
rect -6388 38254 -6386 38306
rect -6386 38254 -6334 38306
rect -6334 38254 -6332 38306
rect -5748 38254 -5746 38306
rect -5746 38254 -5694 38306
rect -5694 38254 -5692 38306
rect -6388 38252 -6332 38254
rect -5748 38252 -5692 38254
rect -5588 38306 -5532 38308
rect -5588 38254 -5586 38306
rect -5586 38254 -5534 38306
rect -5534 38254 -5532 38306
rect -5588 38252 -5532 38254
rect -5428 38306 -5372 38308
rect -5428 38254 -5426 38306
rect -5426 38254 -5374 38306
rect -5374 38254 -5372 38306
rect -5428 38252 -5372 38254
rect -5268 38306 -5212 38308
rect -5268 38254 -5266 38306
rect -5266 38254 -5214 38306
rect -5214 38254 -5212 38306
rect -5268 38252 -5212 38254
rect -5108 38306 -5052 38308
rect -5108 38254 -5106 38306
rect -5106 38254 -5054 38306
rect -5054 38254 -5052 38306
rect -5108 38252 -5052 38254
rect -4948 38306 -4892 38308
rect -4948 38254 -4946 38306
rect -4946 38254 -4894 38306
rect -4894 38254 -4892 38306
rect -4948 38252 -4892 38254
rect -4788 38306 -4732 38308
rect -4148 38306 -4092 38308
rect -4788 38254 -4786 38306
rect -4786 38254 -4734 38306
rect -4734 38254 -4732 38306
rect -4148 38254 -4146 38306
rect -4146 38254 -4094 38306
rect -4094 38254 -4092 38306
rect -4788 38252 -4732 38254
rect -4148 38252 -4092 38254
rect -3988 38306 -3932 38308
rect -3988 38254 -3986 38306
rect -3986 38254 -3934 38306
rect -3934 38254 -3932 38306
rect -3988 38252 -3932 38254
rect -3828 38306 -3772 38308
rect -3828 38254 -3826 38306
rect -3826 38254 -3774 38306
rect -3774 38254 -3772 38306
rect -3828 38252 -3772 38254
rect -3668 38306 -3612 38308
rect -3668 38254 -3666 38306
rect -3666 38254 -3614 38306
rect -3614 38254 -3612 38306
rect -3668 38252 -3612 38254
rect -3508 38306 -3452 38308
rect -3508 38254 -3506 38306
rect -3506 38254 -3454 38306
rect -3454 38254 -3452 38306
rect -3508 38252 -3452 38254
rect -3348 38306 -3292 38308
rect -3348 38254 -3346 38306
rect -3346 38254 -3294 38306
rect -3294 38254 -3292 38306
rect -3348 38252 -3292 38254
rect -3188 38306 -3132 38308
rect -3188 38254 -3186 38306
rect -3186 38254 -3134 38306
rect -3134 38254 -3132 38306
rect -3188 38252 -3132 38254
rect -3028 38306 -2972 38308
rect -3028 38254 -3026 38306
rect -3026 38254 -2974 38306
rect -2974 38254 -2972 38306
rect -3028 38252 -2972 38254
rect -2868 38306 -2812 38308
rect -2868 38254 -2866 38306
rect -2866 38254 -2814 38306
rect -2814 38254 -2812 38306
rect -2868 38252 -2812 38254
rect -2708 38306 -2652 38308
rect -2708 38254 -2706 38306
rect -2706 38254 -2654 38306
rect -2654 38254 -2652 38306
rect -2708 38252 -2652 38254
rect -2548 38306 -2492 38308
rect -2548 38254 -2546 38306
rect -2546 38254 -2494 38306
rect -2494 38254 -2492 38306
rect -2548 38252 -2492 38254
rect -2388 38306 -2332 38308
rect -2388 38254 -2386 38306
rect -2386 38254 -2334 38306
rect -2334 38254 -2332 38306
rect -2388 38252 -2332 38254
rect -2228 38306 -2172 38308
rect -2228 38254 -2226 38306
rect -2226 38254 -2174 38306
rect -2174 38254 -2172 38306
rect -2228 38252 -2172 38254
rect -2068 38306 -2012 38308
rect -2068 38254 -2066 38306
rect -2066 38254 -2014 38306
rect -2014 38254 -2012 38306
rect -2068 38252 -2012 38254
rect -1908 38306 -1852 38308
rect -1908 38254 -1906 38306
rect -1906 38254 -1854 38306
rect -1854 38254 -1852 38306
rect -1908 38252 -1852 38254
rect -1748 38306 -1692 38308
rect -1748 38254 -1746 38306
rect -1746 38254 -1694 38306
rect -1694 38254 -1692 38306
rect -1748 38252 -1692 38254
rect -1588 38306 -1532 38308
rect -1588 38254 -1586 38306
rect -1586 38254 -1534 38306
rect -1534 38254 -1532 38306
rect -1588 38252 -1532 38254
rect -1428 38306 -1372 38308
rect -1428 38254 -1426 38306
rect -1426 38254 -1374 38306
rect -1374 38254 -1372 38306
rect -1428 38252 -1372 38254
rect -1268 38306 -1212 38308
rect -1268 38254 -1266 38306
rect -1266 38254 -1214 38306
rect -1214 38254 -1212 38306
rect -1268 38252 -1212 38254
rect -1108 38306 -1052 38308
rect -1108 38254 -1106 38306
rect -1106 38254 -1054 38306
rect -1054 38254 -1052 38306
rect -1108 38252 -1052 38254
rect -948 38306 -892 38308
rect -948 38254 -946 38306
rect -946 38254 -894 38306
rect -894 38254 -892 38306
rect -948 38252 -892 38254
rect -788 38306 -732 38308
rect -788 38254 -786 38306
rect -786 38254 -734 38306
rect -734 38254 -732 38306
rect -788 38252 -732 38254
rect -628 38306 -572 38308
rect -628 38254 -626 38306
rect -626 38254 -574 38306
rect -574 38254 -572 38306
rect -628 38252 -572 38254
rect -468 38306 -412 38308
rect -468 38254 -466 38306
rect -466 38254 -414 38306
rect -414 38254 -412 38306
rect -468 38252 -412 38254
rect -308 38306 -252 38308
rect -308 38254 -306 38306
rect -306 38254 -254 38306
rect -254 38254 -252 38306
rect -308 38252 -252 38254
rect -148 38306 -92 38308
rect -148 38254 -146 38306
rect -146 38254 -94 38306
rect -94 38254 -92 38306
rect -148 38252 -92 38254
rect 12 38306 68 38308
rect 12 38254 14 38306
rect 14 38254 66 38306
rect 66 38254 68 38306
rect 12 38252 68 38254
rect -6068 38092 -6012 38148
rect -7028 37986 -6972 37988
rect -7028 37934 -7026 37986
rect -7026 37934 -6974 37986
rect -6974 37934 -6972 37986
rect -7028 37932 -6972 37934
rect -6868 37986 -6812 37988
rect -6868 37934 -6866 37986
rect -6866 37934 -6814 37986
rect -6814 37934 -6812 37986
rect -6868 37932 -6812 37934
rect -6708 37986 -6652 37988
rect -6708 37934 -6706 37986
rect -6706 37934 -6654 37986
rect -6654 37934 -6652 37986
rect -6708 37932 -6652 37934
rect -6548 37986 -6492 37988
rect -6548 37934 -6546 37986
rect -6546 37934 -6494 37986
rect -6494 37934 -6492 37986
rect -6548 37932 -6492 37934
rect -6388 37986 -6332 37988
rect -5748 37986 -5692 37988
rect -6388 37934 -6386 37986
rect -6386 37934 -6334 37986
rect -6334 37934 -6332 37986
rect -5748 37934 -5746 37986
rect -5746 37934 -5694 37986
rect -5694 37934 -5692 37986
rect -6388 37932 -6332 37934
rect -5748 37932 -5692 37934
rect -5588 37986 -5532 37988
rect -5588 37934 -5586 37986
rect -5586 37934 -5534 37986
rect -5534 37934 -5532 37986
rect -5588 37932 -5532 37934
rect -5428 37986 -5372 37988
rect -5428 37934 -5426 37986
rect -5426 37934 -5374 37986
rect -5374 37934 -5372 37986
rect -5428 37932 -5372 37934
rect -5268 37986 -5212 37988
rect -5268 37934 -5266 37986
rect -5266 37934 -5214 37986
rect -5214 37934 -5212 37986
rect -5268 37932 -5212 37934
rect -5108 37986 -5052 37988
rect -5108 37934 -5106 37986
rect -5106 37934 -5054 37986
rect -5054 37934 -5052 37986
rect -5108 37932 -5052 37934
rect -4948 37986 -4892 37988
rect -4948 37934 -4946 37986
rect -4946 37934 -4894 37986
rect -4894 37934 -4892 37986
rect -4948 37932 -4892 37934
rect -4788 37986 -4732 37988
rect -4148 37986 -4092 37988
rect -4788 37934 -4786 37986
rect -4786 37934 -4734 37986
rect -4734 37934 -4732 37986
rect -4148 37934 -4146 37986
rect -4146 37934 -4094 37986
rect -4094 37934 -4092 37986
rect -4788 37932 -4732 37934
rect -4148 37932 -4092 37934
rect -3988 37986 -3932 37988
rect -3988 37934 -3986 37986
rect -3986 37934 -3934 37986
rect -3934 37934 -3932 37986
rect -3988 37932 -3932 37934
rect -3828 37986 -3772 37988
rect -3828 37934 -3826 37986
rect -3826 37934 -3774 37986
rect -3774 37934 -3772 37986
rect -3828 37932 -3772 37934
rect -3668 37986 -3612 37988
rect -3668 37934 -3666 37986
rect -3666 37934 -3614 37986
rect -3614 37934 -3612 37986
rect -3668 37932 -3612 37934
rect -3508 37986 -3452 37988
rect -3508 37934 -3506 37986
rect -3506 37934 -3454 37986
rect -3454 37934 -3452 37986
rect -3508 37932 -3452 37934
rect -3348 37986 -3292 37988
rect -3348 37934 -3346 37986
rect -3346 37934 -3294 37986
rect -3294 37934 -3292 37986
rect -3348 37932 -3292 37934
rect -3188 37986 -3132 37988
rect -3188 37934 -3186 37986
rect -3186 37934 -3134 37986
rect -3134 37934 -3132 37986
rect -3188 37932 -3132 37934
rect -3028 37986 -2972 37988
rect -3028 37934 -3026 37986
rect -3026 37934 -2974 37986
rect -2974 37934 -2972 37986
rect -3028 37932 -2972 37934
rect -2868 37986 -2812 37988
rect -2868 37934 -2866 37986
rect -2866 37934 -2814 37986
rect -2814 37934 -2812 37986
rect -2868 37932 -2812 37934
rect -2708 37986 -2652 37988
rect -2708 37934 -2706 37986
rect -2706 37934 -2654 37986
rect -2654 37934 -2652 37986
rect -2708 37932 -2652 37934
rect -2548 37986 -2492 37988
rect -2548 37934 -2546 37986
rect -2546 37934 -2494 37986
rect -2494 37934 -2492 37986
rect -2548 37932 -2492 37934
rect -2388 37986 -2332 37988
rect -2388 37934 -2386 37986
rect -2386 37934 -2334 37986
rect -2334 37934 -2332 37986
rect -2388 37932 -2332 37934
rect -2228 37986 -2172 37988
rect -2228 37934 -2226 37986
rect -2226 37934 -2174 37986
rect -2174 37934 -2172 37986
rect -2228 37932 -2172 37934
rect -2068 37986 -2012 37988
rect -2068 37934 -2066 37986
rect -2066 37934 -2014 37986
rect -2014 37934 -2012 37986
rect -2068 37932 -2012 37934
rect -1908 37986 -1852 37988
rect -1908 37934 -1906 37986
rect -1906 37934 -1854 37986
rect -1854 37934 -1852 37986
rect -1908 37932 -1852 37934
rect -1748 37986 -1692 37988
rect -1748 37934 -1746 37986
rect -1746 37934 -1694 37986
rect -1694 37934 -1692 37986
rect -1748 37932 -1692 37934
rect -1588 37986 -1532 37988
rect -1588 37934 -1586 37986
rect -1586 37934 -1534 37986
rect -1534 37934 -1532 37986
rect -1588 37932 -1532 37934
rect -1428 37986 -1372 37988
rect -1428 37934 -1426 37986
rect -1426 37934 -1374 37986
rect -1374 37934 -1372 37986
rect -1428 37932 -1372 37934
rect -1268 37986 -1212 37988
rect -1268 37934 -1266 37986
rect -1266 37934 -1214 37986
rect -1214 37934 -1212 37986
rect -1268 37932 -1212 37934
rect -1108 37986 -1052 37988
rect -1108 37934 -1106 37986
rect -1106 37934 -1054 37986
rect -1054 37934 -1052 37986
rect -1108 37932 -1052 37934
rect -948 37986 -892 37988
rect -948 37934 -946 37986
rect -946 37934 -894 37986
rect -894 37934 -892 37986
rect -948 37932 -892 37934
rect -788 37986 -732 37988
rect -788 37934 -786 37986
rect -786 37934 -734 37986
rect -734 37934 -732 37986
rect -788 37932 -732 37934
rect -628 37986 -572 37988
rect -628 37934 -626 37986
rect -626 37934 -574 37986
rect -574 37934 -572 37986
rect -628 37932 -572 37934
rect -468 37986 -412 37988
rect -468 37934 -466 37986
rect -466 37934 -414 37986
rect -414 37934 -412 37986
rect -468 37932 -412 37934
rect -308 37986 -252 37988
rect -308 37934 -306 37986
rect -306 37934 -254 37986
rect -254 37934 -252 37986
rect -308 37932 -252 37934
rect -148 37986 -92 37988
rect -148 37934 -146 37986
rect -146 37934 -94 37986
rect -94 37934 -92 37986
rect -148 37932 -92 37934
rect 12 37986 68 37988
rect 12 37934 14 37986
rect 14 37934 66 37986
rect 66 37934 68 37986
rect 12 37932 68 37934
rect -4468 37772 -4412 37828
rect -7028 37666 -6972 37668
rect -7028 37614 -7026 37666
rect -7026 37614 -6974 37666
rect -6974 37614 -6972 37666
rect -7028 37612 -6972 37614
rect -6868 37666 -6812 37668
rect -6868 37614 -6866 37666
rect -6866 37614 -6814 37666
rect -6814 37614 -6812 37666
rect -6868 37612 -6812 37614
rect -6708 37666 -6652 37668
rect -6708 37614 -6706 37666
rect -6706 37614 -6654 37666
rect -6654 37614 -6652 37666
rect -6708 37612 -6652 37614
rect -6548 37666 -6492 37668
rect -6548 37614 -6546 37666
rect -6546 37614 -6494 37666
rect -6494 37614 -6492 37666
rect -6548 37612 -6492 37614
rect -6388 37666 -6332 37668
rect -5748 37666 -5692 37668
rect -6388 37614 -6386 37666
rect -6386 37614 -6334 37666
rect -6334 37614 -6332 37666
rect -5748 37614 -5746 37666
rect -5746 37614 -5694 37666
rect -5694 37614 -5692 37666
rect -6388 37612 -6332 37614
rect -5748 37612 -5692 37614
rect -5588 37666 -5532 37668
rect -5588 37614 -5586 37666
rect -5586 37614 -5534 37666
rect -5534 37614 -5532 37666
rect -5588 37612 -5532 37614
rect -5428 37666 -5372 37668
rect -5428 37614 -5426 37666
rect -5426 37614 -5374 37666
rect -5374 37614 -5372 37666
rect -5428 37612 -5372 37614
rect -5268 37666 -5212 37668
rect -5268 37614 -5266 37666
rect -5266 37614 -5214 37666
rect -5214 37614 -5212 37666
rect -5268 37612 -5212 37614
rect -5108 37666 -5052 37668
rect -5108 37614 -5106 37666
rect -5106 37614 -5054 37666
rect -5054 37614 -5052 37666
rect -5108 37612 -5052 37614
rect -4948 37666 -4892 37668
rect -4948 37614 -4946 37666
rect -4946 37614 -4894 37666
rect -4894 37614 -4892 37666
rect -4948 37612 -4892 37614
rect -4788 37666 -4732 37668
rect -4148 37666 -4092 37668
rect -4788 37614 -4786 37666
rect -4786 37614 -4734 37666
rect -4734 37614 -4732 37666
rect -4148 37614 -4146 37666
rect -4146 37614 -4094 37666
rect -4094 37614 -4092 37666
rect -4788 37612 -4732 37614
rect -4148 37612 -4092 37614
rect -3988 37666 -3932 37668
rect -3988 37614 -3986 37666
rect -3986 37614 -3934 37666
rect -3934 37614 -3932 37666
rect -3988 37612 -3932 37614
rect -3828 37666 -3772 37668
rect -3828 37614 -3826 37666
rect -3826 37614 -3774 37666
rect -3774 37614 -3772 37666
rect -3828 37612 -3772 37614
rect -3668 37666 -3612 37668
rect -3668 37614 -3666 37666
rect -3666 37614 -3614 37666
rect -3614 37614 -3612 37666
rect -3668 37612 -3612 37614
rect -3508 37666 -3452 37668
rect -3508 37614 -3506 37666
rect -3506 37614 -3454 37666
rect -3454 37614 -3452 37666
rect -3508 37612 -3452 37614
rect -3348 37666 -3292 37668
rect -3348 37614 -3346 37666
rect -3346 37614 -3294 37666
rect -3294 37614 -3292 37666
rect -3348 37612 -3292 37614
rect -3188 37666 -3132 37668
rect -3188 37614 -3186 37666
rect -3186 37614 -3134 37666
rect -3134 37614 -3132 37666
rect -3188 37612 -3132 37614
rect -3028 37666 -2972 37668
rect -3028 37614 -3026 37666
rect -3026 37614 -2974 37666
rect -2974 37614 -2972 37666
rect -3028 37612 -2972 37614
rect -2868 37666 -2812 37668
rect -2868 37614 -2866 37666
rect -2866 37614 -2814 37666
rect -2814 37614 -2812 37666
rect -2868 37612 -2812 37614
rect -2708 37666 -2652 37668
rect -2708 37614 -2706 37666
rect -2706 37614 -2654 37666
rect -2654 37614 -2652 37666
rect -2708 37612 -2652 37614
rect -2548 37666 -2492 37668
rect -2548 37614 -2546 37666
rect -2546 37614 -2494 37666
rect -2494 37614 -2492 37666
rect -2548 37612 -2492 37614
rect -2388 37666 -2332 37668
rect -2388 37614 -2386 37666
rect -2386 37614 -2334 37666
rect -2334 37614 -2332 37666
rect -2388 37612 -2332 37614
rect -2228 37666 -2172 37668
rect -2228 37614 -2226 37666
rect -2226 37614 -2174 37666
rect -2174 37614 -2172 37666
rect -2228 37612 -2172 37614
rect -2068 37666 -2012 37668
rect -2068 37614 -2066 37666
rect -2066 37614 -2014 37666
rect -2014 37614 -2012 37666
rect -2068 37612 -2012 37614
rect -1908 37666 -1852 37668
rect -1908 37614 -1906 37666
rect -1906 37614 -1854 37666
rect -1854 37614 -1852 37666
rect -1908 37612 -1852 37614
rect -1748 37666 -1692 37668
rect -1748 37614 -1746 37666
rect -1746 37614 -1694 37666
rect -1694 37614 -1692 37666
rect -1748 37612 -1692 37614
rect -1588 37666 -1532 37668
rect -1588 37614 -1586 37666
rect -1586 37614 -1534 37666
rect -1534 37614 -1532 37666
rect -1588 37612 -1532 37614
rect -1428 37666 -1372 37668
rect -1428 37614 -1426 37666
rect -1426 37614 -1374 37666
rect -1374 37614 -1372 37666
rect -1428 37612 -1372 37614
rect -1268 37666 -1212 37668
rect -1268 37614 -1266 37666
rect -1266 37614 -1214 37666
rect -1214 37614 -1212 37666
rect -1268 37612 -1212 37614
rect -1108 37666 -1052 37668
rect -1108 37614 -1106 37666
rect -1106 37614 -1054 37666
rect -1054 37614 -1052 37666
rect -1108 37612 -1052 37614
rect -948 37666 -892 37668
rect -948 37614 -946 37666
rect -946 37614 -894 37666
rect -894 37614 -892 37666
rect -948 37612 -892 37614
rect -788 37666 -732 37668
rect -788 37614 -786 37666
rect -786 37614 -734 37666
rect -734 37614 -732 37666
rect -788 37612 -732 37614
rect -628 37666 -572 37668
rect -628 37614 -626 37666
rect -626 37614 -574 37666
rect -574 37614 -572 37666
rect -628 37612 -572 37614
rect -468 37666 -412 37668
rect -468 37614 -466 37666
rect -466 37614 -414 37666
rect -414 37614 -412 37666
rect -468 37612 -412 37614
rect -308 37666 -252 37668
rect -308 37614 -306 37666
rect -306 37614 -254 37666
rect -254 37614 -252 37666
rect -308 37612 -252 37614
rect -148 37666 -92 37668
rect -148 37614 -146 37666
rect -146 37614 -94 37666
rect -94 37614 -92 37666
rect -148 37612 -92 37614
rect 12 37666 68 37668
rect 12 37614 14 37666
rect 14 37614 66 37666
rect 66 37614 68 37666
rect 12 37612 68 37614
rect 77052 36892 77108 36948
rect 77372 36892 77428 36948
rect 77212 36732 77268 36788
rect 76732 36626 76788 36628
rect 76732 36574 76734 36626
rect 76734 36574 76786 36626
rect 76786 36574 76788 36626
rect 76732 36572 76788 36574
rect 76892 36626 76948 36628
rect 76892 36574 76894 36626
rect 76894 36574 76946 36626
rect 76946 36574 76948 36626
rect 76892 36572 76948 36574
rect 77052 36572 77108 36628
rect 77372 36572 77428 36628
rect 77212 36412 77268 36468
rect 76732 36306 76788 36308
rect 76732 36254 76734 36306
rect 76734 36254 76786 36306
rect 76786 36254 76788 36306
rect 76732 36252 76788 36254
rect 76892 36306 76948 36308
rect 76892 36254 76894 36306
rect 76894 36254 76946 36306
rect 76946 36254 76948 36306
rect 76892 36252 76948 36254
rect 77052 36252 77108 36308
rect 77372 36252 77428 36308
rect 77052 35932 77108 35988
rect 77372 35932 77428 35988
rect 77212 35772 77268 35828
rect 126732 35692 126948 35908
rect 77052 35612 77108 35668
rect 77372 35612 77428 35668
rect 77052 35452 77108 35508
rect 77372 35452 77428 35508
rect 77052 35292 77108 35348
rect 77372 35292 77428 35348
rect -2548 35266 -2492 35268
rect -2548 35214 -2546 35266
rect -2546 35214 -2494 35266
rect -2494 35214 -2492 35266
rect -2548 35212 -2492 35214
rect -2388 35266 -2332 35268
rect -2388 35214 -2386 35266
rect -2386 35214 -2334 35266
rect -2334 35214 -2332 35266
rect -2388 35212 -2332 35214
rect -2228 35266 -2172 35268
rect -2228 35214 -2226 35266
rect -2226 35214 -2174 35266
rect -2174 35214 -2172 35266
rect -2228 35212 -2172 35214
rect -2068 35266 -2012 35268
rect -2068 35214 -2066 35266
rect -2066 35214 -2014 35266
rect -2014 35214 -2012 35266
rect -2068 35212 -2012 35214
rect -1908 35266 -1852 35268
rect -1908 35214 -1906 35266
rect -1906 35214 -1854 35266
rect -1854 35214 -1852 35266
rect -1908 35212 -1852 35214
rect -1748 35266 -1692 35268
rect -1748 35214 -1746 35266
rect -1746 35214 -1694 35266
rect -1694 35214 -1692 35266
rect -1748 35212 -1692 35214
rect -1588 35266 -1532 35268
rect -1588 35214 -1586 35266
rect -1586 35214 -1534 35266
rect -1534 35214 -1532 35266
rect -1588 35212 -1532 35214
rect -1428 35266 -1372 35268
rect -1428 35214 -1426 35266
rect -1426 35214 -1374 35266
rect -1374 35214 -1372 35266
rect -1428 35212 -1372 35214
rect -1268 35266 -1212 35268
rect -1268 35214 -1266 35266
rect -1266 35214 -1214 35266
rect -1214 35214 -1212 35266
rect -1268 35212 -1212 35214
rect -1108 35266 -1052 35268
rect -1108 35214 -1106 35266
rect -1106 35214 -1054 35266
rect -1054 35214 -1052 35266
rect -1108 35212 -1052 35214
rect -948 35266 -892 35268
rect -948 35214 -946 35266
rect -946 35214 -894 35266
rect -894 35214 -892 35266
rect -948 35212 -892 35214
rect -788 35266 -732 35268
rect -788 35214 -786 35266
rect -786 35214 -734 35266
rect -734 35214 -732 35266
rect -788 35212 -732 35214
rect -628 35266 -572 35268
rect -628 35214 -626 35266
rect -626 35214 -574 35266
rect -574 35214 -572 35266
rect -628 35212 -572 35214
rect -468 35266 -412 35268
rect -468 35214 -466 35266
rect -466 35214 -414 35266
rect -414 35214 -412 35266
rect -468 35212 -412 35214
rect -308 35266 -252 35268
rect -308 35214 -306 35266
rect -306 35214 -254 35266
rect -254 35214 -252 35266
rect -308 35212 -252 35214
rect -148 35266 -92 35268
rect -148 35214 -146 35266
rect -146 35214 -94 35266
rect -94 35214 -92 35266
rect -148 35212 -92 35214
rect 12 35266 68 35268
rect 12 35214 14 35266
rect 14 35214 66 35266
rect 66 35214 68 35266
rect 12 35212 68 35214
rect -2948 34972 -2732 35188
rect 77052 35132 77108 35188
rect 77372 35132 77428 35188
rect 77052 34972 77108 35028
rect 77372 34972 77428 35028
rect -2548 34946 -2492 34948
rect -2548 34894 -2546 34946
rect -2546 34894 -2494 34946
rect -2494 34894 -2492 34946
rect -2548 34892 -2492 34894
rect -2388 34946 -2332 34948
rect -2388 34894 -2386 34946
rect -2386 34894 -2334 34946
rect -2334 34894 -2332 34946
rect -2388 34892 -2332 34894
rect -2228 34946 -2172 34948
rect -2228 34894 -2226 34946
rect -2226 34894 -2174 34946
rect -2174 34894 -2172 34946
rect -2228 34892 -2172 34894
rect -2068 34946 -2012 34948
rect -2068 34894 -2066 34946
rect -2066 34894 -2014 34946
rect -2014 34894 -2012 34946
rect -2068 34892 -2012 34894
rect -1908 34946 -1852 34948
rect -1908 34894 -1906 34946
rect -1906 34894 -1854 34946
rect -1854 34894 -1852 34946
rect -1908 34892 -1852 34894
rect -1748 34946 -1692 34948
rect -1748 34894 -1746 34946
rect -1746 34894 -1694 34946
rect -1694 34894 -1692 34946
rect -1748 34892 -1692 34894
rect -1588 34946 -1532 34948
rect -1588 34894 -1586 34946
rect -1586 34894 -1534 34946
rect -1534 34894 -1532 34946
rect -1588 34892 -1532 34894
rect -1428 34946 -1372 34948
rect -1428 34894 -1426 34946
rect -1426 34894 -1374 34946
rect -1374 34894 -1372 34946
rect -1428 34892 -1372 34894
rect -1268 34946 -1212 34948
rect -1268 34894 -1266 34946
rect -1266 34894 -1214 34946
rect -1214 34894 -1212 34946
rect -1268 34892 -1212 34894
rect -1108 34946 -1052 34948
rect -1108 34894 -1106 34946
rect -1106 34894 -1054 34946
rect -1054 34894 -1052 34946
rect -1108 34892 -1052 34894
rect -948 34946 -892 34948
rect -948 34894 -946 34946
rect -946 34894 -894 34946
rect -894 34894 -892 34946
rect -948 34892 -892 34894
rect -788 34946 -732 34948
rect -788 34894 -786 34946
rect -786 34894 -734 34946
rect -734 34894 -732 34946
rect -788 34892 -732 34894
rect -628 34946 -572 34948
rect -628 34894 -626 34946
rect -626 34894 -574 34946
rect -574 34894 -572 34946
rect -628 34892 -572 34894
rect -468 34946 -412 34948
rect -468 34894 -466 34946
rect -466 34894 -414 34946
rect -414 34894 -412 34946
rect -468 34892 -412 34894
rect -308 34946 -252 34948
rect -308 34894 -306 34946
rect -306 34894 -254 34946
rect -254 34894 -252 34946
rect -308 34892 -252 34894
rect -148 34946 -92 34948
rect -148 34894 -146 34946
rect -146 34894 -94 34946
rect -94 34894 -92 34946
rect -148 34892 -92 34894
rect 12 34946 68 34948
rect 12 34894 14 34946
rect 14 34894 66 34946
rect 66 34894 68 34946
rect 12 34892 68 34894
rect 77212 34812 77268 34868
rect 77052 34652 77108 34708
rect 77372 34652 77428 34708
<< metal3 >>
rect 76880 44468 76960 44480
rect 76880 44412 76892 44468
rect 76948 44412 76960 44468
rect -1440 41832 -1040 41920
rect -1440 41608 -1352 41832
rect -1128 41608 -1040 41832
rect -1440 41520 -1040 41608
rect -960 41908 -880 41920
rect -960 41852 -948 41908
rect -892 41852 -880 41908
rect -960 41588 -880 41852
rect -960 41532 -948 41588
rect -892 41532 -880 41588
rect -960 41520 -880 41532
rect -800 41908 -720 41920
rect -800 41852 -788 41908
rect -732 41852 -720 41908
rect -800 41588 -720 41852
rect -800 41532 -788 41588
rect -732 41532 -720 41588
rect -800 41520 -720 41532
rect -640 41908 -560 41920
rect -640 41852 -628 41908
rect -572 41852 -560 41908
rect -640 41588 -560 41852
rect -640 41532 -628 41588
rect -572 41532 -560 41588
rect -640 41520 -560 41532
rect -480 41908 -400 41920
rect -480 41852 -468 41908
rect -412 41852 -400 41908
rect -480 41588 -400 41852
rect -480 41532 -468 41588
rect -412 41532 -400 41588
rect -480 41520 -400 41532
rect -320 41908 -240 41920
rect -320 41852 -308 41908
rect -252 41852 -240 41908
rect -320 41588 -240 41852
rect -320 41532 -308 41588
rect -252 41532 -240 41588
rect -320 41520 -240 41532
rect -160 41908 -80 41920
rect -160 41852 -148 41908
rect -92 41852 -80 41908
rect -160 41588 -80 41852
rect -160 41532 -148 41588
rect -92 41532 -80 41588
rect -160 41520 -80 41532
rect 0 41908 80 41920
rect 0 41852 12 41908
rect 68 41852 80 41908
rect 0 41588 80 41852
rect 76880 41748 76960 44412
rect 77040 43672 77120 43680
rect 77040 43608 77048 43672
rect 77112 43608 77120 43672
rect 77040 43352 77120 43608
rect 77360 43672 77440 43680
rect 77360 43608 77368 43672
rect 77432 43608 77440 43672
rect 77040 43288 77048 43352
rect 77112 43288 77120 43352
rect 77040 43192 77120 43288
rect 77040 43128 77048 43192
rect 77112 43128 77120 43192
rect 77040 43032 77120 43128
rect 77040 42968 77048 43032
rect 77112 42968 77120 43032
rect 77040 42872 77120 42968
rect 77040 42808 77048 42872
rect 77112 42808 77120 42872
rect 77040 42712 77120 42808
rect 77040 42648 77048 42712
rect 77112 42648 77120 42712
rect 77040 42392 77120 42648
rect 77200 43508 77280 43520
rect 77200 43452 77212 43508
rect 77268 43452 77280 43508
rect 77200 42548 77280 43452
rect 77200 42492 77212 42548
rect 77268 42492 77280 42548
rect 77200 42480 77280 42492
rect 77360 43352 77440 43608
rect 77360 43288 77368 43352
rect 77432 43288 77440 43352
rect 77360 43192 77440 43288
rect 77360 43128 77368 43192
rect 77432 43128 77440 43192
rect 77360 43032 77440 43128
rect 77360 42968 77368 43032
rect 77432 42968 77440 43032
rect 77360 42872 77440 42968
rect 77360 42808 77368 42872
rect 77432 42808 77440 42872
rect 77360 42712 77440 42808
rect 77360 42648 77368 42712
rect 77432 42648 77440 42712
rect 77040 42328 77048 42392
rect 77112 42328 77120 42392
rect 77040 42320 77120 42328
rect 77360 42392 77440 42648
rect 77360 42328 77368 42392
rect 77432 42328 77440 42392
rect 77360 42320 77440 42328
rect 126640 42628 127040 42720
rect 126640 42412 126732 42628
rect 126948 42412 127040 42628
rect 76880 41692 76892 41748
rect 76948 41692 76960 41748
rect 76880 41680 76960 41692
rect 77040 41752 77120 41760
rect 77040 41688 77048 41752
rect 77112 41688 77120 41752
rect 0 41532 12 41588
rect 68 41532 80 41588
rect 0 41520 80 41532
rect 77040 41432 77120 41688
rect 77040 41368 77048 41432
rect 77112 41368 77120 41432
rect 77040 41272 77120 41368
rect 77040 41208 77048 41272
rect 77112 41208 77120 41272
rect 77040 41112 77120 41208
rect 77040 41048 77048 41112
rect 77112 41048 77120 41112
rect 77040 40952 77120 41048
rect 77040 40888 77048 40952
rect 77112 40888 77120 40952
rect 77040 40792 77120 40888
rect 77040 40728 77048 40792
rect 77112 40728 77120 40792
rect 76720 40628 76800 40640
rect 76720 40572 76732 40628
rect 76788 40572 76800 40628
rect 76720 40308 76800 40572
rect 76720 40252 76732 40308
rect 76788 40252 76800 40308
rect 76720 40240 76800 40252
rect 76880 40628 76960 40640
rect 76880 40572 76892 40628
rect 76948 40572 76960 40628
rect 76880 40308 76960 40572
rect 76880 40252 76892 40308
rect 76948 40252 76960 40308
rect 76880 40240 76960 40252
rect 77040 40632 77120 40728
rect 77040 40568 77048 40632
rect 77112 40568 77120 40632
rect 77040 40312 77120 40568
rect 77040 40248 77048 40312
rect 77112 40248 77120 40312
rect 77040 40240 77120 40248
rect 77200 41588 77280 41760
rect 77200 41532 77212 41588
rect 77268 41532 77280 41588
rect 77200 40468 77280 41532
rect 77200 40412 77212 40468
rect 77268 40412 77280 40468
rect 77200 40240 77280 40412
rect 77360 41752 77440 41760
rect 77360 41688 77368 41752
rect 77432 41688 77440 41752
rect 77360 41432 77440 41688
rect 77360 41368 77368 41432
rect 77432 41368 77440 41432
rect 77360 41272 77440 41368
rect 77360 41208 77368 41272
rect 77432 41208 77440 41272
rect 77360 41112 77440 41208
rect 77360 41048 77368 41112
rect 77432 41048 77440 41112
rect 77360 40952 77440 41048
rect 77360 40888 77368 40952
rect 77432 40888 77440 40952
rect 77360 40792 77440 40888
rect 77360 40728 77368 40792
rect 77432 40728 77440 40792
rect 77360 40632 77440 40728
rect 77360 40568 77368 40632
rect 77432 40568 77440 40632
rect 77360 40312 77440 40568
rect 77360 40248 77368 40312
rect 77432 40248 77440 40312
rect 77360 40240 77440 40248
rect 126640 40072 127040 42412
rect 126640 39848 126728 40072
rect 126952 39848 127040 40072
rect 126640 39760 127040 39848
rect 126640 38472 127040 38560
rect -7040 38308 -6960 38320
rect -7040 38252 -7028 38308
rect -6972 38252 -6960 38308
rect -7040 37988 -6960 38252
rect -7040 37932 -7028 37988
rect -6972 37932 -6960 37988
rect -7040 37668 -6960 37932
rect -7040 37612 -7028 37668
rect -6972 37612 -6960 37668
rect -7040 37600 -6960 37612
rect -6880 38308 -6800 38320
rect -6880 38252 -6868 38308
rect -6812 38252 -6800 38308
rect -6880 37988 -6800 38252
rect -6880 37932 -6868 37988
rect -6812 37932 -6800 37988
rect -6880 37668 -6800 37932
rect -6880 37612 -6868 37668
rect -6812 37612 -6800 37668
rect -6880 37600 -6800 37612
rect -6720 38308 -6640 38320
rect -6720 38252 -6708 38308
rect -6652 38252 -6640 38308
rect -6720 37988 -6640 38252
rect -6720 37932 -6708 37988
rect -6652 37932 -6640 37988
rect -6720 37668 -6640 37932
rect -6720 37612 -6708 37668
rect -6652 37612 -6640 37668
rect -6720 37600 -6640 37612
rect -6560 38308 -6480 38320
rect -6560 38252 -6548 38308
rect -6492 38252 -6480 38308
rect -6560 37988 -6480 38252
rect -6560 37932 -6548 37988
rect -6492 37932 -6480 37988
rect -6560 37668 -6480 37932
rect -6560 37612 -6548 37668
rect -6492 37612 -6480 37668
rect -6560 37600 -6480 37612
rect -6400 38308 -6320 38320
rect -6400 38252 -6388 38308
rect -6332 38252 -6320 38308
rect -6400 37988 -6320 38252
rect -6400 37932 -6388 37988
rect -6332 37932 -6320 37988
rect -6400 37668 -6320 37932
rect -6240 38232 -5840 38320
rect -6240 38008 -6152 38232
rect -5928 38008 -5840 38232
rect -6240 37920 -5840 38008
rect -5760 38308 -5680 38320
rect -5760 38252 -5748 38308
rect -5692 38252 -5680 38308
rect -5760 37988 -5680 38252
rect -5760 37932 -5748 37988
rect -5692 37932 -5680 37988
rect -6400 37612 -6388 37668
rect -6332 37612 -6320 37668
rect -6400 37600 -6320 37612
rect -5760 37668 -5680 37932
rect -5760 37612 -5748 37668
rect -5692 37612 -5680 37668
rect -5760 37600 -5680 37612
rect -5600 38308 -5520 38320
rect -5600 38252 -5588 38308
rect -5532 38252 -5520 38308
rect -5600 37988 -5520 38252
rect -5600 37932 -5588 37988
rect -5532 37932 -5520 37988
rect -5600 37668 -5520 37932
rect -5600 37612 -5588 37668
rect -5532 37612 -5520 37668
rect -5600 37600 -5520 37612
rect -5440 38308 -5360 38320
rect -5440 38252 -5428 38308
rect -5372 38252 -5360 38308
rect -5440 37988 -5360 38252
rect -5440 37932 -5428 37988
rect -5372 37932 -5360 37988
rect -5440 37668 -5360 37932
rect -5440 37612 -5428 37668
rect -5372 37612 -5360 37668
rect -5440 37600 -5360 37612
rect -5280 38308 -5200 38320
rect -5280 38252 -5268 38308
rect -5212 38252 -5200 38308
rect -5280 37988 -5200 38252
rect -5280 37932 -5268 37988
rect -5212 37932 -5200 37988
rect -5280 37668 -5200 37932
rect -5280 37612 -5268 37668
rect -5212 37612 -5200 37668
rect -5280 37600 -5200 37612
rect -5120 38308 -5040 38320
rect -5120 38252 -5108 38308
rect -5052 38252 -5040 38308
rect -5120 37988 -5040 38252
rect -5120 37932 -5108 37988
rect -5052 37932 -5040 37988
rect -5120 37668 -5040 37932
rect -5120 37612 -5108 37668
rect -5052 37612 -5040 37668
rect -5120 37600 -5040 37612
rect -4960 38308 -4880 38320
rect -4960 38252 -4948 38308
rect -4892 38252 -4880 38308
rect -4960 37988 -4880 38252
rect -4960 37932 -4948 37988
rect -4892 37932 -4880 37988
rect -4960 37668 -4880 37932
rect -4960 37612 -4948 37668
rect -4892 37612 -4880 37668
rect -4960 37600 -4880 37612
rect -4800 38308 -4720 38320
rect -4800 38252 -4788 38308
rect -4732 38252 -4720 38308
rect -4800 37988 -4720 38252
rect -4160 38308 -4080 38320
rect -4160 38252 -4148 38308
rect -4092 38252 -4080 38308
rect -4800 37932 -4788 37988
rect -4732 37932 -4720 37988
rect -4800 37668 -4720 37932
rect -4800 37612 -4788 37668
rect -4732 37612 -4720 37668
rect -4800 37600 -4720 37612
rect -4640 37912 -4240 38000
rect -4640 37688 -4552 37912
rect -4328 37688 -4240 37912
rect -4640 37600 -4240 37688
rect -4160 37988 -4080 38252
rect -4160 37932 -4148 37988
rect -4092 37932 -4080 37988
rect -4160 37668 -4080 37932
rect -4160 37612 -4148 37668
rect -4092 37612 -4080 37668
rect -4160 37600 -4080 37612
rect -4000 38308 -3920 38320
rect -4000 38252 -3988 38308
rect -3932 38252 -3920 38308
rect -4000 37988 -3920 38252
rect -4000 37932 -3988 37988
rect -3932 37932 -3920 37988
rect -4000 37668 -3920 37932
rect -4000 37612 -3988 37668
rect -3932 37612 -3920 37668
rect -4000 37600 -3920 37612
rect -3840 38308 -3760 38320
rect -3840 38252 -3828 38308
rect -3772 38252 -3760 38308
rect -3840 37988 -3760 38252
rect -3840 37932 -3828 37988
rect -3772 37932 -3760 37988
rect -3840 37668 -3760 37932
rect -3840 37612 -3828 37668
rect -3772 37612 -3760 37668
rect -3840 37600 -3760 37612
rect -3680 38308 -3600 38320
rect -3680 38252 -3668 38308
rect -3612 38252 -3600 38308
rect -3680 37988 -3600 38252
rect -3680 37932 -3668 37988
rect -3612 37932 -3600 37988
rect -3680 37668 -3600 37932
rect -3680 37612 -3668 37668
rect -3612 37612 -3600 37668
rect -3680 37600 -3600 37612
rect -3520 38308 -3440 38320
rect -3520 38252 -3508 38308
rect -3452 38252 -3440 38308
rect -3520 37988 -3440 38252
rect -3520 37932 -3508 37988
rect -3452 37932 -3440 37988
rect -3520 37668 -3440 37932
rect -3520 37612 -3508 37668
rect -3452 37612 -3440 37668
rect -3520 37600 -3440 37612
rect -3360 38308 -3280 38320
rect -3360 38252 -3348 38308
rect -3292 38252 -3280 38308
rect -3360 37988 -3280 38252
rect -3360 37932 -3348 37988
rect -3292 37932 -3280 37988
rect -3360 37668 -3280 37932
rect -3360 37612 -3348 37668
rect -3292 37612 -3280 37668
rect -3360 37600 -3280 37612
rect -3200 38308 -3120 38320
rect -3200 38252 -3188 38308
rect -3132 38252 -3120 38308
rect -3200 37988 -3120 38252
rect -3200 37932 -3188 37988
rect -3132 37932 -3120 37988
rect -3200 37668 -3120 37932
rect -3200 37612 -3188 37668
rect -3132 37612 -3120 37668
rect -3200 37600 -3120 37612
rect -3040 38308 -2960 38320
rect -3040 38252 -3028 38308
rect -2972 38252 -2960 38308
rect -3040 37988 -2960 38252
rect -3040 37932 -3028 37988
rect -2972 37932 -2960 37988
rect -3040 37668 -2960 37932
rect -3040 37612 -3028 37668
rect -2972 37612 -2960 37668
rect -3040 37600 -2960 37612
rect -2880 38308 -2800 38320
rect -2880 38252 -2868 38308
rect -2812 38252 -2800 38308
rect -2880 37988 -2800 38252
rect -2880 37932 -2868 37988
rect -2812 37932 -2800 37988
rect -2880 37668 -2800 37932
rect -2880 37612 -2868 37668
rect -2812 37612 -2800 37668
rect -2880 37600 -2800 37612
rect -2720 38308 -2640 38320
rect -2720 38252 -2708 38308
rect -2652 38252 -2640 38308
rect -2720 37988 -2640 38252
rect -2720 37932 -2708 37988
rect -2652 37932 -2640 37988
rect -2720 37668 -2640 37932
rect -2720 37612 -2708 37668
rect -2652 37612 -2640 37668
rect -2720 37600 -2640 37612
rect -2560 38308 -2480 38320
rect -2560 38252 -2548 38308
rect -2492 38252 -2480 38308
rect -2560 37988 -2480 38252
rect -2560 37932 -2548 37988
rect -2492 37932 -2480 37988
rect -2560 37668 -2480 37932
rect -2560 37612 -2548 37668
rect -2492 37612 -2480 37668
rect -2560 37600 -2480 37612
rect -2400 38308 -2320 38320
rect -2400 38252 -2388 38308
rect -2332 38252 -2320 38308
rect -2400 37988 -2320 38252
rect -2400 37932 -2388 37988
rect -2332 37932 -2320 37988
rect -2400 37668 -2320 37932
rect -2400 37612 -2388 37668
rect -2332 37612 -2320 37668
rect -2400 37600 -2320 37612
rect -2240 38308 -2160 38320
rect -2240 38252 -2228 38308
rect -2172 38252 -2160 38308
rect -2240 37988 -2160 38252
rect -2240 37932 -2228 37988
rect -2172 37932 -2160 37988
rect -2240 37668 -2160 37932
rect -2240 37612 -2228 37668
rect -2172 37612 -2160 37668
rect -2240 37600 -2160 37612
rect -2080 38308 -2000 38320
rect -2080 38252 -2068 38308
rect -2012 38252 -2000 38308
rect -2080 37988 -2000 38252
rect -2080 37932 -2068 37988
rect -2012 37932 -2000 37988
rect -2080 37668 -2000 37932
rect -2080 37612 -2068 37668
rect -2012 37612 -2000 37668
rect -2080 37600 -2000 37612
rect -1920 38308 -1840 38320
rect -1920 38252 -1908 38308
rect -1852 38252 -1840 38308
rect -1920 37988 -1840 38252
rect -1920 37932 -1908 37988
rect -1852 37932 -1840 37988
rect -1920 37668 -1840 37932
rect -1920 37612 -1908 37668
rect -1852 37612 -1840 37668
rect -1920 37600 -1840 37612
rect -1760 38308 -1680 38320
rect -1760 38252 -1748 38308
rect -1692 38252 -1680 38308
rect -1760 37988 -1680 38252
rect -1760 37932 -1748 37988
rect -1692 37932 -1680 37988
rect -1760 37668 -1680 37932
rect -1760 37612 -1748 37668
rect -1692 37612 -1680 37668
rect -1760 37600 -1680 37612
rect -1600 38308 -1520 38320
rect -1600 38252 -1588 38308
rect -1532 38252 -1520 38308
rect -1600 37988 -1520 38252
rect -1600 37932 -1588 37988
rect -1532 37932 -1520 37988
rect -1600 37668 -1520 37932
rect -1600 37612 -1588 37668
rect -1532 37612 -1520 37668
rect -1600 37600 -1520 37612
rect -1440 38308 -1360 38320
rect -1440 38252 -1428 38308
rect -1372 38252 -1360 38308
rect -1440 37988 -1360 38252
rect -1440 37932 -1428 37988
rect -1372 37932 -1360 37988
rect -1440 37668 -1360 37932
rect -1440 37612 -1428 37668
rect -1372 37612 -1360 37668
rect -1440 37600 -1360 37612
rect -1280 38308 -1200 38320
rect -1280 38252 -1268 38308
rect -1212 38252 -1200 38308
rect -1280 37988 -1200 38252
rect -1280 37932 -1268 37988
rect -1212 37932 -1200 37988
rect -1280 37668 -1200 37932
rect -1280 37612 -1268 37668
rect -1212 37612 -1200 37668
rect -1280 37600 -1200 37612
rect -1120 38308 -1040 38320
rect -1120 38252 -1108 38308
rect -1052 38252 -1040 38308
rect -1120 37988 -1040 38252
rect -1120 37932 -1108 37988
rect -1052 37932 -1040 37988
rect -1120 37668 -1040 37932
rect -1120 37612 -1108 37668
rect -1052 37612 -1040 37668
rect -1120 37600 -1040 37612
rect -960 38308 -880 38320
rect -960 38252 -948 38308
rect -892 38252 -880 38308
rect -960 37988 -880 38252
rect -960 37932 -948 37988
rect -892 37932 -880 37988
rect -960 37668 -880 37932
rect -960 37612 -948 37668
rect -892 37612 -880 37668
rect -960 37600 -880 37612
rect -800 38308 -720 38320
rect -800 38252 -788 38308
rect -732 38252 -720 38308
rect -800 37988 -720 38252
rect -800 37932 -788 37988
rect -732 37932 -720 37988
rect -800 37668 -720 37932
rect -800 37612 -788 37668
rect -732 37612 -720 37668
rect -800 37600 -720 37612
rect -640 38308 -560 38320
rect -640 38252 -628 38308
rect -572 38252 -560 38308
rect -640 37988 -560 38252
rect -640 37932 -628 37988
rect -572 37932 -560 37988
rect -640 37668 -560 37932
rect -640 37612 -628 37668
rect -572 37612 -560 37668
rect -640 37600 -560 37612
rect -480 38308 -400 38320
rect -480 38252 -468 38308
rect -412 38252 -400 38308
rect -480 37988 -400 38252
rect -480 37932 -468 37988
rect -412 37932 -400 37988
rect -480 37668 -400 37932
rect -480 37612 -468 37668
rect -412 37612 -400 37668
rect -480 37600 -400 37612
rect -320 38308 -240 38320
rect -320 38252 -308 38308
rect -252 38252 -240 38308
rect -320 37988 -240 38252
rect -320 37932 -308 37988
rect -252 37932 -240 37988
rect -320 37668 -240 37932
rect -320 37612 -308 37668
rect -252 37612 -240 37668
rect -320 37600 -240 37612
rect -160 38308 -80 38320
rect -160 38252 -148 38308
rect -92 38252 -80 38308
rect -160 37988 -80 38252
rect -160 37932 -148 37988
rect -92 37932 -80 37988
rect -160 37668 -80 37932
rect -160 37612 -148 37668
rect -92 37612 -80 37668
rect -160 37600 -80 37612
rect 0 38308 80 38320
rect 0 38252 12 38308
rect 68 38252 80 38308
rect 0 37988 80 38252
rect 0 37932 12 37988
rect 68 37932 80 37988
rect 0 37668 80 37932
rect 0 37612 12 37668
rect 68 37612 80 37668
rect 0 37600 80 37612
rect 126640 38248 126728 38472
rect 126952 38248 127040 38472
rect 77040 36952 77120 36960
rect 77040 36888 77048 36952
rect 77112 36888 77120 36952
rect 76720 36628 76800 36640
rect 76720 36572 76732 36628
rect 76788 36572 76800 36628
rect 76720 36308 76800 36572
rect 76720 36252 76732 36308
rect 76788 36252 76800 36308
rect 76720 36240 76800 36252
rect 76880 36628 76960 36640
rect 76880 36572 76892 36628
rect 76948 36572 76960 36628
rect 76880 36308 76960 36572
rect 76880 36252 76892 36308
rect 76948 36252 76960 36308
rect 76880 36240 76960 36252
rect 77040 36632 77120 36888
rect 77040 36568 77048 36632
rect 77112 36568 77120 36632
rect 77040 36312 77120 36568
rect 77040 36248 77048 36312
rect 77112 36248 77120 36312
rect 77040 36240 77120 36248
rect 77200 36788 77280 36960
rect 77200 36732 77212 36788
rect 77268 36732 77280 36788
rect 77200 36468 77280 36732
rect 77200 36412 77212 36468
rect 77268 36412 77280 36468
rect 77200 36240 77280 36412
rect 77360 36952 77440 36960
rect 77360 36888 77368 36952
rect 77432 36888 77440 36952
rect 77360 36632 77440 36888
rect 77360 36568 77368 36632
rect 77432 36568 77440 36632
rect 77360 36312 77440 36568
rect 77360 36248 77368 36312
rect 77432 36248 77440 36312
rect 77360 36240 77440 36248
rect 77040 35992 77120 36000
rect 77040 35928 77048 35992
rect 77112 35928 77120 35992
rect 77040 35672 77120 35928
rect 77360 35992 77440 36000
rect 77360 35928 77368 35992
rect 77432 35928 77440 35992
rect 77040 35608 77048 35672
rect 77112 35608 77120 35672
rect 77040 35512 77120 35608
rect 77040 35448 77048 35512
rect 77112 35448 77120 35512
rect 77040 35352 77120 35448
rect 77040 35288 77048 35352
rect 77112 35288 77120 35352
rect -3040 35192 -2640 35280
rect -3040 34968 -2952 35192
rect -2728 34968 -2640 35192
rect -3040 34880 -2640 34968
rect -2560 35268 -2480 35280
rect -2560 35212 -2548 35268
rect -2492 35212 -2480 35268
rect -2560 34948 -2480 35212
rect -2560 34892 -2548 34948
rect -2492 34892 -2480 34948
rect -2560 34880 -2480 34892
rect -2400 35268 -2320 35280
rect -2400 35212 -2388 35268
rect -2332 35212 -2320 35268
rect -2400 34948 -2320 35212
rect -2400 34892 -2388 34948
rect -2332 34892 -2320 34948
rect -2400 34880 -2320 34892
rect -2240 35268 -2160 35280
rect -2240 35212 -2228 35268
rect -2172 35212 -2160 35268
rect -2240 34948 -2160 35212
rect -2240 34892 -2228 34948
rect -2172 34892 -2160 34948
rect -2240 34880 -2160 34892
rect -2080 35268 -2000 35280
rect -2080 35212 -2068 35268
rect -2012 35212 -2000 35268
rect -2080 34948 -2000 35212
rect -2080 34892 -2068 34948
rect -2012 34892 -2000 34948
rect -2080 34880 -2000 34892
rect -1920 35268 -1840 35280
rect -1920 35212 -1908 35268
rect -1852 35212 -1840 35268
rect -1920 34948 -1840 35212
rect -1920 34892 -1908 34948
rect -1852 34892 -1840 34948
rect -1920 34880 -1840 34892
rect -1760 35268 -1680 35280
rect -1760 35212 -1748 35268
rect -1692 35212 -1680 35268
rect -1760 34948 -1680 35212
rect -1760 34892 -1748 34948
rect -1692 34892 -1680 34948
rect -1760 34880 -1680 34892
rect -1600 35268 -1520 35280
rect -1600 35212 -1588 35268
rect -1532 35212 -1520 35268
rect -1600 34948 -1520 35212
rect -1600 34892 -1588 34948
rect -1532 34892 -1520 34948
rect -1600 34880 -1520 34892
rect -1440 35268 -1360 35280
rect -1440 35212 -1428 35268
rect -1372 35212 -1360 35268
rect -1440 34948 -1360 35212
rect -1440 34892 -1428 34948
rect -1372 34892 -1360 34948
rect -1440 34880 -1360 34892
rect -1280 35268 -1200 35280
rect -1280 35212 -1268 35268
rect -1212 35212 -1200 35268
rect -1280 34948 -1200 35212
rect -1280 34892 -1268 34948
rect -1212 34892 -1200 34948
rect -1280 34880 -1200 34892
rect -1120 35268 -1040 35280
rect -1120 35212 -1108 35268
rect -1052 35212 -1040 35268
rect -1120 34948 -1040 35212
rect -1120 34892 -1108 34948
rect -1052 34892 -1040 34948
rect -1120 34880 -1040 34892
rect -960 35268 -880 35280
rect -960 35212 -948 35268
rect -892 35212 -880 35268
rect -960 34948 -880 35212
rect -960 34892 -948 34948
rect -892 34892 -880 34948
rect -960 34880 -880 34892
rect -800 35268 -720 35280
rect -800 35212 -788 35268
rect -732 35212 -720 35268
rect -800 34948 -720 35212
rect -800 34892 -788 34948
rect -732 34892 -720 34948
rect -800 34880 -720 34892
rect -640 35268 -560 35280
rect -640 35212 -628 35268
rect -572 35212 -560 35268
rect -640 34948 -560 35212
rect -640 34892 -628 34948
rect -572 34892 -560 34948
rect -640 34880 -560 34892
rect -480 35268 -400 35280
rect -480 35212 -468 35268
rect -412 35212 -400 35268
rect -480 34948 -400 35212
rect -480 34892 -468 34948
rect -412 34892 -400 34948
rect -480 34880 -400 34892
rect -320 35268 -240 35280
rect -320 35212 -308 35268
rect -252 35212 -240 35268
rect -320 34948 -240 35212
rect -320 34892 -308 34948
rect -252 34892 -240 34948
rect -320 34880 -240 34892
rect -160 35268 -80 35280
rect -160 35212 -148 35268
rect -92 35212 -80 35268
rect -160 34948 -80 35212
rect -160 34892 -148 34948
rect -92 34892 -80 34948
rect -160 34880 -80 34892
rect 0 35268 80 35280
rect 0 35212 12 35268
rect 68 35212 80 35268
rect 0 34948 80 35212
rect 0 34892 12 34948
rect 68 34892 80 34948
rect 0 34880 80 34892
rect 77040 35192 77120 35288
rect 77040 35128 77048 35192
rect 77112 35128 77120 35192
rect 77040 35032 77120 35128
rect 77040 34968 77048 35032
rect 77112 34968 77120 35032
rect 77040 34712 77120 34968
rect 77040 34648 77048 34712
rect 77112 34648 77120 34712
rect 77040 34640 77120 34648
rect 77200 35828 77280 35840
rect 77200 35772 77212 35828
rect 77268 35772 77280 35828
rect 77200 34868 77280 35772
rect 77200 34812 77212 34868
rect 77268 34812 77280 34868
rect 77200 34640 77280 34812
rect 77360 35672 77440 35928
rect 77360 35608 77368 35672
rect 77432 35608 77440 35672
rect 77360 35512 77440 35608
rect 126640 35908 127040 38248
rect 126640 35692 126732 35908
rect 126948 35692 127040 35908
rect 126640 35600 127040 35692
rect 77360 35448 77368 35512
rect 77432 35448 77440 35512
rect 77360 35352 77440 35448
rect 77360 35288 77368 35352
rect 77432 35288 77440 35352
rect 77360 35192 77440 35288
rect 77360 35128 77368 35192
rect 77432 35128 77440 35192
rect 77360 35032 77440 35128
rect 77360 34968 77368 35032
rect 77432 34968 77440 35032
rect 77360 34712 77440 34968
rect 77360 34648 77368 34712
rect 77432 34648 77440 34712
rect 77360 34640 77440 34648
<< via3 >>
rect -1352 41828 -1128 41832
rect -1352 41612 -1348 41828
rect -1348 41612 -1132 41828
rect -1132 41612 -1128 41828
rect -1352 41608 -1128 41612
rect 77048 43668 77112 43672
rect 77048 43612 77052 43668
rect 77052 43612 77108 43668
rect 77108 43612 77112 43668
rect 77048 43608 77112 43612
rect 77368 43668 77432 43672
rect 77368 43612 77372 43668
rect 77372 43612 77428 43668
rect 77428 43612 77432 43668
rect 77368 43608 77432 43612
rect 77048 43348 77112 43352
rect 77048 43292 77052 43348
rect 77052 43292 77108 43348
rect 77108 43292 77112 43348
rect 77048 43288 77112 43292
rect 77048 43188 77112 43192
rect 77048 43132 77052 43188
rect 77052 43132 77108 43188
rect 77108 43132 77112 43188
rect 77048 43128 77112 43132
rect 77048 43028 77112 43032
rect 77048 42972 77052 43028
rect 77052 42972 77108 43028
rect 77108 42972 77112 43028
rect 77048 42968 77112 42972
rect 77048 42868 77112 42872
rect 77048 42812 77052 42868
rect 77052 42812 77108 42868
rect 77108 42812 77112 42868
rect 77048 42808 77112 42812
rect 77048 42708 77112 42712
rect 77048 42652 77052 42708
rect 77052 42652 77108 42708
rect 77108 42652 77112 42708
rect 77048 42648 77112 42652
rect 77368 43348 77432 43352
rect 77368 43292 77372 43348
rect 77372 43292 77428 43348
rect 77428 43292 77432 43348
rect 77368 43288 77432 43292
rect 77368 43188 77432 43192
rect 77368 43132 77372 43188
rect 77372 43132 77428 43188
rect 77428 43132 77432 43188
rect 77368 43128 77432 43132
rect 77368 43028 77432 43032
rect 77368 42972 77372 43028
rect 77372 42972 77428 43028
rect 77428 42972 77432 43028
rect 77368 42968 77432 42972
rect 77368 42868 77432 42872
rect 77368 42812 77372 42868
rect 77372 42812 77428 42868
rect 77428 42812 77432 42868
rect 77368 42808 77432 42812
rect 77368 42708 77432 42712
rect 77368 42652 77372 42708
rect 77372 42652 77428 42708
rect 77428 42652 77432 42708
rect 77368 42648 77432 42652
rect 77048 42388 77112 42392
rect 77048 42332 77052 42388
rect 77052 42332 77108 42388
rect 77108 42332 77112 42388
rect 77048 42328 77112 42332
rect 77368 42388 77432 42392
rect 77368 42332 77372 42388
rect 77372 42332 77428 42388
rect 77428 42332 77432 42388
rect 77368 42328 77432 42332
rect 77048 41748 77112 41752
rect 77048 41692 77052 41748
rect 77052 41692 77108 41748
rect 77108 41692 77112 41748
rect 77048 41688 77112 41692
rect 77048 41428 77112 41432
rect 77048 41372 77052 41428
rect 77052 41372 77108 41428
rect 77108 41372 77112 41428
rect 77048 41368 77112 41372
rect 77048 41268 77112 41272
rect 77048 41212 77052 41268
rect 77052 41212 77108 41268
rect 77108 41212 77112 41268
rect 77048 41208 77112 41212
rect 77048 41108 77112 41112
rect 77048 41052 77052 41108
rect 77052 41052 77108 41108
rect 77108 41052 77112 41108
rect 77048 41048 77112 41052
rect 77048 40948 77112 40952
rect 77048 40892 77052 40948
rect 77052 40892 77108 40948
rect 77108 40892 77112 40948
rect 77048 40888 77112 40892
rect 77048 40788 77112 40792
rect 77048 40732 77052 40788
rect 77052 40732 77108 40788
rect 77108 40732 77112 40788
rect 77048 40728 77112 40732
rect 77048 40628 77112 40632
rect 77048 40572 77052 40628
rect 77052 40572 77108 40628
rect 77108 40572 77112 40628
rect 77048 40568 77112 40572
rect 77048 40308 77112 40312
rect 77048 40252 77052 40308
rect 77052 40252 77108 40308
rect 77108 40252 77112 40308
rect 77048 40248 77112 40252
rect 77368 41748 77432 41752
rect 77368 41692 77372 41748
rect 77372 41692 77428 41748
rect 77428 41692 77432 41748
rect 77368 41688 77432 41692
rect 77368 41428 77432 41432
rect 77368 41372 77372 41428
rect 77372 41372 77428 41428
rect 77428 41372 77432 41428
rect 77368 41368 77432 41372
rect 77368 41268 77432 41272
rect 77368 41212 77372 41268
rect 77372 41212 77428 41268
rect 77428 41212 77432 41268
rect 77368 41208 77432 41212
rect 77368 41108 77432 41112
rect 77368 41052 77372 41108
rect 77372 41052 77428 41108
rect 77428 41052 77432 41108
rect 77368 41048 77432 41052
rect 77368 40948 77432 40952
rect 77368 40892 77372 40948
rect 77372 40892 77428 40948
rect 77428 40892 77432 40948
rect 77368 40888 77432 40892
rect 77368 40788 77432 40792
rect 77368 40732 77372 40788
rect 77372 40732 77428 40788
rect 77428 40732 77432 40788
rect 77368 40728 77432 40732
rect 77368 40628 77432 40632
rect 77368 40572 77372 40628
rect 77372 40572 77428 40628
rect 77428 40572 77432 40628
rect 77368 40568 77432 40572
rect 77368 40308 77432 40312
rect 77368 40252 77372 40308
rect 77372 40252 77428 40308
rect 77428 40252 77432 40308
rect 77368 40248 77432 40252
rect 126728 39848 126952 40072
rect -6152 38148 -5928 38232
rect -6152 38092 -6068 38148
rect -6068 38092 -6012 38148
rect -6012 38092 -5928 38148
rect -6152 38008 -5928 38092
rect -4552 37828 -4328 37912
rect -4552 37772 -4468 37828
rect -4468 37772 -4412 37828
rect -4412 37772 -4328 37828
rect -4552 37688 -4328 37772
rect 126728 38248 126952 38472
rect 77048 36948 77112 36952
rect 77048 36892 77052 36948
rect 77052 36892 77108 36948
rect 77108 36892 77112 36948
rect 77048 36888 77112 36892
rect 77048 36628 77112 36632
rect 77048 36572 77052 36628
rect 77052 36572 77108 36628
rect 77108 36572 77112 36628
rect 77048 36568 77112 36572
rect 77048 36308 77112 36312
rect 77048 36252 77052 36308
rect 77052 36252 77108 36308
rect 77108 36252 77112 36308
rect 77048 36248 77112 36252
rect 77368 36948 77432 36952
rect 77368 36892 77372 36948
rect 77372 36892 77428 36948
rect 77428 36892 77432 36948
rect 77368 36888 77432 36892
rect 77368 36628 77432 36632
rect 77368 36572 77372 36628
rect 77372 36572 77428 36628
rect 77428 36572 77432 36628
rect 77368 36568 77432 36572
rect 77368 36308 77432 36312
rect 77368 36252 77372 36308
rect 77372 36252 77428 36308
rect 77428 36252 77432 36308
rect 77368 36248 77432 36252
rect 77048 35988 77112 35992
rect 77048 35932 77052 35988
rect 77052 35932 77108 35988
rect 77108 35932 77112 35988
rect 77048 35928 77112 35932
rect 77368 35988 77432 35992
rect 77368 35932 77372 35988
rect 77372 35932 77428 35988
rect 77428 35932 77432 35988
rect 77368 35928 77432 35932
rect 77048 35668 77112 35672
rect 77048 35612 77052 35668
rect 77052 35612 77108 35668
rect 77108 35612 77112 35668
rect 77048 35608 77112 35612
rect 77048 35508 77112 35512
rect 77048 35452 77052 35508
rect 77052 35452 77108 35508
rect 77108 35452 77112 35508
rect 77048 35448 77112 35452
rect 77048 35348 77112 35352
rect 77048 35292 77052 35348
rect 77052 35292 77108 35348
rect 77108 35292 77112 35348
rect 77048 35288 77112 35292
rect -2952 35188 -2728 35192
rect -2952 34972 -2948 35188
rect -2948 34972 -2732 35188
rect -2732 34972 -2728 35188
rect -2952 34968 -2728 34972
rect 77048 35188 77112 35192
rect 77048 35132 77052 35188
rect 77052 35132 77108 35188
rect 77108 35132 77112 35188
rect 77048 35128 77112 35132
rect 77048 35028 77112 35032
rect 77048 34972 77052 35028
rect 77052 34972 77108 35028
rect 77108 34972 77112 35028
rect 77048 34968 77112 34972
rect 77048 34708 77112 34712
rect 77048 34652 77052 34708
rect 77052 34652 77108 34708
rect 77108 34652 77112 34708
rect 77048 34648 77112 34652
rect 77368 35668 77432 35672
rect 77368 35612 77372 35668
rect 77372 35612 77428 35668
rect 77428 35612 77432 35668
rect 77368 35608 77432 35612
rect 77368 35508 77432 35512
rect 77368 35452 77372 35508
rect 77372 35452 77428 35508
rect 77428 35452 77432 35508
rect 77368 35448 77432 35452
rect 77368 35348 77432 35352
rect 77368 35292 77372 35348
rect 77372 35292 77428 35348
rect 77428 35292 77432 35348
rect 77368 35288 77432 35292
rect 77368 35188 77432 35192
rect 77368 35132 77372 35188
rect 77372 35132 77428 35188
rect 77428 35132 77432 35188
rect 77368 35128 77432 35132
rect 77368 35028 77432 35032
rect 77368 34972 77372 35028
rect 77372 34972 77428 35028
rect 77428 34972 77432 35028
rect 77368 34968 77432 34972
rect 77368 34708 77432 34712
rect 77368 34652 77372 34708
rect 77372 34652 77428 34708
rect 77428 34652 77432 34708
rect 77368 34648 77432 34652
<< metal4 >>
rect 76480 79518 80320 79600
rect 76480 79282 77602 79518
rect 77838 79282 80320 79518
rect 76480 79200 80320 79282
rect 76480 79038 80320 79120
rect 76480 78802 79202 79038
rect 79438 78802 80320 79038
rect 76480 78720 80320 78802
rect 76480 78558 80320 78640
rect 76480 78322 80002 78558
rect 80238 78322 80320 78558
rect 76480 78240 80320 78322
rect 77040 43672 77440 43680
rect 77040 43608 77048 43672
rect 77112 43608 77368 43672
rect 77432 43608 77440 43672
rect 77040 43600 77440 43608
rect 77040 43352 77440 43360
rect 77040 43288 77048 43352
rect 77112 43288 77368 43352
rect 77432 43288 77440 43352
rect 77040 43280 77440 43288
rect 77040 43192 77440 43200
rect 77040 43128 77048 43192
rect 77112 43128 77368 43192
rect 77432 43128 77440 43192
rect 77040 43120 77440 43128
rect 77040 43032 77440 43040
rect 77040 42968 77048 43032
rect 77112 42968 77368 43032
rect 77432 42968 77440 43032
rect 77040 42960 77440 42968
rect 77040 42872 77440 42880
rect 77040 42808 77048 42872
rect 77112 42808 77368 42872
rect 77432 42808 77440 42872
rect 77040 42800 77440 42808
rect 77040 42712 77440 42720
rect 77040 42648 77048 42712
rect 77112 42648 77368 42712
rect 77432 42648 77440 42712
rect 77040 42640 77440 42648
rect 77040 42392 77440 42400
rect 77040 42328 77048 42392
rect 77112 42328 77368 42392
rect 77432 42328 77440 42392
rect 77040 42320 77440 42328
rect -1440 41838 -1040 41920
rect -1440 41602 -1358 41838
rect -1122 41602 -1040 41838
rect 77040 41752 77440 41760
rect 77040 41688 77048 41752
rect 77112 41688 77368 41752
rect 77432 41688 77440 41752
rect 77040 41680 77440 41688
rect -1440 41520 -1040 41602
rect 77040 41432 77440 41440
rect 77040 41368 77048 41432
rect 77112 41368 77368 41432
rect 77432 41368 77440 41432
rect 77040 41360 77440 41368
rect 77040 41272 77440 41280
rect 77040 41208 77048 41272
rect 77112 41208 77368 41272
rect 77432 41208 77440 41272
rect 77040 41200 77440 41208
rect 77040 41112 77440 41120
rect 77040 41048 77048 41112
rect 77112 41048 77368 41112
rect 77432 41048 77440 41112
rect 77040 41040 77440 41048
rect 77040 40952 77440 40960
rect 77040 40888 77048 40952
rect 77112 40888 77368 40952
rect 77432 40888 77440 40952
rect 77040 40880 77440 40888
rect 124400 40878 127440 40960
rect 77040 40792 77440 40800
rect 77040 40728 77048 40792
rect 77112 40728 77368 40792
rect 77432 40728 77440 40792
rect 77040 40720 77440 40728
rect 124400 40642 124482 40878
rect 124718 40642 127440 40878
rect 77040 40632 77440 40640
rect 77040 40568 77048 40632
rect 77112 40568 77368 40632
rect 77432 40568 77440 40632
rect 77040 40560 77440 40568
rect 124400 40560 127440 40642
rect 77040 40312 77440 40320
rect 77040 40248 77048 40312
rect 77112 40248 77368 40312
rect 77432 40248 77440 40312
rect 77040 40240 77440 40248
rect 126640 40072 127440 40160
rect 126640 39848 126728 40072
rect 126952 39848 127440 40072
rect 126640 39760 127440 39848
rect 124400 39278 127440 39360
rect 124400 39042 124482 39278
rect 124718 39042 127440 39278
rect 124400 38960 127440 39042
rect 126640 38472 127440 38560
rect -6240 38238 -5840 38320
rect -6240 38002 -6158 38238
rect -5922 38002 -5840 38238
rect 126640 38248 126728 38472
rect 126952 38248 127440 38472
rect 126640 38160 127440 38248
rect -6240 37920 -5840 38002
rect -4640 37918 -4240 38000
rect -4640 37682 -4558 37918
rect -4322 37682 -4240 37918
rect -4640 37600 -4240 37682
rect 124400 37678 127440 37760
rect 124400 37442 124482 37678
rect 124718 37442 127440 37678
rect 124400 37360 127440 37442
rect 77040 36952 77440 36960
rect 77040 36888 77048 36952
rect 77112 36888 77368 36952
rect 77432 36888 77440 36952
rect 77040 36880 77440 36888
rect 77040 36632 77440 36640
rect 77040 36568 77048 36632
rect 77112 36568 77368 36632
rect 77432 36568 77440 36632
rect 77040 36560 77440 36568
rect 77040 36312 77440 36320
rect 77040 36248 77048 36312
rect 77112 36248 77368 36312
rect 77432 36248 77440 36312
rect 77040 36240 77440 36248
rect 77040 35992 77440 36000
rect 77040 35928 77048 35992
rect 77112 35928 77368 35992
rect 77432 35928 77440 35992
rect 77040 35920 77440 35928
rect 77040 35672 77440 35680
rect 77040 35608 77048 35672
rect 77112 35608 77368 35672
rect 77432 35608 77440 35672
rect 77040 35600 77440 35608
rect 77040 35512 77440 35520
rect 77040 35448 77048 35512
rect 77112 35448 77368 35512
rect 77432 35448 77440 35512
rect 77040 35440 77440 35448
rect 77040 35352 77440 35360
rect 77040 35288 77048 35352
rect 77112 35288 77368 35352
rect 77432 35288 77440 35352
rect 77040 35280 77440 35288
rect -3040 35198 -2640 35280
rect -3040 34962 -2958 35198
rect -2722 34962 -2640 35198
rect 77040 35192 77440 35200
rect 77040 35128 77048 35192
rect 77112 35128 77368 35192
rect 77432 35128 77440 35192
rect 77040 35120 77440 35128
rect -3040 34880 -2640 34962
rect 77040 35032 77440 35040
rect 77040 34968 77048 35032
rect 77112 34968 77368 35032
rect 77432 34968 77440 35032
rect 77040 34960 77440 34968
rect 77040 34712 77440 34720
rect 77040 34648 77048 34712
rect 77112 34648 77368 34712
rect 77432 34648 77440 34712
rect 77040 34640 77440 34648
<< via4 >>
rect 77602 79282 77838 79518
rect 79202 78802 79438 79038
rect 80002 78322 80238 78558
rect -1358 41832 -1122 41838
rect -1358 41608 -1352 41832
rect -1352 41608 -1128 41832
rect -1128 41608 -1122 41832
rect -1358 41602 -1122 41608
rect 124482 40642 124718 40878
rect 124482 39042 124718 39278
rect -6158 38232 -5922 38238
rect -6158 38008 -6152 38232
rect -6152 38008 -5928 38232
rect -5928 38008 -5922 38232
rect -6158 38002 -5922 38008
rect -4558 37912 -4322 37918
rect -4558 37688 -4552 37912
rect -4552 37688 -4328 37912
rect -4328 37688 -4322 37912
rect -4558 37682 -4322 37688
rect 124482 37442 124718 37678
rect -2958 35192 -2722 35198
rect -2958 34968 -2952 35192
rect -2952 34968 -2728 35192
rect -2728 34968 -2722 35192
rect -2958 34962 -2722 34968
<< metal5 >>
rect -7040 37600 -6640 79760
rect -6240 38238 -5840 79760
rect -6240 38002 -6158 38238
rect -5922 38002 -5840 38238
rect -6240 37600 -5840 38002
rect -5440 37600 -5040 79760
rect -4640 37918 -4240 79760
rect -4640 37682 -4558 37918
rect -4322 37682 -4240 37918
rect -4640 37600 -4240 37682
rect -3840 34880 -3440 79760
rect -3040 35198 -2640 79760
rect -3040 34962 -2958 35198
rect -2722 34962 -2640 35198
rect -3040 34880 -2640 34962
rect -2240 34880 -1840 79760
rect -1440 41838 -1040 79760
rect -1440 41602 -1358 41838
rect -1122 41602 -1040 41838
rect -1440 41520 -1040 41602
rect -640 38960 -240 79760
rect 160 79680 560 79760
rect 960 79680 1360 79760
rect 1760 79680 2160 79760
rect 77520 79518 77920 79600
rect 77520 79282 77602 79518
rect 77838 79282 77920 79518
rect 77520 78720 77920 79282
rect 79120 79038 79520 79600
rect 79120 78802 79202 79038
rect 79438 78802 79520 79038
rect 79120 78720 79520 78802
rect 79920 78720 80320 79600
rect 80000 78558 80240 78560
rect 80000 78322 80002 78558
rect 80238 78322 80240 78558
rect 80000 78320 80240 78322
rect 124400 40878 124800 40960
rect 124400 40642 124482 40878
rect 124718 40642 124800 40878
rect 124400 40560 124800 40642
rect 125200 40560 125600 40960
rect 126000 40560 126400 40960
rect 124480 39278 124720 39280
rect 124480 39042 124482 39278
rect 124718 39042 124720 39278
rect 124480 39040 124720 39042
rect 124400 37678 124800 37760
rect 124400 37442 124482 37678
rect 124718 37442 124800 37678
rect 124400 37360 124800 37442
rect 125200 37360 125600 37760
rect 126000 37360 126400 37760
use lna  lna
timestamp 1638148091
transform 1 0 33280 0 1 560
box -33280 -4240 43360 79120
use opamp_pair  buffer
timestamp 1638148091
transform 1 0 80720 0 1 44720
box -3280 -47440 45920 34000
<< labels >>
rlabel metal2 s 76640 40400 76720 40480 4 xp
rlabel metal2 s 76640 36400 76720 36480 4 xm
rlabel metal2 s -80 38080 0 38160 4 ip
port 1 nsew
rlabel metal2 s -80 37760 0 37840 4 im
port 2 nsew
rlabel metal5 s -6240 79680 -5840 79760 4 ip
port 1 nsew
rlabel metal5 s -4640 79680 -4240 79760 4 im
port 2 nsew
rlabel metal4 s 127360 38160 127440 38560 4 om
port 3 nsew
rlabel metal4 s 127360 39760 127440 40160 4 op
port 4 nsew
rlabel metal5 s -3040 79680 -2640 79760 4 fsb
port 5 nsew
rlabel metal5 s -1440 79680 -1040 79760 4 ib
port 6 nsew
rlabel metal5 s 160 79680 560 79760 4 vdda
port 7 nsew
rlabel metal5 s 960 79680 1360 79760 4 gnda
port 8 nsew
rlabel metal5 s 1760 79680 2160 79760 4 vssa
port 9 nsew
<< end >>
