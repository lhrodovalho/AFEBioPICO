**.subckt untitled
x1 net1 net2 net3 net3 n1_2
x2 net2 net2 net1 net3 n1_2
x3 net1 net2 net3 net3 n1_2
x4 net4 net4 net1 net3 n1_2
x5 net5 net2 net3 net3 n1_2
x6 net6 net6 net5 net3 n1_2
x7 net2 net8 net7 net9 p2_1
x8 net7 net24 net9 net9 p2_1
x9 net4 net8 net10 net9 p1_2
x10 net10 net24 net9 net9 p1_2
x11 net6 net8 net11 net9 p1_2
x12 net11 net24 net9 net9 p1_2
x13 net12 net13 net3 net3 n2_1
x14 net19 net13 net12 net3 n2_1
x15 net19 net8 net14 net9 p1_2
x16 net14 net8 net9 net9 p1_2
x17 net15 net4 net3 net3 n1_2
x18 net8 net4 net15 net3 n1_2
x19 net8 net8 net16 net9 p1_2
x20 net16 net25 net9 net9 p1_2
x21 net17 net6 net3 net3 n1_2
x22 net20 net6 net17 net3 n1_2
x23 net20 net8 net18 net9 p1_2
x24 net18 net25 net9 net9 p1_2
x25 net21 net22 net3 net3 n1_2
x26 net22 net22 net21 net3 n1_2
x27 __UNCONNECTED_PIN__0 net8 net23 net9 p1_2
x28 net23 net24 net9 net9 p1_2
x29 net27 net28 net3 net3 n1_2
x30 net24 net27 net28 net3 n1_2
x31 net26 net27 net9 net9 p2_1
x32 net9 net27 net26 net9 p2_1
**.ends

* expanding   symbol:  n1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_2.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_2.sch
.subckt n1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_1
xs X G S B n1_1
.ends


* expanding   symbol:  p2_1.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p2_1.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p2_1.sch
.subckt p2_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xl D G S B p1_1
xr D G S B p1_1
.ends


* expanding   symbol:  p1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_2.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_2.sch
.subckt p1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_1
xd D G X B p1_1
.ends


* expanding   symbol:  n2_1.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n2_1.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n2_1.sch
.subckt n2_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xr D G S B n1_1
xl D G S B n1_1
.ends


* expanding   symbol:  n1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_1.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_1.sch
.subckt n1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8_lvt L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  p1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_1.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_1.sch
.subckt p1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8_lvt L=8 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

** flattened .save nodes
.end
