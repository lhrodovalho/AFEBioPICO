* pseudo-resistor testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "pseudo.spice"
.include "pseudo_bias4x.spice"

vdd vdd 0 1.8
vss vss 0 0.0
ecm cm vss vdd vss 0.5

* DUT
X0 ga da pa cm gb db pb cm cm vss pseudo
*vba ga da 0.2
*vbb gb db 0.1
vp p cm dc 1m ac 1
epa pa cm p cm 1
epb pb cm p cm 1

x1 ib da ga gb db vss dc vss dd vdd vss pseudo_bias4x
ibias ib vss 1n

.save ib ga da db gb pa i(epa) i(epb)

*.option rshunt=1e18
.option gmin=1e-15
.option scale=1e-6
.control

	ac dec 1 1m 1m
	print abs(1/i(epa))

	dc vp -101m 100m 10m
	let ii = abs(i(epa))
	let ri = 1/abs(deriv(ii))
	wrdata pseudo_i.txt ii ri
	plot ylog ii
	plot ylog ri
	let vg = da
	let vd = ga
	plot vd-vg
	wrdata pseudo_v.txt vg vd vd-vg
    
.endc

.end
