* NGSPICE file created from pseudo_bias.ext - technology: sky130A

.subckt p8_1 D G S B SUB
X0 S G D B sky130_fd_pr__pfet_01v8_lvt ad=1.2e+13p pd=5.6e+07u as=1.2e+13p ps=5.6e+07u w=3e+06u l=8e+06u
X1 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X2 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X3 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X4 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X5 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X6 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X7 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
.ends

.subckt p1_8 D G S B SUB
X0 D G a7 B sky130_fd_pr__pfet_01v8_lvt ad=1.5e+12p pd=7e+06u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X1 a6 G a5 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X2 S G a1 B sky130_fd_pr__pfet_01v8_lvt ad=1.5e+12p pd=7e+06u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X3 a6 G a7 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X4 a2 G a3 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X5 a2 G a1 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X6 a4 G a5 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=0p ps=0u w=3e+06u l=8e+06u
X7 a4 G a3 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
.ends

.subckt pseudo_bias ib xa ya xb yb vdda gnda vssa
Xp8_1_0 vdda ib vdda vdda vssa p8_1
Xp8_1_1 ya xa vssa vdda vssa p8_1
Xp8_1_2 ib ib vdda vdda vssa p8_1
Xp8_1_3 yb xb vssa vdda vssa p8_1
Xp8_1_4 vdda ib vdda vdda vssa p8_1
Xp8_1_5 yb xb vssa vdda vssa p8_1
Xp8_1_6 vdda ib vdda vdda vssa p8_1
Xp8_1_7 ib ib vdda vdda vssa p8_1
Xp8_1_8 ya xa vssa vdda vssa p8_1
Xp8_1_9 vdda ib vdda vdda vssa p8_1
Xp1_8_0 ya ib vdda vdda vssa p1_8
Xp1_8_1 yb ib vdda vdda vssa p1_8
Xp1_8_2 yb ib vdda vdda vssa p1_8
Xp1_8_3 ya ib vdda vdda vssa p1_8
C0 gnda xa 125.51fF
C1 gnda ib 125.14fF
C2 gnda yb 81.24fF
C3 gnda xb 79.25fF
C4 gnda vdda 35.96fF
C5 gnda ya 127.58fF
.ends

