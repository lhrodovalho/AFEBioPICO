magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< pwell >>
rect -12906 7734 14906 7866
rect -12906 1466 -12774 7734
rect 14774 1466 14906 7734
rect -12906 1334 14906 1466
<< psubdiff >>
rect -12880 7817 14880 7840
rect -12880 7783 -12719 7817
rect -12685 7783 -12651 7817
rect -12617 7783 -12583 7817
rect -12549 7783 -12515 7817
rect -12481 7783 -12447 7817
rect -12413 7783 -12379 7817
rect -12345 7783 -12311 7817
rect -12277 7783 -12243 7817
rect -12209 7783 -12175 7817
rect -12141 7783 -12107 7817
rect -12073 7783 -12039 7817
rect -12005 7783 -11971 7817
rect -11937 7783 -11903 7817
rect -11869 7783 -11835 7817
rect -11801 7783 -11767 7817
rect -11733 7783 -11699 7817
rect -11665 7783 -11631 7817
rect -11597 7783 -11563 7817
rect -11529 7783 -11495 7817
rect -11461 7783 -11427 7817
rect -11393 7783 -11359 7817
rect -11325 7783 -11291 7817
rect -11257 7783 -11223 7817
rect -11189 7783 -11155 7817
rect -11121 7783 -11087 7817
rect -11053 7783 -11019 7817
rect -10985 7783 -10951 7817
rect -10917 7783 -10883 7817
rect -10849 7783 -10815 7817
rect -10781 7783 -10747 7817
rect -10713 7783 -10679 7817
rect -10645 7783 -10611 7817
rect -10577 7783 -10543 7817
rect -10509 7783 -10475 7817
rect -10441 7783 -10407 7817
rect -10373 7783 -10339 7817
rect -10305 7783 -10271 7817
rect -10237 7783 -10203 7817
rect -10169 7783 -10135 7817
rect -10101 7783 -10067 7817
rect -10033 7783 -9999 7817
rect -9965 7783 -9931 7817
rect -9897 7783 -9863 7817
rect -9829 7783 -9795 7817
rect -9761 7783 -9727 7817
rect -9693 7783 -9659 7817
rect -9625 7783 -9591 7817
rect -9557 7783 -9523 7817
rect -9489 7783 -9455 7817
rect -9421 7783 -9387 7817
rect -9353 7783 -9319 7817
rect -9285 7783 -9251 7817
rect -9217 7783 -9183 7817
rect -9149 7783 -9115 7817
rect -9081 7783 -9047 7817
rect -9013 7783 -8979 7817
rect -8945 7783 -8911 7817
rect -8877 7783 -8843 7817
rect -8809 7783 -8775 7817
rect -8741 7783 -8707 7817
rect -8673 7783 -8639 7817
rect -8605 7783 -8571 7817
rect -8537 7783 -8503 7817
rect -8469 7783 -8435 7817
rect -8401 7783 -8367 7817
rect -8333 7783 -8299 7817
rect -8265 7783 -8231 7817
rect -8197 7783 -8163 7817
rect -8129 7783 -8095 7817
rect -8061 7783 -8027 7817
rect -7993 7783 -7959 7817
rect -7925 7783 -7891 7817
rect -7857 7783 -7823 7817
rect -7789 7783 -7755 7817
rect -7721 7783 -7687 7817
rect -7653 7783 -7619 7817
rect -7585 7783 -7551 7817
rect -7517 7783 -7483 7817
rect -7449 7783 -7415 7817
rect -7381 7783 -7347 7817
rect -7313 7783 -7279 7817
rect -7245 7783 -7211 7817
rect -7177 7783 -7143 7817
rect -7109 7783 -7075 7817
rect -7041 7783 -7007 7817
rect -6973 7783 -6939 7817
rect -6905 7783 -6871 7817
rect -6837 7783 -6803 7817
rect -6769 7783 -6735 7817
rect -6701 7783 -6667 7817
rect -6633 7783 -6599 7817
rect -6565 7783 -6531 7817
rect -6497 7783 -6463 7817
rect -6429 7783 -6395 7817
rect -6361 7783 -6327 7817
rect -6293 7783 -6259 7817
rect -6225 7783 -6191 7817
rect -6157 7783 -6123 7817
rect -6089 7783 -6055 7817
rect -6021 7783 -5987 7817
rect -5953 7783 -5919 7817
rect -5885 7783 -5851 7817
rect -5817 7783 -5783 7817
rect -5749 7783 -5715 7817
rect -5681 7783 -5647 7817
rect -5613 7783 -5579 7817
rect -5545 7783 -5511 7817
rect -5477 7783 -5443 7817
rect -5409 7783 -5375 7817
rect -5341 7783 -5307 7817
rect -5273 7783 -5239 7817
rect -5205 7783 -5171 7817
rect -5137 7783 -5103 7817
rect -5069 7783 -5035 7817
rect -5001 7783 -4967 7817
rect -4933 7783 -4899 7817
rect -4865 7783 -4831 7817
rect -4797 7783 -4763 7817
rect -4729 7783 -4695 7817
rect -4661 7783 -4627 7817
rect -4593 7783 -4559 7817
rect -4525 7783 -4491 7817
rect -4457 7783 -4423 7817
rect -4389 7783 -4355 7817
rect -4321 7783 -4287 7817
rect -4253 7783 -4219 7817
rect -4185 7783 -4151 7817
rect -4117 7783 -4083 7817
rect -4049 7783 -4015 7817
rect -3981 7783 -3947 7817
rect -3913 7783 -3879 7817
rect -3845 7783 -3811 7817
rect -3777 7783 -3743 7817
rect -3709 7783 -3675 7817
rect -3641 7783 -3607 7817
rect -3573 7783 -3539 7817
rect -3505 7783 -3471 7817
rect -3437 7783 -3403 7817
rect -3369 7783 -3335 7817
rect -3301 7783 -3267 7817
rect -3233 7783 -3199 7817
rect -3165 7783 -3131 7817
rect -3097 7783 -3063 7817
rect -3029 7783 -2995 7817
rect -2961 7783 -2927 7817
rect -2893 7783 -2859 7817
rect -2825 7783 -2791 7817
rect -2757 7783 -2723 7817
rect -2689 7783 -2655 7817
rect -2621 7783 -2587 7817
rect -2553 7783 -2519 7817
rect -2485 7783 -2451 7817
rect -2417 7783 -2383 7817
rect -2349 7783 -2315 7817
rect -2281 7783 -2247 7817
rect -2213 7783 -2179 7817
rect -2145 7783 -2111 7817
rect -2077 7783 -2043 7817
rect -2009 7783 -1975 7817
rect -1941 7783 -1907 7817
rect -1873 7783 -1839 7817
rect -1805 7783 -1771 7817
rect -1737 7783 -1703 7817
rect -1669 7783 -1635 7817
rect -1601 7783 -1567 7817
rect -1533 7783 -1499 7817
rect -1465 7783 -1431 7817
rect -1397 7783 -1363 7817
rect -1329 7783 -1295 7817
rect -1261 7783 -1227 7817
rect -1193 7783 -1159 7817
rect -1125 7783 -1091 7817
rect -1057 7783 -1023 7817
rect -989 7783 -955 7817
rect -921 7783 -887 7817
rect -853 7783 -819 7817
rect -785 7783 -751 7817
rect -717 7783 -683 7817
rect -649 7783 -615 7817
rect -581 7783 -547 7817
rect -513 7783 -479 7817
rect -445 7783 -411 7817
rect -377 7783 -343 7817
rect -309 7783 -275 7817
rect -241 7783 -207 7817
rect -173 7783 -139 7817
rect -105 7783 -71 7817
rect -37 7783 -3 7817
rect 31 7783 65 7817
rect 99 7783 133 7817
rect 167 7783 201 7817
rect 235 7783 269 7817
rect 303 7783 337 7817
rect 371 7783 405 7817
rect 439 7783 473 7817
rect 507 7783 541 7817
rect 575 7783 609 7817
rect 643 7783 677 7817
rect 711 7783 745 7817
rect 779 7783 813 7817
rect 847 7783 881 7817
rect 915 7783 949 7817
rect 983 7783 1017 7817
rect 1051 7783 1085 7817
rect 1119 7783 1153 7817
rect 1187 7783 1221 7817
rect 1255 7783 1289 7817
rect 1323 7783 1357 7817
rect 1391 7783 1425 7817
rect 1459 7783 1493 7817
rect 1527 7783 1561 7817
rect 1595 7783 1629 7817
rect 1663 7783 1697 7817
rect 1731 7783 1765 7817
rect 1799 7783 1833 7817
rect 1867 7783 1901 7817
rect 1935 7783 1969 7817
rect 2003 7783 2037 7817
rect 2071 7783 2105 7817
rect 2139 7783 2173 7817
rect 2207 7783 2241 7817
rect 2275 7783 2309 7817
rect 2343 7783 2377 7817
rect 2411 7783 2445 7817
rect 2479 7783 2513 7817
rect 2547 7783 2581 7817
rect 2615 7783 2649 7817
rect 2683 7783 2717 7817
rect 2751 7783 2785 7817
rect 2819 7783 2853 7817
rect 2887 7783 2921 7817
rect 2955 7783 2989 7817
rect 3023 7783 3057 7817
rect 3091 7783 3125 7817
rect 3159 7783 3193 7817
rect 3227 7783 3261 7817
rect 3295 7783 3329 7817
rect 3363 7783 3397 7817
rect 3431 7783 3465 7817
rect 3499 7783 3533 7817
rect 3567 7783 3601 7817
rect 3635 7783 3669 7817
rect 3703 7783 3737 7817
rect 3771 7783 3805 7817
rect 3839 7783 3873 7817
rect 3907 7783 3941 7817
rect 3975 7783 4009 7817
rect 4043 7783 4077 7817
rect 4111 7783 4145 7817
rect 4179 7783 4213 7817
rect 4247 7783 4281 7817
rect 4315 7783 4349 7817
rect 4383 7783 4417 7817
rect 4451 7783 4485 7817
rect 4519 7783 4553 7817
rect 4587 7783 4621 7817
rect 4655 7783 4689 7817
rect 4723 7783 4757 7817
rect 4791 7783 4825 7817
rect 4859 7783 4893 7817
rect 4927 7783 4961 7817
rect 4995 7783 5029 7817
rect 5063 7783 5097 7817
rect 5131 7783 5165 7817
rect 5199 7783 5233 7817
rect 5267 7783 5301 7817
rect 5335 7783 5369 7817
rect 5403 7783 5437 7817
rect 5471 7783 5505 7817
rect 5539 7783 5573 7817
rect 5607 7783 5641 7817
rect 5675 7783 5709 7817
rect 5743 7783 5777 7817
rect 5811 7783 5845 7817
rect 5879 7783 5913 7817
rect 5947 7783 5981 7817
rect 6015 7783 6049 7817
rect 6083 7783 6117 7817
rect 6151 7783 6185 7817
rect 6219 7783 6253 7817
rect 6287 7783 6321 7817
rect 6355 7783 6389 7817
rect 6423 7783 6457 7817
rect 6491 7783 6525 7817
rect 6559 7783 6593 7817
rect 6627 7783 6661 7817
rect 6695 7783 6729 7817
rect 6763 7783 6797 7817
rect 6831 7783 6865 7817
rect 6899 7783 6933 7817
rect 6967 7783 7001 7817
rect 7035 7783 7069 7817
rect 7103 7783 7137 7817
rect 7171 7783 7205 7817
rect 7239 7783 7273 7817
rect 7307 7783 7341 7817
rect 7375 7783 7409 7817
rect 7443 7783 7477 7817
rect 7511 7783 7545 7817
rect 7579 7783 7613 7817
rect 7647 7783 7681 7817
rect 7715 7783 7749 7817
rect 7783 7783 7817 7817
rect 7851 7783 7885 7817
rect 7919 7783 7953 7817
rect 7987 7783 8021 7817
rect 8055 7783 8089 7817
rect 8123 7783 8157 7817
rect 8191 7783 8225 7817
rect 8259 7783 8293 7817
rect 8327 7783 8361 7817
rect 8395 7783 8429 7817
rect 8463 7783 8497 7817
rect 8531 7783 8565 7817
rect 8599 7783 8633 7817
rect 8667 7783 8701 7817
rect 8735 7783 8769 7817
rect 8803 7783 8837 7817
rect 8871 7783 8905 7817
rect 8939 7783 8973 7817
rect 9007 7783 9041 7817
rect 9075 7783 9109 7817
rect 9143 7783 9177 7817
rect 9211 7783 9245 7817
rect 9279 7783 9313 7817
rect 9347 7783 9381 7817
rect 9415 7783 9449 7817
rect 9483 7783 9517 7817
rect 9551 7783 9585 7817
rect 9619 7783 9653 7817
rect 9687 7783 9721 7817
rect 9755 7783 9789 7817
rect 9823 7783 9857 7817
rect 9891 7783 9925 7817
rect 9959 7783 9993 7817
rect 10027 7783 10061 7817
rect 10095 7783 10129 7817
rect 10163 7783 10197 7817
rect 10231 7783 10265 7817
rect 10299 7783 10333 7817
rect 10367 7783 10401 7817
rect 10435 7783 10469 7817
rect 10503 7783 10537 7817
rect 10571 7783 10605 7817
rect 10639 7783 10673 7817
rect 10707 7783 10741 7817
rect 10775 7783 10809 7817
rect 10843 7783 10877 7817
rect 10911 7783 10945 7817
rect 10979 7783 11013 7817
rect 11047 7783 11081 7817
rect 11115 7783 11149 7817
rect 11183 7783 11217 7817
rect 11251 7783 11285 7817
rect 11319 7783 11353 7817
rect 11387 7783 11421 7817
rect 11455 7783 11489 7817
rect 11523 7783 11557 7817
rect 11591 7783 11625 7817
rect 11659 7783 11693 7817
rect 11727 7783 11761 7817
rect 11795 7783 11829 7817
rect 11863 7783 11897 7817
rect 11931 7783 11965 7817
rect 11999 7783 12033 7817
rect 12067 7783 12101 7817
rect 12135 7783 12169 7817
rect 12203 7783 12237 7817
rect 12271 7783 12305 7817
rect 12339 7783 12373 7817
rect 12407 7783 12441 7817
rect 12475 7783 12509 7817
rect 12543 7783 12577 7817
rect 12611 7783 12645 7817
rect 12679 7783 12713 7817
rect 12747 7783 12781 7817
rect 12815 7783 12849 7817
rect 12883 7783 12917 7817
rect 12951 7783 12985 7817
rect 13019 7783 13053 7817
rect 13087 7783 13121 7817
rect 13155 7783 13189 7817
rect 13223 7783 13257 7817
rect 13291 7783 13325 7817
rect 13359 7783 13393 7817
rect 13427 7783 13461 7817
rect 13495 7783 13529 7817
rect 13563 7783 13597 7817
rect 13631 7783 13665 7817
rect 13699 7783 13733 7817
rect 13767 7783 13801 7817
rect 13835 7783 13869 7817
rect 13903 7783 13937 7817
rect 13971 7783 14005 7817
rect 14039 7783 14073 7817
rect 14107 7783 14141 7817
rect 14175 7783 14209 7817
rect 14243 7783 14277 7817
rect 14311 7783 14345 7817
rect 14379 7783 14413 7817
rect 14447 7783 14481 7817
rect 14515 7783 14549 7817
rect 14583 7783 14617 7817
rect 14651 7783 14685 7817
rect 14719 7783 14880 7817
rect -12880 7760 14880 7783
rect -12880 7677 -12800 7760
rect -12880 7643 -12857 7677
rect -12823 7643 -12800 7677
rect -12880 7609 -12800 7643
rect -12880 7575 -12857 7609
rect -12823 7575 -12800 7609
rect -12880 7541 -12800 7575
rect -12880 7507 -12857 7541
rect -12823 7507 -12800 7541
rect -12880 7473 -12800 7507
rect -12880 7439 -12857 7473
rect -12823 7439 -12800 7473
rect -12880 7405 -12800 7439
rect -12880 7371 -12857 7405
rect -12823 7371 -12800 7405
rect -12880 7337 -12800 7371
rect -12880 7303 -12857 7337
rect -12823 7303 -12800 7337
rect -12880 7269 -12800 7303
rect -12880 7235 -12857 7269
rect -12823 7235 -12800 7269
rect -12880 7201 -12800 7235
rect -12880 7167 -12857 7201
rect -12823 7167 -12800 7201
rect -12880 7133 -12800 7167
rect -12880 7099 -12857 7133
rect -12823 7099 -12800 7133
rect -12880 7065 -12800 7099
rect -12880 7031 -12857 7065
rect -12823 7031 -12800 7065
rect -12880 6997 -12800 7031
rect -12880 6963 -12857 6997
rect -12823 6963 -12800 6997
rect -12880 6929 -12800 6963
rect -12880 6895 -12857 6929
rect -12823 6895 -12800 6929
rect -12880 6861 -12800 6895
rect -12880 6827 -12857 6861
rect -12823 6827 -12800 6861
rect -12880 6793 -12800 6827
rect -12880 6759 -12857 6793
rect -12823 6759 -12800 6793
rect -12880 6725 -12800 6759
rect -12880 6691 -12857 6725
rect -12823 6691 -12800 6725
rect -12880 6657 -12800 6691
rect -12880 6623 -12857 6657
rect -12823 6623 -12800 6657
rect -12880 6589 -12800 6623
rect -12880 6555 -12857 6589
rect -12823 6555 -12800 6589
rect -12880 6521 -12800 6555
rect -12880 6487 -12857 6521
rect -12823 6487 -12800 6521
rect -12880 6453 -12800 6487
rect -12880 6419 -12857 6453
rect -12823 6419 -12800 6453
rect -12880 6385 -12800 6419
rect -12880 6351 -12857 6385
rect -12823 6351 -12800 6385
rect -12880 6317 -12800 6351
rect -12880 6283 -12857 6317
rect -12823 6283 -12800 6317
rect -12880 6249 -12800 6283
rect -12880 6215 -12857 6249
rect -12823 6215 -12800 6249
rect -12880 6181 -12800 6215
rect -12880 6147 -12857 6181
rect -12823 6147 -12800 6181
rect -12880 6113 -12800 6147
rect -12880 6079 -12857 6113
rect -12823 6079 -12800 6113
rect -12880 6045 -12800 6079
rect -12880 6011 -12857 6045
rect -12823 6011 -12800 6045
rect -12880 5977 -12800 6011
rect -12880 5943 -12857 5977
rect -12823 5943 -12800 5977
rect -12880 5909 -12800 5943
rect -12880 5875 -12857 5909
rect -12823 5875 -12800 5909
rect -12880 5841 -12800 5875
rect -12880 5807 -12857 5841
rect -12823 5807 -12800 5841
rect -12880 5773 -12800 5807
rect -12880 5739 -12857 5773
rect -12823 5739 -12800 5773
rect -12880 5705 -12800 5739
rect -12880 5671 -12857 5705
rect -12823 5671 -12800 5705
rect -12880 5637 -12800 5671
rect -12880 5603 -12857 5637
rect -12823 5603 -12800 5637
rect -12880 5569 -12800 5603
rect -12880 5535 -12857 5569
rect -12823 5535 -12800 5569
rect -12880 5501 -12800 5535
rect -12880 5467 -12857 5501
rect -12823 5467 -12800 5501
rect -12880 5433 -12800 5467
rect -12880 5399 -12857 5433
rect -12823 5399 -12800 5433
rect -12880 5365 -12800 5399
rect -12880 5331 -12857 5365
rect -12823 5331 -12800 5365
rect -12880 5297 -12800 5331
rect -12880 5263 -12857 5297
rect -12823 5263 -12800 5297
rect -12880 5229 -12800 5263
rect -12880 5195 -12857 5229
rect -12823 5195 -12800 5229
rect -12880 5161 -12800 5195
rect -12880 5127 -12857 5161
rect -12823 5127 -12800 5161
rect -12880 5093 -12800 5127
rect -12880 5059 -12857 5093
rect -12823 5059 -12800 5093
rect -12880 5025 -12800 5059
rect -12880 4991 -12857 5025
rect -12823 4991 -12800 5025
rect -12880 4957 -12800 4991
rect -12880 4923 -12857 4957
rect -12823 4923 -12800 4957
rect -12880 4889 -12800 4923
rect -12880 4855 -12857 4889
rect -12823 4855 -12800 4889
rect -12880 4821 -12800 4855
rect -12880 4787 -12857 4821
rect -12823 4787 -12800 4821
rect -12880 4753 -12800 4787
rect -12880 4719 -12857 4753
rect -12823 4719 -12800 4753
rect -12880 4685 -12800 4719
rect -12880 4651 -12857 4685
rect -12823 4651 -12800 4685
rect -12880 4617 -12800 4651
rect -12880 4583 -12857 4617
rect -12823 4583 -12800 4617
rect -12880 4549 -12800 4583
rect -12880 4515 -12857 4549
rect -12823 4515 -12800 4549
rect -12880 4481 -12800 4515
rect -12880 4447 -12857 4481
rect -12823 4447 -12800 4481
rect -12880 4413 -12800 4447
rect -12880 4379 -12857 4413
rect -12823 4379 -12800 4413
rect -12880 4345 -12800 4379
rect -12880 4311 -12857 4345
rect -12823 4311 -12800 4345
rect -12880 4277 -12800 4311
rect -12880 4243 -12857 4277
rect -12823 4243 -12800 4277
rect -12880 4209 -12800 4243
rect -12880 4175 -12857 4209
rect -12823 4175 -12800 4209
rect -12880 4141 -12800 4175
rect -12880 4107 -12857 4141
rect -12823 4107 -12800 4141
rect -12880 4073 -12800 4107
rect -12880 4039 -12857 4073
rect -12823 4039 -12800 4073
rect -12880 4005 -12800 4039
rect -12880 3971 -12857 4005
rect -12823 3971 -12800 4005
rect -12880 3937 -12800 3971
rect -12880 3903 -12857 3937
rect -12823 3903 -12800 3937
rect -12880 3869 -12800 3903
rect -12880 3835 -12857 3869
rect -12823 3835 -12800 3869
rect -12880 3801 -12800 3835
rect -12880 3767 -12857 3801
rect -12823 3767 -12800 3801
rect -12880 3733 -12800 3767
rect -12880 3699 -12857 3733
rect -12823 3699 -12800 3733
rect -12880 3665 -12800 3699
rect -12880 3631 -12857 3665
rect -12823 3631 -12800 3665
rect -12880 3597 -12800 3631
rect -12880 3563 -12857 3597
rect -12823 3563 -12800 3597
rect -12880 3529 -12800 3563
rect -12880 3495 -12857 3529
rect -12823 3495 -12800 3529
rect -12880 3461 -12800 3495
rect -12880 3427 -12857 3461
rect -12823 3427 -12800 3461
rect -12880 3393 -12800 3427
rect -12880 3359 -12857 3393
rect -12823 3359 -12800 3393
rect -12880 3325 -12800 3359
rect -12880 3291 -12857 3325
rect -12823 3291 -12800 3325
rect -12880 3257 -12800 3291
rect -12880 3223 -12857 3257
rect -12823 3223 -12800 3257
rect -12880 3189 -12800 3223
rect -12880 3155 -12857 3189
rect -12823 3155 -12800 3189
rect -12880 3121 -12800 3155
rect -12880 3087 -12857 3121
rect -12823 3087 -12800 3121
rect -12880 3053 -12800 3087
rect -12880 3019 -12857 3053
rect -12823 3019 -12800 3053
rect -12880 2985 -12800 3019
rect -12880 2951 -12857 2985
rect -12823 2951 -12800 2985
rect -12880 2917 -12800 2951
rect -12880 2883 -12857 2917
rect -12823 2883 -12800 2917
rect -12880 2849 -12800 2883
rect -12880 2815 -12857 2849
rect -12823 2815 -12800 2849
rect -12880 2781 -12800 2815
rect -12880 2747 -12857 2781
rect -12823 2747 -12800 2781
rect -12880 2713 -12800 2747
rect -12880 2679 -12857 2713
rect -12823 2679 -12800 2713
rect -12880 2645 -12800 2679
rect -12880 2611 -12857 2645
rect -12823 2611 -12800 2645
rect -12880 2577 -12800 2611
rect -12880 2543 -12857 2577
rect -12823 2543 -12800 2577
rect -12880 2509 -12800 2543
rect -12880 2475 -12857 2509
rect -12823 2475 -12800 2509
rect -12880 2441 -12800 2475
rect -12880 2407 -12857 2441
rect -12823 2407 -12800 2441
rect -12880 2373 -12800 2407
rect -12880 2339 -12857 2373
rect -12823 2339 -12800 2373
rect -12880 2305 -12800 2339
rect -12880 2271 -12857 2305
rect -12823 2271 -12800 2305
rect -12880 2237 -12800 2271
rect -12880 2203 -12857 2237
rect -12823 2203 -12800 2237
rect -12880 2169 -12800 2203
rect -12880 2135 -12857 2169
rect -12823 2135 -12800 2169
rect -12880 2101 -12800 2135
rect -12880 2067 -12857 2101
rect -12823 2067 -12800 2101
rect -12880 2033 -12800 2067
rect -12880 1999 -12857 2033
rect -12823 1999 -12800 2033
rect -12880 1965 -12800 1999
rect -12880 1931 -12857 1965
rect -12823 1931 -12800 1965
rect -12880 1897 -12800 1931
rect -12880 1863 -12857 1897
rect -12823 1863 -12800 1897
rect -12880 1829 -12800 1863
rect -12880 1795 -12857 1829
rect -12823 1795 -12800 1829
rect -12880 1761 -12800 1795
rect -12880 1727 -12857 1761
rect -12823 1727 -12800 1761
rect -12880 1693 -12800 1727
rect -12880 1659 -12857 1693
rect -12823 1659 -12800 1693
rect -12880 1625 -12800 1659
rect -12880 1591 -12857 1625
rect -12823 1591 -12800 1625
rect -12880 1557 -12800 1591
rect -12880 1523 -12857 1557
rect -12823 1523 -12800 1557
rect -12880 1440 -12800 1523
rect 14800 7677 14880 7760
rect 14800 7643 14823 7677
rect 14857 7643 14880 7677
rect 14800 7609 14880 7643
rect 14800 7575 14823 7609
rect 14857 7575 14880 7609
rect 14800 7541 14880 7575
rect 14800 7507 14823 7541
rect 14857 7507 14880 7541
rect 14800 7473 14880 7507
rect 14800 7439 14823 7473
rect 14857 7439 14880 7473
rect 14800 7405 14880 7439
rect 14800 7371 14823 7405
rect 14857 7371 14880 7405
rect 14800 7337 14880 7371
rect 14800 7303 14823 7337
rect 14857 7303 14880 7337
rect 14800 7269 14880 7303
rect 14800 7235 14823 7269
rect 14857 7235 14880 7269
rect 14800 7201 14880 7235
rect 14800 7167 14823 7201
rect 14857 7167 14880 7201
rect 14800 7133 14880 7167
rect 14800 7099 14823 7133
rect 14857 7099 14880 7133
rect 14800 7065 14880 7099
rect 14800 7031 14823 7065
rect 14857 7031 14880 7065
rect 14800 6997 14880 7031
rect 14800 6963 14823 6997
rect 14857 6963 14880 6997
rect 14800 6929 14880 6963
rect 14800 6895 14823 6929
rect 14857 6895 14880 6929
rect 14800 6861 14880 6895
rect 14800 6827 14823 6861
rect 14857 6827 14880 6861
rect 14800 6793 14880 6827
rect 14800 6759 14823 6793
rect 14857 6759 14880 6793
rect 14800 6725 14880 6759
rect 14800 6691 14823 6725
rect 14857 6691 14880 6725
rect 14800 6657 14880 6691
rect 14800 6623 14823 6657
rect 14857 6623 14880 6657
rect 14800 6589 14880 6623
rect 14800 6555 14823 6589
rect 14857 6555 14880 6589
rect 14800 6521 14880 6555
rect 14800 6487 14823 6521
rect 14857 6487 14880 6521
rect 14800 6453 14880 6487
rect 14800 6419 14823 6453
rect 14857 6419 14880 6453
rect 14800 6385 14880 6419
rect 14800 6351 14823 6385
rect 14857 6351 14880 6385
rect 14800 6317 14880 6351
rect 14800 6283 14823 6317
rect 14857 6283 14880 6317
rect 14800 6249 14880 6283
rect 14800 6215 14823 6249
rect 14857 6215 14880 6249
rect 14800 6181 14880 6215
rect 14800 6147 14823 6181
rect 14857 6147 14880 6181
rect 14800 6113 14880 6147
rect 14800 6079 14823 6113
rect 14857 6079 14880 6113
rect 14800 6045 14880 6079
rect 14800 6011 14823 6045
rect 14857 6011 14880 6045
rect 14800 5977 14880 6011
rect 14800 5943 14823 5977
rect 14857 5943 14880 5977
rect 14800 5909 14880 5943
rect 14800 5875 14823 5909
rect 14857 5875 14880 5909
rect 14800 5841 14880 5875
rect 14800 5807 14823 5841
rect 14857 5807 14880 5841
rect 14800 5773 14880 5807
rect 14800 5739 14823 5773
rect 14857 5739 14880 5773
rect 14800 5705 14880 5739
rect 14800 5671 14823 5705
rect 14857 5671 14880 5705
rect 14800 5637 14880 5671
rect 14800 5603 14823 5637
rect 14857 5603 14880 5637
rect 14800 5569 14880 5603
rect 14800 5535 14823 5569
rect 14857 5535 14880 5569
rect 14800 5501 14880 5535
rect 14800 5467 14823 5501
rect 14857 5467 14880 5501
rect 14800 5433 14880 5467
rect 14800 5399 14823 5433
rect 14857 5399 14880 5433
rect 14800 5365 14880 5399
rect 14800 5331 14823 5365
rect 14857 5331 14880 5365
rect 14800 5297 14880 5331
rect 14800 5263 14823 5297
rect 14857 5263 14880 5297
rect 14800 5229 14880 5263
rect 14800 5195 14823 5229
rect 14857 5195 14880 5229
rect 14800 5161 14880 5195
rect 14800 5127 14823 5161
rect 14857 5127 14880 5161
rect 14800 5093 14880 5127
rect 14800 5059 14823 5093
rect 14857 5059 14880 5093
rect 14800 5025 14880 5059
rect 14800 4991 14823 5025
rect 14857 4991 14880 5025
rect 14800 4957 14880 4991
rect 14800 4923 14823 4957
rect 14857 4923 14880 4957
rect 14800 4889 14880 4923
rect 14800 4855 14823 4889
rect 14857 4855 14880 4889
rect 14800 4821 14880 4855
rect 14800 4787 14823 4821
rect 14857 4787 14880 4821
rect 14800 4753 14880 4787
rect 14800 4719 14823 4753
rect 14857 4719 14880 4753
rect 14800 4685 14880 4719
rect 14800 4651 14823 4685
rect 14857 4651 14880 4685
rect 14800 4617 14880 4651
rect 14800 4583 14823 4617
rect 14857 4583 14880 4617
rect 14800 4549 14880 4583
rect 14800 4515 14823 4549
rect 14857 4515 14880 4549
rect 14800 4481 14880 4515
rect 14800 4447 14823 4481
rect 14857 4447 14880 4481
rect 14800 4413 14880 4447
rect 14800 4379 14823 4413
rect 14857 4379 14880 4413
rect 14800 4345 14880 4379
rect 14800 4311 14823 4345
rect 14857 4311 14880 4345
rect 14800 4277 14880 4311
rect 14800 4243 14823 4277
rect 14857 4243 14880 4277
rect 14800 4209 14880 4243
rect 14800 4175 14823 4209
rect 14857 4175 14880 4209
rect 14800 4141 14880 4175
rect 14800 4107 14823 4141
rect 14857 4107 14880 4141
rect 14800 4073 14880 4107
rect 14800 4039 14823 4073
rect 14857 4039 14880 4073
rect 14800 4005 14880 4039
rect 14800 3971 14823 4005
rect 14857 3971 14880 4005
rect 14800 3937 14880 3971
rect 14800 3903 14823 3937
rect 14857 3903 14880 3937
rect 14800 3869 14880 3903
rect 14800 3835 14823 3869
rect 14857 3835 14880 3869
rect 14800 3801 14880 3835
rect 14800 3767 14823 3801
rect 14857 3767 14880 3801
rect 14800 3733 14880 3767
rect 14800 3699 14823 3733
rect 14857 3699 14880 3733
rect 14800 3665 14880 3699
rect 14800 3631 14823 3665
rect 14857 3631 14880 3665
rect 14800 3597 14880 3631
rect 14800 3563 14823 3597
rect 14857 3563 14880 3597
rect 14800 3529 14880 3563
rect 14800 3495 14823 3529
rect 14857 3495 14880 3529
rect 14800 3461 14880 3495
rect 14800 3427 14823 3461
rect 14857 3427 14880 3461
rect 14800 3393 14880 3427
rect 14800 3359 14823 3393
rect 14857 3359 14880 3393
rect 14800 3325 14880 3359
rect 14800 3291 14823 3325
rect 14857 3291 14880 3325
rect 14800 3257 14880 3291
rect 14800 3223 14823 3257
rect 14857 3223 14880 3257
rect 14800 3189 14880 3223
rect 14800 3155 14823 3189
rect 14857 3155 14880 3189
rect 14800 3121 14880 3155
rect 14800 3087 14823 3121
rect 14857 3087 14880 3121
rect 14800 3053 14880 3087
rect 14800 3019 14823 3053
rect 14857 3019 14880 3053
rect 14800 2985 14880 3019
rect 14800 2951 14823 2985
rect 14857 2951 14880 2985
rect 14800 2917 14880 2951
rect 14800 2883 14823 2917
rect 14857 2883 14880 2917
rect 14800 2849 14880 2883
rect 14800 2815 14823 2849
rect 14857 2815 14880 2849
rect 14800 2781 14880 2815
rect 14800 2747 14823 2781
rect 14857 2747 14880 2781
rect 14800 2713 14880 2747
rect 14800 2679 14823 2713
rect 14857 2679 14880 2713
rect 14800 2645 14880 2679
rect 14800 2611 14823 2645
rect 14857 2611 14880 2645
rect 14800 2577 14880 2611
rect 14800 2543 14823 2577
rect 14857 2543 14880 2577
rect 14800 2509 14880 2543
rect 14800 2475 14823 2509
rect 14857 2475 14880 2509
rect 14800 2441 14880 2475
rect 14800 2407 14823 2441
rect 14857 2407 14880 2441
rect 14800 2373 14880 2407
rect 14800 2339 14823 2373
rect 14857 2339 14880 2373
rect 14800 2305 14880 2339
rect 14800 2271 14823 2305
rect 14857 2271 14880 2305
rect 14800 2237 14880 2271
rect 14800 2203 14823 2237
rect 14857 2203 14880 2237
rect 14800 2169 14880 2203
rect 14800 2135 14823 2169
rect 14857 2135 14880 2169
rect 14800 2101 14880 2135
rect 14800 2067 14823 2101
rect 14857 2067 14880 2101
rect 14800 2033 14880 2067
rect 14800 1999 14823 2033
rect 14857 1999 14880 2033
rect 14800 1965 14880 1999
rect 14800 1931 14823 1965
rect 14857 1931 14880 1965
rect 14800 1897 14880 1931
rect 14800 1863 14823 1897
rect 14857 1863 14880 1897
rect 14800 1829 14880 1863
rect 14800 1795 14823 1829
rect 14857 1795 14880 1829
rect 14800 1761 14880 1795
rect 14800 1727 14823 1761
rect 14857 1727 14880 1761
rect 14800 1693 14880 1727
rect 14800 1659 14823 1693
rect 14857 1659 14880 1693
rect 14800 1625 14880 1659
rect 14800 1591 14823 1625
rect 14857 1591 14880 1625
rect 14800 1557 14880 1591
rect 14800 1523 14823 1557
rect 14857 1523 14880 1557
rect 14800 1440 14880 1523
rect -12880 1417 14880 1440
rect -12880 1383 -12719 1417
rect -12685 1383 -12651 1417
rect -12617 1383 -12583 1417
rect -12549 1383 -12515 1417
rect -12481 1383 -12447 1417
rect -12413 1383 -12379 1417
rect -12345 1383 -12311 1417
rect -12277 1383 -12243 1417
rect -12209 1383 -12175 1417
rect -12141 1383 -12107 1417
rect -12073 1383 -12039 1417
rect -12005 1383 -11971 1417
rect -11937 1383 -11903 1417
rect -11869 1383 -11835 1417
rect -11801 1383 -11767 1417
rect -11733 1383 -11699 1417
rect -11665 1383 -11631 1417
rect -11597 1383 -11563 1417
rect -11529 1383 -11495 1417
rect -11461 1383 -11427 1417
rect -11393 1383 -11359 1417
rect -11325 1383 -11291 1417
rect -11257 1383 -11223 1417
rect -11189 1383 -11155 1417
rect -11121 1383 -11087 1417
rect -11053 1383 -11019 1417
rect -10985 1383 -10951 1417
rect -10917 1383 -10883 1417
rect -10849 1383 -10815 1417
rect -10781 1383 -10747 1417
rect -10713 1383 -10679 1417
rect -10645 1383 -10611 1417
rect -10577 1383 -10543 1417
rect -10509 1383 -10475 1417
rect -10441 1383 -10407 1417
rect -10373 1383 -10339 1417
rect -10305 1383 -10271 1417
rect -10237 1383 -10203 1417
rect -10169 1383 -10135 1417
rect -10101 1383 -10067 1417
rect -10033 1383 -9999 1417
rect -9965 1383 -9931 1417
rect -9897 1383 -9863 1417
rect -9829 1383 -9795 1417
rect -9761 1383 -9727 1417
rect -9693 1383 -9659 1417
rect -9625 1383 -9591 1417
rect -9557 1383 -9523 1417
rect -9489 1383 -9455 1417
rect -9421 1383 -9387 1417
rect -9353 1383 -9319 1417
rect -9285 1383 -9251 1417
rect -9217 1383 -9183 1417
rect -9149 1383 -9115 1417
rect -9081 1383 -9047 1417
rect -9013 1383 -8979 1417
rect -8945 1383 -8911 1417
rect -8877 1383 -8843 1417
rect -8809 1383 -8775 1417
rect -8741 1383 -8707 1417
rect -8673 1383 -8639 1417
rect -8605 1383 -8571 1417
rect -8537 1383 -8503 1417
rect -8469 1383 -8435 1417
rect -8401 1383 -8367 1417
rect -8333 1383 -8299 1417
rect -8265 1383 -8231 1417
rect -8197 1383 -8163 1417
rect -8129 1383 -8095 1417
rect -8061 1383 -8027 1417
rect -7993 1383 -7959 1417
rect -7925 1383 -7891 1417
rect -7857 1383 -7823 1417
rect -7789 1383 -7755 1417
rect -7721 1383 -7687 1417
rect -7653 1383 -7619 1417
rect -7585 1383 -7551 1417
rect -7517 1383 -7483 1417
rect -7449 1383 -7415 1417
rect -7381 1383 -7347 1417
rect -7313 1383 -7279 1417
rect -7245 1383 -7211 1417
rect -7177 1383 -7143 1417
rect -7109 1383 -7075 1417
rect -7041 1383 -7007 1417
rect -6973 1383 -6939 1417
rect -6905 1383 -6871 1417
rect -6837 1383 -6803 1417
rect -6769 1383 -6735 1417
rect -6701 1383 -6667 1417
rect -6633 1383 -6599 1417
rect -6565 1383 -6531 1417
rect -6497 1383 -6463 1417
rect -6429 1383 -6395 1417
rect -6361 1383 -6327 1417
rect -6293 1383 -6259 1417
rect -6225 1383 -6191 1417
rect -6157 1383 -6123 1417
rect -6089 1383 -6055 1417
rect -6021 1383 -5987 1417
rect -5953 1383 -5919 1417
rect -5885 1383 -5851 1417
rect -5817 1383 -5783 1417
rect -5749 1383 -5715 1417
rect -5681 1383 -5647 1417
rect -5613 1383 -5579 1417
rect -5545 1383 -5511 1417
rect -5477 1383 -5443 1417
rect -5409 1383 -5375 1417
rect -5341 1383 -5307 1417
rect -5273 1383 -5239 1417
rect -5205 1383 -5171 1417
rect -5137 1383 -5103 1417
rect -5069 1383 -5035 1417
rect -5001 1383 -4967 1417
rect -4933 1383 -4899 1417
rect -4865 1383 -4831 1417
rect -4797 1383 -4763 1417
rect -4729 1383 -4695 1417
rect -4661 1383 -4627 1417
rect -4593 1383 -4559 1417
rect -4525 1383 -4491 1417
rect -4457 1383 -4423 1417
rect -4389 1383 -4355 1417
rect -4321 1383 -4287 1417
rect -4253 1383 -4219 1417
rect -4185 1383 -4151 1417
rect -4117 1383 -4083 1417
rect -4049 1383 -4015 1417
rect -3981 1383 -3947 1417
rect -3913 1383 -3879 1417
rect -3845 1383 -3811 1417
rect -3777 1383 -3743 1417
rect -3709 1383 -3675 1417
rect -3641 1383 -3607 1417
rect -3573 1383 -3539 1417
rect -3505 1383 -3471 1417
rect -3437 1383 -3403 1417
rect -3369 1383 -3335 1417
rect -3301 1383 -3267 1417
rect -3233 1383 -3199 1417
rect -3165 1383 -3131 1417
rect -3097 1383 -3063 1417
rect -3029 1383 -2995 1417
rect -2961 1383 -2927 1417
rect -2893 1383 -2859 1417
rect -2825 1383 -2791 1417
rect -2757 1383 -2723 1417
rect -2689 1383 -2655 1417
rect -2621 1383 -2587 1417
rect -2553 1383 -2519 1417
rect -2485 1383 -2451 1417
rect -2417 1383 -2383 1417
rect -2349 1383 -2315 1417
rect -2281 1383 -2247 1417
rect -2213 1383 -2179 1417
rect -2145 1383 -2111 1417
rect -2077 1383 -2043 1417
rect -2009 1383 -1975 1417
rect -1941 1383 -1907 1417
rect -1873 1383 -1839 1417
rect -1805 1383 -1771 1417
rect -1737 1383 -1703 1417
rect -1669 1383 -1635 1417
rect -1601 1383 -1567 1417
rect -1533 1383 -1499 1417
rect -1465 1383 -1431 1417
rect -1397 1383 -1363 1417
rect -1329 1383 -1295 1417
rect -1261 1383 -1227 1417
rect -1193 1383 -1159 1417
rect -1125 1383 -1091 1417
rect -1057 1383 -1023 1417
rect -989 1383 -955 1417
rect -921 1383 -887 1417
rect -853 1383 -819 1417
rect -785 1383 -751 1417
rect -717 1383 -683 1417
rect -649 1383 -615 1417
rect -581 1383 -547 1417
rect -513 1383 -479 1417
rect -445 1383 -411 1417
rect -377 1383 -343 1417
rect -309 1383 -275 1417
rect -241 1383 -207 1417
rect -173 1383 -139 1417
rect -105 1383 -71 1417
rect -37 1383 -3 1417
rect 31 1383 65 1417
rect 99 1383 133 1417
rect 167 1383 201 1417
rect 235 1383 269 1417
rect 303 1383 337 1417
rect 371 1383 405 1417
rect 439 1383 473 1417
rect 507 1383 541 1417
rect 575 1383 609 1417
rect 643 1383 677 1417
rect 711 1383 745 1417
rect 779 1383 813 1417
rect 847 1383 881 1417
rect 915 1383 949 1417
rect 983 1383 1017 1417
rect 1051 1383 1085 1417
rect 1119 1383 1153 1417
rect 1187 1383 1221 1417
rect 1255 1383 1289 1417
rect 1323 1383 1357 1417
rect 1391 1383 1425 1417
rect 1459 1383 1493 1417
rect 1527 1383 1561 1417
rect 1595 1383 1629 1417
rect 1663 1383 1697 1417
rect 1731 1383 1765 1417
rect 1799 1383 1833 1417
rect 1867 1383 1901 1417
rect 1935 1383 1969 1417
rect 2003 1383 2037 1417
rect 2071 1383 2105 1417
rect 2139 1383 2173 1417
rect 2207 1383 2241 1417
rect 2275 1383 2309 1417
rect 2343 1383 2377 1417
rect 2411 1383 2445 1417
rect 2479 1383 2513 1417
rect 2547 1383 2581 1417
rect 2615 1383 2649 1417
rect 2683 1383 2717 1417
rect 2751 1383 2785 1417
rect 2819 1383 2853 1417
rect 2887 1383 2921 1417
rect 2955 1383 2989 1417
rect 3023 1383 3057 1417
rect 3091 1383 3125 1417
rect 3159 1383 3193 1417
rect 3227 1383 3261 1417
rect 3295 1383 3329 1417
rect 3363 1383 3397 1417
rect 3431 1383 3465 1417
rect 3499 1383 3533 1417
rect 3567 1383 3601 1417
rect 3635 1383 3669 1417
rect 3703 1383 3737 1417
rect 3771 1383 3805 1417
rect 3839 1383 3873 1417
rect 3907 1383 3941 1417
rect 3975 1383 4009 1417
rect 4043 1383 4077 1417
rect 4111 1383 4145 1417
rect 4179 1383 4213 1417
rect 4247 1383 4281 1417
rect 4315 1383 4349 1417
rect 4383 1383 4417 1417
rect 4451 1383 4485 1417
rect 4519 1383 4553 1417
rect 4587 1383 4621 1417
rect 4655 1383 4689 1417
rect 4723 1383 4757 1417
rect 4791 1383 4825 1417
rect 4859 1383 4893 1417
rect 4927 1383 4961 1417
rect 4995 1383 5029 1417
rect 5063 1383 5097 1417
rect 5131 1383 5165 1417
rect 5199 1383 5233 1417
rect 5267 1383 5301 1417
rect 5335 1383 5369 1417
rect 5403 1383 5437 1417
rect 5471 1383 5505 1417
rect 5539 1383 5573 1417
rect 5607 1383 5641 1417
rect 5675 1383 5709 1417
rect 5743 1383 5777 1417
rect 5811 1383 5845 1417
rect 5879 1383 5913 1417
rect 5947 1383 5981 1417
rect 6015 1383 6049 1417
rect 6083 1383 6117 1417
rect 6151 1383 6185 1417
rect 6219 1383 6253 1417
rect 6287 1383 6321 1417
rect 6355 1383 6389 1417
rect 6423 1383 6457 1417
rect 6491 1383 6525 1417
rect 6559 1383 6593 1417
rect 6627 1383 6661 1417
rect 6695 1383 6729 1417
rect 6763 1383 6797 1417
rect 6831 1383 6865 1417
rect 6899 1383 6933 1417
rect 6967 1383 7001 1417
rect 7035 1383 7069 1417
rect 7103 1383 7137 1417
rect 7171 1383 7205 1417
rect 7239 1383 7273 1417
rect 7307 1383 7341 1417
rect 7375 1383 7409 1417
rect 7443 1383 7477 1417
rect 7511 1383 7545 1417
rect 7579 1383 7613 1417
rect 7647 1383 7681 1417
rect 7715 1383 7749 1417
rect 7783 1383 7817 1417
rect 7851 1383 7885 1417
rect 7919 1383 7953 1417
rect 7987 1383 8021 1417
rect 8055 1383 8089 1417
rect 8123 1383 8157 1417
rect 8191 1383 8225 1417
rect 8259 1383 8293 1417
rect 8327 1383 8361 1417
rect 8395 1383 8429 1417
rect 8463 1383 8497 1417
rect 8531 1383 8565 1417
rect 8599 1383 8633 1417
rect 8667 1383 8701 1417
rect 8735 1383 8769 1417
rect 8803 1383 8837 1417
rect 8871 1383 8905 1417
rect 8939 1383 8973 1417
rect 9007 1383 9041 1417
rect 9075 1383 9109 1417
rect 9143 1383 9177 1417
rect 9211 1383 9245 1417
rect 9279 1383 9313 1417
rect 9347 1383 9381 1417
rect 9415 1383 9449 1417
rect 9483 1383 9517 1417
rect 9551 1383 9585 1417
rect 9619 1383 9653 1417
rect 9687 1383 9721 1417
rect 9755 1383 9789 1417
rect 9823 1383 9857 1417
rect 9891 1383 9925 1417
rect 9959 1383 9993 1417
rect 10027 1383 10061 1417
rect 10095 1383 10129 1417
rect 10163 1383 10197 1417
rect 10231 1383 10265 1417
rect 10299 1383 10333 1417
rect 10367 1383 10401 1417
rect 10435 1383 10469 1417
rect 10503 1383 10537 1417
rect 10571 1383 10605 1417
rect 10639 1383 10673 1417
rect 10707 1383 10741 1417
rect 10775 1383 10809 1417
rect 10843 1383 10877 1417
rect 10911 1383 10945 1417
rect 10979 1383 11013 1417
rect 11047 1383 11081 1417
rect 11115 1383 11149 1417
rect 11183 1383 11217 1417
rect 11251 1383 11285 1417
rect 11319 1383 11353 1417
rect 11387 1383 11421 1417
rect 11455 1383 11489 1417
rect 11523 1383 11557 1417
rect 11591 1383 11625 1417
rect 11659 1383 11693 1417
rect 11727 1383 11761 1417
rect 11795 1383 11829 1417
rect 11863 1383 11897 1417
rect 11931 1383 11965 1417
rect 11999 1383 12033 1417
rect 12067 1383 12101 1417
rect 12135 1383 12169 1417
rect 12203 1383 12237 1417
rect 12271 1383 12305 1417
rect 12339 1383 12373 1417
rect 12407 1383 12441 1417
rect 12475 1383 12509 1417
rect 12543 1383 12577 1417
rect 12611 1383 12645 1417
rect 12679 1383 12713 1417
rect 12747 1383 12781 1417
rect 12815 1383 12849 1417
rect 12883 1383 12917 1417
rect 12951 1383 12985 1417
rect 13019 1383 13053 1417
rect 13087 1383 13121 1417
rect 13155 1383 13189 1417
rect 13223 1383 13257 1417
rect 13291 1383 13325 1417
rect 13359 1383 13393 1417
rect 13427 1383 13461 1417
rect 13495 1383 13529 1417
rect 13563 1383 13597 1417
rect 13631 1383 13665 1417
rect 13699 1383 13733 1417
rect 13767 1383 13801 1417
rect 13835 1383 13869 1417
rect 13903 1383 13937 1417
rect 13971 1383 14005 1417
rect 14039 1383 14073 1417
rect 14107 1383 14141 1417
rect 14175 1383 14209 1417
rect 14243 1383 14277 1417
rect 14311 1383 14345 1417
rect 14379 1383 14413 1417
rect 14447 1383 14481 1417
rect 14515 1383 14549 1417
rect 14583 1383 14617 1417
rect 14651 1383 14685 1417
rect 14719 1383 14880 1417
rect -12880 1360 14880 1383
<< psubdiffcont >>
rect -12719 7783 -12685 7817
rect -12651 7783 -12617 7817
rect -12583 7783 -12549 7817
rect -12515 7783 -12481 7817
rect -12447 7783 -12413 7817
rect -12379 7783 -12345 7817
rect -12311 7783 -12277 7817
rect -12243 7783 -12209 7817
rect -12175 7783 -12141 7817
rect -12107 7783 -12073 7817
rect -12039 7783 -12005 7817
rect -11971 7783 -11937 7817
rect -11903 7783 -11869 7817
rect -11835 7783 -11801 7817
rect -11767 7783 -11733 7817
rect -11699 7783 -11665 7817
rect -11631 7783 -11597 7817
rect -11563 7783 -11529 7817
rect -11495 7783 -11461 7817
rect -11427 7783 -11393 7817
rect -11359 7783 -11325 7817
rect -11291 7783 -11257 7817
rect -11223 7783 -11189 7817
rect -11155 7783 -11121 7817
rect -11087 7783 -11053 7817
rect -11019 7783 -10985 7817
rect -10951 7783 -10917 7817
rect -10883 7783 -10849 7817
rect -10815 7783 -10781 7817
rect -10747 7783 -10713 7817
rect -10679 7783 -10645 7817
rect -10611 7783 -10577 7817
rect -10543 7783 -10509 7817
rect -10475 7783 -10441 7817
rect -10407 7783 -10373 7817
rect -10339 7783 -10305 7817
rect -10271 7783 -10237 7817
rect -10203 7783 -10169 7817
rect -10135 7783 -10101 7817
rect -10067 7783 -10033 7817
rect -9999 7783 -9965 7817
rect -9931 7783 -9897 7817
rect -9863 7783 -9829 7817
rect -9795 7783 -9761 7817
rect -9727 7783 -9693 7817
rect -9659 7783 -9625 7817
rect -9591 7783 -9557 7817
rect -9523 7783 -9489 7817
rect -9455 7783 -9421 7817
rect -9387 7783 -9353 7817
rect -9319 7783 -9285 7817
rect -9251 7783 -9217 7817
rect -9183 7783 -9149 7817
rect -9115 7783 -9081 7817
rect -9047 7783 -9013 7817
rect -8979 7783 -8945 7817
rect -8911 7783 -8877 7817
rect -8843 7783 -8809 7817
rect -8775 7783 -8741 7817
rect -8707 7783 -8673 7817
rect -8639 7783 -8605 7817
rect -8571 7783 -8537 7817
rect -8503 7783 -8469 7817
rect -8435 7783 -8401 7817
rect -8367 7783 -8333 7817
rect -8299 7783 -8265 7817
rect -8231 7783 -8197 7817
rect -8163 7783 -8129 7817
rect -8095 7783 -8061 7817
rect -8027 7783 -7993 7817
rect -7959 7783 -7925 7817
rect -7891 7783 -7857 7817
rect -7823 7783 -7789 7817
rect -7755 7783 -7721 7817
rect -7687 7783 -7653 7817
rect -7619 7783 -7585 7817
rect -7551 7783 -7517 7817
rect -7483 7783 -7449 7817
rect -7415 7783 -7381 7817
rect -7347 7783 -7313 7817
rect -7279 7783 -7245 7817
rect -7211 7783 -7177 7817
rect -7143 7783 -7109 7817
rect -7075 7783 -7041 7817
rect -7007 7783 -6973 7817
rect -6939 7783 -6905 7817
rect -6871 7783 -6837 7817
rect -6803 7783 -6769 7817
rect -6735 7783 -6701 7817
rect -6667 7783 -6633 7817
rect -6599 7783 -6565 7817
rect -6531 7783 -6497 7817
rect -6463 7783 -6429 7817
rect -6395 7783 -6361 7817
rect -6327 7783 -6293 7817
rect -6259 7783 -6225 7817
rect -6191 7783 -6157 7817
rect -6123 7783 -6089 7817
rect -6055 7783 -6021 7817
rect -5987 7783 -5953 7817
rect -5919 7783 -5885 7817
rect -5851 7783 -5817 7817
rect -5783 7783 -5749 7817
rect -5715 7783 -5681 7817
rect -5647 7783 -5613 7817
rect -5579 7783 -5545 7817
rect -5511 7783 -5477 7817
rect -5443 7783 -5409 7817
rect -5375 7783 -5341 7817
rect -5307 7783 -5273 7817
rect -5239 7783 -5205 7817
rect -5171 7783 -5137 7817
rect -5103 7783 -5069 7817
rect -5035 7783 -5001 7817
rect -4967 7783 -4933 7817
rect -4899 7783 -4865 7817
rect -4831 7783 -4797 7817
rect -4763 7783 -4729 7817
rect -4695 7783 -4661 7817
rect -4627 7783 -4593 7817
rect -4559 7783 -4525 7817
rect -4491 7783 -4457 7817
rect -4423 7783 -4389 7817
rect -4355 7783 -4321 7817
rect -4287 7783 -4253 7817
rect -4219 7783 -4185 7817
rect -4151 7783 -4117 7817
rect -4083 7783 -4049 7817
rect -4015 7783 -3981 7817
rect -3947 7783 -3913 7817
rect -3879 7783 -3845 7817
rect -3811 7783 -3777 7817
rect -3743 7783 -3709 7817
rect -3675 7783 -3641 7817
rect -3607 7783 -3573 7817
rect -3539 7783 -3505 7817
rect -3471 7783 -3437 7817
rect -3403 7783 -3369 7817
rect -3335 7783 -3301 7817
rect -3267 7783 -3233 7817
rect -3199 7783 -3165 7817
rect -3131 7783 -3097 7817
rect -3063 7783 -3029 7817
rect -2995 7783 -2961 7817
rect -2927 7783 -2893 7817
rect -2859 7783 -2825 7817
rect -2791 7783 -2757 7817
rect -2723 7783 -2689 7817
rect -2655 7783 -2621 7817
rect -2587 7783 -2553 7817
rect -2519 7783 -2485 7817
rect -2451 7783 -2417 7817
rect -2383 7783 -2349 7817
rect -2315 7783 -2281 7817
rect -2247 7783 -2213 7817
rect -2179 7783 -2145 7817
rect -2111 7783 -2077 7817
rect -2043 7783 -2009 7817
rect -1975 7783 -1941 7817
rect -1907 7783 -1873 7817
rect -1839 7783 -1805 7817
rect -1771 7783 -1737 7817
rect -1703 7783 -1669 7817
rect -1635 7783 -1601 7817
rect -1567 7783 -1533 7817
rect -1499 7783 -1465 7817
rect -1431 7783 -1397 7817
rect -1363 7783 -1329 7817
rect -1295 7783 -1261 7817
rect -1227 7783 -1193 7817
rect -1159 7783 -1125 7817
rect -1091 7783 -1057 7817
rect -1023 7783 -989 7817
rect -955 7783 -921 7817
rect -887 7783 -853 7817
rect -819 7783 -785 7817
rect -751 7783 -717 7817
rect -683 7783 -649 7817
rect -615 7783 -581 7817
rect -547 7783 -513 7817
rect -479 7783 -445 7817
rect -411 7783 -377 7817
rect -343 7783 -309 7817
rect -275 7783 -241 7817
rect -207 7783 -173 7817
rect -139 7783 -105 7817
rect -71 7783 -37 7817
rect -3 7783 31 7817
rect 65 7783 99 7817
rect 133 7783 167 7817
rect 201 7783 235 7817
rect 269 7783 303 7817
rect 337 7783 371 7817
rect 405 7783 439 7817
rect 473 7783 507 7817
rect 541 7783 575 7817
rect 609 7783 643 7817
rect 677 7783 711 7817
rect 745 7783 779 7817
rect 813 7783 847 7817
rect 881 7783 915 7817
rect 949 7783 983 7817
rect 1017 7783 1051 7817
rect 1085 7783 1119 7817
rect 1153 7783 1187 7817
rect 1221 7783 1255 7817
rect 1289 7783 1323 7817
rect 1357 7783 1391 7817
rect 1425 7783 1459 7817
rect 1493 7783 1527 7817
rect 1561 7783 1595 7817
rect 1629 7783 1663 7817
rect 1697 7783 1731 7817
rect 1765 7783 1799 7817
rect 1833 7783 1867 7817
rect 1901 7783 1935 7817
rect 1969 7783 2003 7817
rect 2037 7783 2071 7817
rect 2105 7783 2139 7817
rect 2173 7783 2207 7817
rect 2241 7783 2275 7817
rect 2309 7783 2343 7817
rect 2377 7783 2411 7817
rect 2445 7783 2479 7817
rect 2513 7783 2547 7817
rect 2581 7783 2615 7817
rect 2649 7783 2683 7817
rect 2717 7783 2751 7817
rect 2785 7783 2819 7817
rect 2853 7783 2887 7817
rect 2921 7783 2955 7817
rect 2989 7783 3023 7817
rect 3057 7783 3091 7817
rect 3125 7783 3159 7817
rect 3193 7783 3227 7817
rect 3261 7783 3295 7817
rect 3329 7783 3363 7817
rect 3397 7783 3431 7817
rect 3465 7783 3499 7817
rect 3533 7783 3567 7817
rect 3601 7783 3635 7817
rect 3669 7783 3703 7817
rect 3737 7783 3771 7817
rect 3805 7783 3839 7817
rect 3873 7783 3907 7817
rect 3941 7783 3975 7817
rect 4009 7783 4043 7817
rect 4077 7783 4111 7817
rect 4145 7783 4179 7817
rect 4213 7783 4247 7817
rect 4281 7783 4315 7817
rect 4349 7783 4383 7817
rect 4417 7783 4451 7817
rect 4485 7783 4519 7817
rect 4553 7783 4587 7817
rect 4621 7783 4655 7817
rect 4689 7783 4723 7817
rect 4757 7783 4791 7817
rect 4825 7783 4859 7817
rect 4893 7783 4927 7817
rect 4961 7783 4995 7817
rect 5029 7783 5063 7817
rect 5097 7783 5131 7817
rect 5165 7783 5199 7817
rect 5233 7783 5267 7817
rect 5301 7783 5335 7817
rect 5369 7783 5403 7817
rect 5437 7783 5471 7817
rect 5505 7783 5539 7817
rect 5573 7783 5607 7817
rect 5641 7783 5675 7817
rect 5709 7783 5743 7817
rect 5777 7783 5811 7817
rect 5845 7783 5879 7817
rect 5913 7783 5947 7817
rect 5981 7783 6015 7817
rect 6049 7783 6083 7817
rect 6117 7783 6151 7817
rect 6185 7783 6219 7817
rect 6253 7783 6287 7817
rect 6321 7783 6355 7817
rect 6389 7783 6423 7817
rect 6457 7783 6491 7817
rect 6525 7783 6559 7817
rect 6593 7783 6627 7817
rect 6661 7783 6695 7817
rect 6729 7783 6763 7817
rect 6797 7783 6831 7817
rect 6865 7783 6899 7817
rect 6933 7783 6967 7817
rect 7001 7783 7035 7817
rect 7069 7783 7103 7817
rect 7137 7783 7171 7817
rect 7205 7783 7239 7817
rect 7273 7783 7307 7817
rect 7341 7783 7375 7817
rect 7409 7783 7443 7817
rect 7477 7783 7511 7817
rect 7545 7783 7579 7817
rect 7613 7783 7647 7817
rect 7681 7783 7715 7817
rect 7749 7783 7783 7817
rect 7817 7783 7851 7817
rect 7885 7783 7919 7817
rect 7953 7783 7987 7817
rect 8021 7783 8055 7817
rect 8089 7783 8123 7817
rect 8157 7783 8191 7817
rect 8225 7783 8259 7817
rect 8293 7783 8327 7817
rect 8361 7783 8395 7817
rect 8429 7783 8463 7817
rect 8497 7783 8531 7817
rect 8565 7783 8599 7817
rect 8633 7783 8667 7817
rect 8701 7783 8735 7817
rect 8769 7783 8803 7817
rect 8837 7783 8871 7817
rect 8905 7783 8939 7817
rect 8973 7783 9007 7817
rect 9041 7783 9075 7817
rect 9109 7783 9143 7817
rect 9177 7783 9211 7817
rect 9245 7783 9279 7817
rect 9313 7783 9347 7817
rect 9381 7783 9415 7817
rect 9449 7783 9483 7817
rect 9517 7783 9551 7817
rect 9585 7783 9619 7817
rect 9653 7783 9687 7817
rect 9721 7783 9755 7817
rect 9789 7783 9823 7817
rect 9857 7783 9891 7817
rect 9925 7783 9959 7817
rect 9993 7783 10027 7817
rect 10061 7783 10095 7817
rect 10129 7783 10163 7817
rect 10197 7783 10231 7817
rect 10265 7783 10299 7817
rect 10333 7783 10367 7817
rect 10401 7783 10435 7817
rect 10469 7783 10503 7817
rect 10537 7783 10571 7817
rect 10605 7783 10639 7817
rect 10673 7783 10707 7817
rect 10741 7783 10775 7817
rect 10809 7783 10843 7817
rect 10877 7783 10911 7817
rect 10945 7783 10979 7817
rect 11013 7783 11047 7817
rect 11081 7783 11115 7817
rect 11149 7783 11183 7817
rect 11217 7783 11251 7817
rect 11285 7783 11319 7817
rect 11353 7783 11387 7817
rect 11421 7783 11455 7817
rect 11489 7783 11523 7817
rect 11557 7783 11591 7817
rect 11625 7783 11659 7817
rect 11693 7783 11727 7817
rect 11761 7783 11795 7817
rect 11829 7783 11863 7817
rect 11897 7783 11931 7817
rect 11965 7783 11999 7817
rect 12033 7783 12067 7817
rect 12101 7783 12135 7817
rect 12169 7783 12203 7817
rect 12237 7783 12271 7817
rect 12305 7783 12339 7817
rect 12373 7783 12407 7817
rect 12441 7783 12475 7817
rect 12509 7783 12543 7817
rect 12577 7783 12611 7817
rect 12645 7783 12679 7817
rect 12713 7783 12747 7817
rect 12781 7783 12815 7817
rect 12849 7783 12883 7817
rect 12917 7783 12951 7817
rect 12985 7783 13019 7817
rect 13053 7783 13087 7817
rect 13121 7783 13155 7817
rect 13189 7783 13223 7817
rect 13257 7783 13291 7817
rect 13325 7783 13359 7817
rect 13393 7783 13427 7817
rect 13461 7783 13495 7817
rect 13529 7783 13563 7817
rect 13597 7783 13631 7817
rect 13665 7783 13699 7817
rect 13733 7783 13767 7817
rect 13801 7783 13835 7817
rect 13869 7783 13903 7817
rect 13937 7783 13971 7817
rect 14005 7783 14039 7817
rect 14073 7783 14107 7817
rect 14141 7783 14175 7817
rect 14209 7783 14243 7817
rect 14277 7783 14311 7817
rect 14345 7783 14379 7817
rect 14413 7783 14447 7817
rect 14481 7783 14515 7817
rect 14549 7783 14583 7817
rect 14617 7783 14651 7817
rect 14685 7783 14719 7817
rect -12857 7643 -12823 7677
rect -12857 7575 -12823 7609
rect -12857 7507 -12823 7541
rect -12857 7439 -12823 7473
rect -12857 7371 -12823 7405
rect -12857 7303 -12823 7337
rect -12857 7235 -12823 7269
rect -12857 7167 -12823 7201
rect -12857 7099 -12823 7133
rect -12857 7031 -12823 7065
rect -12857 6963 -12823 6997
rect -12857 6895 -12823 6929
rect -12857 6827 -12823 6861
rect -12857 6759 -12823 6793
rect -12857 6691 -12823 6725
rect -12857 6623 -12823 6657
rect -12857 6555 -12823 6589
rect -12857 6487 -12823 6521
rect -12857 6419 -12823 6453
rect -12857 6351 -12823 6385
rect -12857 6283 -12823 6317
rect -12857 6215 -12823 6249
rect -12857 6147 -12823 6181
rect -12857 6079 -12823 6113
rect -12857 6011 -12823 6045
rect -12857 5943 -12823 5977
rect -12857 5875 -12823 5909
rect -12857 5807 -12823 5841
rect -12857 5739 -12823 5773
rect -12857 5671 -12823 5705
rect -12857 5603 -12823 5637
rect -12857 5535 -12823 5569
rect -12857 5467 -12823 5501
rect -12857 5399 -12823 5433
rect -12857 5331 -12823 5365
rect -12857 5263 -12823 5297
rect -12857 5195 -12823 5229
rect -12857 5127 -12823 5161
rect -12857 5059 -12823 5093
rect -12857 4991 -12823 5025
rect -12857 4923 -12823 4957
rect -12857 4855 -12823 4889
rect -12857 4787 -12823 4821
rect -12857 4719 -12823 4753
rect -12857 4651 -12823 4685
rect -12857 4583 -12823 4617
rect -12857 4515 -12823 4549
rect -12857 4447 -12823 4481
rect -12857 4379 -12823 4413
rect -12857 4311 -12823 4345
rect -12857 4243 -12823 4277
rect -12857 4175 -12823 4209
rect -12857 4107 -12823 4141
rect -12857 4039 -12823 4073
rect -12857 3971 -12823 4005
rect -12857 3903 -12823 3937
rect -12857 3835 -12823 3869
rect -12857 3767 -12823 3801
rect -12857 3699 -12823 3733
rect -12857 3631 -12823 3665
rect -12857 3563 -12823 3597
rect -12857 3495 -12823 3529
rect -12857 3427 -12823 3461
rect -12857 3359 -12823 3393
rect -12857 3291 -12823 3325
rect -12857 3223 -12823 3257
rect -12857 3155 -12823 3189
rect -12857 3087 -12823 3121
rect -12857 3019 -12823 3053
rect -12857 2951 -12823 2985
rect -12857 2883 -12823 2917
rect -12857 2815 -12823 2849
rect -12857 2747 -12823 2781
rect -12857 2679 -12823 2713
rect -12857 2611 -12823 2645
rect -12857 2543 -12823 2577
rect -12857 2475 -12823 2509
rect -12857 2407 -12823 2441
rect -12857 2339 -12823 2373
rect -12857 2271 -12823 2305
rect -12857 2203 -12823 2237
rect -12857 2135 -12823 2169
rect -12857 2067 -12823 2101
rect -12857 1999 -12823 2033
rect -12857 1931 -12823 1965
rect -12857 1863 -12823 1897
rect -12857 1795 -12823 1829
rect -12857 1727 -12823 1761
rect -12857 1659 -12823 1693
rect -12857 1591 -12823 1625
rect -12857 1523 -12823 1557
rect 14823 7643 14857 7677
rect 14823 7575 14857 7609
rect 14823 7507 14857 7541
rect 14823 7439 14857 7473
rect 14823 7371 14857 7405
rect 14823 7303 14857 7337
rect 14823 7235 14857 7269
rect 14823 7167 14857 7201
rect 14823 7099 14857 7133
rect 14823 7031 14857 7065
rect 14823 6963 14857 6997
rect 14823 6895 14857 6929
rect 14823 6827 14857 6861
rect 14823 6759 14857 6793
rect 14823 6691 14857 6725
rect 14823 6623 14857 6657
rect 14823 6555 14857 6589
rect 14823 6487 14857 6521
rect 14823 6419 14857 6453
rect 14823 6351 14857 6385
rect 14823 6283 14857 6317
rect 14823 6215 14857 6249
rect 14823 6147 14857 6181
rect 14823 6079 14857 6113
rect 14823 6011 14857 6045
rect 14823 5943 14857 5977
rect 14823 5875 14857 5909
rect 14823 5807 14857 5841
rect 14823 5739 14857 5773
rect 14823 5671 14857 5705
rect 14823 5603 14857 5637
rect 14823 5535 14857 5569
rect 14823 5467 14857 5501
rect 14823 5399 14857 5433
rect 14823 5331 14857 5365
rect 14823 5263 14857 5297
rect 14823 5195 14857 5229
rect 14823 5127 14857 5161
rect 14823 5059 14857 5093
rect 14823 4991 14857 5025
rect 14823 4923 14857 4957
rect 14823 4855 14857 4889
rect 14823 4787 14857 4821
rect 14823 4719 14857 4753
rect 14823 4651 14857 4685
rect 14823 4583 14857 4617
rect 14823 4515 14857 4549
rect 14823 4447 14857 4481
rect 14823 4379 14857 4413
rect 14823 4311 14857 4345
rect 14823 4243 14857 4277
rect 14823 4175 14857 4209
rect 14823 4107 14857 4141
rect 14823 4039 14857 4073
rect 14823 3971 14857 4005
rect 14823 3903 14857 3937
rect 14823 3835 14857 3869
rect 14823 3767 14857 3801
rect 14823 3699 14857 3733
rect 14823 3631 14857 3665
rect 14823 3563 14857 3597
rect 14823 3495 14857 3529
rect 14823 3427 14857 3461
rect 14823 3359 14857 3393
rect 14823 3291 14857 3325
rect 14823 3223 14857 3257
rect 14823 3155 14857 3189
rect 14823 3087 14857 3121
rect 14823 3019 14857 3053
rect 14823 2951 14857 2985
rect 14823 2883 14857 2917
rect 14823 2815 14857 2849
rect 14823 2747 14857 2781
rect 14823 2679 14857 2713
rect 14823 2611 14857 2645
rect 14823 2543 14857 2577
rect 14823 2475 14857 2509
rect 14823 2407 14857 2441
rect 14823 2339 14857 2373
rect 14823 2271 14857 2305
rect 14823 2203 14857 2237
rect 14823 2135 14857 2169
rect 14823 2067 14857 2101
rect 14823 1999 14857 2033
rect 14823 1931 14857 1965
rect 14823 1863 14857 1897
rect 14823 1795 14857 1829
rect 14823 1727 14857 1761
rect 14823 1659 14857 1693
rect 14823 1591 14857 1625
rect 14823 1523 14857 1557
rect -12719 1383 -12685 1417
rect -12651 1383 -12617 1417
rect -12583 1383 -12549 1417
rect -12515 1383 -12481 1417
rect -12447 1383 -12413 1417
rect -12379 1383 -12345 1417
rect -12311 1383 -12277 1417
rect -12243 1383 -12209 1417
rect -12175 1383 -12141 1417
rect -12107 1383 -12073 1417
rect -12039 1383 -12005 1417
rect -11971 1383 -11937 1417
rect -11903 1383 -11869 1417
rect -11835 1383 -11801 1417
rect -11767 1383 -11733 1417
rect -11699 1383 -11665 1417
rect -11631 1383 -11597 1417
rect -11563 1383 -11529 1417
rect -11495 1383 -11461 1417
rect -11427 1383 -11393 1417
rect -11359 1383 -11325 1417
rect -11291 1383 -11257 1417
rect -11223 1383 -11189 1417
rect -11155 1383 -11121 1417
rect -11087 1383 -11053 1417
rect -11019 1383 -10985 1417
rect -10951 1383 -10917 1417
rect -10883 1383 -10849 1417
rect -10815 1383 -10781 1417
rect -10747 1383 -10713 1417
rect -10679 1383 -10645 1417
rect -10611 1383 -10577 1417
rect -10543 1383 -10509 1417
rect -10475 1383 -10441 1417
rect -10407 1383 -10373 1417
rect -10339 1383 -10305 1417
rect -10271 1383 -10237 1417
rect -10203 1383 -10169 1417
rect -10135 1383 -10101 1417
rect -10067 1383 -10033 1417
rect -9999 1383 -9965 1417
rect -9931 1383 -9897 1417
rect -9863 1383 -9829 1417
rect -9795 1383 -9761 1417
rect -9727 1383 -9693 1417
rect -9659 1383 -9625 1417
rect -9591 1383 -9557 1417
rect -9523 1383 -9489 1417
rect -9455 1383 -9421 1417
rect -9387 1383 -9353 1417
rect -9319 1383 -9285 1417
rect -9251 1383 -9217 1417
rect -9183 1383 -9149 1417
rect -9115 1383 -9081 1417
rect -9047 1383 -9013 1417
rect -8979 1383 -8945 1417
rect -8911 1383 -8877 1417
rect -8843 1383 -8809 1417
rect -8775 1383 -8741 1417
rect -8707 1383 -8673 1417
rect -8639 1383 -8605 1417
rect -8571 1383 -8537 1417
rect -8503 1383 -8469 1417
rect -8435 1383 -8401 1417
rect -8367 1383 -8333 1417
rect -8299 1383 -8265 1417
rect -8231 1383 -8197 1417
rect -8163 1383 -8129 1417
rect -8095 1383 -8061 1417
rect -8027 1383 -7993 1417
rect -7959 1383 -7925 1417
rect -7891 1383 -7857 1417
rect -7823 1383 -7789 1417
rect -7755 1383 -7721 1417
rect -7687 1383 -7653 1417
rect -7619 1383 -7585 1417
rect -7551 1383 -7517 1417
rect -7483 1383 -7449 1417
rect -7415 1383 -7381 1417
rect -7347 1383 -7313 1417
rect -7279 1383 -7245 1417
rect -7211 1383 -7177 1417
rect -7143 1383 -7109 1417
rect -7075 1383 -7041 1417
rect -7007 1383 -6973 1417
rect -6939 1383 -6905 1417
rect -6871 1383 -6837 1417
rect -6803 1383 -6769 1417
rect -6735 1383 -6701 1417
rect -6667 1383 -6633 1417
rect -6599 1383 -6565 1417
rect -6531 1383 -6497 1417
rect -6463 1383 -6429 1417
rect -6395 1383 -6361 1417
rect -6327 1383 -6293 1417
rect -6259 1383 -6225 1417
rect -6191 1383 -6157 1417
rect -6123 1383 -6089 1417
rect -6055 1383 -6021 1417
rect -5987 1383 -5953 1417
rect -5919 1383 -5885 1417
rect -5851 1383 -5817 1417
rect -5783 1383 -5749 1417
rect -5715 1383 -5681 1417
rect -5647 1383 -5613 1417
rect -5579 1383 -5545 1417
rect -5511 1383 -5477 1417
rect -5443 1383 -5409 1417
rect -5375 1383 -5341 1417
rect -5307 1383 -5273 1417
rect -5239 1383 -5205 1417
rect -5171 1383 -5137 1417
rect -5103 1383 -5069 1417
rect -5035 1383 -5001 1417
rect -4967 1383 -4933 1417
rect -4899 1383 -4865 1417
rect -4831 1383 -4797 1417
rect -4763 1383 -4729 1417
rect -4695 1383 -4661 1417
rect -4627 1383 -4593 1417
rect -4559 1383 -4525 1417
rect -4491 1383 -4457 1417
rect -4423 1383 -4389 1417
rect -4355 1383 -4321 1417
rect -4287 1383 -4253 1417
rect -4219 1383 -4185 1417
rect -4151 1383 -4117 1417
rect -4083 1383 -4049 1417
rect -4015 1383 -3981 1417
rect -3947 1383 -3913 1417
rect -3879 1383 -3845 1417
rect -3811 1383 -3777 1417
rect -3743 1383 -3709 1417
rect -3675 1383 -3641 1417
rect -3607 1383 -3573 1417
rect -3539 1383 -3505 1417
rect -3471 1383 -3437 1417
rect -3403 1383 -3369 1417
rect -3335 1383 -3301 1417
rect -3267 1383 -3233 1417
rect -3199 1383 -3165 1417
rect -3131 1383 -3097 1417
rect -3063 1383 -3029 1417
rect -2995 1383 -2961 1417
rect -2927 1383 -2893 1417
rect -2859 1383 -2825 1417
rect -2791 1383 -2757 1417
rect -2723 1383 -2689 1417
rect -2655 1383 -2621 1417
rect -2587 1383 -2553 1417
rect -2519 1383 -2485 1417
rect -2451 1383 -2417 1417
rect -2383 1383 -2349 1417
rect -2315 1383 -2281 1417
rect -2247 1383 -2213 1417
rect -2179 1383 -2145 1417
rect -2111 1383 -2077 1417
rect -2043 1383 -2009 1417
rect -1975 1383 -1941 1417
rect -1907 1383 -1873 1417
rect -1839 1383 -1805 1417
rect -1771 1383 -1737 1417
rect -1703 1383 -1669 1417
rect -1635 1383 -1601 1417
rect -1567 1383 -1533 1417
rect -1499 1383 -1465 1417
rect -1431 1383 -1397 1417
rect -1363 1383 -1329 1417
rect -1295 1383 -1261 1417
rect -1227 1383 -1193 1417
rect -1159 1383 -1125 1417
rect -1091 1383 -1057 1417
rect -1023 1383 -989 1417
rect -955 1383 -921 1417
rect -887 1383 -853 1417
rect -819 1383 -785 1417
rect -751 1383 -717 1417
rect -683 1383 -649 1417
rect -615 1383 -581 1417
rect -547 1383 -513 1417
rect -479 1383 -445 1417
rect -411 1383 -377 1417
rect -343 1383 -309 1417
rect -275 1383 -241 1417
rect -207 1383 -173 1417
rect -139 1383 -105 1417
rect -71 1383 -37 1417
rect -3 1383 31 1417
rect 65 1383 99 1417
rect 133 1383 167 1417
rect 201 1383 235 1417
rect 269 1383 303 1417
rect 337 1383 371 1417
rect 405 1383 439 1417
rect 473 1383 507 1417
rect 541 1383 575 1417
rect 609 1383 643 1417
rect 677 1383 711 1417
rect 745 1383 779 1417
rect 813 1383 847 1417
rect 881 1383 915 1417
rect 949 1383 983 1417
rect 1017 1383 1051 1417
rect 1085 1383 1119 1417
rect 1153 1383 1187 1417
rect 1221 1383 1255 1417
rect 1289 1383 1323 1417
rect 1357 1383 1391 1417
rect 1425 1383 1459 1417
rect 1493 1383 1527 1417
rect 1561 1383 1595 1417
rect 1629 1383 1663 1417
rect 1697 1383 1731 1417
rect 1765 1383 1799 1417
rect 1833 1383 1867 1417
rect 1901 1383 1935 1417
rect 1969 1383 2003 1417
rect 2037 1383 2071 1417
rect 2105 1383 2139 1417
rect 2173 1383 2207 1417
rect 2241 1383 2275 1417
rect 2309 1383 2343 1417
rect 2377 1383 2411 1417
rect 2445 1383 2479 1417
rect 2513 1383 2547 1417
rect 2581 1383 2615 1417
rect 2649 1383 2683 1417
rect 2717 1383 2751 1417
rect 2785 1383 2819 1417
rect 2853 1383 2887 1417
rect 2921 1383 2955 1417
rect 2989 1383 3023 1417
rect 3057 1383 3091 1417
rect 3125 1383 3159 1417
rect 3193 1383 3227 1417
rect 3261 1383 3295 1417
rect 3329 1383 3363 1417
rect 3397 1383 3431 1417
rect 3465 1383 3499 1417
rect 3533 1383 3567 1417
rect 3601 1383 3635 1417
rect 3669 1383 3703 1417
rect 3737 1383 3771 1417
rect 3805 1383 3839 1417
rect 3873 1383 3907 1417
rect 3941 1383 3975 1417
rect 4009 1383 4043 1417
rect 4077 1383 4111 1417
rect 4145 1383 4179 1417
rect 4213 1383 4247 1417
rect 4281 1383 4315 1417
rect 4349 1383 4383 1417
rect 4417 1383 4451 1417
rect 4485 1383 4519 1417
rect 4553 1383 4587 1417
rect 4621 1383 4655 1417
rect 4689 1383 4723 1417
rect 4757 1383 4791 1417
rect 4825 1383 4859 1417
rect 4893 1383 4927 1417
rect 4961 1383 4995 1417
rect 5029 1383 5063 1417
rect 5097 1383 5131 1417
rect 5165 1383 5199 1417
rect 5233 1383 5267 1417
rect 5301 1383 5335 1417
rect 5369 1383 5403 1417
rect 5437 1383 5471 1417
rect 5505 1383 5539 1417
rect 5573 1383 5607 1417
rect 5641 1383 5675 1417
rect 5709 1383 5743 1417
rect 5777 1383 5811 1417
rect 5845 1383 5879 1417
rect 5913 1383 5947 1417
rect 5981 1383 6015 1417
rect 6049 1383 6083 1417
rect 6117 1383 6151 1417
rect 6185 1383 6219 1417
rect 6253 1383 6287 1417
rect 6321 1383 6355 1417
rect 6389 1383 6423 1417
rect 6457 1383 6491 1417
rect 6525 1383 6559 1417
rect 6593 1383 6627 1417
rect 6661 1383 6695 1417
rect 6729 1383 6763 1417
rect 6797 1383 6831 1417
rect 6865 1383 6899 1417
rect 6933 1383 6967 1417
rect 7001 1383 7035 1417
rect 7069 1383 7103 1417
rect 7137 1383 7171 1417
rect 7205 1383 7239 1417
rect 7273 1383 7307 1417
rect 7341 1383 7375 1417
rect 7409 1383 7443 1417
rect 7477 1383 7511 1417
rect 7545 1383 7579 1417
rect 7613 1383 7647 1417
rect 7681 1383 7715 1417
rect 7749 1383 7783 1417
rect 7817 1383 7851 1417
rect 7885 1383 7919 1417
rect 7953 1383 7987 1417
rect 8021 1383 8055 1417
rect 8089 1383 8123 1417
rect 8157 1383 8191 1417
rect 8225 1383 8259 1417
rect 8293 1383 8327 1417
rect 8361 1383 8395 1417
rect 8429 1383 8463 1417
rect 8497 1383 8531 1417
rect 8565 1383 8599 1417
rect 8633 1383 8667 1417
rect 8701 1383 8735 1417
rect 8769 1383 8803 1417
rect 8837 1383 8871 1417
rect 8905 1383 8939 1417
rect 8973 1383 9007 1417
rect 9041 1383 9075 1417
rect 9109 1383 9143 1417
rect 9177 1383 9211 1417
rect 9245 1383 9279 1417
rect 9313 1383 9347 1417
rect 9381 1383 9415 1417
rect 9449 1383 9483 1417
rect 9517 1383 9551 1417
rect 9585 1383 9619 1417
rect 9653 1383 9687 1417
rect 9721 1383 9755 1417
rect 9789 1383 9823 1417
rect 9857 1383 9891 1417
rect 9925 1383 9959 1417
rect 9993 1383 10027 1417
rect 10061 1383 10095 1417
rect 10129 1383 10163 1417
rect 10197 1383 10231 1417
rect 10265 1383 10299 1417
rect 10333 1383 10367 1417
rect 10401 1383 10435 1417
rect 10469 1383 10503 1417
rect 10537 1383 10571 1417
rect 10605 1383 10639 1417
rect 10673 1383 10707 1417
rect 10741 1383 10775 1417
rect 10809 1383 10843 1417
rect 10877 1383 10911 1417
rect 10945 1383 10979 1417
rect 11013 1383 11047 1417
rect 11081 1383 11115 1417
rect 11149 1383 11183 1417
rect 11217 1383 11251 1417
rect 11285 1383 11319 1417
rect 11353 1383 11387 1417
rect 11421 1383 11455 1417
rect 11489 1383 11523 1417
rect 11557 1383 11591 1417
rect 11625 1383 11659 1417
rect 11693 1383 11727 1417
rect 11761 1383 11795 1417
rect 11829 1383 11863 1417
rect 11897 1383 11931 1417
rect 11965 1383 11999 1417
rect 12033 1383 12067 1417
rect 12101 1383 12135 1417
rect 12169 1383 12203 1417
rect 12237 1383 12271 1417
rect 12305 1383 12339 1417
rect 12373 1383 12407 1417
rect 12441 1383 12475 1417
rect 12509 1383 12543 1417
rect 12577 1383 12611 1417
rect 12645 1383 12679 1417
rect 12713 1383 12747 1417
rect 12781 1383 12815 1417
rect 12849 1383 12883 1417
rect 12917 1383 12951 1417
rect 12985 1383 13019 1417
rect 13053 1383 13087 1417
rect 13121 1383 13155 1417
rect 13189 1383 13223 1417
rect 13257 1383 13291 1417
rect 13325 1383 13359 1417
rect 13393 1383 13427 1417
rect 13461 1383 13495 1417
rect 13529 1383 13563 1417
rect 13597 1383 13631 1417
rect 13665 1383 13699 1417
rect 13733 1383 13767 1417
rect 13801 1383 13835 1417
rect 13869 1383 13903 1417
rect 13937 1383 13971 1417
rect 14005 1383 14039 1417
rect 14073 1383 14107 1417
rect 14141 1383 14175 1417
rect 14209 1383 14243 1417
rect 14277 1383 14311 1417
rect 14345 1383 14379 1417
rect 14413 1383 14447 1417
rect 14481 1383 14515 1417
rect 14549 1383 14583 1417
rect 14617 1383 14651 1417
rect 14685 1383 14719 1417
<< locali >>
rect -12880 7817 14880 7840
rect -12880 7783 -12719 7817
rect -12685 7783 -12651 7817
rect -12617 7783 -12583 7817
rect -12549 7783 -12515 7817
rect -12481 7783 -12447 7817
rect -12413 7783 -12379 7817
rect -12345 7783 -12311 7817
rect -12277 7783 -12243 7817
rect -12209 7783 -12175 7817
rect -12141 7783 -12107 7817
rect -12073 7783 -12039 7817
rect -12005 7783 -11971 7817
rect -11937 7783 -11903 7817
rect -11869 7783 -11835 7817
rect -11801 7783 -11767 7817
rect -11733 7783 -11699 7817
rect -11665 7783 -11631 7817
rect -11597 7783 -11563 7817
rect -11529 7783 -11495 7817
rect -11461 7783 -11427 7817
rect -11393 7783 -11359 7817
rect -11325 7783 -11291 7817
rect -11257 7783 -11223 7817
rect -11189 7783 -11155 7817
rect -11121 7783 -11087 7817
rect -11053 7783 -11019 7817
rect -10985 7783 -10951 7817
rect -10917 7783 -10883 7817
rect -10849 7783 -10815 7817
rect -10781 7783 -10747 7817
rect -10713 7783 -10679 7817
rect -10645 7783 -10611 7817
rect -10577 7783 -10543 7817
rect -10509 7783 -10475 7817
rect -10441 7783 -10407 7817
rect -10373 7783 -10339 7817
rect -10305 7783 -10271 7817
rect -10237 7783 -10203 7817
rect -10169 7783 -10135 7817
rect -10101 7783 -10067 7817
rect -10033 7783 -9999 7817
rect -9965 7783 -9931 7817
rect -9897 7783 -9863 7817
rect -9829 7783 -9795 7817
rect -9761 7783 -9727 7817
rect -9693 7783 -9659 7817
rect -9625 7783 -9591 7817
rect -9557 7783 -9523 7817
rect -9489 7783 -9455 7817
rect -9421 7783 -9387 7817
rect -9353 7783 -9319 7817
rect -9285 7783 -9251 7817
rect -9217 7783 -9183 7817
rect -9149 7783 -9115 7817
rect -9081 7783 -9047 7817
rect -9013 7783 -8979 7817
rect -8945 7783 -8911 7817
rect -8877 7783 -8843 7817
rect -8809 7783 -8775 7817
rect -8741 7783 -8707 7817
rect -8673 7783 -8639 7817
rect -8605 7783 -8571 7817
rect -8537 7783 -8503 7817
rect -8469 7783 -8435 7817
rect -8401 7783 -8367 7817
rect -8333 7783 -8299 7817
rect -8265 7783 -8231 7817
rect -8197 7783 -8163 7817
rect -8129 7783 -8095 7817
rect -8061 7783 -8027 7817
rect -7993 7783 -7959 7817
rect -7925 7783 -7891 7817
rect -7857 7783 -7823 7817
rect -7789 7783 -7755 7817
rect -7721 7783 -7687 7817
rect -7653 7783 -7619 7817
rect -7585 7783 -7551 7817
rect -7517 7783 -7483 7817
rect -7449 7783 -7415 7817
rect -7381 7783 -7347 7817
rect -7313 7783 -7279 7817
rect -7245 7783 -7211 7817
rect -7177 7783 -7143 7817
rect -7109 7783 -7075 7817
rect -7041 7783 -7007 7817
rect -6973 7783 -6939 7817
rect -6905 7783 -6871 7817
rect -6837 7783 -6803 7817
rect -6769 7783 -6735 7817
rect -6701 7783 -6667 7817
rect -6633 7783 -6599 7817
rect -6565 7783 -6531 7817
rect -6497 7783 -6463 7817
rect -6429 7783 -6395 7817
rect -6361 7783 -6327 7817
rect -6293 7783 -6259 7817
rect -6225 7783 -6191 7817
rect -6157 7783 -6123 7817
rect -6089 7783 -6055 7817
rect -6021 7783 -5987 7817
rect -5953 7783 -5919 7817
rect -5885 7783 -5851 7817
rect -5817 7783 -5783 7817
rect -5749 7783 -5715 7817
rect -5681 7783 -5647 7817
rect -5613 7783 -5579 7817
rect -5545 7783 -5511 7817
rect -5477 7783 -5443 7817
rect -5409 7783 -5375 7817
rect -5341 7783 -5307 7817
rect -5273 7783 -5239 7817
rect -5205 7783 -5171 7817
rect -5137 7783 -5103 7817
rect -5069 7783 -5035 7817
rect -5001 7783 -4967 7817
rect -4933 7783 -4899 7817
rect -4865 7783 -4831 7817
rect -4797 7783 -4763 7817
rect -4729 7783 -4695 7817
rect -4661 7783 -4627 7817
rect -4593 7783 -4559 7817
rect -4525 7783 -4491 7817
rect -4457 7783 -4423 7817
rect -4389 7783 -4355 7817
rect -4321 7783 -4287 7817
rect -4253 7783 -4219 7817
rect -4185 7783 -4151 7817
rect -4117 7783 -4083 7817
rect -4049 7783 -4015 7817
rect -3981 7783 -3947 7817
rect -3913 7783 -3879 7817
rect -3845 7783 -3811 7817
rect -3777 7783 -3743 7817
rect -3709 7783 -3675 7817
rect -3641 7783 -3607 7817
rect -3573 7783 -3539 7817
rect -3505 7783 -3471 7817
rect -3437 7783 -3403 7817
rect -3369 7783 -3335 7817
rect -3301 7783 -3267 7817
rect -3233 7783 -3199 7817
rect -3165 7783 -3131 7817
rect -3097 7783 -3063 7817
rect -3029 7783 -2995 7817
rect -2961 7783 -2927 7817
rect -2893 7783 -2859 7817
rect -2825 7783 -2791 7817
rect -2757 7783 -2723 7817
rect -2689 7783 -2655 7817
rect -2621 7783 -2587 7817
rect -2553 7783 -2519 7817
rect -2485 7783 -2451 7817
rect -2417 7783 -2383 7817
rect -2349 7783 -2315 7817
rect -2281 7783 -2247 7817
rect -2213 7783 -2179 7817
rect -2145 7783 -2111 7817
rect -2077 7783 -2043 7817
rect -2009 7783 -1975 7817
rect -1941 7783 -1907 7817
rect -1873 7783 -1839 7817
rect -1805 7783 -1771 7817
rect -1737 7783 -1703 7817
rect -1669 7783 -1635 7817
rect -1601 7783 -1567 7817
rect -1533 7783 -1499 7817
rect -1465 7783 -1431 7817
rect -1397 7783 -1363 7817
rect -1329 7783 -1295 7817
rect -1261 7783 -1227 7817
rect -1193 7783 -1159 7817
rect -1125 7783 -1091 7817
rect -1057 7783 -1023 7817
rect -989 7783 -955 7817
rect -921 7783 -887 7817
rect -853 7783 -819 7817
rect -785 7783 -751 7817
rect -717 7783 -683 7817
rect -649 7783 -615 7817
rect -581 7783 -547 7817
rect -513 7783 -479 7817
rect -445 7783 -411 7817
rect -377 7783 -343 7817
rect -309 7783 -275 7817
rect -241 7783 -207 7817
rect -173 7783 -139 7817
rect -105 7783 -71 7817
rect -37 7783 -3 7817
rect 31 7783 65 7817
rect 99 7783 133 7817
rect 167 7783 201 7817
rect 235 7783 269 7817
rect 303 7783 337 7817
rect 371 7783 405 7817
rect 439 7783 473 7817
rect 507 7783 541 7817
rect 575 7783 609 7817
rect 643 7783 677 7817
rect 711 7783 745 7817
rect 779 7783 813 7817
rect 847 7783 881 7817
rect 915 7783 949 7817
rect 983 7783 1017 7817
rect 1051 7783 1085 7817
rect 1119 7783 1153 7817
rect 1187 7783 1221 7817
rect 1255 7783 1289 7817
rect 1323 7783 1357 7817
rect 1391 7783 1425 7817
rect 1459 7783 1493 7817
rect 1527 7783 1561 7817
rect 1595 7783 1629 7817
rect 1663 7783 1697 7817
rect 1731 7783 1765 7817
rect 1799 7783 1833 7817
rect 1867 7783 1901 7817
rect 1935 7783 1969 7817
rect 2003 7783 2037 7817
rect 2071 7783 2105 7817
rect 2139 7783 2173 7817
rect 2207 7783 2241 7817
rect 2275 7783 2309 7817
rect 2343 7783 2377 7817
rect 2411 7783 2445 7817
rect 2479 7783 2513 7817
rect 2547 7783 2581 7817
rect 2615 7783 2649 7817
rect 2683 7783 2717 7817
rect 2751 7783 2785 7817
rect 2819 7783 2853 7817
rect 2887 7783 2921 7817
rect 2955 7783 2989 7817
rect 3023 7783 3057 7817
rect 3091 7783 3125 7817
rect 3159 7783 3193 7817
rect 3227 7783 3261 7817
rect 3295 7783 3329 7817
rect 3363 7783 3397 7817
rect 3431 7783 3465 7817
rect 3499 7783 3533 7817
rect 3567 7783 3601 7817
rect 3635 7783 3669 7817
rect 3703 7783 3737 7817
rect 3771 7783 3805 7817
rect 3839 7783 3873 7817
rect 3907 7783 3941 7817
rect 3975 7783 4009 7817
rect 4043 7783 4077 7817
rect 4111 7783 4145 7817
rect 4179 7783 4213 7817
rect 4247 7783 4281 7817
rect 4315 7783 4349 7817
rect 4383 7783 4417 7817
rect 4451 7783 4485 7817
rect 4519 7783 4553 7817
rect 4587 7783 4621 7817
rect 4655 7783 4689 7817
rect 4723 7783 4757 7817
rect 4791 7783 4825 7817
rect 4859 7783 4893 7817
rect 4927 7783 4961 7817
rect 4995 7783 5029 7817
rect 5063 7783 5097 7817
rect 5131 7783 5165 7817
rect 5199 7783 5233 7817
rect 5267 7783 5301 7817
rect 5335 7783 5369 7817
rect 5403 7783 5437 7817
rect 5471 7783 5505 7817
rect 5539 7783 5573 7817
rect 5607 7783 5641 7817
rect 5675 7783 5709 7817
rect 5743 7783 5777 7817
rect 5811 7783 5845 7817
rect 5879 7783 5913 7817
rect 5947 7783 5981 7817
rect 6015 7783 6049 7817
rect 6083 7783 6117 7817
rect 6151 7783 6185 7817
rect 6219 7783 6253 7817
rect 6287 7783 6321 7817
rect 6355 7783 6389 7817
rect 6423 7783 6457 7817
rect 6491 7783 6525 7817
rect 6559 7783 6593 7817
rect 6627 7783 6661 7817
rect 6695 7783 6729 7817
rect 6763 7783 6797 7817
rect 6831 7783 6865 7817
rect 6899 7783 6933 7817
rect 6967 7783 7001 7817
rect 7035 7783 7069 7817
rect 7103 7783 7137 7817
rect 7171 7783 7205 7817
rect 7239 7783 7273 7817
rect 7307 7783 7341 7817
rect 7375 7783 7409 7817
rect 7443 7783 7477 7817
rect 7511 7783 7545 7817
rect 7579 7783 7613 7817
rect 7647 7783 7681 7817
rect 7715 7783 7749 7817
rect 7783 7783 7817 7817
rect 7851 7783 7885 7817
rect 7919 7783 7953 7817
rect 7987 7783 8021 7817
rect 8055 7783 8089 7817
rect 8123 7783 8157 7817
rect 8191 7783 8225 7817
rect 8259 7783 8293 7817
rect 8327 7783 8361 7817
rect 8395 7783 8429 7817
rect 8463 7783 8497 7817
rect 8531 7783 8565 7817
rect 8599 7783 8633 7817
rect 8667 7783 8701 7817
rect 8735 7783 8769 7817
rect 8803 7783 8837 7817
rect 8871 7783 8905 7817
rect 8939 7783 8973 7817
rect 9007 7783 9041 7817
rect 9075 7783 9109 7817
rect 9143 7783 9177 7817
rect 9211 7783 9245 7817
rect 9279 7783 9313 7817
rect 9347 7783 9381 7817
rect 9415 7783 9449 7817
rect 9483 7783 9517 7817
rect 9551 7783 9585 7817
rect 9619 7783 9653 7817
rect 9687 7783 9721 7817
rect 9755 7783 9789 7817
rect 9823 7783 9857 7817
rect 9891 7783 9925 7817
rect 9959 7783 9993 7817
rect 10027 7783 10061 7817
rect 10095 7783 10129 7817
rect 10163 7783 10197 7817
rect 10231 7783 10265 7817
rect 10299 7783 10333 7817
rect 10367 7783 10401 7817
rect 10435 7783 10469 7817
rect 10503 7783 10537 7817
rect 10571 7783 10605 7817
rect 10639 7783 10673 7817
rect 10707 7783 10741 7817
rect 10775 7783 10809 7817
rect 10843 7783 10877 7817
rect 10911 7783 10945 7817
rect 10979 7783 11013 7817
rect 11047 7783 11081 7817
rect 11115 7783 11149 7817
rect 11183 7783 11217 7817
rect 11251 7783 11285 7817
rect 11319 7783 11353 7817
rect 11387 7783 11421 7817
rect 11455 7783 11489 7817
rect 11523 7783 11557 7817
rect 11591 7783 11625 7817
rect 11659 7783 11693 7817
rect 11727 7783 11761 7817
rect 11795 7783 11829 7817
rect 11863 7783 11897 7817
rect 11931 7783 11965 7817
rect 11999 7783 12033 7817
rect 12067 7783 12101 7817
rect 12135 7783 12169 7817
rect 12203 7783 12237 7817
rect 12271 7783 12305 7817
rect 12339 7783 12373 7817
rect 12407 7783 12441 7817
rect 12475 7783 12509 7817
rect 12543 7783 12577 7817
rect 12611 7783 12645 7817
rect 12679 7783 12713 7817
rect 12747 7783 12781 7817
rect 12815 7783 12849 7817
rect 12883 7783 12917 7817
rect 12951 7783 12985 7817
rect 13019 7783 13053 7817
rect 13087 7783 13121 7817
rect 13155 7783 13189 7817
rect 13223 7783 13257 7817
rect 13291 7783 13325 7817
rect 13359 7783 13393 7817
rect 13427 7783 13461 7817
rect 13495 7783 13529 7817
rect 13563 7783 13597 7817
rect 13631 7783 13665 7817
rect 13699 7783 13733 7817
rect 13767 7783 13801 7817
rect 13835 7783 13869 7817
rect 13903 7783 13937 7817
rect 13971 7783 14005 7817
rect 14039 7783 14073 7817
rect 14107 7783 14141 7817
rect 14175 7783 14209 7817
rect 14243 7783 14277 7817
rect 14311 7783 14345 7817
rect 14379 7783 14413 7817
rect 14447 7783 14481 7817
rect 14515 7783 14549 7817
rect 14583 7783 14617 7817
rect 14651 7783 14685 7817
rect 14719 7783 14880 7817
rect -12880 7760 14880 7783
rect -12880 7677 -12800 7760
rect -12880 7643 -12857 7677
rect -12823 7643 -12800 7677
rect -12880 7609 -12800 7643
rect -12880 7575 -12857 7609
rect -12823 7575 -12800 7609
rect -12880 7541 -12800 7575
rect -12880 7507 -12857 7541
rect -12823 7507 -12800 7541
rect -12880 7473 -12800 7507
rect -12880 7439 -12857 7473
rect -12823 7439 -12800 7473
rect -12880 7405 -12800 7439
rect -12880 7371 -12857 7405
rect -12823 7371 -12800 7405
rect -12880 7337 -12800 7371
rect -12880 7303 -12857 7337
rect -12823 7303 -12800 7337
rect -12880 7269 -12800 7303
rect -12880 7235 -12857 7269
rect -12823 7235 -12800 7269
rect -12880 7201 -12800 7235
rect -12880 7167 -12857 7201
rect -12823 7167 -12800 7201
rect -12880 7133 -12800 7167
rect -12880 7099 -12857 7133
rect -12823 7099 -12800 7133
rect -12880 7065 -12800 7099
rect -12880 7031 -12857 7065
rect -12823 7031 -12800 7065
rect -12880 6997 -12800 7031
rect -12880 6963 -12857 6997
rect -12823 6963 -12800 6997
rect -12880 6929 -12800 6963
rect -12880 6895 -12857 6929
rect -12823 6895 -12800 6929
rect -12880 6861 -12800 6895
rect -12880 6827 -12857 6861
rect -12823 6827 -12800 6861
rect -12880 6793 -12800 6827
rect -12880 6759 -12857 6793
rect -12823 6759 -12800 6793
rect -12880 6725 -12800 6759
rect -12880 6691 -12857 6725
rect -12823 6691 -12800 6725
rect -12880 6657 -12800 6691
rect -12880 6623 -12857 6657
rect -12823 6623 -12800 6657
rect -12880 6589 -12800 6623
rect -12880 6555 -12857 6589
rect -12823 6555 -12800 6589
rect -12880 6521 -12800 6555
rect -12880 6487 -12857 6521
rect -12823 6487 -12800 6521
rect -12880 6453 -12800 6487
rect -12880 6419 -12857 6453
rect -12823 6419 -12800 6453
rect -12880 6385 -12800 6419
rect -12880 6351 -12857 6385
rect -12823 6351 -12800 6385
rect -12880 6317 -12800 6351
rect -12880 6283 -12857 6317
rect -12823 6283 -12800 6317
rect -12880 6249 -12800 6283
rect -12880 6215 -12857 6249
rect -12823 6215 -12800 6249
rect -12880 6181 -12800 6215
rect -12880 6147 -12857 6181
rect -12823 6147 -12800 6181
rect -12880 6113 -12800 6147
rect -12880 6079 -12857 6113
rect -12823 6079 -12800 6113
rect -12880 6045 -12800 6079
rect -12880 6011 -12857 6045
rect -12823 6011 -12800 6045
rect -12880 5977 -12800 6011
rect -12880 5943 -12857 5977
rect -12823 5943 -12800 5977
rect -12880 5909 -12800 5943
rect -12880 5875 -12857 5909
rect -12823 5875 -12800 5909
rect -12880 5841 -12800 5875
rect -12880 5807 -12857 5841
rect -12823 5807 -12800 5841
rect -12880 5773 -12800 5807
rect -12880 5739 -12857 5773
rect -12823 5739 -12800 5773
rect -12880 5705 -12800 5739
rect -12880 5671 -12857 5705
rect -12823 5671 -12800 5705
rect -12880 5637 -12800 5671
rect -12880 5603 -12857 5637
rect -12823 5603 -12800 5637
rect -12880 5569 -12800 5603
rect -12880 5535 -12857 5569
rect -12823 5535 -12800 5569
rect -12880 5501 -12800 5535
rect -12880 5467 -12857 5501
rect -12823 5467 -12800 5501
rect -12880 5433 -12800 5467
rect -12880 5399 -12857 5433
rect -12823 5399 -12800 5433
rect -12880 5365 -12800 5399
rect -12880 5331 -12857 5365
rect -12823 5331 -12800 5365
rect -12880 5297 -12800 5331
rect -12880 5263 -12857 5297
rect -12823 5263 -12800 5297
rect -12880 5229 -12800 5263
rect -12880 5195 -12857 5229
rect -12823 5195 -12800 5229
rect -12880 5161 -12800 5195
rect -12880 5127 -12857 5161
rect -12823 5127 -12800 5161
rect -12880 5093 -12800 5127
rect -12880 5059 -12857 5093
rect -12823 5059 -12800 5093
rect -12880 5025 -12800 5059
rect -12880 4991 -12857 5025
rect -12823 4991 -12800 5025
rect -12880 4957 -12800 4991
rect -12880 4923 -12857 4957
rect -12823 4923 -12800 4957
rect -12880 4889 -12800 4923
rect -12880 4855 -12857 4889
rect -12823 4855 -12800 4889
rect -12880 4821 -12800 4855
rect -12880 4787 -12857 4821
rect -12823 4787 -12800 4821
rect -12880 4753 -12800 4787
rect -12880 4719 -12857 4753
rect -12823 4719 -12800 4753
rect -12880 4685 -12800 4719
rect -12880 4651 -12857 4685
rect -12823 4651 -12800 4685
rect -12880 4617 -12800 4651
rect -12880 4583 -12857 4617
rect -12823 4583 -12800 4617
rect -12880 4549 -12800 4583
rect -12880 4515 -12857 4549
rect -12823 4515 -12800 4549
rect -12880 4481 -12800 4515
rect -12880 4447 -12857 4481
rect -12823 4447 -12800 4481
rect -12880 4413 -12800 4447
rect -12880 4379 -12857 4413
rect -12823 4379 -12800 4413
rect -12880 4345 -12800 4379
rect -12880 4311 -12857 4345
rect -12823 4311 -12800 4345
rect -12880 4277 -12800 4311
rect -12880 4243 -12857 4277
rect -12823 4243 -12800 4277
rect -12880 4209 -12800 4243
rect -12880 4175 -12857 4209
rect -12823 4175 -12800 4209
rect -12880 4141 -12800 4175
rect -12880 4107 -12857 4141
rect -12823 4107 -12800 4141
rect -12880 4073 -12800 4107
rect -12880 4039 -12857 4073
rect -12823 4039 -12800 4073
rect -12880 4005 -12800 4039
rect -12880 3971 -12857 4005
rect -12823 3971 -12800 4005
rect -12880 3937 -12800 3971
rect -12880 3903 -12857 3937
rect -12823 3903 -12800 3937
rect -12880 3869 -12800 3903
rect -12880 3835 -12857 3869
rect -12823 3835 -12800 3869
rect -12880 3801 -12800 3835
rect -12880 3767 -12857 3801
rect -12823 3767 -12800 3801
rect -12880 3733 -12800 3767
rect -12880 3699 -12857 3733
rect -12823 3699 -12800 3733
rect -12880 3665 -12800 3699
rect -12880 3631 -12857 3665
rect -12823 3631 -12800 3665
rect -12880 3597 -12800 3631
rect -12880 3563 -12857 3597
rect -12823 3563 -12800 3597
rect -12880 3529 -12800 3563
rect -12880 3495 -12857 3529
rect -12823 3495 -12800 3529
rect -12880 3461 -12800 3495
rect -12880 3427 -12857 3461
rect -12823 3427 -12800 3461
rect -12880 3393 -12800 3427
rect -12880 3359 -12857 3393
rect -12823 3359 -12800 3393
rect -12880 3325 -12800 3359
rect -12880 3291 -12857 3325
rect -12823 3291 -12800 3325
rect -12880 3257 -12800 3291
rect -12880 3223 -12857 3257
rect -12823 3223 -12800 3257
rect -12880 3189 -12800 3223
rect -12880 3155 -12857 3189
rect -12823 3155 -12800 3189
rect -12880 3121 -12800 3155
rect -12880 3087 -12857 3121
rect -12823 3087 -12800 3121
rect -12880 3053 -12800 3087
rect -12880 3019 -12857 3053
rect -12823 3019 -12800 3053
rect -12880 2985 -12800 3019
rect -12880 2951 -12857 2985
rect -12823 2951 -12800 2985
rect -12880 2917 -12800 2951
rect -12880 2883 -12857 2917
rect -12823 2883 -12800 2917
rect -12880 2849 -12800 2883
rect -12880 2815 -12857 2849
rect -12823 2815 -12800 2849
rect -12880 2781 -12800 2815
rect -12880 2747 -12857 2781
rect -12823 2747 -12800 2781
rect -12880 2713 -12800 2747
rect -12880 2679 -12857 2713
rect -12823 2679 -12800 2713
rect -12880 2645 -12800 2679
rect -12880 2611 -12857 2645
rect -12823 2611 -12800 2645
rect -12880 2577 -12800 2611
rect -12880 2543 -12857 2577
rect -12823 2543 -12800 2577
rect -12880 2509 -12800 2543
rect -12880 2475 -12857 2509
rect -12823 2475 -12800 2509
rect -12880 2441 -12800 2475
rect -12880 2407 -12857 2441
rect -12823 2407 -12800 2441
rect -12880 2373 -12800 2407
rect -12880 2339 -12857 2373
rect -12823 2339 -12800 2373
rect -12880 2305 -12800 2339
rect -12880 2271 -12857 2305
rect -12823 2271 -12800 2305
rect -12880 2237 -12800 2271
rect -12880 2203 -12857 2237
rect -12823 2203 -12800 2237
rect -12880 2169 -12800 2203
rect -12880 2135 -12857 2169
rect -12823 2135 -12800 2169
rect -12880 2101 -12800 2135
rect -12880 2067 -12857 2101
rect -12823 2067 -12800 2101
rect -12880 2033 -12800 2067
rect -12880 1999 -12857 2033
rect -12823 1999 -12800 2033
rect -12880 1965 -12800 1999
rect -12880 1931 -12857 1965
rect -12823 1931 -12800 1965
rect -12880 1897 -12800 1931
rect -12880 1863 -12857 1897
rect -12823 1863 -12800 1897
rect -12880 1829 -12800 1863
rect -12880 1795 -12857 1829
rect -12823 1795 -12800 1829
rect -12880 1761 -12800 1795
rect -12880 1727 -12857 1761
rect -12823 1727 -12800 1761
rect -12880 1693 -12800 1727
rect -12880 1659 -12857 1693
rect -12823 1659 -12800 1693
rect -12880 1625 -12800 1659
rect -12880 1591 -12857 1625
rect -12823 1591 -12800 1625
rect -12880 1557 -12800 1591
rect -12880 1523 -12857 1557
rect -12823 1523 -12800 1557
rect -12880 1440 -12800 1523
rect 14800 7677 14880 7760
rect 14800 7643 14823 7677
rect 14857 7643 14880 7677
rect 14800 7609 14880 7643
rect 14800 7575 14823 7609
rect 14857 7575 14880 7609
rect 14800 7541 14880 7575
rect 14800 7507 14823 7541
rect 14857 7507 14880 7541
rect 14800 7473 14880 7507
rect 14800 7439 14823 7473
rect 14857 7439 14880 7473
rect 14800 7405 14880 7439
rect 14800 7371 14823 7405
rect 14857 7371 14880 7405
rect 14800 7337 14880 7371
rect 14800 7303 14823 7337
rect 14857 7303 14880 7337
rect 14800 7269 14880 7303
rect 14800 7235 14823 7269
rect 14857 7235 14880 7269
rect 14800 7201 14880 7235
rect 14800 7167 14823 7201
rect 14857 7167 14880 7201
rect 14800 7133 14880 7167
rect 14800 7099 14823 7133
rect 14857 7099 14880 7133
rect 14800 7065 14880 7099
rect 14800 7031 14823 7065
rect 14857 7031 14880 7065
rect 14800 6997 14880 7031
rect 14800 6963 14823 6997
rect 14857 6963 14880 6997
rect 14800 6929 14880 6963
rect 14800 6895 14823 6929
rect 14857 6895 14880 6929
rect 14800 6861 14880 6895
rect 14800 6827 14823 6861
rect 14857 6827 14880 6861
rect 14800 6793 14880 6827
rect 14800 6759 14823 6793
rect 14857 6759 14880 6793
rect 14800 6725 14880 6759
rect 14800 6691 14823 6725
rect 14857 6691 14880 6725
rect 14800 6657 14880 6691
rect 14800 6623 14823 6657
rect 14857 6623 14880 6657
rect 14800 6589 14880 6623
rect 14800 6555 14823 6589
rect 14857 6555 14880 6589
rect 14800 6521 14880 6555
rect 14800 6487 14823 6521
rect 14857 6487 14880 6521
rect 14800 6453 14880 6487
rect 14800 6419 14823 6453
rect 14857 6419 14880 6453
rect 14800 6385 14880 6419
rect 14800 6351 14823 6385
rect 14857 6351 14880 6385
rect 14800 6317 14880 6351
rect 14800 6283 14823 6317
rect 14857 6283 14880 6317
rect 14800 6249 14880 6283
rect 14800 6215 14823 6249
rect 14857 6215 14880 6249
rect 14800 6181 14880 6215
rect 14800 6147 14823 6181
rect 14857 6147 14880 6181
rect 14800 6113 14880 6147
rect 14800 6079 14823 6113
rect 14857 6079 14880 6113
rect 14800 6045 14880 6079
rect 14800 6011 14823 6045
rect 14857 6011 14880 6045
rect 14800 5977 14880 6011
rect 14800 5943 14823 5977
rect 14857 5943 14880 5977
rect 14800 5909 14880 5943
rect 14800 5875 14823 5909
rect 14857 5875 14880 5909
rect 14800 5841 14880 5875
rect 14800 5807 14823 5841
rect 14857 5807 14880 5841
rect 14800 5773 14880 5807
rect 14800 5739 14823 5773
rect 14857 5739 14880 5773
rect 14800 5705 14880 5739
rect 14800 5671 14823 5705
rect 14857 5671 14880 5705
rect 14800 5637 14880 5671
rect 14800 5603 14823 5637
rect 14857 5603 14880 5637
rect 14800 5569 14880 5603
rect 14800 5535 14823 5569
rect 14857 5535 14880 5569
rect 14800 5501 14880 5535
rect 14800 5467 14823 5501
rect 14857 5467 14880 5501
rect 14800 5433 14880 5467
rect 14800 5399 14823 5433
rect 14857 5399 14880 5433
rect 14800 5365 14880 5399
rect 14800 5331 14823 5365
rect 14857 5331 14880 5365
rect 14800 5297 14880 5331
rect 14800 5263 14823 5297
rect 14857 5263 14880 5297
rect 14800 5229 14880 5263
rect 14800 5195 14823 5229
rect 14857 5195 14880 5229
rect 14800 5161 14880 5195
rect 14800 5127 14823 5161
rect 14857 5127 14880 5161
rect 14800 5093 14880 5127
rect 14800 5059 14823 5093
rect 14857 5059 14880 5093
rect 14800 5025 14880 5059
rect 14800 4991 14823 5025
rect 14857 4991 14880 5025
rect 14800 4957 14880 4991
rect 14800 4923 14823 4957
rect 14857 4923 14880 4957
rect 14800 4889 14880 4923
rect 14800 4855 14823 4889
rect 14857 4855 14880 4889
rect 14800 4821 14880 4855
rect 14800 4787 14823 4821
rect 14857 4787 14880 4821
rect 14800 4753 14880 4787
rect 14800 4719 14823 4753
rect 14857 4719 14880 4753
rect 14800 4685 14880 4719
rect 14800 4651 14823 4685
rect 14857 4651 14880 4685
rect 14800 4617 14880 4651
rect 14800 4583 14823 4617
rect 14857 4583 14880 4617
rect 14800 4549 14880 4583
rect 14800 4515 14823 4549
rect 14857 4515 14880 4549
rect 14800 4481 14880 4515
rect 14800 4447 14823 4481
rect 14857 4447 14880 4481
rect 14800 4413 14880 4447
rect 14800 4379 14823 4413
rect 14857 4379 14880 4413
rect 14800 4345 14880 4379
rect 14800 4311 14823 4345
rect 14857 4311 14880 4345
rect 14800 4277 14880 4311
rect 14800 4243 14823 4277
rect 14857 4243 14880 4277
rect 14800 4209 14880 4243
rect 14800 4175 14823 4209
rect 14857 4175 14880 4209
rect 14800 4141 14880 4175
rect 14800 4107 14823 4141
rect 14857 4107 14880 4141
rect 14800 4073 14880 4107
rect 14800 4039 14823 4073
rect 14857 4039 14880 4073
rect 14800 4005 14880 4039
rect 14800 3971 14823 4005
rect 14857 3971 14880 4005
rect 14800 3937 14880 3971
rect 14800 3903 14823 3937
rect 14857 3903 14880 3937
rect 14800 3869 14880 3903
rect 14800 3835 14823 3869
rect 14857 3835 14880 3869
rect 14800 3801 14880 3835
rect 14800 3767 14823 3801
rect 14857 3767 14880 3801
rect 14800 3733 14880 3767
rect 14800 3699 14823 3733
rect 14857 3699 14880 3733
rect 14800 3665 14880 3699
rect 14800 3631 14823 3665
rect 14857 3631 14880 3665
rect 14800 3597 14880 3631
rect 14800 3563 14823 3597
rect 14857 3563 14880 3597
rect 14800 3529 14880 3563
rect 14800 3495 14823 3529
rect 14857 3495 14880 3529
rect 14800 3461 14880 3495
rect 14800 3427 14823 3461
rect 14857 3427 14880 3461
rect 14800 3393 14880 3427
rect 14800 3359 14823 3393
rect 14857 3359 14880 3393
rect 14800 3325 14880 3359
rect 14800 3291 14823 3325
rect 14857 3291 14880 3325
rect 14800 3257 14880 3291
rect 14800 3223 14823 3257
rect 14857 3223 14880 3257
rect 14800 3189 14880 3223
rect 14800 3155 14823 3189
rect 14857 3155 14880 3189
rect 14800 3121 14880 3155
rect 14800 3087 14823 3121
rect 14857 3087 14880 3121
rect 14800 3053 14880 3087
rect 14800 3019 14823 3053
rect 14857 3019 14880 3053
rect 14800 2985 14880 3019
rect 14800 2951 14823 2985
rect 14857 2951 14880 2985
rect 14800 2917 14880 2951
rect 14800 2883 14823 2917
rect 14857 2883 14880 2917
rect 14800 2849 14880 2883
rect 14800 2815 14823 2849
rect 14857 2815 14880 2849
rect 14800 2781 14880 2815
rect 14800 2747 14823 2781
rect 14857 2747 14880 2781
rect 14800 2713 14880 2747
rect 14800 2679 14823 2713
rect 14857 2679 14880 2713
rect 14800 2645 14880 2679
rect 14800 2611 14823 2645
rect 14857 2611 14880 2645
rect 14800 2577 14880 2611
rect 14800 2543 14823 2577
rect 14857 2543 14880 2577
rect 14800 2509 14880 2543
rect 14800 2475 14823 2509
rect 14857 2475 14880 2509
rect 14800 2441 14880 2475
rect 14800 2407 14823 2441
rect 14857 2407 14880 2441
rect 14800 2373 14880 2407
rect 14800 2339 14823 2373
rect 14857 2339 14880 2373
rect 14800 2305 14880 2339
rect 14800 2271 14823 2305
rect 14857 2271 14880 2305
rect 14800 2237 14880 2271
rect 14800 2203 14823 2237
rect 14857 2203 14880 2237
rect 14800 2169 14880 2203
rect 14800 2135 14823 2169
rect 14857 2135 14880 2169
rect 14800 2101 14880 2135
rect 14800 2067 14823 2101
rect 14857 2067 14880 2101
rect 14800 2033 14880 2067
rect 14800 1999 14823 2033
rect 14857 1999 14880 2033
rect 14800 1965 14880 1999
rect 14800 1931 14823 1965
rect 14857 1931 14880 1965
rect 14800 1897 14880 1931
rect 14800 1863 14823 1897
rect 14857 1863 14880 1897
rect 14800 1829 14880 1863
rect 14800 1795 14823 1829
rect 14857 1795 14880 1829
rect 14800 1761 14880 1795
rect 14800 1727 14823 1761
rect 14857 1727 14880 1761
rect 14800 1693 14880 1727
rect 14800 1659 14823 1693
rect 14857 1659 14880 1693
rect 14800 1625 14880 1659
rect 14800 1591 14823 1625
rect 14857 1591 14880 1625
rect 14800 1557 14880 1591
rect 14800 1523 14823 1557
rect 14857 1523 14880 1557
rect 14800 1440 14880 1523
rect -12880 1417 14880 1440
rect -12880 1383 -12719 1417
rect -12685 1383 -12651 1417
rect -12617 1383 -12583 1417
rect -12549 1383 -12515 1417
rect -12481 1383 -12447 1417
rect -12413 1383 -12379 1417
rect -12345 1383 -12311 1417
rect -12277 1383 -12243 1417
rect -12209 1383 -12175 1417
rect -12141 1383 -12107 1417
rect -12073 1383 -12039 1417
rect -12005 1383 -11971 1417
rect -11937 1383 -11903 1417
rect -11869 1383 -11835 1417
rect -11801 1383 -11767 1417
rect -11733 1383 -11699 1417
rect -11665 1383 -11631 1417
rect -11597 1383 -11563 1417
rect -11529 1383 -11495 1417
rect -11461 1383 -11427 1417
rect -11393 1383 -11359 1417
rect -11325 1383 -11291 1417
rect -11257 1383 -11223 1417
rect -11189 1383 -11155 1417
rect -11121 1383 -11087 1417
rect -11053 1383 -11019 1417
rect -10985 1383 -10951 1417
rect -10917 1383 -10883 1417
rect -10849 1383 -10815 1417
rect -10781 1383 -10747 1417
rect -10713 1383 -10679 1417
rect -10645 1383 -10611 1417
rect -10577 1383 -10543 1417
rect -10509 1383 -10475 1417
rect -10441 1383 -10407 1417
rect -10373 1383 -10339 1417
rect -10305 1383 -10271 1417
rect -10237 1383 -10203 1417
rect -10169 1383 -10135 1417
rect -10101 1383 -10067 1417
rect -10033 1383 -9999 1417
rect -9965 1383 -9931 1417
rect -9897 1383 -9863 1417
rect -9829 1383 -9795 1417
rect -9761 1383 -9727 1417
rect -9693 1383 -9659 1417
rect -9625 1383 -9591 1417
rect -9557 1383 -9523 1417
rect -9489 1383 -9455 1417
rect -9421 1383 -9387 1417
rect -9353 1383 -9319 1417
rect -9285 1383 -9251 1417
rect -9217 1383 -9183 1417
rect -9149 1383 -9115 1417
rect -9081 1383 -9047 1417
rect -9013 1383 -8979 1417
rect -8945 1383 -8911 1417
rect -8877 1383 -8843 1417
rect -8809 1383 -8775 1417
rect -8741 1383 -8707 1417
rect -8673 1383 -8639 1417
rect -8605 1383 -8571 1417
rect -8537 1383 -8503 1417
rect -8469 1383 -8435 1417
rect -8401 1383 -8367 1417
rect -8333 1383 -8299 1417
rect -8265 1383 -8231 1417
rect -8197 1383 -8163 1417
rect -8129 1383 -8095 1417
rect -8061 1383 -8027 1417
rect -7993 1383 -7959 1417
rect -7925 1383 -7891 1417
rect -7857 1383 -7823 1417
rect -7789 1383 -7755 1417
rect -7721 1383 -7687 1417
rect -7653 1383 -7619 1417
rect -7585 1383 -7551 1417
rect -7517 1383 -7483 1417
rect -7449 1383 -7415 1417
rect -7381 1383 -7347 1417
rect -7313 1383 -7279 1417
rect -7245 1383 -7211 1417
rect -7177 1383 -7143 1417
rect -7109 1383 -7075 1417
rect -7041 1383 -7007 1417
rect -6973 1383 -6939 1417
rect -6905 1383 -6871 1417
rect -6837 1383 -6803 1417
rect -6769 1383 -6735 1417
rect -6701 1383 -6667 1417
rect -6633 1383 -6599 1417
rect -6565 1383 -6531 1417
rect -6497 1383 -6463 1417
rect -6429 1383 -6395 1417
rect -6361 1383 -6327 1417
rect -6293 1383 -6259 1417
rect -6225 1383 -6191 1417
rect -6157 1383 -6123 1417
rect -6089 1383 -6055 1417
rect -6021 1383 -5987 1417
rect -5953 1383 -5919 1417
rect -5885 1383 -5851 1417
rect -5817 1383 -5783 1417
rect -5749 1383 -5715 1417
rect -5681 1383 -5647 1417
rect -5613 1383 -5579 1417
rect -5545 1383 -5511 1417
rect -5477 1383 -5443 1417
rect -5409 1383 -5375 1417
rect -5341 1383 -5307 1417
rect -5273 1383 -5239 1417
rect -5205 1383 -5171 1417
rect -5137 1383 -5103 1417
rect -5069 1383 -5035 1417
rect -5001 1383 -4967 1417
rect -4933 1383 -4899 1417
rect -4865 1383 -4831 1417
rect -4797 1383 -4763 1417
rect -4729 1383 -4695 1417
rect -4661 1383 -4627 1417
rect -4593 1383 -4559 1417
rect -4525 1383 -4491 1417
rect -4457 1383 -4423 1417
rect -4389 1383 -4355 1417
rect -4321 1383 -4287 1417
rect -4253 1383 -4219 1417
rect -4185 1383 -4151 1417
rect -4117 1383 -4083 1417
rect -4049 1383 -4015 1417
rect -3981 1383 -3947 1417
rect -3913 1383 -3879 1417
rect -3845 1383 -3811 1417
rect -3777 1383 -3743 1417
rect -3709 1383 -3675 1417
rect -3641 1383 -3607 1417
rect -3573 1383 -3539 1417
rect -3505 1383 -3471 1417
rect -3437 1383 -3403 1417
rect -3369 1383 -3335 1417
rect -3301 1383 -3267 1417
rect -3233 1383 -3199 1417
rect -3165 1383 -3131 1417
rect -3097 1383 -3063 1417
rect -3029 1383 -2995 1417
rect -2961 1383 -2927 1417
rect -2893 1383 -2859 1417
rect -2825 1383 -2791 1417
rect -2757 1383 -2723 1417
rect -2689 1383 -2655 1417
rect -2621 1383 -2587 1417
rect -2553 1383 -2519 1417
rect -2485 1383 -2451 1417
rect -2417 1383 -2383 1417
rect -2349 1383 -2315 1417
rect -2281 1383 -2247 1417
rect -2213 1383 -2179 1417
rect -2145 1383 -2111 1417
rect -2077 1383 -2043 1417
rect -2009 1383 -1975 1417
rect -1941 1383 -1907 1417
rect -1873 1383 -1839 1417
rect -1805 1383 -1771 1417
rect -1737 1383 -1703 1417
rect -1669 1383 -1635 1417
rect -1601 1383 -1567 1417
rect -1533 1383 -1499 1417
rect -1465 1383 -1431 1417
rect -1397 1383 -1363 1417
rect -1329 1383 -1295 1417
rect -1261 1383 -1227 1417
rect -1193 1383 -1159 1417
rect -1125 1383 -1091 1417
rect -1057 1383 -1023 1417
rect -989 1383 -955 1417
rect -921 1383 -887 1417
rect -853 1383 -819 1417
rect -785 1383 -751 1417
rect -717 1383 -683 1417
rect -649 1383 -615 1417
rect -581 1383 -547 1417
rect -513 1383 -479 1417
rect -445 1383 -411 1417
rect -377 1383 -343 1417
rect -309 1383 -275 1417
rect -241 1383 -207 1417
rect -173 1383 -139 1417
rect -105 1383 -71 1417
rect -37 1383 -3 1417
rect 31 1383 65 1417
rect 99 1383 133 1417
rect 167 1383 201 1417
rect 235 1383 269 1417
rect 303 1383 337 1417
rect 371 1383 405 1417
rect 439 1383 473 1417
rect 507 1383 541 1417
rect 575 1383 609 1417
rect 643 1383 677 1417
rect 711 1383 745 1417
rect 779 1383 813 1417
rect 847 1383 881 1417
rect 915 1383 949 1417
rect 983 1383 1017 1417
rect 1051 1383 1085 1417
rect 1119 1383 1153 1417
rect 1187 1383 1221 1417
rect 1255 1383 1289 1417
rect 1323 1383 1357 1417
rect 1391 1383 1425 1417
rect 1459 1383 1493 1417
rect 1527 1383 1561 1417
rect 1595 1383 1629 1417
rect 1663 1383 1697 1417
rect 1731 1383 1765 1417
rect 1799 1383 1833 1417
rect 1867 1383 1901 1417
rect 1935 1383 1969 1417
rect 2003 1383 2037 1417
rect 2071 1383 2105 1417
rect 2139 1383 2173 1417
rect 2207 1383 2241 1417
rect 2275 1383 2309 1417
rect 2343 1383 2377 1417
rect 2411 1383 2445 1417
rect 2479 1383 2513 1417
rect 2547 1383 2581 1417
rect 2615 1383 2649 1417
rect 2683 1383 2717 1417
rect 2751 1383 2785 1417
rect 2819 1383 2853 1417
rect 2887 1383 2921 1417
rect 2955 1383 2989 1417
rect 3023 1383 3057 1417
rect 3091 1383 3125 1417
rect 3159 1383 3193 1417
rect 3227 1383 3261 1417
rect 3295 1383 3329 1417
rect 3363 1383 3397 1417
rect 3431 1383 3465 1417
rect 3499 1383 3533 1417
rect 3567 1383 3601 1417
rect 3635 1383 3669 1417
rect 3703 1383 3737 1417
rect 3771 1383 3805 1417
rect 3839 1383 3873 1417
rect 3907 1383 3941 1417
rect 3975 1383 4009 1417
rect 4043 1383 4077 1417
rect 4111 1383 4145 1417
rect 4179 1383 4213 1417
rect 4247 1383 4281 1417
rect 4315 1383 4349 1417
rect 4383 1383 4417 1417
rect 4451 1383 4485 1417
rect 4519 1383 4553 1417
rect 4587 1383 4621 1417
rect 4655 1383 4689 1417
rect 4723 1383 4757 1417
rect 4791 1383 4825 1417
rect 4859 1383 4893 1417
rect 4927 1383 4961 1417
rect 4995 1383 5029 1417
rect 5063 1383 5097 1417
rect 5131 1383 5165 1417
rect 5199 1383 5233 1417
rect 5267 1383 5301 1417
rect 5335 1383 5369 1417
rect 5403 1383 5437 1417
rect 5471 1383 5505 1417
rect 5539 1383 5573 1417
rect 5607 1383 5641 1417
rect 5675 1383 5709 1417
rect 5743 1383 5777 1417
rect 5811 1383 5845 1417
rect 5879 1383 5913 1417
rect 5947 1383 5981 1417
rect 6015 1383 6049 1417
rect 6083 1383 6117 1417
rect 6151 1383 6185 1417
rect 6219 1383 6253 1417
rect 6287 1383 6321 1417
rect 6355 1383 6389 1417
rect 6423 1383 6457 1417
rect 6491 1383 6525 1417
rect 6559 1383 6593 1417
rect 6627 1383 6661 1417
rect 6695 1383 6729 1417
rect 6763 1383 6797 1417
rect 6831 1383 6865 1417
rect 6899 1383 6933 1417
rect 6967 1383 7001 1417
rect 7035 1383 7069 1417
rect 7103 1383 7137 1417
rect 7171 1383 7205 1417
rect 7239 1383 7273 1417
rect 7307 1383 7341 1417
rect 7375 1383 7409 1417
rect 7443 1383 7477 1417
rect 7511 1383 7545 1417
rect 7579 1383 7613 1417
rect 7647 1383 7681 1417
rect 7715 1383 7749 1417
rect 7783 1383 7817 1417
rect 7851 1383 7885 1417
rect 7919 1383 7953 1417
rect 7987 1383 8021 1417
rect 8055 1383 8089 1417
rect 8123 1383 8157 1417
rect 8191 1383 8225 1417
rect 8259 1383 8293 1417
rect 8327 1383 8361 1417
rect 8395 1383 8429 1417
rect 8463 1383 8497 1417
rect 8531 1383 8565 1417
rect 8599 1383 8633 1417
rect 8667 1383 8701 1417
rect 8735 1383 8769 1417
rect 8803 1383 8837 1417
rect 8871 1383 8905 1417
rect 8939 1383 8973 1417
rect 9007 1383 9041 1417
rect 9075 1383 9109 1417
rect 9143 1383 9177 1417
rect 9211 1383 9245 1417
rect 9279 1383 9313 1417
rect 9347 1383 9381 1417
rect 9415 1383 9449 1417
rect 9483 1383 9517 1417
rect 9551 1383 9585 1417
rect 9619 1383 9653 1417
rect 9687 1383 9721 1417
rect 9755 1383 9789 1417
rect 9823 1383 9857 1417
rect 9891 1383 9925 1417
rect 9959 1383 9993 1417
rect 10027 1383 10061 1417
rect 10095 1383 10129 1417
rect 10163 1383 10197 1417
rect 10231 1383 10265 1417
rect 10299 1383 10333 1417
rect 10367 1383 10401 1417
rect 10435 1383 10469 1417
rect 10503 1383 10537 1417
rect 10571 1383 10605 1417
rect 10639 1383 10673 1417
rect 10707 1383 10741 1417
rect 10775 1383 10809 1417
rect 10843 1383 10877 1417
rect 10911 1383 10945 1417
rect 10979 1383 11013 1417
rect 11047 1383 11081 1417
rect 11115 1383 11149 1417
rect 11183 1383 11217 1417
rect 11251 1383 11285 1417
rect 11319 1383 11353 1417
rect 11387 1383 11421 1417
rect 11455 1383 11489 1417
rect 11523 1383 11557 1417
rect 11591 1383 11625 1417
rect 11659 1383 11693 1417
rect 11727 1383 11761 1417
rect 11795 1383 11829 1417
rect 11863 1383 11897 1417
rect 11931 1383 11965 1417
rect 11999 1383 12033 1417
rect 12067 1383 12101 1417
rect 12135 1383 12169 1417
rect 12203 1383 12237 1417
rect 12271 1383 12305 1417
rect 12339 1383 12373 1417
rect 12407 1383 12441 1417
rect 12475 1383 12509 1417
rect 12543 1383 12577 1417
rect 12611 1383 12645 1417
rect 12679 1383 12713 1417
rect 12747 1383 12781 1417
rect 12815 1383 12849 1417
rect 12883 1383 12917 1417
rect 12951 1383 12985 1417
rect 13019 1383 13053 1417
rect 13087 1383 13121 1417
rect 13155 1383 13189 1417
rect 13223 1383 13257 1417
rect 13291 1383 13325 1417
rect 13359 1383 13393 1417
rect 13427 1383 13461 1417
rect 13495 1383 13529 1417
rect 13563 1383 13597 1417
rect 13631 1383 13665 1417
rect 13699 1383 13733 1417
rect 13767 1383 13801 1417
rect 13835 1383 13869 1417
rect 13903 1383 13937 1417
rect 13971 1383 14005 1417
rect 14039 1383 14073 1417
rect 14107 1383 14141 1417
rect 14175 1383 14209 1417
rect 14243 1383 14277 1417
rect 14311 1383 14345 1417
rect 14379 1383 14413 1417
rect 14447 1383 14481 1417
rect 14515 1383 14549 1417
rect 14583 1383 14617 1417
rect 14651 1383 14685 1417
rect 14719 1383 14880 1417
rect -12880 1360 14880 1383
<< metal3 >>
rect -12720 7672 -12640 7680
rect -12720 7608 -12712 7672
rect -12648 7608 -12640 7672
rect -12720 7352 -12640 7608
rect -12720 7288 -12712 7352
rect -12648 7288 -12640 7352
rect -12720 7032 -12640 7288
rect -12720 6968 -12712 7032
rect -12648 6968 -12640 7032
rect -12720 6880 -12640 6968
rect -12560 7672 -12480 7680
rect -12560 7608 -12552 7672
rect -12488 7608 -12480 7672
rect -12560 7352 -12480 7608
rect -12560 7288 -12552 7352
rect -12488 7288 -12480 7352
rect -12560 7032 -12480 7288
rect -12560 6968 -12552 7032
rect -12488 6968 -12480 7032
rect -12560 6880 -12480 6968
rect -12400 7672 -12320 7680
rect -12400 7608 -12392 7672
rect -12328 7608 -12320 7672
rect -12400 7352 -12320 7608
rect 14320 7672 14400 7680
rect 14320 7608 14328 7672
rect 14392 7608 14400 7672
rect -12400 7288 -12392 7352
rect -12328 7288 -12320 7352
rect -12400 7032 -12320 7288
rect -11040 7512 -10960 7520
rect -11040 7448 -11032 7512
rect -10968 7448 -10960 7512
rect -12400 6968 -12392 7032
rect -12328 6968 -12320 7032
rect -12400 6880 -12320 6968
rect -12720 4720 -12320 6880
rect -12240 7032 -12160 7040
rect -12240 6968 -12232 7032
rect -12168 6968 -12160 7032
rect -12240 4720 -12160 6968
rect -11040 6880 -10960 7448
rect -8640 7512 -8560 7520
rect -8640 7448 -8632 7512
rect -8568 7448 -8560 7512
rect -9840 7032 -9760 7040
rect -9840 6968 -9832 7032
rect -9768 6968 -9760 7032
rect -12080 4720 -9920 6880
rect -9840 4720 -9760 6968
rect -8640 6880 -8560 7448
rect -6240 7512 -6160 7520
rect -6240 7448 -6232 7512
rect -6168 7448 -6160 7512
rect -7440 7032 -7360 7040
rect -7440 6968 -7432 7032
rect -7368 6968 -7360 7032
rect -9680 4720 -7520 6880
rect -7440 4720 -7360 6968
rect -6240 6880 -6160 7448
rect -3840 7512 -3760 7520
rect -3840 7448 -3832 7512
rect -3768 7448 -3760 7512
rect -5040 7032 -4960 7040
rect -5040 6968 -5032 7032
rect -4968 6968 -4960 7032
rect -7280 4720 -5120 6880
rect -5040 4720 -4960 6968
rect -3840 6880 -3760 7448
rect -1440 7512 -1360 7520
rect -1440 7448 -1432 7512
rect -1368 7448 -1360 7512
rect -2640 7032 -2560 7040
rect -2640 6968 -2632 7032
rect -2568 6968 -2560 7032
rect -4880 4720 -2720 6880
rect -2640 4720 -2560 6968
rect -1440 6880 -1360 7448
rect 3360 7512 3440 7520
rect 3360 7448 3368 7512
rect 3432 7448 3440 7512
rect 960 7192 1040 7200
rect 960 7128 968 7192
rect 1032 7128 1040 7192
rect -240 7032 -160 7040
rect -240 6968 -232 7032
rect -168 6968 -160 7032
rect -2480 4720 -320 6880
rect -240 4720 -160 6968
rect 960 6880 1040 7128
rect 2160 7032 2240 7040
rect 2160 6968 2168 7032
rect 2232 6968 2240 7032
rect -80 4720 2080 6880
rect 2160 4720 2240 6968
rect 3360 6880 3440 7448
rect 5760 7512 5840 7520
rect 5760 7448 5768 7512
rect 5832 7448 5840 7512
rect 4560 7032 4640 7040
rect 4560 6968 4568 7032
rect 4632 6968 4640 7032
rect 2320 4720 4480 6880
rect 4560 4720 4640 6968
rect 5760 6880 5840 7448
rect 8160 7512 8240 7520
rect 8160 7448 8168 7512
rect 8232 7448 8240 7512
rect 6960 7032 7040 7040
rect 6960 6968 6968 7032
rect 7032 6968 7040 7032
rect 4720 4720 6880 6880
rect 6960 4720 7040 6968
rect 8160 6880 8240 7448
rect 10560 7512 10640 7520
rect 10560 7448 10568 7512
rect 10632 7448 10640 7512
rect 9360 7032 9440 7040
rect 9360 6968 9368 7032
rect 9432 6968 9440 7032
rect 7120 4720 9280 6880
rect 9360 4720 9440 6968
rect 10560 6880 10640 7448
rect 12960 7512 13040 7520
rect 12960 7448 12968 7512
rect 13032 7448 13040 7512
rect 11760 7032 11840 7040
rect 11760 6968 11768 7032
rect 11832 6968 11840 7032
rect 9520 4720 11680 6880
rect 11760 4720 11840 6968
rect 12960 6880 13040 7448
rect 14320 7352 14400 7608
rect 14320 7288 14328 7352
rect 14392 7288 14400 7352
rect 14160 7032 14240 7040
rect 14160 6968 14168 7032
rect 14232 6968 14240 7032
rect 11920 4720 14080 6880
rect 14160 4720 14240 6968
rect 14320 7032 14400 7288
rect 14320 6968 14328 7032
rect 14392 6968 14400 7032
rect 14320 6880 14400 6968
rect 14480 7672 14560 7680
rect 14480 7608 14488 7672
rect 14552 7608 14560 7672
rect 14480 7352 14560 7608
rect 14480 7288 14488 7352
rect 14552 7288 14560 7352
rect 14480 7032 14560 7288
rect 14480 6968 14488 7032
rect 14552 6968 14560 7032
rect 14480 6880 14560 6968
rect 14640 7672 14720 7680
rect 14640 7608 14648 7672
rect 14712 7608 14720 7672
rect 14640 7352 14720 7608
rect 14640 7288 14648 7352
rect 14712 7288 14720 7352
rect 14640 7032 14720 7288
rect 14640 6968 14648 7032
rect 14712 6968 14720 7032
rect 14640 6880 14720 6968
rect 14320 4720 14720 6880
rect -12720 4480 -12640 4720
rect -12560 4480 -12480 4720
rect -12400 4480 -12320 4720
rect 14320 4480 14400 4720
rect 14480 4480 14560 4720
rect 14640 4480 14720 4720
rect -12720 2320 -12320 4480
rect -12720 2232 -12640 2320
rect -12720 2168 -12712 2232
rect -12648 2168 -12640 2232
rect -12720 1912 -12640 2168
rect -12720 1848 -12712 1912
rect -12648 1848 -12640 1912
rect -12720 1592 -12640 1848
rect -12720 1528 -12712 1592
rect -12648 1528 -12640 1592
rect -12720 1520 -12640 1528
rect -12560 2232 -12480 2320
rect -12560 2168 -12552 2232
rect -12488 2168 -12480 2232
rect -12560 1912 -12480 2168
rect -12560 1848 -12552 1912
rect -12488 1848 -12480 1912
rect -12560 1592 -12480 1848
rect -12560 1528 -12552 1592
rect -12488 1528 -12480 1592
rect -12560 1520 -12480 1528
rect -12400 2232 -12320 2320
rect -12400 2168 -12392 2232
rect -12328 2168 -12320 2232
rect -12400 1912 -12320 2168
rect -12240 2232 -12160 4480
rect -12080 2320 -9920 4480
rect -12240 2168 -12232 2232
rect -12168 2168 -12160 2232
rect -12240 2160 -12160 2168
rect -12400 1848 -12392 1912
rect -12328 1848 -12320 1912
rect -12400 1592 -12320 1848
rect -11040 1752 -10960 2320
rect -9840 2232 -9760 4480
rect -9680 2320 -7520 4480
rect -9840 2168 -9832 2232
rect -9768 2168 -9760 2232
rect -9840 2160 -9760 2168
rect -11040 1688 -11032 1752
rect -10968 1688 -10960 1752
rect -11040 1680 -10960 1688
rect -8640 1752 -8560 2320
rect -7440 2232 -7360 4480
rect -7280 2320 -5120 4480
rect -7440 2168 -7432 2232
rect -7368 2168 -7360 2232
rect -7440 2160 -7360 2168
rect -8640 1688 -8632 1752
rect -8568 1688 -8560 1752
rect -8640 1680 -8560 1688
rect -6240 1752 -6160 2320
rect -5040 2232 -4960 4480
rect -4880 2320 -2720 4480
rect -5040 2168 -5032 2232
rect -4968 2168 -4960 2232
rect -5040 2160 -4960 2168
rect -6240 1688 -6232 1752
rect -6168 1688 -6160 1752
rect -6240 1680 -6160 1688
rect -3840 1752 -3760 2320
rect -2640 2232 -2560 4480
rect -2480 2320 -320 4480
rect -2640 2168 -2632 2232
rect -2568 2168 -2560 2232
rect -2640 2160 -2560 2168
rect -3840 1688 -3832 1752
rect -3768 1688 -3760 1752
rect -3840 1680 -3760 1688
rect -1440 1752 -1360 2320
rect -240 2232 -160 4480
rect -80 2320 2080 4480
rect -240 2168 -232 2232
rect -168 2168 -160 2232
rect -240 2160 -160 2168
rect 960 2072 1040 2320
rect 2160 2232 2240 4480
rect 2320 2320 4480 4480
rect 2160 2168 2168 2232
rect 2232 2168 2240 2232
rect 2160 2160 2240 2168
rect 960 2008 968 2072
rect 1032 2008 1040 2072
rect 960 2000 1040 2008
rect -1440 1688 -1432 1752
rect -1368 1688 -1360 1752
rect -1440 1680 -1360 1688
rect 3360 1752 3440 2320
rect 4560 2232 4640 4480
rect 4720 2320 6880 4480
rect 4560 2168 4568 2232
rect 4632 2168 4640 2232
rect 4560 2160 4640 2168
rect 3360 1688 3368 1752
rect 3432 1688 3440 1752
rect 3360 1680 3440 1688
rect 5760 1752 5840 2320
rect 6960 2232 7040 4480
rect 7120 2320 9280 4480
rect 6960 2168 6968 2232
rect 7032 2168 7040 2232
rect 6960 2160 7040 2168
rect 5760 1688 5768 1752
rect 5832 1688 5840 1752
rect 5760 1680 5840 1688
rect 8160 1752 8240 2320
rect 9360 2232 9440 4480
rect 9520 2320 11680 4480
rect 9360 2168 9368 2232
rect 9432 2168 9440 2232
rect 9360 2160 9440 2168
rect 8160 1688 8168 1752
rect 8232 1688 8240 1752
rect 8160 1680 8240 1688
rect 10560 1752 10640 2320
rect 11760 2232 11840 4480
rect 11920 2320 14080 4480
rect 11760 2168 11768 2232
rect 11832 2168 11840 2232
rect 11760 2160 11840 2168
rect 10560 1688 10568 1752
rect 10632 1688 10640 1752
rect 10560 1680 10640 1688
rect 12960 1752 13040 2320
rect 14160 2232 14240 4480
rect 14160 2168 14168 2232
rect 14232 2168 14240 2232
rect 14160 2160 14240 2168
rect 14320 2320 14720 4480
rect 14320 2232 14400 2320
rect 14320 2168 14328 2232
rect 14392 2168 14400 2232
rect 12960 1688 12968 1752
rect 13032 1688 13040 1752
rect 12960 1680 13040 1688
rect 14320 1912 14400 2168
rect 14320 1848 14328 1912
rect 14392 1848 14400 1912
rect -12400 1528 -12392 1592
rect -12328 1528 -12320 1592
rect -12400 1520 -12320 1528
rect 14320 1592 14400 1848
rect 14320 1528 14328 1592
rect 14392 1528 14400 1592
rect 14320 1520 14400 1528
rect 14480 2232 14560 2320
rect 14480 2168 14488 2232
rect 14552 2168 14560 2232
rect 14480 1912 14560 2168
rect 14480 1848 14488 1912
rect 14552 1848 14560 1912
rect 14480 1592 14560 1848
rect 14480 1528 14488 1592
rect 14552 1528 14560 1592
rect 14480 1520 14560 1528
rect 14640 2232 14720 2320
rect 14640 2168 14648 2232
rect 14712 2168 14720 2232
rect 14640 1912 14720 2168
rect 14640 1848 14648 1912
rect 14712 1848 14720 1912
rect 14640 1592 14720 1848
rect 14640 1528 14648 1592
rect 14712 1528 14720 1592
rect 14640 1520 14720 1528
<< via3 >>
rect -12712 7608 -12648 7672
rect -12712 7288 -12648 7352
rect -12712 6968 -12648 7032
rect -12552 7608 -12488 7672
rect -12552 7288 -12488 7352
rect -12552 6968 -12488 7032
rect -12392 7608 -12328 7672
rect 14328 7608 14392 7672
rect -12392 7288 -12328 7352
rect -11032 7448 -10968 7512
rect -12392 6968 -12328 7032
rect -12232 6968 -12168 7032
rect -8632 7448 -8568 7512
rect -9832 6968 -9768 7032
rect -6232 7448 -6168 7512
rect -7432 6968 -7368 7032
rect -3832 7448 -3768 7512
rect -5032 6968 -4968 7032
rect -1432 7448 -1368 7512
rect -2632 6968 -2568 7032
rect 3368 7448 3432 7512
rect 968 7128 1032 7192
rect -232 6968 -168 7032
rect 2168 6968 2232 7032
rect 5768 7448 5832 7512
rect 4568 6968 4632 7032
rect 8168 7448 8232 7512
rect 6968 6968 7032 7032
rect 10568 7448 10632 7512
rect 9368 6968 9432 7032
rect 12968 7448 13032 7512
rect 11768 6968 11832 7032
rect 14328 7288 14392 7352
rect 14168 6968 14232 7032
rect 14328 6968 14392 7032
rect 14488 7608 14552 7672
rect 14488 7288 14552 7352
rect 14488 6968 14552 7032
rect 14648 7608 14712 7672
rect 14648 7288 14712 7352
rect 14648 6968 14712 7032
rect -12712 2168 -12648 2232
rect -12712 1848 -12648 1912
rect -12712 1528 -12648 1592
rect -12552 2168 -12488 2232
rect -12552 1848 -12488 1912
rect -12552 1528 -12488 1592
rect -12392 2168 -12328 2232
rect -12232 2168 -12168 2232
rect -12392 1848 -12328 1912
rect -9832 2168 -9768 2232
rect -11032 1688 -10968 1752
rect -7432 2168 -7368 2232
rect -8632 1688 -8568 1752
rect -5032 2168 -4968 2232
rect -6232 1688 -6168 1752
rect -2632 2168 -2568 2232
rect -3832 1688 -3768 1752
rect -232 2168 -168 2232
rect 2168 2168 2232 2232
rect 968 2008 1032 2072
rect -1432 1688 -1368 1752
rect 4568 2168 4632 2232
rect 3368 1688 3432 1752
rect 6968 2168 7032 2232
rect 5768 1688 5832 1752
rect 9368 2168 9432 2232
rect 8168 1688 8232 1752
rect 11768 2168 11832 2232
rect 10568 1688 10632 1752
rect 14168 2168 14232 2232
rect 14328 2168 14392 2232
rect 12968 1688 13032 1752
rect 14328 1848 14392 1912
rect -12392 1528 -12328 1592
rect 14328 1528 14392 1592
rect 14488 2168 14552 2232
rect 14488 1848 14552 1912
rect 14488 1528 14552 1592
rect 14648 2168 14712 2232
rect 14648 1848 14712 1912
rect 14648 1528 14712 1592
<< mimcap >>
rect -12640 6712 -12400 6800
rect -12640 4888 -12552 6712
rect -12488 4888 -12400 6712
rect -12640 4800 -12400 4888
rect -12000 6712 -10000 6800
rect -12000 4888 -11912 6712
rect -10088 4888 -10000 6712
rect -12000 4800 -10000 4888
rect -9600 6712 -7600 6800
rect -9600 4888 -9512 6712
rect -7688 4888 -7600 6712
rect -9600 4800 -7600 4888
rect -7200 6712 -5200 6800
rect -7200 4888 -7112 6712
rect -5288 4888 -5200 6712
rect -7200 4800 -5200 4888
rect -4800 6712 -2800 6800
rect -4800 4888 -4712 6712
rect -2888 4888 -2800 6712
rect -4800 4800 -2800 4888
rect -2400 6712 -400 6800
rect -2400 4888 -2312 6712
rect -488 4888 -400 6712
rect -2400 4800 -400 4888
rect 0 6712 2000 6800
rect 0 4888 88 6712
rect 1912 4888 2000 6712
rect 0 4800 2000 4888
rect 2400 6712 4400 6800
rect 2400 4888 2488 6712
rect 4312 4888 4400 6712
rect 2400 4800 4400 4888
rect 4800 6712 6800 6800
rect 4800 4888 4888 6712
rect 6712 4888 6800 6712
rect 4800 4800 6800 4888
rect 7200 6712 9200 6800
rect 7200 4888 7288 6712
rect 9112 4888 9200 6712
rect 7200 4800 9200 4888
rect 9600 6712 11600 6800
rect 9600 4888 9688 6712
rect 11512 4888 11600 6712
rect 9600 4800 11600 4888
rect 12000 6712 14000 6800
rect 12000 4888 12088 6712
rect 13912 4888 14000 6712
rect 12000 4800 14000 4888
rect 14400 6712 14640 6800
rect 14400 4888 14488 6712
rect 14552 4888 14640 6712
rect 14400 4800 14640 4888
rect -12640 4312 -12400 4400
rect -12640 2488 -12552 4312
rect -12488 2488 -12400 4312
rect -12640 2400 -12400 2488
rect -12000 4312 -10000 4400
rect -12000 2488 -11912 4312
rect -10088 2488 -10000 4312
rect -12000 2400 -10000 2488
rect -9600 4312 -7600 4400
rect -9600 2488 -9512 4312
rect -7688 2488 -7600 4312
rect -9600 2400 -7600 2488
rect -7200 4312 -5200 4400
rect -7200 2488 -7112 4312
rect -5288 2488 -5200 4312
rect -7200 2400 -5200 2488
rect -4800 4312 -2800 4400
rect -4800 2488 -4712 4312
rect -2888 2488 -2800 4312
rect -4800 2400 -2800 2488
rect -2400 4312 -400 4400
rect -2400 2488 -2312 4312
rect -488 2488 -400 4312
rect -2400 2400 -400 2488
rect 0 4312 2000 4400
rect 0 2488 88 4312
rect 1912 2488 2000 4312
rect 0 2400 2000 2488
rect 2400 4312 4400 4400
rect 2400 2488 2488 4312
rect 4312 2488 4400 4312
rect 2400 2400 4400 2488
rect 4800 4312 6800 4400
rect 4800 2488 4888 4312
rect 6712 2488 6800 4312
rect 4800 2400 6800 2488
rect 7200 4312 9200 4400
rect 7200 2488 7288 4312
rect 9112 2488 9200 4312
rect 7200 2400 9200 2488
rect 9600 4312 11600 4400
rect 9600 2488 9688 4312
rect 11512 2488 11600 4312
rect 9600 2400 11600 2488
rect 12000 4312 14000 4400
rect 12000 2488 12088 4312
rect 13912 2488 14000 4312
rect 12000 2400 14000 2488
rect 14400 4312 14640 4400
rect 14400 2488 14488 4312
rect 14552 2488 14640 4312
rect 14400 2400 14640 2488
<< mimcapcontact >>
rect -12552 4888 -12488 6712
rect -11912 4888 -10088 6712
rect -9512 4888 -7688 6712
rect -7112 4888 -5288 6712
rect -4712 4888 -2888 6712
rect -2312 4888 -488 6712
rect 88 4888 1912 6712
rect 2488 4888 4312 6712
rect 4888 4888 6712 6712
rect 7288 4888 9112 6712
rect 9688 4888 11512 6712
rect 12088 4888 13912 6712
rect 14488 4888 14552 6712
rect -12552 2488 -12488 4312
rect -11912 2488 -10088 4312
rect -9512 2488 -7688 4312
rect -7112 2488 -5288 4312
rect -4712 2488 -2888 4312
rect -2312 2488 -488 4312
rect 88 2488 1912 4312
rect 2488 2488 4312 4312
rect 4888 2488 6712 4312
rect 7288 2488 9112 4312
rect 9688 2488 11512 4312
rect 12088 2488 13912 4312
rect 14488 2488 14552 4312
<< metal4 >>
rect -12720 7672 14880 7680
rect -12720 7608 -12712 7672
rect -12648 7608 -12552 7672
rect -12488 7608 -12392 7672
rect -12328 7608 14328 7672
rect 14392 7608 14488 7672
rect 14552 7608 14648 7672
rect 14712 7608 14880 7672
rect -12720 7600 14880 7608
rect -12720 7512 14880 7520
rect -12720 7448 -11032 7512
rect -10968 7448 -8632 7512
rect -8568 7448 -6232 7512
rect -6168 7448 -3832 7512
rect -3768 7448 -1432 7512
rect -1368 7448 3368 7512
rect 3432 7448 5768 7512
rect 5832 7448 8168 7512
rect 8232 7448 10568 7512
rect 10632 7448 12968 7512
rect 13032 7448 14880 7512
rect -12720 7440 14880 7448
rect -12720 7352 14880 7360
rect -12720 7288 -12712 7352
rect -12648 7288 -12552 7352
rect -12488 7288 -12392 7352
rect -12328 7288 14328 7352
rect 14392 7288 14488 7352
rect 14552 7288 14648 7352
rect 14712 7288 14880 7352
rect -12720 7280 14880 7288
rect -12720 7192 14880 7200
rect -12720 7128 968 7192
rect 1032 7128 14880 7192
rect -12720 7120 14880 7128
rect -12720 7032 14880 7040
rect -12720 6968 -12712 7032
rect -12648 6968 -12552 7032
rect -12488 6968 -12392 7032
rect -12328 6968 -12232 7032
rect -12168 6968 -9832 7032
rect -9768 6968 -7432 7032
rect -7368 6968 -5032 7032
rect -4968 6968 -2632 7032
rect -2568 6968 -232 7032
rect -168 6968 2168 7032
rect 2232 6968 4568 7032
rect 4632 6968 6968 7032
rect 7032 6968 9368 7032
rect 9432 6968 11768 7032
rect 11832 6968 14168 7032
rect 14232 6968 14328 7032
rect 14392 6968 14488 7032
rect 14552 6968 14648 7032
rect 14712 6968 14880 7032
rect -12720 6960 14880 6968
rect -12720 6880 -12640 6960
rect -12560 6880 -12480 6960
rect -12400 6880 -12320 6960
rect -12720 6712 -12320 6880
rect -12720 4888 -12552 6712
rect -12488 4888 -12320 6712
rect -12720 4720 -12320 4888
rect -12240 4720 -12160 6960
rect -12080 6712 -9920 6880
rect -12080 4888 -11912 6712
rect -10088 4888 -9920 6712
rect -12080 4720 -9920 4888
rect -9840 4720 -9760 6960
rect -9680 6712 -7520 6880
rect -9680 4888 -9512 6712
rect -7688 4888 -7520 6712
rect -9680 4720 -7520 4888
rect -7440 4720 -7360 6960
rect -7280 6712 -5120 6880
rect -7280 4888 -7112 6712
rect -5288 4888 -5120 6712
rect -7280 4720 -5120 4888
rect -5040 4720 -4960 6960
rect -4880 6712 -2720 6880
rect -4880 4888 -4712 6712
rect -2888 4888 -2720 6712
rect -4880 4720 -2720 4888
rect -2640 4720 -2560 6960
rect -2480 6712 -320 6880
rect -2480 4888 -2312 6712
rect -488 4888 -320 6712
rect -2480 4720 -320 4888
rect -240 4720 -160 6960
rect -80 6712 2080 6880
rect -80 4888 88 6712
rect 1912 4888 2080 6712
rect -80 4720 2080 4888
rect 2160 4720 2240 6960
rect 2320 6712 4480 6880
rect 2320 4888 2488 6712
rect 4312 4888 4480 6712
rect 2320 4720 4480 4888
rect 4560 4720 4640 6960
rect 4720 6712 6880 6880
rect 4720 4888 4888 6712
rect 6712 4888 6880 6712
rect 4720 4720 6880 4888
rect 6960 4720 7040 6960
rect 7120 6712 9280 6880
rect 7120 4888 7288 6712
rect 9112 4888 9280 6712
rect 7120 4720 9280 4888
rect 9360 4720 9440 6960
rect 9520 6712 11680 6880
rect 9520 4888 9688 6712
rect 11512 4888 11680 6712
rect 9520 4720 11680 4888
rect 11760 4720 11840 6960
rect 11920 6712 14080 6880
rect 11920 4888 12088 6712
rect 13912 4888 14080 6712
rect 11920 4720 14080 4888
rect 14160 4720 14240 6960
rect 14320 6880 14400 6960
rect 14480 6880 14560 6960
rect 14640 6880 14720 6960
rect 14320 6712 14720 6880
rect 14320 4888 14488 6712
rect 14552 4888 14720 6712
rect 14320 4720 14720 4888
rect -12080 4640 -12000 4720
rect -11920 4640 -11840 4720
rect -11760 4640 -11680 4720
rect -11600 4640 -11520 4720
rect -11440 4640 -11360 4720
rect -11280 4640 -11200 4720
rect -11120 4640 -11040 4720
rect -10960 4640 -10880 4720
rect -10800 4640 -10720 4720
rect -10640 4640 -10560 4720
rect -10480 4640 -10400 4720
rect -10320 4640 -10240 4720
rect -10160 4640 -10080 4720
rect -10000 4640 -9920 4720
rect -9680 4640 -9600 4720
rect -9520 4640 -9440 4720
rect -9360 4640 -9280 4720
rect -9200 4640 -9120 4720
rect -9040 4640 -8960 4720
rect -8880 4640 -8800 4720
rect -8720 4640 -8640 4720
rect -8560 4640 -8480 4720
rect -8400 4640 -8320 4720
rect -8240 4640 -8160 4720
rect -8080 4640 -8000 4720
rect -7920 4640 -7840 4720
rect -7760 4640 -7680 4720
rect -7600 4640 -7520 4720
rect -7280 4640 -7200 4720
rect -7120 4640 -7040 4720
rect -6960 4640 -6880 4720
rect -6800 4640 -6720 4720
rect -6640 4640 -6560 4720
rect -6480 4640 -6400 4720
rect -6320 4640 -6240 4720
rect -6160 4640 -6080 4720
rect -6000 4640 -5920 4720
rect -5840 4640 -5760 4720
rect -5680 4640 -5600 4720
rect -5520 4640 -5440 4720
rect -5360 4640 -5280 4720
rect -5200 4640 -5120 4720
rect -4880 4640 -4800 4720
rect -4720 4640 -4640 4720
rect -4560 4640 -4480 4720
rect -4400 4640 -4320 4720
rect -4240 4640 -4160 4720
rect -4080 4640 -4000 4720
rect -3920 4640 -3840 4720
rect -3760 4640 -3680 4720
rect -3600 4640 -3520 4720
rect -3440 4640 -3360 4720
rect -3280 4640 -3200 4720
rect -3120 4640 -3040 4720
rect -2960 4640 -2880 4720
rect -2800 4640 -2720 4720
rect -2480 4640 -2400 4720
rect -2320 4640 -2240 4720
rect -2160 4640 -2080 4720
rect -2000 4640 -1920 4720
rect -1840 4640 -1760 4720
rect -1680 4640 -1600 4720
rect -1520 4640 -1440 4720
rect -1360 4640 -1280 4720
rect -1200 4640 -1120 4720
rect -1040 4640 -960 4720
rect -880 4640 -800 4720
rect -720 4640 -640 4720
rect -560 4640 -480 4720
rect -400 4640 -320 4720
rect -80 4640 0 4720
rect 80 4640 160 4720
rect 240 4640 320 4720
rect 400 4640 480 4720
rect 560 4640 640 4720
rect 720 4640 800 4720
rect 880 4640 960 4720
rect 1040 4640 1120 4720
rect 1200 4640 1280 4720
rect 1360 4640 1440 4720
rect 1520 4640 1600 4720
rect 1680 4640 1760 4720
rect 1840 4640 1920 4720
rect 2000 4640 2080 4720
rect 2320 4640 2400 4720
rect 2480 4640 2560 4720
rect 2640 4640 2720 4720
rect 2800 4640 2880 4720
rect 2960 4640 3040 4720
rect 3120 4640 3200 4720
rect 3280 4640 3360 4720
rect 3440 4640 3520 4720
rect 3600 4640 3680 4720
rect 3760 4640 3840 4720
rect 3920 4640 4000 4720
rect 4080 4640 4160 4720
rect 4240 4640 4320 4720
rect 4400 4640 4480 4720
rect 4720 4640 4800 4720
rect 4880 4640 4960 4720
rect 5040 4640 5120 4720
rect 5200 4640 5280 4720
rect 5360 4640 5440 4720
rect 5520 4640 5600 4720
rect 5680 4640 5760 4720
rect 5840 4640 5920 4720
rect 6000 4640 6080 4720
rect 6160 4640 6240 4720
rect 6320 4640 6400 4720
rect 6480 4640 6560 4720
rect 6640 4640 6720 4720
rect 6800 4640 6880 4720
rect 7120 4640 7200 4720
rect 7280 4640 7360 4720
rect 7440 4640 7520 4720
rect 7600 4640 7680 4720
rect 7760 4640 7840 4720
rect 7920 4640 8000 4720
rect 8080 4640 8160 4720
rect 8240 4640 8320 4720
rect 8400 4640 8480 4720
rect 8560 4640 8640 4720
rect 8720 4640 8800 4720
rect 8880 4640 8960 4720
rect 9040 4640 9120 4720
rect 9200 4640 9280 4720
rect 9520 4640 9600 4720
rect 9680 4640 9760 4720
rect 9840 4640 9920 4720
rect 10000 4640 10080 4720
rect 10160 4640 10240 4720
rect 10320 4640 10400 4720
rect 10480 4640 10560 4720
rect 10640 4640 10720 4720
rect 10800 4640 10880 4720
rect 10960 4640 11040 4720
rect 11120 4640 11200 4720
rect 11280 4640 11360 4720
rect 11440 4640 11520 4720
rect 11600 4640 11680 4720
rect 11920 4640 12000 4720
rect 12080 4640 12160 4720
rect 12240 4640 12320 4720
rect 12400 4640 12480 4720
rect 12560 4640 12640 4720
rect 12720 4640 12800 4720
rect 12880 4640 12960 4720
rect 13040 4640 13120 4720
rect 13200 4640 13280 4720
rect 13360 4640 13440 4720
rect 13520 4640 13600 4720
rect 13680 4640 13760 4720
rect 13840 4640 13920 4720
rect 14000 4640 14080 4720
rect -12800 4560 14880 4640
rect -12080 4480 -12000 4560
rect -11920 4480 -11840 4560
rect -11760 4480 -11680 4560
rect -11600 4480 -11520 4560
rect -11440 4480 -11360 4560
rect -11280 4480 -11200 4560
rect -11120 4480 -11040 4560
rect -10960 4480 -10880 4560
rect -10800 4480 -10720 4560
rect -10640 4480 -10560 4560
rect -10480 4480 -10400 4560
rect -10320 4480 -10240 4560
rect -10160 4480 -10080 4560
rect -10000 4480 -9920 4560
rect -9680 4480 -9600 4560
rect -9520 4480 -9440 4560
rect -9360 4480 -9280 4560
rect -9200 4480 -9120 4560
rect -9040 4480 -8960 4560
rect -8880 4480 -8800 4560
rect -8720 4480 -8640 4560
rect -8560 4480 -8480 4560
rect -8400 4480 -8320 4560
rect -8240 4480 -8160 4560
rect -8080 4480 -8000 4560
rect -7920 4480 -7840 4560
rect -7760 4480 -7680 4560
rect -7600 4480 -7520 4560
rect -7280 4480 -7200 4560
rect -7120 4480 -7040 4560
rect -6960 4480 -6880 4560
rect -6800 4480 -6720 4560
rect -6640 4480 -6560 4560
rect -6480 4480 -6400 4560
rect -6320 4480 -6240 4560
rect -6160 4480 -6080 4560
rect -6000 4480 -5920 4560
rect -5840 4480 -5760 4560
rect -5680 4480 -5600 4560
rect -5520 4480 -5440 4560
rect -5360 4480 -5280 4560
rect -5200 4480 -5120 4560
rect -4880 4480 -4800 4560
rect -4720 4480 -4640 4560
rect -4560 4480 -4480 4560
rect -4400 4480 -4320 4560
rect -4240 4480 -4160 4560
rect -4080 4480 -4000 4560
rect -3920 4480 -3840 4560
rect -3760 4480 -3680 4560
rect -3600 4480 -3520 4560
rect -3440 4480 -3360 4560
rect -3280 4480 -3200 4560
rect -3120 4480 -3040 4560
rect -2960 4480 -2880 4560
rect -2800 4480 -2720 4560
rect -2480 4480 -2400 4560
rect -2320 4480 -2240 4560
rect -2160 4480 -2080 4560
rect -2000 4480 -1920 4560
rect -1840 4480 -1760 4560
rect -1680 4480 -1600 4560
rect -1520 4480 -1440 4560
rect -1360 4480 -1280 4560
rect -1200 4480 -1120 4560
rect -1040 4480 -960 4560
rect -880 4480 -800 4560
rect -720 4480 -640 4560
rect -560 4480 -480 4560
rect -400 4480 -320 4560
rect -80 4480 0 4560
rect 80 4480 160 4560
rect 240 4480 320 4560
rect 400 4480 480 4560
rect 560 4480 640 4560
rect 720 4480 800 4560
rect 880 4480 960 4560
rect 1040 4480 1120 4560
rect 1200 4480 1280 4560
rect 1360 4480 1440 4560
rect 1520 4480 1600 4560
rect 1680 4480 1760 4560
rect 1840 4480 1920 4560
rect 2000 4480 2080 4560
rect 2320 4480 2400 4560
rect 2480 4480 2560 4560
rect 2640 4480 2720 4560
rect 2800 4480 2880 4560
rect 2960 4480 3040 4560
rect 3120 4480 3200 4560
rect 3280 4480 3360 4560
rect 3440 4480 3520 4560
rect 3600 4480 3680 4560
rect 3760 4480 3840 4560
rect 3920 4480 4000 4560
rect 4080 4480 4160 4560
rect 4240 4480 4320 4560
rect 4400 4480 4480 4560
rect 4720 4480 4800 4560
rect 4880 4480 4960 4560
rect 5040 4480 5120 4560
rect 5200 4480 5280 4560
rect 5360 4480 5440 4560
rect 5520 4480 5600 4560
rect 5680 4480 5760 4560
rect 5840 4480 5920 4560
rect 6000 4480 6080 4560
rect 6160 4480 6240 4560
rect 6320 4480 6400 4560
rect 6480 4480 6560 4560
rect 6640 4480 6720 4560
rect 6800 4480 6880 4560
rect 7120 4480 7200 4560
rect 7280 4480 7360 4560
rect 7440 4480 7520 4560
rect 7600 4480 7680 4560
rect 7760 4480 7840 4560
rect 7920 4480 8000 4560
rect 8080 4480 8160 4560
rect 8240 4480 8320 4560
rect 8400 4480 8480 4560
rect 8560 4480 8640 4560
rect 8720 4480 8800 4560
rect 8880 4480 8960 4560
rect 9040 4480 9120 4560
rect 9200 4480 9280 4560
rect 9520 4480 9600 4560
rect 9680 4480 9760 4560
rect 9840 4480 9920 4560
rect 10000 4480 10080 4560
rect 10160 4480 10240 4560
rect 10320 4480 10400 4560
rect 10480 4480 10560 4560
rect 10640 4480 10720 4560
rect 10800 4480 10880 4560
rect 10960 4480 11040 4560
rect 11120 4480 11200 4560
rect 11280 4480 11360 4560
rect 11440 4480 11520 4560
rect 11600 4480 11680 4560
rect 11920 4480 12000 4560
rect 12080 4480 12160 4560
rect 12240 4480 12320 4560
rect 12400 4480 12480 4560
rect 12560 4480 12640 4560
rect 12720 4480 12800 4560
rect 12880 4480 12960 4560
rect 13040 4480 13120 4560
rect 13200 4480 13280 4560
rect 13360 4480 13440 4560
rect 13520 4480 13600 4560
rect 13680 4480 13760 4560
rect 13840 4480 13920 4560
rect 14000 4480 14080 4560
rect -12720 4312 -12320 4480
rect -12720 2488 -12552 4312
rect -12488 2488 -12320 4312
rect -12720 2320 -12320 2488
rect -12720 2240 -12640 2320
rect -12560 2240 -12480 2320
rect -12400 2240 -12320 2320
rect -12240 2240 -12160 4480
rect -12080 4312 -9920 4480
rect -12080 2488 -11912 4312
rect -10088 2488 -9920 4312
rect -12080 2320 -9920 2488
rect -9840 2240 -9760 4480
rect -9680 4312 -7520 4480
rect -9680 2488 -9512 4312
rect -7688 2488 -7520 4312
rect -9680 2320 -7520 2488
rect -7440 2240 -7360 4480
rect -7280 4312 -5120 4480
rect -7280 2488 -7112 4312
rect -5288 2488 -5120 4312
rect -7280 2320 -5120 2488
rect -5040 2240 -4960 4480
rect -4880 4312 -2720 4480
rect -4880 2488 -4712 4312
rect -2888 2488 -2720 4312
rect -4880 2320 -2720 2488
rect -2640 2240 -2560 4480
rect -2480 4312 -320 4480
rect -2480 2488 -2312 4312
rect -488 2488 -320 4312
rect -2480 2320 -320 2488
rect -240 2240 -160 4480
rect -80 4312 2080 4480
rect -80 2488 88 4312
rect 1912 2488 2080 4312
rect -80 2320 2080 2488
rect 2160 2240 2240 4480
rect 2320 4312 4480 4480
rect 2320 2488 2488 4312
rect 4312 2488 4480 4312
rect 2320 2320 4480 2488
rect 4560 2240 4640 4480
rect 4720 4312 6880 4480
rect 4720 2488 4888 4312
rect 6712 2488 6880 4312
rect 4720 2320 6880 2488
rect 6960 2240 7040 4480
rect 7120 4312 9280 4480
rect 7120 2488 7288 4312
rect 9112 2488 9280 4312
rect 7120 2320 9280 2488
rect 9360 2240 9440 4480
rect 9520 4312 11680 4480
rect 9520 2488 9688 4312
rect 11512 2488 11680 4312
rect 9520 2320 11680 2488
rect 11760 2240 11840 4480
rect 11920 4312 14080 4480
rect 11920 2488 12088 4312
rect 13912 2488 14080 4312
rect 11920 2320 14080 2488
rect 14160 2240 14240 4480
rect 14320 4312 14720 4480
rect 14320 2488 14488 4312
rect 14552 2488 14720 4312
rect 14320 2320 14720 2488
rect 14320 2240 14400 2320
rect 14480 2240 14560 2320
rect 14640 2240 14720 2320
rect -12800 2232 14880 2240
rect -12800 2168 -12712 2232
rect -12648 2168 -12552 2232
rect -12488 2168 -12392 2232
rect -12328 2168 -12232 2232
rect -12168 2168 -9832 2232
rect -9768 2168 -7432 2232
rect -7368 2168 -5032 2232
rect -4968 2168 -2632 2232
rect -2568 2168 -232 2232
rect -168 2168 2168 2232
rect 2232 2168 4568 2232
rect 4632 2168 6968 2232
rect 7032 2168 9368 2232
rect 9432 2168 11768 2232
rect 11832 2168 14168 2232
rect 14232 2168 14328 2232
rect 14392 2168 14488 2232
rect 14552 2168 14648 2232
rect 14712 2168 14880 2232
rect -12800 2160 14880 2168
rect -12800 2072 14880 2080
rect -12800 2008 968 2072
rect 1032 2008 14880 2072
rect -12800 2000 14880 2008
rect -12800 1912 14880 1920
rect -12800 1848 -12712 1912
rect -12648 1848 -12552 1912
rect -12488 1848 -12392 1912
rect -12328 1848 14328 1912
rect 14392 1848 14488 1912
rect 14552 1848 14648 1912
rect 14712 1848 14880 1912
rect -12800 1840 14880 1848
rect -12800 1752 14880 1760
rect -12800 1688 -11032 1752
rect -10968 1688 -8632 1752
rect -8568 1688 -6232 1752
rect -6168 1688 -3832 1752
rect -3768 1688 -1432 1752
rect -1368 1688 3368 1752
rect 3432 1688 5768 1752
rect 5832 1688 8168 1752
rect 8232 1688 10568 1752
rect 10632 1688 12968 1752
rect 13032 1688 14880 1752
rect -12800 1680 14880 1688
rect -12800 1592 14880 1600
rect -12800 1528 -12712 1592
rect -12648 1528 -12552 1592
rect -12488 1528 -12392 1592
rect -12328 1528 14328 1592
rect 14392 1528 14488 1592
rect 14552 1528 14648 1592
rect 14712 1528 14880 1592
rect -12800 1520 14880 1528
<< labels >>
rlabel metal4 s 14800 4560 14880 4640 4 a
port 1 nsew
rlabel metal4 s 14800 7120 14880 7200 4 b1
port 2 nsew
rlabel metal4 s 14800 2000 14880 2080 4 b2
port 3 nsew
rlabel metal4 s 14800 7440 14880 7520 4 c1
port 4 nsew
rlabel metal4 s 14800 1680 14880 1760 4 c2
port 5 nsew
rlabel metal4 s 14800 7280 14880 7360 4 gnda
port 6 nsew
rlabel locali s 14800 1360 14880 1440 4 vssa
port 7 nsew
<< end >>
