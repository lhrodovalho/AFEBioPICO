* NGSPICE file created from opamp_coreb.ext - technology: sky130A

.subckt opamp_coreb gpa dpa gpb gn xn vdda vssa
X0 dpb gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X1 dpb gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X2 n2 gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X3 xp gpa p5 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X4 dpb gpb dpa dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.875e+12p pd=4.625e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X5 dpb gpb dpa dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.875e+12p pd=4.625e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X6 dpb gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X7 n7 gn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.5e+11p ps=2.55e+06u w=1e+06u l=2e+06u
X8 xp gpa dpa vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X9 dpa gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X10 xn gn dpb vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X11 vdda gpa p8 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.95e+12p pd=5.05e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X12 dpa gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X13 dpa gpb dpb dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.875e+12p ps=4.625e+06u w=3e+06u l=2e+06u
X14 xn gn n7 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X15 p7 gpa vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.95e+12p ps=5.05e+06u w=3e+06u l=2e+06u
X16 xn gn dpb vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X17 xn gn n5 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X18 dpa gpb dpb dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.875e+12p ps=4.625e+06u w=3e+06u l=2e+06u
X19 dpa gpb dpb dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.875e+12p ps=4.625e+06u w=3e+06u l=2e+06u
X20 p1 gpa vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.95e+12p ps=5.05e+06u w=3e+06u l=2e+06u
X21 xp gpa dpa vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X22 dpa gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X23 dpb gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X24 xn gn dpb vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X25 n6 gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X26 dpb gpb dpa dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.875e+12p pd=4.625e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X27 dpb gpb dpa dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.875e+12p pd=4.625e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X28 dpb gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X29 n1 gn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.5e+11p ps=2.55e+06u w=1e+06u l=2e+06u
X30 n4 gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X31 xp gpa p3 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X32 dpa gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X33 xp gpa dpa vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X34 p2 gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X35 p8 gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X36 dpb gpb dpa dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.875e+12p pd=4.625e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X37 xp gpa dpa vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X38 dpa gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X39 dpb gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X40 vssa gn n2 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.5e+11p pd=2.55e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X41 vssa gn n6 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.5e+11p pd=2.55e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X42 p5 gpa vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.95e+12p ps=5.05e+06u w=3e+06u l=2e+06u
X43 xp gpa dpa vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X44 dpa gpb dpb dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.875e+12p ps=4.625e+06u w=3e+06u l=2e+06u
X45 xp gpa p1 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X46 dpa gpb dpb dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.875e+12p ps=4.625e+06u w=3e+06u l=2e+06u
X47 xn gn dpb vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X48 vssa gn n4 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.5e+11p pd=2.55e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X49 xn gn dpb vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X50 dpa gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X51 xp gpa dpa vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X52 dpb gpb dpa dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.875e+12p pd=4.625e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X53 dpa gpb dpb dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.875e+12p ps=4.625e+06u w=3e+06u l=2e+06u
X54 n5 gn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.5e+11p ps=2.55e+06u w=1e+06u l=2e+06u
X55 p3 gpa vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.95e+12p ps=5.05e+06u w=3e+06u l=2e+06u
X56 vdda gpa p6 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.95e+12p pd=5.05e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X57 dpb gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X58 n3 gn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.5e+11p ps=2.55e+06u w=1e+06u l=2e+06u
X59 dpb gpb dpa dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.875e+12p pd=4.625e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X60 dpb gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X61 n8 gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X62 vdda gpa p2 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.95e+12p pd=5.05e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X63 p6 gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X64 xp gpa dpa vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X65 xn gn n3 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X66 vdda gpa p4 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.95e+12p pd=5.05e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X67 xn gn dpb vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X68 vssa gn n8 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.5e+11p pd=2.55e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X69 dpb gpb dpa dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.875e+12p pd=4.625e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X70 xn gn dpb vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X71 p4 gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X72 xp gpa dpa vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X73 dpa gpb dpb dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.875e+12p ps=4.625e+06u w=3e+06u l=2e+06u
X74 xn gn dpb vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X75 xp gpa p7 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X76 dpa gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X77 dpa gpb dpb dpa sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.875e+12p ps=4.625e+06u w=3e+06u l=2e+06u
X78 dpa gpa xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X79 xn gn n1 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
.ends

