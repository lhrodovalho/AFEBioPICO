* operational amplifier buffer testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "../mag/ota.spice"

* supply voltages
vdda vdda 0 1.8
vssa vssa 0 0.0
egnda gnda vssa vdda vssa 0.5

* input signals
vin in gnda dc 0 ac 1 SINE(0 0.4 1 0 0 0)
IB ib vss 5n


* DUT
Xdut out in out ib vdda gnda vssa ota
CL out gnda 1p

.save v(in) v(out) v(ib) v(Xdut.x) i(vdda)
.option gmin=1e-15
.control

	op
	print ib i(vdda)
	
	ac dec 10 1m 1Meg
	wrdata ../data/ota_tb_buf_ac.txt vdb(out) phase(out)*180/PI
	plot vdb(out)
	plot phase(out)*180/PI
		
	tran 10m 5 1
	wrdata ../data/ota_tb_buf_tran.txt v(in) v(out) i(vdda)
	plot v(in) v(out)

.endc

.end
