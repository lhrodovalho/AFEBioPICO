magic
tech sky130A
timestamp 1634680784
<< nwell >>
rect -2870 -3290 -2820 -460
rect 23500 -3290 23550 -460
rect -2870 -12540 -2820 -9710
rect 23500 -12540 23550 -9710
rect -2870 -15850 -2820 -13020
rect 23500 -15850 23550 -13020
rect -2870 -25100 -2820 -22270
rect 23500 -25100 23550 -22270
<< pwell >>
rect -2910 -440 -2820 -410
rect 23500 -440 23590 -410
rect -2920 -5150 -2810 -5120
rect 23500 -5150 23600 -5120
rect -2920 -6280 -2890 -5150
rect 23570 -6280 23600 -5150
rect -2920 -7850 -2890 -6720
rect 23570 -7850 23600 -6720
rect -2920 -7880 -2810 -7850
rect 23500 -7880 23600 -7850
rect -2910 -12590 -2820 -12560
rect 23500 -12590 23590 -12560
rect -2910 -13000 -2820 -12970
rect 23500 -13000 23590 -12970
rect -2920 -17710 -2810 -17680
rect 23500 -17710 23600 -17680
rect -2920 -18840 -2890 -17710
rect 23570 -18840 23600 -17710
rect -2920 -20410 -2890 -19280
rect 23570 -20410 23600 -19280
rect -2920 -20440 -2810 -20410
rect 23500 -20440 23600 -20410
rect -2910 -25150 -2820 -25120
rect 23500 -25150 23590 -25120
<< psubdiff >>
rect -2920 -440 -2820 -410
rect 23500 -440 23600 -410
rect -2920 -3310 -2890 -440
rect 23570 -3310 23600 -440
rect -2920 -3340 -1810 -3310
rect 10270 -3340 10410 -3310
rect 22490 -3340 23600 -3310
rect -2920 -5120 -2890 -3340
rect 23570 -5120 23600 -3340
rect -2920 -5150 -2810 -5120
rect 23500 -5150 23600 -5120
rect -2920 -6280 -2890 -5150
rect 23570 -6280 23600 -5150
rect -2920 -6310 23600 -6280
rect -2920 -6720 23600 -6690
rect -2920 -7850 -2890 -6720
rect 23570 -7850 23600 -6720
rect -2920 -7880 -2810 -7850
rect 23500 -7880 23600 -7850
rect -2920 -9660 -2890 -7880
rect 23570 -9660 23600 -7880
rect -2920 -9690 -1810 -9660
rect 10270 -9690 10410 -9660
rect 22490 -9690 23600 -9660
rect -2920 -12560 -2890 -9690
rect 23570 -12560 23600 -9690
rect -2920 -12590 -2820 -12560
rect 23500 -12590 23600 -12560
rect -2920 -13000 -2820 -12970
rect 23500 -13000 23600 -12970
rect -2920 -15870 -2890 -13000
rect 23570 -15870 23600 -13000
rect -2920 -15900 -1810 -15870
rect 10270 -15900 10410 -15870
rect 22490 -15900 23600 -15870
rect -2920 -17680 -2890 -15900
rect 23570 -17680 23600 -15900
rect -2920 -17710 -2810 -17680
rect 23500 -17710 23600 -17680
rect -2920 -18840 -2890 -17710
rect 23570 -18840 23600 -17710
rect -2920 -18870 23600 -18840
rect -2920 -19280 23600 -19250
rect -2920 -20410 -2890 -19280
rect 23570 -20410 23600 -19280
rect -2920 -20440 -2810 -20410
rect 23500 -20440 23600 -20410
rect -2920 -22220 -2890 -20440
rect 23570 -22220 23600 -20440
rect -2920 -22250 -1810 -22220
rect 10270 -22250 10410 -22220
rect 22490 -22250 23600 -22220
rect -2920 -25120 -2890 -22250
rect 23570 -25120 23600 -22250
rect -2920 -25150 -2820 -25120
rect 23500 -25150 23600 -25120
rect -2920 -25440 -2890 -25150
rect -2920 -25470 -2880 -25440
rect 21100 -25470 21130 -25440
rect -2920 -28490 -2890 -25470
rect -2920 -28520 -2880 -28490
rect 21100 -28520 21130 -28490
<< psubdiffcont >>
rect -1810 -3340 10270 -3310
rect 10410 -3340 22490 -3310
rect -1810 -9690 10270 -9660
rect 10410 -9690 22490 -9660
rect -1810 -15900 10270 -15870
rect 10410 -15900 22490 -15870
rect -1810 -22250 10270 -22220
rect 10410 -22250 22490 -22220
rect -2880 -25470 21100 -25440
rect -2880 -28520 21100 -28490
<< locali >>
rect -6280 -4120 -6110 -220
rect -6080 -4120 -5910 -220
rect -5880 -4120 -5710 -220
rect -5680 -4120 -5510 -220
rect -5480 -4120 -5310 -220
rect -5280 -4120 -5110 -220
rect -5080 -4120 -4710 -220
rect -4680 -4120 -4510 -220
rect -4480 -4120 -4310 -220
rect -4280 -4120 -4110 -220
rect -4080 -4120 -3910 -220
rect -3880 -4120 -3710 -220
rect -3680 -3400 -3510 -220
rect -2920 -440 -2820 -410
rect 23500 -440 23600 -410
rect -2920 -3310 -2890 -440
rect -1010 -480 -960 -470
rect -2850 -3270 -2820 -480
rect -1010 -510 -1000 -480
rect -970 -510 -960 -480
rect -1010 -520 -960 -510
rect 21640 -480 21690 -470
rect 21640 -510 21650 -480
rect 21680 -510 21690 -480
rect 21640 -520 21690 -510
rect 23500 -3270 23530 -480
rect 23570 -3310 23600 -440
rect -2920 -3340 -1850 -3310
rect -1820 -3340 -1810 -3310
rect 10270 -3340 10410 -3310
rect 22490 -3340 22500 -3310
rect 22530 -3340 23600 -3310
rect -3680 -3490 23560 -3400
rect -3680 -3520 -3510 -3490
rect -3680 -3610 23560 -3520
rect -3680 -3640 -3510 -3610
rect -3680 -3730 23560 -3640
rect -3680 -3760 -3510 -3730
rect -3680 -3850 23560 -3760
rect -3680 -3880 -3510 -3850
rect -3680 -3970 23560 -3880
rect -3680 -4000 -3510 -3970
rect -3680 -4090 23560 -4000
rect -3680 -4120 -3510 -4090
rect -6280 -4160 24420 -4120
rect -6280 -4300 24270 -4160
rect 24410 -4300 24420 -4160
rect -6280 -4340 24420 -4300
rect -6280 -8660 -6110 -4340
rect -6080 -8660 -5910 -4340
rect -5880 -8660 -5710 -4340
rect -5680 -8660 -5510 -4340
rect -5480 -8660 -5310 -4340
rect -5280 -8660 -5110 -4340
rect -5080 -8660 -4710 -4340
rect -4680 -8660 -4510 -4340
rect -4480 -8660 -4310 -4340
rect -4280 -8660 -4110 -4340
rect -4080 -8660 -3910 -4340
rect -3880 -8660 -3710 -4340
rect -3680 -4370 -3510 -4340
rect -3680 -4460 23560 -4370
rect -3680 -4490 -3510 -4460
rect -3680 -4580 23560 -4490
rect -3680 -4610 -3510 -4580
rect -3680 -4700 23560 -4610
rect -3680 -4730 -3510 -4700
rect -3680 -4820 23560 -4730
rect -3680 -4850 -3510 -4820
rect -3680 -4940 23560 -4850
rect -3680 -4970 -3510 -4940
rect -3680 -5060 23560 -4970
rect -3680 -7940 -3510 -5060
rect -2920 -5150 -2810 -5120
rect 23500 -5150 23600 -5120
rect -2920 -6280 -2890 -5150
rect -1860 -6280 -1810 -6270
rect 22490 -6280 22540 -6270
rect 23570 -6280 23600 -5150
rect -2920 -6310 -1850 -6280
rect -1820 -6310 22500 -6280
rect 22530 -6310 23600 -6280
rect -1860 -6320 -1810 -6310
rect 22490 -6320 22540 -6310
rect -1860 -6690 -1810 -6680
rect 22490 -6690 22540 -6680
rect -2920 -6720 -1850 -6690
rect -1820 -6720 22500 -6690
rect 22530 -6720 23600 -6690
rect -2920 -7850 -2890 -6720
rect -1860 -6730 -1810 -6720
rect 22490 -6730 22540 -6720
rect 23570 -7850 23600 -6720
rect -2920 -7880 -2810 -7850
rect 23500 -7880 23600 -7850
rect -3680 -8030 23560 -7940
rect -3680 -8060 -3510 -8030
rect -3680 -8150 23560 -8060
rect -3680 -8180 -3510 -8150
rect -3680 -8270 23560 -8180
rect -3680 -8300 -3510 -8270
rect -3680 -8390 23560 -8300
rect -3680 -8420 -3510 -8390
rect -3680 -8510 23560 -8420
rect -3680 -8540 -3510 -8510
rect -3680 -8630 23560 -8540
rect -3680 -8660 -3510 -8630
rect -6280 -8700 24420 -8660
rect -6280 -8840 24270 -8700
rect 24410 -8840 24420 -8700
rect -6280 -8880 24420 -8840
rect -6280 -16680 -6110 -8880
rect -6080 -16680 -5910 -8880
rect -5880 -16680 -5710 -8880
rect -5680 -16680 -5510 -8880
rect -5480 -16680 -5310 -8880
rect -5280 -16680 -5110 -8880
rect -5080 -16680 -4710 -8880
rect -4680 -16680 -4510 -8880
rect -4480 -16680 -4310 -8880
rect -4280 -16680 -4110 -8880
rect -4080 -16680 -3910 -8880
rect -3880 -16680 -3710 -8880
rect -3680 -8910 -3510 -8880
rect -3680 -9000 23560 -8910
rect -3680 -9030 -3510 -9000
rect -3680 -9120 23560 -9030
rect -3680 -9150 -3510 -9120
rect -3680 -9240 23560 -9150
rect -3680 -9270 -3510 -9240
rect -3680 -9360 23560 -9270
rect -3680 -9390 -3510 -9360
rect -3680 -9480 23560 -9390
rect -3680 -9510 -3510 -9480
rect -3680 -9600 23560 -9510
rect -3680 -15960 -3510 -9600
rect -2920 -9690 -1850 -9660
rect -1820 -9690 -1810 -9660
rect 10270 -9690 10410 -9660
rect 22490 -9690 22500 -9660
rect 22530 -9690 23600 -9660
rect -2920 -12560 -2890 -9690
rect -2850 -12520 -2820 -9730
rect -1010 -12490 -960 -12480
rect -1010 -12520 -1000 -12490
rect -970 -12520 -960 -12490
rect -1010 -12530 -960 -12520
rect 21640 -12490 21690 -12480
rect 21640 -12520 21650 -12490
rect 21680 -12520 21690 -12490
rect 23500 -12520 23530 -9730
rect 21640 -12530 21690 -12520
rect 23570 -12560 23600 -9690
rect -2920 -12590 -2820 -12560
rect 23500 -12590 23600 -12560
rect -2920 -13000 -2820 -12970
rect 23500 -13000 23600 -12970
rect -2920 -15870 -2890 -13000
rect -1010 -13040 -960 -13030
rect -2850 -15830 -2820 -13040
rect -1010 -13070 -1000 -13040
rect -970 -13070 -960 -13040
rect -1010 -13080 -960 -13070
rect 21640 -13040 21690 -13030
rect 21640 -13070 21650 -13040
rect 21680 -13070 21690 -13040
rect 21640 -13080 21690 -13070
rect 23500 -15830 23530 -13040
rect 23570 -15870 23600 -13000
rect -2920 -15900 -1850 -15870
rect -1820 -15900 -1810 -15870
rect 10270 -15900 10410 -15870
rect 22490 -15900 22500 -15870
rect 22530 -15900 23600 -15870
rect -3680 -16050 23560 -15960
rect -3680 -16080 -3510 -16050
rect -3680 -16170 23560 -16080
rect -3680 -16200 -3510 -16170
rect -3680 -16290 23560 -16200
rect -3680 -16320 -3510 -16290
rect -3680 -16410 23560 -16320
rect -3680 -16440 -3510 -16410
rect -3680 -16530 23560 -16440
rect -3680 -16560 -3510 -16530
rect -3680 -16650 23560 -16560
rect -3680 -16680 -3510 -16650
rect -6280 -16720 24420 -16680
rect -6280 -16860 24270 -16720
rect 24410 -16860 24420 -16720
rect -6280 -16900 24420 -16860
rect -6280 -21220 -6110 -16900
rect -6080 -21220 -5910 -16900
rect -5880 -21220 -5710 -16900
rect -5680 -21220 -5510 -16900
rect -5480 -21220 -5310 -16900
rect -5280 -21220 -5110 -16900
rect -5080 -21220 -4710 -16900
rect -4680 -21220 -4510 -16900
rect -4480 -21220 -4310 -16900
rect -4280 -21220 -4110 -16900
rect -4080 -21220 -3910 -16900
rect -3880 -21220 -3710 -16900
rect -3680 -16930 -3510 -16900
rect -3680 -17020 23560 -16930
rect -3680 -17050 -3510 -17020
rect -3680 -17140 23560 -17050
rect -3680 -17170 -3510 -17140
rect -3680 -17260 23560 -17170
rect -3680 -17290 -3510 -17260
rect -3680 -17380 23560 -17290
rect -3680 -17410 -3510 -17380
rect -3680 -17500 23560 -17410
rect -3680 -17530 -3510 -17500
rect -3680 -17620 23560 -17530
rect -3680 -20500 -3510 -17620
rect -2920 -17710 -2810 -17680
rect 23500 -17710 23600 -17680
rect -2920 -18840 -2890 -17710
rect -1860 -18840 -1810 -18830
rect 22490 -18840 22540 -18830
rect 23570 -18840 23600 -17710
rect -2920 -18870 -1850 -18840
rect -1820 -18870 22500 -18840
rect 22530 -18870 23600 -18840
rect -1860 -18880 -1810 -18870
rect 22490 -18880 22540 -18870
rect -1860 -19250 -1810 -19240
rect 22490 -19250 22540 -19240
rect -2920 -19280 -1850 -19250
rect -1820 -19280 22500 -19250
rect 22530 -19280 23600 -19250
rect -2920 -20410 -2890 -19280
rect -1860 -19290 -1810 -19280
rect 22490 -19290 22540 -19280
rect 23570 -20410 23600 -19280
rect -2920 -20440 -2810 -20410
rect 23500 -20440 23600 -20410
rect -3680 -20590 23560 -20500
rect -3680 -20620 -3510 -20590
rect -3680 -20710 23560 -20620
rect -3680 -20740 -3510 -20710
rect -3680 -20830 23560 -20740
rect -3680 -20860 -3510 -20830
rect -3680 -20950 23560 -20860
rect -3680 -20980 -3510 -20950
rect -3680 -21070 23560 -20980
rect -3680 -21100 -3510 -21070
rect -3680 -21190 23560 -21100
rect -3680 -21220 -3510 -21190
rect -6280 -21260 24420 -21220
rect -6280 -21400 24270 -21260
rect 24410 -21400 24420 -21260
rect -6280 -21440 24420 -21400
rect -6280 -28520 -6110 -21440
rect -6080 -28520 -5910 -21440
rect -5880 -28520 -5710 -21440
rect -5680 -28520 -5510 -21440
rect -5480 -28520 -5310 -21440
rect -5280 -28520 -5110 -21440
rect -5080 -28520 -4710 -21440
rect -4680 -28520 -4510 -21440
rect -4480 -28520 -4310 -21440
rect -4280 -28520 -4110 -21440
rect -4080 -28520 -3910 -21440
rect -3880 -28520 -3710 -21440
rect -3680 -21470 -3510 -21440
rect -3680 -21560 23560 -21470
rect -3680 -21590 -3510 -21560
rect -3680 -21680 23560 -21590
rect -3680 -21710 -3510 -21680
rect -3680 -21800 23560 -21710
rect -3680 -21830 -3510 -21800
rect -3680 -21920 23560 -21830
rect -3680 -21950 -3510 -21920
rect -3680 -22040 23560 -21950
rect -3680 -22070 -3510 -22040
rect -3680 -22160 23560 -22070
rect -3680 -28520 -3510 -22160
rect -2920 -22250 -1850 -22220
rect -1820 -22250 -1810 -22220
rect 10270 -22250 10410 -22220
rect 22490 -22250 22500 -22220
rect 22530 -22250 23600 -22220
rect -2920 -25120 -2890 -22250
rect -2850 -25080 -2820 -22290
rect -1010 -25050 -960 -25040
rect -1010 -25080 -1000 -25050
rect -970 -25080 -960 -25050
rect -1010 -25090 -960 -25080
rect 21640 -25050 21690 -25040
rect 21640 -25080 21650 -25050
rect 21680 -25080 21690 -25050
rect 23500 -25080 23530 -22290
rect 21640 -25090 21690 -25080
rect 23570 -25120 23600 -22250
rect -2920 -25150 -2820 -25120
rect 23500 -25150 23600 -25120
rect -2920 -25440 -2890 -25150
rect -2920 -25470 -2880 -25440
rect 21100 -25470 21130 -25440
rect -2920 -28490 -2890 -25470
rect -2920 -28520 -2880 -28490
rect 21100 -28520 21130 -28490
<< viali >>
rect -1000 -510 -970 -480
rect 21650 -510 21680 -480
rect -1850 -3340 -1820 -3310
rect 22500 -3340 22530 -3310
rect 24270 -4300 24410 -4160
rect -1850 -6310 -1820 -6280
rect 22500 -6310 22530 -6280
rect -1850 -6720 -1820 -6690
rect 22500 -6720 22530 -6690
rect 24270 -8840 24410 -8700
rect -1850 -9690 -1820 -9660
rect 22500 -9690 22530 -9660
rect -1000 -12520 -970 -12490
rect 21650 -12520 21680 -12490
rect -1000 -13070 -970 -13040
rect 21650 -13070 21680 -13040
rect -1850 -15900 -1820 -15870
rect 22500 -15900 22530 -15870
rect 24270 -16860 24410 -16720
rect -1850 -18870 -1820 -18840
rect 22500 -18870 22530 -18840
rect -1850 -19280 -1820 -19250
rect 22500 -19280 22530 -19250
rect 24270 -21400 24410 -21260
rect -1850 -22250 -1820 -22220
rect 22500 -22250 22530 -22220
rect -1000 -25080 -970 -25050
rect 21650 -25080 21680 -25050
<< metal1 >>
rect -6310 -3360 -6280 -220
rect -6110 -3360 -6080 -220
rect -5910 -3360 -5880 -220
rect -5710 -3360 -5680 -220
rect -5510 -3360 -5480 -220
rect -5310 -3360 -5280 -220
rect -5110 -3360 -5080 -220
rect -4710 -3360 -4680 -220
rect -4510 -3360 -4480 -220
rect -4310 -3360 -4280 -220
rect -4110 -3360 -4080 -220
rect -3910 -3360 -3880 -220
rect -3710 -3360 -3680 -220
rect -3510 -3360 -3480 -220
rect -2790 -230 -2760 -220
rect -2790 -3360 -2760 -370
rect -1940 -230 -1910 -220
rect -1940 -390 -1910 -370
rect -1000 -230 -970 -220
rect -1000 -390 -970 -370
rect 880 -230 910 -220
rect 880 -450 910 -370
rect 1820 -230 1850 -220
rect 1820 -450 1850 -370
rect 3700 -230 3730 -220
rect 3700 -390 3730 -370
rect 5580 -230 5610 -220
rect 5580 -390 5610 -370
rect 7460 -230 7490 -220
rect 7460 -390 7490 -370
rect 10280 -230 10310 -220
rect 10280 -390 10310 -370
rect 10370 -230 10400 -220
rect 10370 -390 10400 -370
rect 13190 -230 13220 -220
rect 13190 -390 13220 -370
rect 15070 -230 15100 -220
rect 15070 -390 15100 -370
rect 16950 -230 16980 -220
rect 16950 -390 16980 -370
rect 18830 -230 18860 -220
rect 18830 -450 18860 -370
rect 19770 -230 19800 -220
rect 19770 -450 19800 -370
rect 21650 -230 21680 -220
rect 21650 -390 21680 -370
rect 22590 -230 22620 -220
rect 22590 -390 22620 -370
rect 23440 -230 23470 -220
rect -1010 -480 -960 -470
rect -1010 -510 -1000 -480
rect -970 -510 -960 -480
rect -1010 -520 -960 -510
rect 21640 -480 21690 -470
rect 21640 -510 21650 -480
rect 21680 -510 21690 -480
rect 21640 -520 21690 -510
rect 23440 -540 23470 -370
rect -1860 -3310 -1810 -3300
rect -1860 -3340 -1850 -3310
rect -1820 -3340 -1810 -3310
rect -1860 -3350 -1810 -3340
rect -6320 -3370 -6270 -3360
rect -6320 -3400 -6310 -3370
rect -6280 -3400 -6270 -3370
rect -6320 -3410 -6270 -3400
rect -6120 -3370 -6070 -3360
rect -6120 -3400 -6110 -3370
rect -6080 -3400 -6070 -3370
rect -6120 -3410 -6070 -3400
rect -5920 -3370 -5870 -3360
rect -5920 -3400 -5910 -3370
rect -5880 -3400 -5870 -3370
rect -5920 -3410 -5870 -3400
rect -5720 -3370 -5670 -3360
rect -5720 -3400 -5710 -3370
rect -5680 -3400 -5670 -3370
rect -5720 -3410 -5670 -3400
rect -5520 -3370 -5470 -3360
rect -5520 -3400 -5510 -3370
rect -5480 -3400 -5470 -3370
rect -5520 -3410 -5470 -3400
rect -5320 -3370 -5270 -3360
rect -5320 -3400 -5310 -3370
rect -5280 -3400 -5270 -3370
rect -5320 -3410 -5270 -3400
rect -5120 -3370 -5070 -3360
rect -5120 -3400 -5110 -3370
rect -5080 -3400 -5070 -3370
rect -5120 -3410 -5070 -3400
rect -4720 -3370 -4670 -3360
rect -4720 -3400 -4710 -3370
rect -4680 -3400 -4670 -3370
rect -4720 -3410 -4670 -3400
rect -4520 -3370 -4470 -3360
rect -4520 -3400 -4510 -3370
rect -4480 -3400 -4470 -3370
rect -4520 -3410 -4470 -3400
rect -4320 -3370 -4270 -3360
rect -4320 -3400 -4310 -3370
rect -4280 -3400 -4270 -3370
rect -4320 -3410 -4270 -3400
rect -4120 -3370 -4070 -3360
rect -4120 -3400 -4110 -3370
rect -4080 -3400 -4070 -3370
rect -4120 -3410 -4070 -3400
rect -3920 -3370 -3870 -3360
rect -3920 -3400 -3910 -3370
rect -3880 -3400 -3870 -3370
rect -3920 -3410 -3870 -3400
rect -3720 -3370 -3670 -3360
rect -3720 -3400 -3710 -3370
rect -3680 -3400 -3670 -3370
rect -3720 -3410 -3670 -3400
rect -3520 -3370 -3470 -3360
rect -3520 -3400 -3510 -3370
rect -3480 -3400 -3470 -3370
rect -3520 -3410 -3470 -3400
rect -6310 -3480 -6280 -3410
rect -6320 -3490 -6270 -3480
rect -6320 -3520 -6310 -3490
rect -6280 -3520 -6270 -3490
rect -6320 -3530 -6270 -3520
rect -6310 -3600 -6280 -3530
rect -6320 -3610 -6270 -3600
rect -6320 -3640 -6310 -3610
rect -6280 -3640 -6270 -3610
rect -6320 -3650 -6270 -3640
rect -6310 -3720 -6280 -3650
rect -6320 -3730 -6270 -3720
rect -6320 -3760 -6310 -3730
rect -6280 -3760 -6270 -3730
rect -6320 -3770 -6270 -3760
rect -6310 -3840 -6280 -3770
rect -6320 -3850 -6270 -3840
rect -6320 -3880 -6310 -3850
rect -6280 -3880 -6270 -3850
rect -6320 -3890 -6270 -3880
rect -6310 -3960 -6280 -3890
rect -6320 -3970 -6270 -3960
rect -6320 -4000 -6310 -3970
rect -6280 -4000 -6270 -3970
rect -6320 -4010 -6270 -4000
rect -6310 -4080 -6280 -4010
rect -6320 -4090 -6270 -4080
rect -6320 -4120 -6310 -4090
rect -6280 -4120 -6270 -4090
rect -6320 -4130 -6270 -4120
rect -6310 -4330 -6280 -4130
rect -6320 -4340 -6270 -4330
rect -6320 -4370 -6310 -4340
rect -6280 -4370 -6270 -4340
rect -6320 -4380 -6270 -4370
rect -6310 -4450 -6280 -4380
rect -6320 -4460 -6270 -4450
rect -6320 -4490 -6310 -4460
rect -6280 -4490 -6270 -4460
rect -6320 -4500 -6270 -4490
rect -6310 -4570 -6280 -4500
rect -6320 -4580 -6270 -4570
rect -6320 -4610 -6310 -4580
rect -6280 -4610 -6270 -4580
rect -6320 -4620 -6270 -4610
rect -6310 -4690 -6280 -4620
rect -6320 -4700 -6270 -4690
rect -6320 -4730 -6310 -4700
rect -6280 -4730 -6270 -4700
rect -6320 -4740 -6270 -4730
rect -6310 -4810 -6280 -4740
rect -6320 -4820 -6270 -4810
rect -6320 -4850 -6310 -4820
rect -6280 -4850 -6270 -4820
rect -6320 -4860 -6270 -4850
rect -6310 -4930 -6280 -4860
rect -6320 -4940 -6270 -4930
rect -6320 -4970 -6310 -4940
rect -6280 -4970 -6270 -4940
rect -6320 -4980 -6270 -4970
rect -6310 -5050 -6280 -4980
rect -6110 -5050 -6080 -3410
rect -5910 -5050 -5880 -3410
rect -5710 -5050 -5680 -3410
rect -5510 -5050 -5480 -3410
rect -5310 -5050 -5280 -3410
rect -5110 -5050 -5080 -3410
rect -4710 -5050 -4680 -3410
rect -4510 -5050 -4480 -3410
rect -4310 -5050 -4280 -3410
rect -4110 -5050 -4080 -3410
rect -3910 -5050 -3880 -3410
rect -3710 -5050 -3680 -3410
rect -3510 -5050 -3480 -3410
rect -2670 -3430 -2640 -3360
rect -2670 -3470 -2640 -3460
rect -2060 -5000 -2030 -4990
rect -6320 -5060 -6270 -5050
rect -6320 -5090 -6310 -5060
rect -6280 -5090 -6270 -5060
rect -6320 -5100 -6270 -5090
rect -6120 -5060 -6070 -5050
rect -6120 -5090 -6110 -5060
rect -6080 -5090 -6070 -5060
rect -6120 -5100 -6070 -5090
rect -5920 -5060 -5870 -5050
rect -5920 -5090 -5910 -5060
rect -5880 -5090 -5870 -5060
rect -5920 -5100 -5870 -5090
rect -5720 -5060 -5670 -5050
rect -5720 -5090 -5710 -5060
rect -5680 -5090 -5670 -5060
rect -5720 -5100 -5670 -5090
rect -5520 -5060 -5470 -5050
rect -5520 -5090 -5510 -5060
rect -5480 -5090 -5470 -5060
rect -5520 -5100 -5470 -5090
rect -5320 -5060 -5270 -5050
rect -5320 -5090 -5310 -5060
rect -5280 -5090 -5270 -5060
rect -5320 -5100 -5270 -5090
rect -5120 -5060 -5070 -5050
rect -5120 -5090 -5110 -5060
rect -5080 -5090 -5070 -5060
rect -5120 -5100 -5070 -5090
rect -4720 -5060 -4670 -5050
rect -4720 -5090 -4710 -5060
rect -4680 -5090 -4670 -5060
rect -4720 -5100 -4670 -5090
rect -4520 -5060 -4470 -5050
rect -4520 -5090 -4510 -5060
rect -4480 -5090 -4470 -5060
rect -4520 -5100 -4470 -5090
rect -4320 -5060 -4270 -5050
rect -4320 -5090 -4310 -5060
rect -4280 -5090 -4270 -5060
rect -4320 -5100 -4270 -5090
rect -4120 -5060 -4070 -5050
rect -4120 -5090 -4110 -5060
rect -4080 -5090 -4070 -5060
rect -4120 -5100 -4070 -5090
rect -3920 -5060 -3870 -5050
rect -3920 -5090 -3910 -5060
rect -3880 -5090 -3870 -5060
rect -3920 -5100 -3870 -5090
rect -3720 -5060 -3670 -5050
rect -3720 -5090 -3710 -5060
rect -3680 -5090 -3670 -5060
rect -3720 -5100 -3670 -5090
rect -3520 -5060 -3470 -5050
rect -3520 -5090 -3510 -5060
rect -3480 -5090 -3470 -5060
rect -3520 -5100 -3470 -5090
rect -6310 -7900 -6280 -5100
rect -6110 -7900 -6080 -5100
rect -5910 -7900 -5880 -5100
rect -5710 -7900 -5680 -5100
rect -5510 -7900 -5480 -5100
rect -5310 -7900 -5280 -5100
rect -5110 -7900 -5080 -5100
rect -4710 -7900 -4680 -5100
rect -4510 -7900 -4480 -5100
rect -4310 -7900 -4280 -5100
rect -4110 -7900 -4080 -5100
rect -3910 -7900 -3880 -5100
rect -3710 -7900 -3680 -5100
rect -3510 -7900 -3480 -5100
rect -2790 -6350 -2760 -5100
rect -2060 -5110 -2030 -5030
rect -2790 -6510 -2760 -6490
rect -2790 -7900 -2760 -6650
rect -1940 -6350 -1910 -5100
rect -1850 -6270 -1820 -3350
rect -1730 -3430 -1700 -3360
rect -1730 -3470 -1700 -3460
rect -1000 -3430 -970 -3360
rect -1000 -3470 -970 -3460
rect -910 -3550 -880 -3360
rect -910 -3590 -880 -3580
rect -790 -3550 -760 -3360
rect -60 -3430 -30 -3150
rect 1820 -3160 1850 -3150
rect -60 -3470 -30 -3460
rect 150 -3430 180 -3360
rect 150 -3470 180 -3460
rect -790 -3590 -760 -3580
rect 760 -4880 790 -4870
rect -1120 -5000 -1090 -4990
rect -1120 -5100 -1090 -5030
rect -910 -5000 -880 -4990
rect -910 -5100 -880 -5030
rect -180 -5000 -150 -4990
rect -180 -5100 -150 -5030
rect 30 -5000 60 -4990
rect 30 -5240 60 -5030
rect 760 -5100 790 -4910
rect 880 -4880 910 -3360
rect 1090 -3430 1120 -3360
rect 1090 -3470 1120 -3460
rect 1820 -3670 1850 -3360
rect 1820 -3710 1850 -3700
rect 1910 -3670 1940 -3360
rect 1910 -3710 1940 -3700
rect 2030 -3790 2060 -3360
rect 2030 -3830 2060 -3820
rect 880 -5100 910 -4910
rect 970 -4030 1000 -4020
rect 970 -5100 1000 -4060
rect 1910 -4030 1940 -4020
rect 1700 -4520 1730 -4510
rect 1700 -5100 1730 -4550
rect 1910 -5240 1940 -4060
rect 2760 -4030 2790 -3150
rect 2970 -3430 3000 -3360
rect 2970 -3470 3000 -3460
rect 3700 -3670 3730 -3360
rect 3700 -3710 3730 -3700
rect 3790 -3670 3820 -3360
rect 3790 -3710 3820 -3700
rect 3910 -3910 3940 -3350
rect 3910 -3950 3940 -3940
rect 2760 -4070 2790 -4060
rect 2850 -4400 2880 -4390
rect 2640 -4520 2670 -4510
rect 2640 -5100 2670 -4550
rect 2760 -4520 2790 -4510
rect 2760 -5100 2790 -4550
rect 2850 -5100 2880 -4430
rect 3790 -4400 3820 -4390
rect 3580 -4520 3610 -4510
rect 3580 -5100 3610 -4550
rect 3790 -5240 3820 -4430
rect 4640 -4400 4670 -3150
rect 4850 -3430 4880 -3360
rect 4850 -3470 4880 -3460
rect 4640 -4440 4670 -4430
rect 4730 -4400 4760 -4390
rect 4520 -4520 4550 -4510
rect 4520 -5100 4550 -4550
rect 4640 -4760 4670 -4750
rect 4640 -5100 4670 -4790
rect 4730 -5100 4760 -4430
rect 5460 -4520 5490 -4510
rect 5460 -5100 5490 -4550
rect 5580 -4520 5610 -3360
rect 5670 -3670 5700 -3360
rect 5670 -3710 5700 -3700
rect 5790 -3910 5820 -3360
rect 5790 -3950 5820 -3940
rect 5580 -4560 5610 -4550
rect 5670 -4400 5700 -4390
rect 5670 -5240 5700 -4430
rect 6520 -4400 6550 -3150
rect 6730 -3430 6760 -3360
rect 6730 -3470 6760 -3460
rect 6520 -4440 6550 -4430
rect 6610 -4030 6640 -4020
rect 6400 -4520 6430 -4510
rect 6400 -5100 6430 -4550
rect 6520 -4760 6550 -4750
rect 6520 -5100 6550 -4790
rect 6610 -5100 6640 -4060
rect 7340 -4520 7370 -4510
rect 7340 -5100 7370 -4550
rect 7460 -4640 7490 -3360
rect 7550 -3670 7580 -3360
rect 7550 -3710 7580 -3700
rect 7670 -3790 7700 -3360
rect 7670 -3830 7700 -3820
rect 7460 -4680 7490 -4670
rect 7550 -4030 7580 -4020
rect 7550 -5240 7580 -4060
rect 8400 -4030 8430 -3150
rect 8400 -4070 8430 -4060
rect 8280 -4520 8310 -4510
rect 8280 -5100 8310 -4550
rect 8400 -4520 8430 -4510
rect 8400 -5100 8430 -4550
rect 8490 -4640 8520 -3360
rect 8610 -3550 8640 -3360
rect 8610 -3590 8640 -3580
rect 8490 -5240 8520 -4670
rect 9340 -4760 9370 -3150
rect 9220 -4880 9250 -4870
rect 9220 -5100 9250 -4910
rect 9340 -5100 9370 -4790
rect 9430 -4160 9460 -4150
rect 9430 -5100 9460 -4300
rect 9550 -4640 9580 -3350
rect 10280 -4160 10310 -2570
rect 10280 -4310 10310 -4300
rect 10370 -4160 10400 -3360
rect 10370 -4310 10400 -4300
rect 9550 -4680 9580 -4670
rect 11100 -4640 11130 -3360
rect 11100 -4680 11130 -4670
rect 11220 -4160 11250 -4150
rect 10160 -4760 10190 -4750
rect 10160 -5100 10190 -4790
rect 10490 -4760 10520 -4750
rect 10490 -5100 10520 -4790
rect 11220 -5100 11250 -4300
rect 11310 -4760 11340 -3150
rect 12040 -3550 12070 -3360
rect 12040 -3590 12070 -3580
rect 11310 -5100 11340 -4790
rect 12160 -4640 12190 -3360
rect 12250 -4030 12280 -3150
rect 12980 -3790 13010 -3360
rect 13100 -3670 13130 -3360
rect 13100 -3710 13130 -3700
rect 12980 -3830 13010 -3820
rect 12250 -4070 12280 -4060
rect 13100 -4030 13130 -4020
rect 11430 -4880 11460 -4870
rect 11430 -5100 11460 -4910
rect 12160 -5240 12190 -4670
rect 12250 -4520 12280 -4510
rect 12250 -5100 12280 -4550
rect 12370 -4520 12400 -4510
rect 12370 -5100 12400 -4550
rect 13100 -5240 13130 -4060
rect 13190 -4640 13220 -3360
rect 13920 -3430 13950 -3360
rect 13920 -3470 13950 -3460
rect 14040 -4030 14070 -4020
rect 13190 -4680 13220 -4670
rect 13310 -4520 13340 -4510
rect 13310 -5100 13340 -4550
rect 14040 -5100 14070 -4060
rect 14130 -4400 14160 -3150
rect 14860 -3910 14890 -3360
rect 14980 -3670 15010 -3360
rect 14980 -3710 15010 -3700
rect 14860 -3950 14890 -3940
rect 14130 -4440 14160 -4430
rect 14980 -4400 15010 -4390
rect 14250 -4520 14280 -4510
rect 14130 -4760 14160 -4750
rect 14130 -5100 14160 -4790
rect 14250 -5100 14280 -4550
rect 14980 -5240 15010 -4430
rect 15070 -4520 15100 -3360
rect 15800 -3430 15830 -3360
rect 15800 -3470 15830 -3460
rect 15920 -4400 15950 -4390
rect 15070 -4560 15100 -4550
rect 15190 -4520 15220 -4510
rect 15190 -5100 15220 -4550
rect 15920 -5100 15950 -4430
rect 16010 -4400 16040 -3150
rect 16740 -3910 16770 -3350
rect 16860 -3670 16890 -3360
rect 16860 -3710 16890 -3700
rect 16950 -3670 16980 -3360
rect 17680 -3430 17710 -3360
rect 17680 -3470 17710 -3460
rect 16950 -3710 16980 -3700
rect 16740 -3950 16770 -3940
rect 17890 -4030 17920 -3150
rect 18830 -3160 18860 -3150
rect 18620 -3790 18650 -3360
rect 18740 -3670 18770 -3360
rect 18740 -3710 18770 -3700
rect 18830 -3670 18860 -3360
rect 19560 -3430 19590 -3360
rect 19560 -3470 19590 -3460
rect 18830 -3710 18860 -3700
rect 18620 -3830 18650 -3820
rect 17890 -4070 17920 -4060
rect 18740 -4030 18770 -4020
rect 16010 -4440 16040 -4430
rect 16860 -4400 16890 -4390
rect 16130 -4520 16160 -4510
rect 16010 -4760 16040 -4750
rect 16010 -5100 16040 -4790
rect 16130 -5100 16160 -4550
rect 16860 -5240 16890 -4430
rect 17800 -4400 17830 -4390
rect 17070 -4520 17100 -4510
rect 17070 -5100 17100 -4550
rect 17800 -5100 17830 -4430
rect 17890 -4520 17920 -4510
rect 17890 -5100 17920 -4550
rect 18010 -4520 18040 -4510
rect 18010 -5100 18040 -4550
rect 18740 -5240 18770 -4060
rect 19680 -4030 19710 -4020
rect 18950 -4520 18980 -4510
rect 18950 -5100 18980 -4550
rect 19680 -5100 19710 -4060
rect 19770 -4880 19800 -3360
rect 20500 -3430 20530 -3360
rect 20500 -3470 20530 -3460
rect 20710 -3430 20740 -3150
rect 22490 -3310 22540 -3300
rect 22490 -3340 22500 -3310
rect 22530 -3340 22540 -3310
rect 22490 -3350 22540 -3340
rect 20710 -3470 20740 -3460
rect 21440 -3550 21470 -3360
rect 21440 -3590 21470 -3580
rect 21560 -3550 21590 -3360
rect 21650 -3430 21680 -3360
rect 21650 -3470 21680 -3460
rect 22380 -3430 22410 -3360
rect 22380 -3470 22410 -3460
rect 21560 -3590 21590 -3580
rect 19770 -5100 19800 -4910
rect 19890 -4880 19920 -4870
rect 19890 -5100 19920 -4910
rect 20620 -5000 20650 -4990
rect 20620 -5240 20650 -5030
rect 20830 -5000 20860 -4990
rect 20830 -5100 20860 -5030
rect 21560 -5000 21590 -4990
rect 21560 -5100 21590 -5030
rect 21770 -5000 21800 -4990
rect 21770 -5100 21800 -5030
rect 22500 -6270 22530 -3350
rect 23320 -3430 23350 -3330
rect 23320 -3470 23350 -3460
rect 24260 -4160 24420 -4150
rect 24260 -4300 24270 -4160
rect 24410 -4300 24420 -4160
rect 24260 -4310 24420 -4300
rect 22710 -5000 22740 -4990
rect 22710 -5100 22740 -5030
rect -1860 -6280 -1810 -6270
rect -1860 -6310 -1850 -6280
rect -1820 -6310 -1810 -6280
rect -1860 -6320 -1810 -6310
rect 22490 -6280 22540 -6270
rect 22490 -6310 22500 -6280
rect 22530 -6310 22540 -6280
rect 22490 -6320 22540 -6310
rect -1940 -6510 -1910 -6490
rect -6320 -7910 -6270 -7900
rect -6320 -7940 -6310 -7910
rect -6280 -7940 -6270 -7910
rect -6320 -7950 -6270 -7940
rect -6120 -7910 -6070 -7900
rect -6120 -7940 -6110 -7910
rect -6080 -7940 -6070 -7910
rect -6120 -7950 -6070 -7940
rect -5920 -7910 -5870 -7900
rect -5920 -7940 -5910 -7910
rect -5880 -7940 -5870 -7910
rect -5920 -7950 -5870 -7940
rect -5720 -7910 -5670 -7900
rect -5720 -7940 -5710 -7910
rect -5680 -7940 -5670 -7910
rect -5720 -7950 -5670 -7940
rect -5520 -7910 -5470 -7900
rect -5520 -7940 -5510 -7910
rect -5480 -7940 -5470 -7910
rect -5520 -7950 -5470 -7940
rect -5320 -7910 -5270 -7900
rect -5320 -7940 -5310 -7910
rect -5280 -7940 -5270 -7910
rect -5320 -7950 -5270 -7940
rect -5120 -7910 -5070 -7900
rect -5120 -7940 -5110 -7910
rect -5080 -7940 -5070 -7910
rect -5120 -7950 -5070 -7940
rect -4720 -7910 -4670 -7900
rect -4720 -7940 -4710 -7910
rect -4680 -7940 -4670 -7910
rect -4720 -7950 -4670 -7940
rect -4520 -7910 -4470 -7900
rect -4520 -7940 -4510 -7910
rect -4480 -7940 -4470 -7910
rect -4520 -7950 -4470 -7940
rect -4320 -7910 -4270 -7900
rect -4320 -7940 -4310 -7910
rect -4280 -7940 -4270 -7910
rect -4320 -7950 -4270 -7940
rect -4120 -7910 -4070 -7900
rect -4120 -7940 -4110 -7910
rect -4080 -7940 -4070 -7910
rect -4120 -7950 -4070 -7940
rect -3920 -7910 -3870 -7900
rect -3920 -7940 -3910 -7910
rect -3880 -7940 -3870 -7910
rect -3920 -7950 -3870 -7940
rect -3720 -7910 -3670 -7900
rect -3720 -7940 -3710 -7910
rect -3680 -7940 -3670 -7910
rect -3720 -7950 -3670 -7940
rect -3520 -7910 -3470 -7900
rect -3520 -7940 -3510 -7910
rect -3480 -7940 -3470 -7910
rect -3520 -7950 -3470 -7940
rect -6310 -8020 -6280 -7950
rect -6320 -8030 -6270 -8020
rect -6320 -8060 -6310 -8030
rect -6280 -8060 -6270 -8030
rect -6320 -8070 -6270 -8060
rect -6310 -8140 -6280 -8070
rect -6320 -8150 -6270 -8140
rect -6320 -8180 -6310 -8150
rect -6280 -8180 -6270 -8150
rect -6320 -8190 -6270 -8180
rect -6310 -8260 -6280 -8190
rect -6320 -8270 -6270 -8260
rect -6320 -8300 -6310 -8270
rect -6280 -8300 -6270 -8270
rect -6320 -8310 -6270 -8300
rect -6310 -8380 -6280 -8310
rect -6320 -8390 -6270 -8380
rect -6320 -8420 -6310 -8390
rect -6280 -8420 -6270 -8390
rect -6320 -8430 -6270 -8420
rect -6310 -8500 -6280 -8430
rect -6320 -8510 -6270 -8500
rect -6320 -8540 -6310 -8510
rect -6280 -8540 -6270 -8510
rect -6320 -8550 -6270 -8540
rect -6310 -8620 -6280 -8550
rect -6320 -8630 -6270 -8620
rect -6320 -8660 -6310 -8630
rect -6280 -8660 -6270 -8630
rect -6320 -8670 -6270 -8660
rect -6310 -8870 -6280 -8670
rect -6320 -8880 -6270 -8870
rect -6320 -8910 -6310 -8880
rect -6280 -8910 -6270 -8880
rect -6320 -8920 -6270 -8910
rect -6310 -8990 -6280 -8920
rect -6320 -9000 -6270 -8990
rect -6320 -9030 -6310 -9000
rect -6280 -9030 -6270 -9000
rect -6320 -9040 -6270 -9030
rect -6310 -9110 -6280 -9040
rect -6320 -9120 -6270 -9110
rect -6320 -9150 -6310 -9120
rect -6280 -9150 -6270 -9120
rect -6320 -9160 -6270 -9150
rect -6310 -9230 -6280 -9160
rect -6320 -9240 -6270 -9230
rect -6320 -9270 -6310 -9240
rect -6280 -9270 -6270 -9240
rect -6320 -9280 -6270 -9270
rect -6310 -9350 -6280 -9280
rect -6320 -9360 -6270 -9350
rect -6320 -9390 -6310 -9360
rect -6280 -9390 -6270 -9360
rect -6320 -9400 -6270 -9390
rect -6310 -9470 -6280 -9400
rect -6320 -9480 -6270 -9470
rect -6320 -9510 -6310 -9480
rect -6280 -9510 -6270 -9480
rect -6320 -9520 -6270 -9510
rect -6310 -9590 -6280 -9520
rect -6110 -9590 -6080 -7950
rect -5910 -9590 -5880 -7950
rect -5710 -9590 -5680 -7950
rect -5510 -9590 -5480 -7950
rect -5310 -9590 -5280 -7950
rect -5110 -9590 -5080 -7950
rect -4710 -9590 -4680 -7950
rect -4510 -9590 -4480 -7950
rect -4310 -9590 -4280 -7950
rect -4110 -9590 -4080 -7950
rect -3910 -9590 -3880 -7950
rect -3710 -9590 -3680 -7950
rect -3510 -9590 -3480 -7950
rect -2060 -7970 -2030 -7890
rect -1940 -7900 -1910 -6650
rect -1850 -6350 -1820 -6320
rect -1850 -6510 -1820 -6490
rect -1850 -6680 -1820 -6650
rect -910 -6350 -880 -6330
rect -910 -6510 -880 -6490
rect -910 -6670 -880 -6650
rect 970 -6350 1000 -6330
rect 970 -6510 1000 -6490
rect 970 -6670 1000 -6650
rect 2850 -6350 2880 -6330
rect 2850 -6510 2880 -6490
rect 2850 -6670 2880 -6650
rect 4730 -6350 4760 -6330
rect 4730 -6510 4760 -6490
rect 4730 -6670 4760 -6650
rect 6610 -6350 6640 -6330
rect 6610 -6510 6640 -6490
rect 6610 -6670 6640 -6650
rect 9430 -6350 9460 -6330
rect 9430 -6510 9460 -6490
rect 9430 -6670 9460 -6650
rect 11220 -6350 11250 -6330
rect 11220 -6510 11250 -6490
rect 11220 -6670 11250 -6650
rect 14040 -6350 14070 -6330
rect 14040 -6510 14070 -6490
rect 14040 -6670 14070 -6650
rect 15920 -6350 15950 -6330
rect 15920 -6510 15950 -6490
rect 15920 -6670 15950 -6650
rect 17800 -6350 17830 -6330
rect 17800 -6510 17830 -6490
rect 17800 -6670 17830 -6650
rect 19680 -6350 19710 -6330
rect 19680 -6510 19710 -6490
rect 19680 -6670 19710 -6650
rect 21560 -6350 21590 -6330
rect 21560 -6510 21590 -6490
rect 21560 -6670 21590 -6650
rect 22500 -6350 22530 -6320
rect 22500 -6510 22530 -6490
rect 22500 -6680 22530 -6650
rect 22590 -6350 22620 -6250
rect 22590 -6510 22620 -6490
rect -1860 -6690 -1810 -6680
rect -1860 -6720 -1850 -6690
rect -1820 -6720 -1810 -6690
rect -1860 -6730 -1810 -6720
rect 22490 -6690 22540 -6680
rect 22490 -6720 22500 -6690
rect 22530 -6720 22540 -6690
rect 22490 -6730 22540 -6720
rect -2060 -8010 -2030 -8000
rect -2670 -9540 -2640 -9530
rect -6320 -9600 -6270 -9590
rect -6320 -9630 -6310 -9600
rect -6280 -9630 -6270 -9600
rect -6320 -9640 -6270 -9630
rect -6120 -9600 -6070 -9590
rect -6120 -9630 -6110 -9600
rect -6080 -9630 -6070 -9600
rect -6120 -9640 -6070 -9630
rect -5920 -9600 -5870 -9590
rect -5920 -9630 -5910 -9600
rect -5880 -9630 -5870 -9600
rect -5920 -9640 -5870 -9630
rect -5720 -9600 -5670 -9590
rect -5720 -9630 -5710 -9600
rect -5680 -9630 -5670 -9600
rect -5720 -9640 -5670 -9630
rect -5520 -9600 -5470 -9590
rect -5520 -9630 -5510 -9600
rect -5480 -9630 -5470 -9600
rect -5520 -9640 -5470 -9630
rect -5320 -9600 -5270 -9590
rect -5320 -9630 -5310 -9600
rect -5280 -9630 -5270 -9600
rect -5320 -9640 -5270 -9630
rect -5120 -9600 -5070 -9590
rect -5120 -9630 -5110 -9600
rect -5080 -9630 -5070 -9600
rect -5120 -9640 -5070 -9630
rect -4720 -9600 -4670 -9590
rect -4720 -9630 -4710 -9600
rect -4680 -9630 -4670 -9600
rect -4720 -9640 -4670 -9630
rect -4520 -9600 -4470 -9590
rect -4520 -9630 -4510 -9600
rect -4480 -9630 -4470 -9600
rect -4520 -9640 -4470 -9630
rect -4320 -9600 -4270 -9590
rect -4320 -9630 -4310 -9600
rect -4280 -9630 -4270 -9600
rect -4320 -9640 -4270 -9630
rect -4120 -9600 -4070 -9590
rect -4120 -9630 -4110 -9600
rect -4080 -9630 -4070 -9600
rect -4120 -9640 -4070 -9630
rect -3920 -9600 -3870 -9590
rect -3920 -9630 -3910 -9600
rect -3880 -9630 -3870 -9600
rect -3920 -9640 -3870 -9630
rect -3720 -9600 -3670 -9590
rect -3720 -9630 -3710 -9600
rect -3680 -9630 -3670 -9600
rect -3720 -9640 -3670 -9630
rect -3520 -9600 -3470 -9590
rect -3520 -9630 -3510 -9600
rect -3480 -9630 -3470 -9600
rect -3520 -9640 -3470 -9630
rect -2670 -9640 -2640 -9570
rect -6310 -15920 -6280 -9640
rect -6110 -15920 -6080 -9640
rect -5910 -15920 -5880 -9640
rect -5710 -15920 -5680 -9640
rect -5510 -15920 -5480 -9640
rect -5310 -15920 -5280 -9640
rect -5110 -15920 -5080 -9640
rect -4710 -15920 -4680 -9640
rect -4510 -15920 -4480 -9640
rect -4310 -15920 -4280 -9640
rect -4110 -15920 -4080 -9640
rect -3910 -15920 -3880 -9640
rect -3710 -15920 -3680 -9640
rect -3510 -15920 -3480 -9640
rect -2790 -12630 -2760 -9640
rect -1850 -9650 -1820 -6730
rect -1120 -7970 -1090 -7900
rect -1120 -8010 -1090 -8000
rect -910 -7970 -880 -7900
rect -910 -8010 -880 -8000
rect -180 -7970 -150 -7900
rect -180 -8010 -150 -8000
rect 30 -7970 60 -7760
rect 30 -8010 60 -8000
rect 760 -8090 790 -7900
rect 760 -8130 790 -8120
rect 880 -8090 910 -7900
rect -910 -9420 -880 -9410
rect -1730 -9540 -1700 -9530
rect -1730 -9640 -1700 -9570
rect -1000 -9540 -970 -9530
rect -1000 -9640 -970 -9570
rect -910 -9640 -880 -9450
rect -790 -9420 -760 -9410
rect -790 -9640 -760 -9450
rect -60 -9540 -30 -9530
rect -1860 -9660 -1810 -9650
rect -1860 -9690 -1850 -9660
rect -1820 -9690 -1810 -9660
rect -1860 -9700 -1810 -9690
rect -60 -9850 -30 -9570
rect 150 -9540 180 -9530
rect 150 -9640 180 -9570
rect 880 -9640 910 -8120
rect 970 -8940 1000 -7900
rect 1700 -8450 1730 -7900
rect 1700 -8490 1730 -8480
rect 970 -8980 1000 -8970
rect 1910 -8940 1940 -7760
rect 2640 -8450 2670 -7900
rect 2640 -8490 2670 -8480
rect 2760 -8450 2790 -7900
rect 2760 -8490 2790 -8480
rect 2850 -8570 2880 -7900
rect 3580 -8450 3610 -7900
rect 3580 -8490 3610 -8480
rect 2850 -8610 2880 -8600
rect 3790 -8570 3820 -7760
rect 4520 -8450 4550 -7900
rect 4640 -8210 4670 -7900
rect 4640 -8250 4670 -8240
rect 4520 -8490 4550 -8480
rect 3790 -8610 3820 -8600
rect 4640 -8570 4670 -8560
rect 1910 -8980 1940 -8970
rect 2760 -8940 2790 -8930
rect 2030 -9180 2060 -9170
rect 1820 -9300 1850 -9290
rect 1090 -9540 1120 -9530
rect 1090 -9640 1120 -9570
rect 1820 -9640 1850 -9330
rect 1910 -9300 1940 -9290
rect 1910 -9640 1940 -9330
rect 2030 -9640 2060 -9210
rect 1820 -9850 1850 -9840
rect 2760 -9850 2790 -8970
rect 3910 -9060 3940 -9050
rect 3700 -9300 3730 -9290
rect 2970 -9540 3000 -9530
rect 2970 -9640 3000 -9570
rect 3700 -9640 3730 -9330
rect 3790 -9300 3820 -9290
rect 3790 -9640 3820 -9330
rect 3910 -9650 3940 -9090
rect 4640 -9850 4670 -8600
rect 4730 -8570 4760 -7900
rect 5460 -8450 5490 -7900
rect 5460 -8490 5490 -8480
rect 5580 -8450 5610 -8440
rect 4730 -8610 4760 -8600
rect 4850 -9540 4880 -9530
rect 4850 -9640 4880 -9570
rect 5580 -9640 5610 -8480
rect 5670 -8570 5700 -7760
rect 6400 -8450 6430 -7900
rect 6520 -8210 6550 -7900
rect 6520 -8250 6550 -8240
rect 6400 -8490 6430 -8480
rect 5670 -8610 5700 -8600
rect 6520 -8570 6550 -8560
rect 5790 -9060 5820 -9050
rect 5670 -9300 5700 -9290
rect 5670 -9640 5700 -9330
rect 5790 -9640 5820 -9090
rect 6520 -9850 6550 -8600
rect 6610 -8940 6640 -7900
rect 7340 -8450 7370 -7900
rect 7340 -8490 7370 -8480
rect 7460 -8330 7490 -8320
rect 6610 -8980 6640 -8970
rect 6730 -9540 6760 -9530
rect 6730 -9640 6760 -9570
rect 7460 -9640 7490 -8360
rect 7550 -8940 7580 -7760
rect 8280 -8450 8310 -7900
rect 8280 -8490 8310 -8480
rect 8400 -8450 8430 -7900
rect 8400 -8490 8430 -8480
rect 8490 -8330 8520 -7760
rect 9220 -8090 9250 -7900
rect 9220 -8130 9250 -8120
rect 7550 -8980 7580 -8970
rect 8400 -8940 8430 -8930
rect 7670 -9180 7700 -9170
rect 7550 -9300 7580 -9290
rect 7550 -9640 7580 -9330
rect 7670 -9640 7700 -9210
rect 8400 -9850 8430 -8970
rect 8490 -9640 8520 -8360
rect 9340 -8210 9370 -7900
rect 8610 -9420 8640 -9410
rect 8610 -9640 8640 -9450
rect 9340 -9850 9370 -8240
rect 9430 -8700 9460 -7900
rect 10160 -8210 10190 -7900
rect 10160 -8250 10190 -8240
rect 10490 -8210 10520 -7900
rect 10490 -8250 10520 -8240
rect 9430 -8850 9460 -8840
rect 9550 -8330 9580 -8320
rect 9550 -9650 9580 -8360
rect 11100 -8330 11130 -8320
rect 10280 -8700 10310 -8690
rect 10280 -10430 10310 -8840
rect 10370 -8700 10400 -8690
rect 10370 -9640 10400 -8840
rect 11100 -9640 11130 -8360
rect 11220 -8700 11250 -7900
rect 11220 -8850 11250 -8840
rect 11310 -8210 11340 -7900
rect 11430 -8090 11460 -7900
rect 11430 -8130 11460 -8120
rect 11310 -9850 11340 -8240
rect 12160 -8330 12190 -7760
rect 12040 -9420 12070 -9410
rect 12040 -9640 12070 -9450
rect 12160 -9640 12190 -8360
rect 12250 -8450 12280 -7900
rect 12250 -8490 12280 -8480
rect 12370 -8450 12400 -7900
rect 12370 -8490 12400 -8480
rect 12250 -8940 12280 -8930
rect 12250 -9850 12280 -8970
rect 13100 -8940 13130 -7760
rect 13100 -8980 13130 -8970
rect 13190 -8330 13220 -8320
rect 12980 -9180 13010 -9170
rect 12980 -9640 13010 -9210
rect 13100 -9300 13130 -9290
rect 13100 -9640 13130 -9330
rect 13190 -9640 13220 -8360
rect 13310 -8450 13340 -7900
rect 13310 -8490 13340 -8480
rect 14040 -8940 14070 -7900
rect 14130 -8210 14160 -7900
rect 14130 -8250 14160 -8240
rect 14250 -8450 14280 -7900
rect 14250 -8490 14280 -8480
rect 14040 -8980 14070 -8970
rect 14130 -8570 14160 -8560
rect 13920 -9540 13950 -9530
rect 13920 -9640 13950 -9570
rect 14130 -9850 14160 -8600
rect 14980 -8570 15010 -7760
rect 14980 -8610 15010 -8600
rect 15070 -8450 15100 -8440
rect 14860 -9060 14890 -9050
rect 14860 -9640 14890 -9090
rect 14980 -9300 15010 -9290
rect 14980 -9640 15010 -9330
rect 15070 -9640 15100 -8480
rect 15190 -8450 15220 -7900
rect 15190 -8490 15220 -8480
rect 15920 -8570 15950 -7900
rect 16010 -8210 16040 -7900
rect 16010 -8250 16040 -8240
rect 16130 -8450 16160 -7900
rect 16130 -8490 16160 -8480
rect 15920 -8610 15950 -8600
rect 16010 -8570 16040 -8560
rect 15800 -9540 15830 -9530
rect 15800 -9640 15830 -9570
rect 16010 -9850 16040 -8600
rect 16860 -8570 16890 -7760
rect 17070 -8450 17100 -7900
rect 17070 -8490 17100 -8480
rect 16860 -8610 16890 -8600
rect 17800 -8570 17830 -7900
rect 17890 -8450 17920 -7900
rect 17890 -8490 17920 -8480
rect 18010 -8450 18040 -7900
rect 18010 -8490 18040 -8480
rect 17800 -8610 17830 -8600
rect 17890 -8940 17920 -8930
rect 16740 -9060 16770 -9050
rect 16740 -9650 16770 -9090
rect 16860 -9300 16890 -9290
rect 16860 -9640 16890 -9330
rect 16950 -9300 16980 -9290
rect 16950 -9640 16980 -9330
rect 17680 -9540 17710 -9530
rect 17680 -9640 17710 -9570
rect 17890 -9850 17920 -8970
rect 18740 -8940 18770 -7760
rect 18950 -8450 18980 -7900
rect 18950 -8490 18980 -8480
rect 18740 -8980 18770 -8970
rect 19680 -8940 19710 -7900
rect 19680 -8980 19710 -8970
rect 19770 -8090 19800 -7900
rect 18620 -9180 18650 -9170
rect 18620 -9640 18650 -9210
rect 18740 -9300 18770 -9290
rect 18740 -9640 18770 -9330
rect 18830 -9300 18860 -9290
rect 18830 -9640 18860 -9330
rect 19560 -9540 19590 -9530
rect 19560 -9640 19590 -9570
rect 19770 -9640 19800 -8120
rect 19890 -8090 19920 -7900
rect 20620 -7970 20650 -7760
rect 20620 -8010 20650 -8000
rect 20830 -7970 20860 -7900
rect 20830 -8010 20860 -8000
rect 21560 -7970 21590 -7900
rect 21560 -8010 21590 -8000
rect 21770 -7970 21800 -7900
rect 21770 -8010 21800 -8000
rect 19890 -8130 19920 -8120
rect 21440 -9420 21470 -9410
rect 20500 -9540 20530 -9530
rect 20500 -9640 20530 -9570
rect 20710 -9540 20740 -9530
rect 18830 -9850 18860 -9840
rect 20710 -9850 20740 -9570
rect 21440 -9640 21470 -9450
rect 21560 -9420 21590 -9410
rect 21560 -9640 21590 -9450
rect 21650 -9540 21680 -9530
rect 21650 -9640 21680 -9570
rect 22380 -9540 22410 -9530
rect 22380 -9640 22410 -9570
rect 22500 -9650 22530 -6730
rect 22590 -6750 22620 -6650
rect 23440 -6350 23470 -6330
rect 23440 -6510 23470 -6490
rect 23440 -6670 23470 -6650
rect 22710 -7970 22740 -7900
rect 22710 -8010 22740 -8000
rect 24260 -8700 24420 -8690
rect 24260 -8840 24270 -8700
rect 24410 -8840 24420 -8700
rect 24260 -8850 24420 -8840
rect 23320 -9540 23350 -9530
rect 22490 -9660 22540 -9650
rect 22490 -9690 22500 -9660
rect 22530 -9690 22540 -9660
rect 23320 -9670 23350 -9570
rect 22490 -9700 22540 -9690
rect -1010 -12490 -960 -12480
rect -1010 -12520 -1000 -12490
rect -970 -12520 -960 -12490
rect -1010 -12530 -960 -12520
rect 21640 -12490 21690 -12480
rect 21640 -12520 21650 -12490
rect 21680 -12520 21690 -12490
rect 21640 -12530 21690 -12520
rect -2790 -12790 -2760 -12770
rect -2790 -15920 -2760 -12930
rect -1940 -12630 -1910 -12610
rect -1940 -12790 -1910 -12770
rect -1940 -12950 -1910 -12930
rect -1000 -12630 -970 -12610
rect -1000 -12790 -970 -12770
rect -1000 -12950 -970 -12930
rect 880 -12630 910 -12550
rect 880 -12790 910 -12770
rect 880 -13010 910 -12930
rect 1820 -12630 1850 -12550
rect 1820 -12790 1850 -12770
rect 1820 -13010 1850 -12930
rect 3700 -12630 3730 -12610
rect 3700 -12790 3730 -12770
rect 3700 -12950 3730 -12930
rect 5580 -12630 5610 -12610
rect 5580 -12790 5610 -12770
rect 5580 -12950 5610 -12930
rect 7460 -12630 7490 -12610
rect 7460 -12790 7490 -12770
rect 7460 -12950 7490 -12930
rect 10280 -12630 10310 -12610
rect 10280 -12790 10310 -12770
rect 10280 -12950 10310 -12930
rect 10370 -12630 10400 -12610
rect 10370 -12790 10400 -12770
rect 10370 -12950 10400 -12930
rect 13190 -12630 13220 -12610
rect 13190 -12790 13220 -12770
rect 13190 -12950 13220 -12930
rect 15070 -12630 15100 -12610
rect 15070 -12790 15100 -12770
rect 15070 -12950 15100 -12930
rect 16950 -12630 16980 -12610
rect 16950 -12790 16980 -12770
rect 16950 -12950 16980 -12930
rect 18830 -12630 18860 -12550
rect 18830 -12790 18860 -12770
rect 18830 -13010 18860 -12930
rect 19770 -12630 19800 -12550
rect 19770 -12790 19800 -12770
rect 19770 -13010 19800 -12930
rect 21650 -12630 21680 -12610
rect 21650 -12790 21680 -12770
rect 21650 -12950 21680 -12930
rect 22590 -12630 22620 -12610
rect 22590 -12790 22620 -12770
rect 22590 -12950 22620 -12930
rect 23440 -12630 23470 -12460
rect 23440 -12790 23470 -12770
rect -1010 -13040 -960 -13030
rect -1010 -13070 -1000 -13040
rect -970 -13070 -960 -13040
rect -1010 -13080 -960 -13070
rect 21640 -13040 21690 -13030
rect 21640 -13070 21650 -13040
rect 21680 -13070 21690 -13040
rect 21640 -13080 21690 -13070
rect 23440 -13100 23470 -12930
rect -1860 -15870 -1810 -15860
rect -1860 -15900 -1850 -15870
rect -1820 -15900 -1810 -15870
rect -1860 -15910 -1810 -15900
rect -6320 -15930 -6270 -15920
rect -6320 -15960 -6310 -15930
rect -6280 -15960 -6270 -15930
rect -6320 -15970 -6270 -15960
rect -6120 -15930 -6070 -15920
rect -6120 -15960 -6110 -15930
rect -6080 -15960 -6070 -15930
rect -6120 -15970 -6070 -15960
rect -5920 -15930 -5870 -15920
rect -5920 -15960 -5910 -15930
rect -5880 -15960 -5870 -15930
rect -5920 -15970 -5870 -15960
rect -5720 -15930 -5670 -15920
rect -5720 -15960 -5710 -15930
rect -5680 -15960 -5670 -15930
rect -5720 -15970 -5670 -15960
rect -5520 -15930 -5470 -15920
rect -5520 -15960 -5510 -15930
rect -5480 -15960 -5470 -15930
rect -5520 -15970 -5470 -15960
rect -5320 -15930 -5270 -15920
rect -5320 -15960 -5310 -15930
rect -5280 -15960 -5270 -15930
rect -5320 -15970 -5270 -15960
rect -5120 -15930 -5070 -15920
rect -5120 -15960 -5110 -15930
rect -5080 -15960 -5070 -15930
rect -5120 -15970 -5070 -15960
rect -4720 -15930 -4670 -15920
rect -4720 -15960 -4710 -15930
rect -4680 -15960 -4670 -15930
rect -4720 -15970 -4670 -15960
rect -4520 -15930 -4470 -15920
rect -4520 -15960 -4510 -15930
rect -4480 -15960 -4470 -15930
rect -4520 -15970 -4470 -15960
rect -4320 -15930 -4270 -15920
rect -4320 -15960 -4310 -15930
rect -4280 -15960 -4270 -15930
rect -4320 -15970 -4270 -15960
rect -4120 -15930 -4070 -15920
rect -4120 -15960 -4110 -15930
rect -4080 -15960 -4070 -15930
rect -4120 -15970 -4070 -15960
rect -3920 -15930 -3870 -15920
rect -3920 -15960 -3910 -15930
rect -3880 -15960 -3870 -15930
rect -3920 -15970 -3870 -15960
rect -3720 -15930 -3670 -15920
rect -3720 -15960 -3710 -15930
rect -3680 -15960 -3670 -15930
rect -3720 -15970 -3670 -15960
rect -3520 -15930 -3470 -15920
rect -3520 -15960 -3510 -15930
rect -3480 -15960 -3470 -15930
rect -3520 -15970 -3470 -15960
rect -6310 -16040 -6280 -15970
rect -6320 -16050 -6270 -16040
rect -6320 -16080 -6310 -16050
rect -6280 -16080 -6270 -16050
rect -6320 -16090 -6270 -16080
rect -6310 -16160 -6280 -16090
rect -6320 -16170 -6270 -16160
rect -6320 -16200 -6310 -16170
rect -6280 -16200 -6270 -16170
rect -6320 -16210 -6270 -16200
rect -6310 -16280 -6280 -16210
rect -6320 -16290 -6270 -16280
rect -6320 -16320 -6310 -16290
rect -6280 -16320 -6270 -16290
rect -6320 -16330 -6270 -16320
rect -6310 -16400 -6280 -16330
rect -6320 -16410 -6270 -16400
rect -6320 -16440 -6310 -16410
rect -6280 -16440 -6270 -16410
rect -6320 -16450 -6270 -16440
rect -6310 -16520 -6280 -16450
rect -6320 -16530 -6270 -16520
rect -6320 -16560 -6310 -16530
rect -6280 -16560 -6270 -16530
rect -6320 -16570 -6270 -16560
rect -6310 -16640 -6280 -16570
rect -6320 -16650 -6270 -16640
rect -6320 -16680 -6310 -16650
rect -6280 -16680 -6270 -16650
rect -6320 -16690 -6270 -16680
rect -6310 -16890 -6280 -16690
rect -6320 -16900 -6270 -16890
rect -6320 -16930 -6310 -16900
rect -6280 -16930 -6270 -16900
rect -6320 -16940 -6270 -16930
rect -6310 -17010 -6280 -16940
rect -6320 -17020 -6270 -17010
rect -6320 -17050 -6310 -17020
rect -6280 -17050 -6270 -17020
rect -6320 -17060 -6270 -17050
rect -6310 -17130 -6280 -17060
rect -6320 -17140 -6270 -17130
rect -6320 -17170 -6310 -17140
rect -6280 -17170 -6270 -17140
rect -6320 -17180 -6270 -17170
rect -6310 -17250 -6280 -17180
rect -6320 -17260 -6270 -17250
rect -6320 -17290 -6310 -17260
rect -6280 -17290 -6270 -17260
rect -6320 -17300 -6270 -17290
rect -6310 -17370 -6280 -17300
rect -6320 -17380 -6270 -17370
rect -6320 -17410 -6310 -17380
rect -6280 -17410 -6270 -17380
rect -6320 -17420 -6270 -17410
rect -6310 -17490 -6280 -17420
rect -6320 -17500 -6270 -17490
rect -6320 -17530 -6310 -17500
rect -6280 -17530 -6270 -17500
rect -6320 -17540 -6270 -17530
rect -6310 -17610 -6280 -17540
rect -6110 -17610 -6080 -15970
rect -5910 -17610 -5880 -15970
rect -5710 -17610 -5680 -15970
rect -5510 -17610 -5480 -15970
rect -5310 -17610 -5280 -15970
rect -5110 -17610 -5080 -15970
rect -4710 -17610 -4680 -15970
rect -4510 -17610 -4480 -15970
rect -4310 -17610 -4280 -15970
rect -4110 -17610 -4080 -15970
rect -3910 -17610 -3880 -15970
rect -3710 -17610 -3680 -15970
rect -3510 -17610 -3480 -15970
rect -2670 -15990 -2640 -15920
rect -2670 -16030 -2640 -16020
rect -2060 -17560 -2030 -17550
rect -6320 -17620 -6270 -17610
rect -6320 -17650 -6310 -17620
rect -6280 -17650 -6270 -17620
rect -6320 -17660 -6270 -17650
rect -6120 -17620 -6070 -17610
rect -6120 -17650 -6110 -17620
rect -6080 -17650 -6070 -17620
rect -6120 -17660 -6070 -17650
rect -5920 -17620 -5870 -17610
rect -5920 -17650 -5910 -17620
rect -5880 -17650 -5870 -17620
rect -5920 -17660 -5870 -17650
rect -5720 -17620 -5670 -17610
rect -5720 -17650 -5710 -17620
rect -5680 -17650 -5670 -17620
rect -5720 -17660 -5670 -17650
rect -5520 -17620 -5470 -17610
rect -5520 -17650 -5510 -17620
rect -5480 -17650 -5470 -17620
rect -5520 -17660 -5470 -17650
rect -5320 -17620 -5270 -17610
rect -5320 -17650 -5310 -17620
rect -5280 -17650 -5270 -17620
rect -5320 -17660 -5270 -17650
rect -5120 -17620 -5070 -17610
rect -5120 -17650 -5110 -17620
rect -5080 -17650 -5070 -17620
rect -5120 -17660 -5070 -17650
rect -4720 -17620 -4670 -17610
rect -4720 -17650 -4710 -17620
rect -4680 -17650 -4670 -17620
rect -4720 -17660 -4670 -17650
rect -4520 -17620 -4470 -17610
rect -4520 -17650 -4510 -17620
rect -4480 -17650 -4470 -17620
rect -4520 -17660 -4470 -17650
rect -4320 -17620 -4270 -17610
rect -4320 -17650 -4310 -17620
rect -4280 -17650 -4270 -17620
rect -4320 -17660 -4270 -17650
rect -4120 -17620 -4070 -17610
rect -4120 -17650 -4110 -17620
rect -4080 -17650 -4070 -17620
rect -4120 -17660 -4070 -17650
rect -3920 -17620 -3870 -17610
rect -3920 -17650 -3910 -17620
rect -3880 -17650 -3870 -17620
rect -3920 -17660 -3870 -17650
rect -3720 -17620 -3670 -17610
rect -3720 -17650 -3710 -17620
rect -3680 -17650 -3670 -17620
rect -3720 -17660 -3670 -17650
rect -3520 -17620 -3470 -17610
rect -3520 -17650 -3510 -17620
rect -3480 -17650 -3470 -17620
rect -3520 -17660 -3470 -17650
rect -6310 -20460 -6280 -17660
rect -6110 -20460 -6080 -17660
rect -5910 -20460 -5880 -17660
rect -5710 -20460 -5680 -17660
rect -5510 -20460 -5480 -17660
rect -5310 -20460 -5280 -17660
rect -5110 -20460 -5080 -17660
rect -4710 -20460 -4680 -17660
rect -4510 -20460 -4480 -17660
rect -4310 -20460 -4280 -17660
rect -4110 -20460 -4080 -17660
rect -3910 -20460 -3880 -17660
rect -3710 -20460 -3680 -17660
rect -3510 -20460 -3480 -17660
rect -2790 -18910 -2760 -17660
rect -2060 -17670 -2030 -17590
rect -2790 -19070 -2760 -19050
rect -2790 -20460 -2760 -19210
rect -1940 -18910 -1910 -17660
rect -1850 -18830 -1820 -15910
rect -1730 -15990 -1700 -15920
rect -1730 -16030 -1700 -16020
rect -1000 -15990 -970 -15920
rect -1000 -16030 -970 -16020
rect -910 -16110 -880 -15920
rect -910 -16150 -880 -16140
rect -790 -16110 -760 -15920
rect -60 -15990 -30 -15710
rect 1820 -15720 1850 -15710
rect -60 -16030 -30 -16020
rect 150 -15990 180 -15920
rect 150 -16030 180 -16020
rect -790 -16150 -760 -16140
rect 760 -17440 790 -17430
rect -1120 -17560 -1090 -17550
rect -1120 -17660 -1090 -17590
rect -910 -17560 -880 -17550
rect -910 -17660 -880 -17590
rect -180 -17560 -150 -17550
rect -180 -17660 -150 -17590
rect 30 -17560 60 -17550
rect 30 -17800 60 -17590
rect 760 -17660 790 -17470
rect 880 -17440 910 -15920
rect 1090 -15990 1120 -15920
rect 1090 -16030 1120 -16020
rect 1820 -16230 1850 -15920
rect 1820 -16270 1850 -16260
rect 1910 -16230 1940 -15920
rect 1910 -16270 1940 -16260
rect 2030 -16350 2060 -15920
rect 2030 -16390 2060 -16380
rect 880 -17660 910 -17470
rect 970 -16590 1000 -16580
rect 970 -17660 1000 -16620
rect 1910 -16590 1940 -16580
rect 1700 -17080 1730 -17070
rect 1700 -17660 1730 -17110
rect 1910 -17800 1940 -16620
rect 2760 -16590 2790 -15710
rect 2970 -15990 3000 -15920
rect 2970 -16030 3000 -16020
rect 3700 -16230 3730 -15920
rect 3700 -16270 3730 -16260
rect 3790 -16230 3820 -15920
rect 3790 -16270 3820 -16260
rect 3910 -16470 3940 -15910
rect 3910 -16510 3940 -16500
rect 2760 -16630 2790 -16620
rect 2850 -16960 2880 -16950
rect 2640 -17080 2670 -17070
rect 2640 -17660 2670 -17110
rect 2760 -17080 2790 -17070
rect 2760 -17660 2790 -17110
rect 2850 -17660 2880 -16990
rect 3790 -16960 3820 -16950
rect 3580 -17080 3610 -17070
rect 3580 -17660 3610 -17110
rect 3790 -17800 3820 -16990
rect 4640 -16960 4670 -15710
rect 4850 -15990 4880 -15920
rect 4850 -16030 4880 -16020
rect 4640 -17000 4670 -16990
rect 4730 -16960 4760 -16950
rect 4520 -17080 4550 -17070
rect 4520 -17660 4550 -17110
rect 4640 -17320 4670 -17310
rect 4640 -17660 4670 -17350
rect 4730 -17660 4760 -16990
rect 5460 -17080 5490 -17070
rect 5460 -17660 5490 -17110
rect 5580 -17080 5610 -15920
rect 5670 -16230 5700 -15920
rect 5670 -16270 5700 -16260
rect 5790 -16470 5820 -15920
rect 5790 -16510 5820 -16500
rect 5580 -17120 5610 -17110
rect 5670 -16960 5700 -16950
rect 5670 -17800 5700 -16990
rect 6520 -16960 6550 -15710
rect 6730 -15990 6760 -15920
rect 6730 -16030 6760 -16020
rect 6520 -17000 6550 -16990
rect 6610 -16590 6640 -16580
rect 6400 -17080 6430 -17070
rect 6400 -17660 6430 -17110
rect 6520 -17320 6550 -17310
rect 6520 -17660 6550 -17350
rect 6610 -17660 6640 -16620
rect 7340 -17080 7370 -17070
rect 7340 -17660 7370 -17110
rect 7460 -17200 7490 -15920
rect 7550 -16230 7580 -15920
rect 7550 -16270 7580 -16260
rect 7670 -16350 7700 -15920
rect 7670 -16390 7700 -16380
rect 7460 -17240 7490 -17230
rect 7550 -16590 7580 -16580
rect 7550 -17800 7580 -16620
rect 8400 -16590 8430 -15710
rect 8400 -16630 8430 -16620
rect 8280 -17080 8310 -17070
rect 8280 -17660 8310 -17110
rect 8400 -17080 8430 -17070
rect 8400 -17660 8430 -17110
rect 8490 -17200 8520 -15920
rect 8610 -16110 8640 -15920
rect 8610 -16150 8640 -16140
rect 8490 -17800 8520 -17230
rect 9340 -17320 9370 -15710
rect 9220 -17440 9250 -17430
rect 9220 -17660 9250 -17470
rect 9340 -17660 9370 -17350
rect 9430 -16720 9460 -16710
rect 9430 -17660 9460 -16860
rect 9550 -17200 9580 -15910
rect 10280 -16720 10310 -15130
rect 10280 -16870 10310 -16860
rect 10370 -16720 10400 -15920
rect 10370 -16870 10400 -16860
rect 9550 -17240 9580 -17230
rect 11100 -17200 11130 -15920
rect 11100 -17240 11130 -17230
rect 11220 -16720 11250 -16710
rect 10160 -17320 10190 -17310
rect 10160 -17660 10190 -17350
rect 10490 -17320 10520 -17310
rect 10490 -17660 10520 -17350
rect 11220 -17660 11250 -16860
rect 11310 -17320 11340 -15710
rect 12040 -16110 12070 -15920
rect 12040 -16150 12070 -16140
rect 11310 -17660 11340 -17350
rect 12160 -17200 12190 -15920
rect 12250 -16590 12280 -15710
rect 12980 -16350 13010 -15920
rect 13100 -16230 13130 -15920
rect 13100 -16270 13130 -16260
rect 12980 -16390 13010 -16380
rect 12250 -16630 12280 -16620
rect 13100 -16590 13130 -16580
rect 11430 -17440 11460 -17430
rect 11430 -17660 11460 -17470
rect 12160 -17800 12190 -17230
rect 12250 -17080 12280 -17070
rect 12250 -17660 12280 -17110
rect 12370 -17080 12400 -17070
rect 12370 -17660 12400 -17110
rect 13100 -17800 13130 -16620
rect 13190 -17200 13220 -15920
rect 13920 -15990 13950 -15920
rect 13920 -16030 13950 -16020
rect 14040 -16590 14070 -16580
rect 13190 -17240 13220 -17230
rect 13310 -17080 13340 -17070
rect 13310 -17660 13340 -17110
rect 14040 -17660 14070 -16620
rect 14130 -16960 14160 -15710
rect 14860 -16470 14890 -15920
rect 14980 -16230 15010 -15920
rect 14980 -16270 15010 -16260
rect 14860 -16510 14890 -16500
rect 14130 -17000 14160 -16990
rect 14980 -16960 15010 -16950
rect 14250 -17080 14280 -17070
rect 14130 -17320 14160 -17310
rect 14130 -17660 14160 -17350
rect 14250 -17660 14280 -17110
rect 14980 -17800 15010 -16990
rect 15070 -17080 15100 -15920
rect 15800 -15990 15830 -15920
rect 15800 -16030 15830 -16020
rect 15920 -16960 15950 -16950
rect 15070 -17120 15100 -17110
rect 15190 -17080 15220 -17070
rect 15190 -17660 15220 -17110
rect 15920 -17660 15950 -16990
rect 16010 -16960 16040 -15710
rect 16740 -16470 16770 -15910
rect 16860 -16230 16890 -15920
rect 16860 -16270 16890 -16260
rect 16950 -16230 16980 -15920
rect 17680 -15990 17710 -15920
rect 17680 -16030 17710 -16020
rect 16950 -16270 16980 -16260
rect 16740 -16510 16770 -16500
rect 17890 -16590 17920 -15710
rect 18830 -15720 18860 -15710
rect 18620 -16350 18650 -15920
rect 18740 -16230 18770 -15920
rect 18740 -16270 18770 -16260
rect 18830 -16230 18860 -15920
rect 19560 -15990 19590 -15920
rect 19560 -16030 19590 -16020
rect 18830 -16270 18860 -16260
rect 18620 -16390 18650 -16380
rect 17890 -16630 17920 -16620
rect 18740 -16590 18770 -16580
rect 16010 -17000 16040 -16990
rect 16860 -16960 16890 -16950
rect 16130 -17080 16160 -17070
rect 16010 -17320 16040 -17310
rect 16010 -17660 16040 -17350
rect 16130 -17660 16160 -17110
rect 16860 -17800 16890 -16990
rect 17800 -16960 17830 -16950
rect 17070 -17080 17100 -17070
rect 17070 -17660 17100 -17110
rect 17800 -17660 17830 -16990
rect 17890 -17080 17920 -17070
rect 17890 -17660 17920 -17110
rect 18010 -17080 18040 -17070
rect 18010 -17660 18040 -17110
rect 18740 -17800 18770 -16620
rect 19680 -16590 19710 -16580
rect 18950 -17080 18980 -17070
rect 18950 -17660 18980 -17110
rect 19680 -17660 19710 -16620
rect 19770 -17440 19800 -15920
rect 20500 -15990 20530 -15920
rect 20500 -16030 20530 -16020
rect 20710 -15990 20740 -15710
rect 22490 -15870 22540 -15860
rect 22490 -15900 22500 -15870
rect 22530 -15900 22540 -15870
rect 22490 -15910 22540 -15900
rect 20710 -16030 20740 -16020
rect 21440 -16110 21470 -15920
rect 21440 -16150 21470 -16140
rect 21560 -16110 21590 -15920
rect 21650 -15990 21680 -15920
rect 21650 -16030 21680 -16020
rect 22380 -15990 22410 -15920
rect 22380 -16030 22410 -16020
rect 21560 -16150 21590 -16140
rect 19770 -17660 19800 -17470
rect 19890 -17440 19920 -17430
rect 19890 -17660 19920 -17470
rect 20620 -17560 20650 -17550
rect 20620 -17800 20650 -17590
rect 20830 -17560 20860 -17550
rect 20830 -17660 20860 -17590
rect 21560 -17560 21590 -17550
rect 21560 -17660 21590 -17590
rect 21770 -17560 21800 -17550
rect 21770 -17660 21800 -17590
rect 22500 -18830 22530 -15910
rect 23320 -15990 23350 -15890
rect 23320 -16030 23350 -16020
rect 24260 -16720 24420 -16710
rect 24260 -16860 24270 -16720
rect 24410 -16860 24420 -16720
rect 24260 -16870 24420 -16860
rect 22710 -17560 22740 -17550
rect 22710 -17660 22740 -17590
rect -1860 -18840 -1810 -18830
rect -1860 -18870 -1850 -18840
rect -1820 -18870 -1810 -18840
rect -1860 -18880 -1810 -18870
rect 22490 -18840 22540 -18830
rect 22490 -18870 22500 -18840
rect 22530 -18870 22540 -18840
rect 22490 -18880 22540 -18870
rect -1940 -19070 -1910 -19050
rect -6320 -20470 -6270 -20460
rect -6320 -20500 -6310 -20470
rect -6280 -20500 -6270 -20470
rect -6320 -20510 -6270 -20500
rect -6120 -20470 -6070 -20460
rect -6120 -20500 -6110 -20470
rect -6080 -20500 -6070 -20470
rect -6120 -20510 -6070 -20500
rect -5920 -20470 -5870 -20460
rect -5920 -20500 -5910 -20470
rect -5880 -20500 -5870 -20470
rect -5920 -20510 -5870 -20500
rect -5720 -20470 -5670 -20460
rect -5720 -20500 -5710 -20470
rect -5680 -20500 -5670 -20470
rect -5720 -20510 -5670 -20500
rect -5520 -20470 -5470 -20460
rect -5520 -20500 -5510 -20470
rect -5480 -20500 -5470 -20470
rect -5520 -20510 -5470 -20500
rect -5320 -20470 -5270 -20460
rect -5320 -20500 -5310 -20470
rect -5280 -20500 -5270 -20470
rect -5320 -20510 -5270 -20500
rect -5120 -20470 -5070 -20460
rect -5120 -20500 -5110 -20470
rect -5080 -20500 -5070 -20470
rect -5120 -20510 -5070 -20500
rect -4720 -20470 -4670 -20460
rect -4720 -20500 -4710 -20470
rect -4680 -20500 -4670 -20470
rect -4720 -20510 -4670 -20500
rect -4520 -20470 -4470 -20460
rect -4520 -20500 -4510 -20470
rect -4480 -20500 -4470 -20470
rect -4520 -20510 -4470 -20500
rect -4320 -20470 -4270 -20460
rect -4320 -20500 -4310 -20470
rect -4280 -20500 -4270 -20470
rect -4320 -20510 -4270 -20500
rect -4120 -20470 -4070 -20460
rect -4120 -20500 -4110 -20470
rect -4080 -20500 -4070 -20470
rect -4120 -20510 -4070 -20500
rect -3920 -20470 -3870 -20460
rect -3920 -20500 -3910 -20470
rect -3880 -20500 -3870 -20470
rect -3920 -20510 -3870 -20500
rect -3720 -20470 -3670 -20460
rect -3720 -20500 -3710 -20470
rect -3680 -20500 -3670 -20470
rect -3720 -20510 -3670 -20500
rect -3520 -20470 -3470 -20460
rect -3520 -20500 -3510 -20470
rect -3480 -20500 -3470 -20470
rect -3520 -20510 -3470 -20500
rect -6310 -20580 -6280 -20510
rect -6320 -20590 -6270 -20580
rect -6320 -20620 -6310 -20590
rect -6280 -20620 -6270 -20590
rect -6320 -20630 -6270 -20620
rect -6310 -20700 -6280 -20630
rect -6320 -20710 -6270 -20700
rect -6320 -20740 -6310 -20710
rect -6280 -20740 -6270 -20710
rect -6320 -20750 -6270 -20740
rect -6310 -20820 -6280 -20750
rect -6320 -20830 -6270 -20820
rect -6320 -20860 -6310 -20830
rect -6280 -20860 -6270 -20830
rect -6320 -20870 -6270 -20860
rect -6310 -20940 -6280 -20870
rect -6320 -20950 -6270 -20940
rect -6320 -20980 -6310 -20950
rect -6280 -20980 -6270 -20950
rect -6320 -20990 -6270 -20980
rect -6310 -21060 -6280 -20990
rect -6320 -21070 -6270 -21060
rect -6320 -21100 -6310 -21070
rect -6280 -21100 -6270 -21070
rect -6320 -21110 -6270 -21100
rect -6310 -21180 -6280 -21110
rect -6320 -21190 -6270 -21180
rect -6320 -21220 -6310 -21190
rect -6280 -21220 -6270 -21190
rect -6320 -21230 -6270 -21220
rect -6310 -21430 -6280 -21230
rect -6320 -21440 -6270 -21430
rect -6320 -21470 -6310 -21440
rect -6280 -21470 -6270 -21440
rect -6320 -21480 -6270 -21470
rect -6310 -21550 -6280 -21480
rect -6320 -21560 -6270 -21550
rect -6320 -21590 -6310 -21560
rect -6280 -21590 -6270 -21560
rect -6320 -21600 -6270 -21590
rect -6310 -21670 -6280 -21600
rect -6320 -21680 -6270 -21670
rect -6320 -21710 -6310 -21680
rect -6280 -21710 -6270 -21680
rect -6320 -21720 -6270 -21710
rect -6310 -21790 -6280 -21720
rect -6320 -21800 -6270 -21790
rect -6320 -21830 -6310 -21800
rect -6280 -21830 -6270 -21800
rect -6320 -21840 -6270 -21830
rect -6310 -21910 -6280 -21840
rect -6320 -21920 -6270 -21910
rect -6320 -21950 -6310 -21920
rect -6280 -21950 -6270 -21920
rect -6320 -21960 -6270 -21950
rect -6310 -22030 -6280 -21960
rect -6320 -22040 -6270 -22030
rect -6320 -22070 -6310 -22040
rect -6280 -22070 -6270 -22040
rect -6320 -22080 -6270 -22070
rect -6310 -22150 -6280 -22080
rect -6110 -22150 -6080 -20510
rect -5910 -22150 -5880 -20510
rect -5710 -22150 -5680 -20510
rect -5510 -22150 -5480 -20510
rect -5310 -22150 -5280 -20510
rect -5110 -22150 -5080 -20510
rect -4710 -22150 -4680 -20510
rect -4510 -22150 -4480 -20510
rect -4310 -22150 -4280 -20510
rect -4110 -22150 -4080 -20510
rect -3910 -22150 -3880 -20510
rect -3710 -22150 -3680 -20510
rect -3510 -22150 -3480 -20510
rect -2060 -20530 -2030 -20450
rect -1940 -20460 -1910 -19210
rect -1850 -18910 -1820 -18880
rect -1850 -19070 -1820 -19050
rect -1850 -19240 -1820 -19210
rect -910 -18910 -880 -18890
rect -910 -19070 -880 -19050
rect -910 -19230 -880 -19210
rect 970 -18910 1000 -18890
rect 970 -19070 1000 -19050
rect 970 -19230 1000 -19210
rect 2850 -18910 2880 -18890
rect 2850 -19070 2880 -19050
rect 2850 -19230 2880 -19210
rect 4730 -18910 4760 -18890
rect 4730 -19070 4760 -19050
rect 4730 -19230 4760 -19210
rect 6610 -18910 6640 -18890
rect 6610 -19070 6640 -19050
rect 6610 -19230 6640 -19210
rect 9430 -18910 9460 -18890
rect 9430 -19070 9460 -19050
rect 9430 -19230 9460 -19210
rect 11220 -18910 11250 -18890
rect 11220 -19070 11250 -19050
rect 11220 -19230 11250 -19210
rect 14040 -18910 14070 -18890
rect 14040 -19070 14070 -19050
rect 14040 -19230 14070 -19210
rect 15920 -18910 15950 -18890
rect 15920 -19070 15950 -19050
rect 15920 -19230 15950 -19210
rect 17800 -18910 17830 -18890
rect 17800 -19070 17830 -19050
rect 17800 -19230 17830 -19210
rect 19680 -18910 19710 -18890
rect 19680 -19070 19710 -19050
rect 19680 -19230 19710 -19210
rect 21560 -18910 21590 -18890
rect 21560 -19070 21590 -19050
rect 21560 -19230 21590 -19210
rect 22500 -18910 22530 -18880
rect 22500 -19070 22530 -19050
rect 22500 -19240 22530 -19210
rect 22590 -18910 22620 -18810
rect 22590 -19070 22620 -19050
rect -1860 -19250 -1810 -19240
rect -1860 -19280 -1850 -19250
rect -1820 -19280 -1810 -19250
rect -1860 -19290 -1810 -19280
rect 22490 -19250 22540 -19240
rect 22490 -19280 22500 -19250
rect 22530 -19280 22540 -19250
rect 22490 -19290 22540 -19280
rect -2060 -20570 -2030 -20560
rect -2670 -22100 -2640 -22090
rect -6320 -22160 -6270 -22150
rect -6320 -22190 -6310 -22160
rect -6280 -22190 -6270 -22160
rect -6320 -22200 -6270 -22190
rect -6120 -22160 -6070 -22150
rect -6120 -22190 -6110 -22160
rect -6080 -22190 -6070 -22160
rect -6120 -22200 -6070 -22190
rect -5920 -22160 -5870 -22150
rect -5920 -22190 -5910 -22160
rect -5880 -22190 -5870 -22160
rect -5920 -22200 -5870 -22190
rect -5720 -22160 -5670 -22150
rect -5720 -22190 -5710 -22160
rect -5680 -22190 -5670 -22160
rect -5720 -22200 -5670 -22190
rect -5520 -22160 -5470 -22150
rect -5520 -22190 -5510 -22160
rect -5480 -22190 -5470 -22160
rect -5520 -22200 -5470 -22190
rect -5320 -22160 -5270 -22150
rect -5320 -22190 -5310 -22160
rect -5280 -22190 -5270 -22160
rect -5320 -22200 -5270 -22190
rect -5120 -22160 -5070 -22150
rect -5120 -22190 -5110 -22160
rect -5080 -22190 -5070 -22160
rect -5120 -22200 -5070 -22190
rect -4720 -22160 -4670 -22150
rect -4720 -22190 -4710 -22160
rect -4680 -22190 -4670 -22160
rect -4720 -22200 -4670 -22190
rect -4520 -22160 -4470 -22150
rect -4520 -22190 -4510 -22160
rect -4480 -22190 -4470 -22160
rect -4520 -22200 -4470 -22190
rect -4320 -22160 -4270 -22150
rect -4320 -22190 -4310 -22160
rect -4280 -22190 -4270 -22160
rect -4320 -22200 -4270 -22190
rect -4120 -22160 -4070 -22150
rect -4120 -22190 -4110 -22160
rect -4080 -22190 -4070 -22160
rect -4120 -22200 -4070 -22190
rect -3920 -22160 -3870 -22150
rect -3920 -22190 -3910 -22160
rect -3880 -22190 -3870 -22160
rect -3920 -22200 -3870 -22190
rect -3720 -22160 -3670 -22150
rect -3720 -22190 -3710 -22160
rect -3680 -22190 -3670 -22160
rect -3720 -22200 -3670 -22190
rect -3520 -22160 -3470 -22150
rect -3520 -22190 -3510 -22160
rect -3480 -22190 -3470 -22160
rect -3520 -22200 -3470 -22190
rect -2670 -22200 -2640 -22130
rect -6310 -28520 -6280 -22200
rect -6110 -28520 -6080 -22200
rect -5910 -28520 -5880 -22200
rect -5710 -28520 -5680 -22200
rect -5510 -28520 -5480 -22200
rect -5310 -28520 -5280 -22200
rect -5110 -28520 -5080 -22200
rect -4710 -28520 -4680 -22200
rect -4510 -28520 -4480 -22200
rect -4310 -28520 -4280 -22200
rect -4110 -28520 -4080 -22200
rect -3910 -28520 -3880 -22200
rect -3710 -28520 -3680 -22200
rect -3510 -28520 -3480 -22200
rect -2790 -25190 -2760 -22200
rect -1850 -22210 -1820 -19290
rect -1120 -20530 -1090 -20460
rect -1120 -20570 -1090 -20560
rect -910 -20530 -880 -20460
rect -910 -20570 -880 -20560
rect -180 -20530 -150 -20460
rect -180 -20570 -150 -20560
rect 30 -20530 60 -20320
rect 30 -20570 60 -20560
rect 760 -20650 790 -20460
rect 760 -20690 790 -20680
rect 880 -20650 910 -20460
rect -910 -21980 -880 -21970
rect -1730 -22100 -1700 -22090
rect -1730 -22200 -1700 -22130
rect -1000 -22100 -970 -22090
rect -1000 -22200 -970 -22130
rect -910 -22200 -880 -22010
rect -790 -21980 -760 -21970
rect -790 -22200 -760 -22010
rect -60 -22100 -30 -22090
rect -1860 -22220 -1810 -22210
rect -1860 -22250 -1850 -22220
rect -1820 -22250 -1810 -22220
rect -1860 -22260 -1810 -22250
rect -60 -22410 -30 -22130
rect 150 -22100 180 -22090
rect 150 -22200 180 -22130
rect 880 -22200 910 -20680
rect 970 -21500 1000 -20460
rect 1700 -21010 1730 -20460
rect 1700 -21050 1730 -21040
rect 970 -21540 1000 -21530
rect 1910 -21500 1940 -20320
rect 2640 -21010 2670 -20460
rect 2640 -21050 2670 -21040
rect 2760 -21010 2790 -20460
rect 2760 -21050 2790 -21040
rect 2850 -21130 2880 -20460
rect 3580 -21010 3610 -20460
rect 3580 -21050 3610 -21040
rect 2850 -21170 2880 -21160
rect 3790 -21130 3820 -20320
rect 4520 -21010 4550 -20460
rect 4640 -20770 4670 -20460
rect 4640 -20810 4670 -20800
rect 4520 -21050 4550 -21040
rect 3790 -21170 3820 -21160
rect 4640 -21130 4670 -21120
rect 1910 -21540 1940 -21530
rect 2760 -21500 2790 -21490
rect 2030 -21740 2060 -21730
rect 1820 -21860 1850 -21850
rect 1090 -22100 1120 -22090
rect 1090 -22200 1120 -22130
rect 1820 -22200 1850 -21890
rect 1910 -21860 1940 -21850
rect 1910 -22200 1940 -21890
rect 2030 -22200 2060 -21770
rect 1820 -22410 1850 -22400
rect 2760 -22410 2790 -21530
rect 3910 -21620 3940 -21610
rect 3700 -21860 3730 -21850
rect 2970 -22100 3000 -22090
rect 2970 -22200 3000 -22130
rect 3700 -22200 3730 -21890
rect 3790 -21860 3820 -21850
rect 3790 -22200 3820 -21890
rect 3910 -22210 3940 -21650
rect 4640 -22410 4670 -21160
rect 4730 -21130 4760 -20460
rect 5460 -21010 5490 -20460
rect 5460 -21050 5490 -21040
rect 5580 -21010 5610 -21000
rect 4730 -21170 4760 -21160
rect 4850 -22100 4880 -22090
rect 4850 -22200 4880 -22130
rect 5580 -22200 5610 -21040
rect 5670 -21130 5700 -20320
rect 6400 -21010 6430 -20460
rect 6520 -20770 6550 -20460
rect 6520 -20810 6550 -20800
rect 6400 -21050 6430 -21040
rect 5670 -21170 5700 -21160
rect 6520 -21130 6550 -21120
rect 5790 -21620 5820 -21610
rect 5670 -21860 5700 -21850
rect 5670 -22200 5700 -21890
rect 5790 -22200 5820 -21650
rect 6520 -22410 6550 -21160
rect 6610 -21500 6640 -20460
rect 7340 -21010 7370 -20460
rect 7340 -21050 7370 -21040
rect 7460 -20890 7490 -20880
rect 6610 -21540 6640 -21530
rect 6730 -22100 6760 -22090
rect 6730 -22200 6760 -22130
rect 7460 -22200 7490 -20920
rect 7550 -21500 7580 -20320
rect 8280 -21010 8310 -20460
rect 8280 -21050 8310 -21040
rect 8400 -21010 8430 -20460
rect 8400 -21050 8430 -21040
rect 8490 -20890 8520 -20320
rect 9220 -20650 9250 -20460
rect 9220 -20690 9250 -20680
rect 7550 -21540 7580 -21530
rect 8400 -21500 8430 -21490
rect 7670 -21740 7700 -21730
rect 7550 -21860 7580 -21850
rect 7550 -22200 7580 -21890
rect 7670 -22200 7700 -21770
rect 8400 -22410 8430 -21530
rect 8490 -22200 8520 -20920
rect 9340 -20770 9370 -20460
rect 8610 -21980 8640 -21970
rect 8610 -22200 8640 -22010
rect 9340 -22410 9370 -20800
rect 9430 -21260 9460 -20460
rect 10160 -20770 10190 -20460
rect 10160 -20810 10190 -20800
rect 10490 -20770 10520 -20460
rect 10490 -20810 10520 -20800
rect 9430 -21410 9460 -21400
rect 9550 -20890 9580 -20880
rect 9550 -22210 9580 -20920
rect 11100 -20890 11130 -20880
rect 10280 -21260 10310 -21250
rect 10280 -22990 10310 -21400
rect 10370 -21260 10400 -21250
rect 10370 -22200 10400 -21400
rect 11100 -22200 11130 -20920
rect 11220 -21260 11250 -20460
rect 11220 -21410 11250 -21400
rect 11310 -20770 11340 -20460
rect 11430 -20650 11460 -20460
rect 11430 -20690 11460 -20680
rect 11310 -22410 11340 -20800
rect 12160 -20890 12190 -20320
rect 12040 -21980 12070 -21970
rect 12040 -22200 12070 -22010
rect 12160 -22200 12190 -20920
rect 12250 -21010 12280 -20460
rect 12250 -21050 12280 -21040
rect 12370 -21010 12400 -20460
rect 12370 -21050 12400 -21040
rect 12250 -21500 12280 -21490
rect 12250 -22410 12280 -21530
rect 13100 -21500 13130 -20320
rect 13100 -21540 13130 -21530
rect 13190 -20890 13220 -20880
rect 12980 -21740 13010 -21730
rect 12980 -22200 13010 -21770
rect 13100 -21860 13130 -21850
rect 13100 -22200 13130 -21890
rect 13190 -22200 13220 -20920
rect 13310 -21010 13340 -20460
rect 13310 -21050 13340 -21040
rect 14040 -21500 14070 -20460
rect 14130 -20770 14160 -20460
rect 14130 -20810 14160 -20800
rect 14250 -21010 14280 -20460
rect 14250 -21050 14280 -21040
rect 14040 -21540 14070 -21530
rect 14130 -21130 14160 -21120
rect 13920 -22100 13950 -22090
rect 13920 -22200 13950 -22130
rect 14130 -22410 14160 -21160
rect 14980 -21130 15010 -20320
rect 14980 -21170 15010 -21160
rect 15070 -21010 15100 -21000
rect 14860 -21620 14890 -21610
rect 14860 -22200 14890 -21650
rect 14980 -21860 15010 -21850
rect 14980 -22200 15010 -21890
rect 15070 -22200 15100 -21040
rect 15190 -21010 15220 -20460
rect 15190 -21050 15220 -21040
rect 15920 -21130 15950 -20460
rect 16010 -20770 16040 -20460
rect 16010 -20810 16040 -20800
rect 16130 -21010 16160 -20460
rect 16130 -21050 16160 -21040
rect 15920 -21170 15950 -21160
rect 16010 -21130 16040 -21120
rect 15800 -22100 15830 -22090
rect 15800 -22200 15830 -22130
rect 16010 -22410 16040 -21160
rect 16860 -21130 16890 -20320
rect 17070 -21010 17100 -20460
rect 17070 -21050 17100 -21040
rect 16860 -21170 16890 -21160
rect 17800 -21130 17830 -20460
rect 17890 -21010 17920 -20460
rect 17890 -21050 17920 -21040
rect 18010 -21010 18040 -20460
rect 18010 -21050 18040 -21040
rect 17800 -21170 17830 -21160
rect 17890 -21500 17920 -21490
rect 16740 -21620 16770 -21610
rect 16740 -22210 16770 -21650
rect 16860 -21860 16890 -21850
rect 16860 -22200 16890 -21890
rect 16950 -21860 16980 -21850
rect 16950 -22200 16980 -21890
rect 17680 -22100 17710 -22090
rect 17680 -22200 17710 -22130
rect 17890 -22410 17920 -21530
rect 18740 -21500 18770 -20320
rect 18950 -21010 18980 -20460
rect 18950 -21050 18980 -21040
rect 18740 -21540 18770 -21530
rect 19680 -21500 19710 -20460
rect 19680 -21540 19710 -21530
rect 19770 -20650 19800 -20460
rect 18620 -21740 18650 -21730
rect 18620 -22200 18650 -21770
rect 18740 -21860 18770 -21850
rect 18740 -22200 18770 -21890
rect 18830 -21860 18860 -21850
rect 18830 -22200 18860 -21890
rect 19560 -22100 19590 -22090
rect 19560 -22200 19590 -22130
rect 19770 -22200 19800 -20680
rect 19890 -20650 19920 -20460
rect 20620 -20530 20650 -20320
rect 20620 -20570 20650 -20560
rect 20830 -20530 20860 -20460
rect 20830 -20570 20860 -20560
rect 21560 -20530 21590 -20460
rect 21560 -20570 21590 -20560
rect 21770 -20530 21800 -20460
rect 21770 -20570 21800 -20560
rect 19890 -20690 19920 -20680
rect 21440 -21980 21470 -21970
rect 20500 -22100 20530 -22090
rect 20500 -22200 20530 -22130
rect 20710 -22100 20740 -22090
rect 18830 -22410 18860 -22400
rect 20710 -22410 20740 -22130
rect 21440 -22200 21470 -22010
rect 21560 -21980 21590 -21970
rect 21560 -22200 21590 -22010
rect 21650 -22100 21680 -22090
rect 21650 -22200 21680 -22130
rect 22380 -22100 22410 -22090
rect 22380 -22200 22410 -22130
rect 22500 -22210 22530 -19290
rect 22590 -19310 22620 -19210
rect 23440 -18910 23470 -18890
rect 23440 -19070 23470 -19050
rect 23440 -19230 23470 -19210
rect 22710 -20530 22740 -20460
rect 22710 -20570 22740 -20560
rect 24260 -21260 24420 -21250
rect 24260 -21400 24270 -21260
rect 24410 -21400 24420 -21260
rect 24260 -21410 24420 -21400
rect 23320 -22100 23350 -22090
rect 22490 -22220 22540 -22210
rect 22490 -22250 22500 -22220
rect 22530 -22250 22540 -22220
rect 23320 -22230 23350 -22130
rect 22490 -22260 22540 -22250
rect -1010 -25050 -960 -25040
rect -1010 -25080 -1000 -25050
rect -970 -25080 -960 -25050
rect -1010 -25090 -960 -25080
rect 21640 -25050 21690 -25040
rect 21640 -25080 21650 -25050
rect 21680 -25080 21690 -25050
rect 21640 -25090 21690 -25080
rect -2790 -25340 -2760 -25330
rect -1940 -25190 -1910 -25170
rect -1940 -25340 -1910 -25330
rect -1000 -25190 -970 -25170
rect -1000 -25340 -970 -25330
rect 880 -25190 910 -25110
rect 880 -25340 910 -25330
rect 1820 -25190 1850 -25110
rect 1820 -25340 1850 -25330
rect 3700 -25190 3730 -25170
rect 3700 -25340 3730 -25330
rect 5580 -25190 5610 -25170
rect 5580 -25340 5610 -25330
rect 7460 -25190 7490 -25170
rect 7460 -25340 7490 -25330
rect 10280 -25190 10310 -25170
rect 10280 -25340 10310 -25330
rect 10370 -25190 10400 -25170
rect 10370 -25340 10400 -25330
rect 13190 -25190 13220 -25170
rect 13190 -25340 13220 -25330
rect 15070 -25190 15100 -25170
rect 15070 -25340 15100 -25330
rect 16950 -25190 16980 -25170
rect 16950 -25340 16980 -25330
rect 18830 -25190 18860 -25110
rect 18830 -25340 18860 -25330
rect 19770 -25190 19800 -25110
rect 19770 -25340 19800 -25330
rect 21650 -25190 21680 -25170
rect 21650 -25340 21680 -25330
rect 22590 -25190 22620 -25170
rect 22590 -25340 22620 -25330
rect 23440 -25190 23470 -25020
rect 23440 -25340 23470 -25330
<< via1 >>
rect -2790 -370 -2760 -230
rect -1940 -370 -1910 -230
rect -1000 -370 -970 -230
rect 880 -370 910 -230
rect 1820 -370 1850 -230
rect 3700 -370 3730 -230
rect 5580 -370 5610 -230
rect 7460 -370 7490 -230
rect 10280 -370 10310 -230
rect 10370 -370 10400 -230
rect 13190 -370 13220 -230
rect 15070 -370 15100 -230
rect 16950 -370 16980 -230
rect 18830 -370 18860 -230
rect 19770 -370 19800 -230
rect 21650 -370 21680 -230
rect 22590 -370 22620 -230
rect 23440 -370 23470 -230
rect -6310 -3400 -6280 -3370
rect -6110 -3400 -6080 -3370
rect -5910 -3400 -5880 -3370
rect -5710 -3400 -5680 -3370
rect -5510 -3400 -5480 -3370
rect -5310 -3400 -5280 -3370
rect -5110 -3400 -5080 -3370
rect -4710 -3400 -4680 -3370
rect -4510 -3400 -4480 -3370
rect -4310 -3400 -4280 -3370
rect -4110 -3400 -4080 -3370
rect -3910 -3400 -3880 -3370
rect -3710 -3400 -3680 -3370
rect -3510 -3400 -3480 -3370
rect -6310 -3520 -6280 -3490
rect -6310 -3640 -6280 -3610
rect -6310 -3760 -6280 -3730
rect -6310 -3880 -6280 -3850
rect -6310 -4000 -6280 -3970
rect -6310 -4120 -6280 -4090
rect -6310 -4370 -6280 -4340
rect -6310 -4490 -6280 -4460
rect -6310 -4610 -6280 -4580
rect -6310 -4730 -6280 -4700
rect -6310 -4850 -6280 -4820
rect -6310 -4970 -6280 -4940
rect -2670 -3460 -2640 -3430
rect -2060 -5030 -2030 -5000
rect -6310 -5090 -6280 -5060
rect -6110 -5090 -6080 -5060
rect -5910 -5090 -5880 -5060
rect -5710 -5090 -5680 -5060
rect -5510 -5090 -5480 -5060
rect -5310 -5090 -5280 -5060
rect -5110 -5090 -5080 -5060
rect -4710 -5090 -4680 -5060
rect -4510 -5090 -4480 -5060
rect -4310 -5090 -4280 -5060
rect -4110 -5090 -4080 -5060
rect -3910 -5090 -3880 -5060
rect -3710 -5090 -3680 -5060
rect -3510 -5090 -3480 -5060
rect -2790 -6490 -2760 -6350
rect -2790 -6650 -2760 -6510
rect -1730 -3460 -1700 -3430
rect -1000 -3460 -970 -3430
rect -910 -3580 -880 -3550
rect -60 -3460 -30 -3430
rect 150 -3460 180 -3430
rect -790 -3580 -760 -3550
rect 760 -4910 790 -4880
rect -1120 -5030 -1090 -5000
rect -910 -5030 -880 -5000
rect -180 -5030 -150 -5000
rect 30 -5030 60 -5000
rect 1090 -3460 1120 -3430
rect 1820 -3700 1850 -3670
rect 1910 -3700 1940 -3670
rect 2030 -3820 2060 -3790
rect 880 -4910 910 -4880
rect 970 -4060 1000 -4030
rect 1910 -4060 1940 -4030
rect 1700 -4550 1730 -4520
rect 2970 -3460 3000 -3430
rect 3700 -3700 3730 -3670
rect 3790 -3700 3820 -3670
rect 3910 -3940 3940 -3910
rect 2760 -4060 2790 -4030
rect 2850 -4430 2880 -4400
rect 2640 -4550 2670 -4520
rect 2760 -4550 2790 -4520
rect 3790 -4430 3820 -4400
rect 3580 -4550 3610 -4520
rect 4850 -3460 4880 -3430
rect 4640 -4430 4670 -4400
rect 4730 -4430 4760 -4400
rect 4520 -4550 4550 -4520
rect 4640 -4790 4670 -4760
rect 5460 -4550 5490 -4520
rect 5670 -3700 5700 -3670
rect 5790 -3940 5820 -3910
rect 5580 -4550 5610 -4520
rect 5670 -4430 5700 -4400
rect 6730 -3460 6760 -3430
rect 6520 -4430 6550 -4400
rect 6610 -4060 6640 -4030
rect 6400 -4550 6430 -4520
rect 6520 -4790 6550 -4760
rect 7340 -4550 7370 -4520
rect 7550 -3700 7580 -3670
rect 7670 -3820 7700 -3790
rect 7460 -4670 7490 -4640
rect 7550 -4060 7580 -4030
rect 8400 -4060 8430 -4030
rect 8280 -4550 8310 -4520
rect 8400 -4550 8430 -4520
rect 8610 -3580 8640 -3550
rect 8490 -4670 8520 -4640
rect 9340 -4790 9370 -4760
rect 9220 -4910 9250 -4880
rect 9430 -4300 9460 -4160
rect 10280 -4300 10310 -4160
rect 10370 -4300 10400 -4160
rect 9550 -4670 9580 -4640
rect 11100 -4670 11130 -4640
rect 11220 -4300 11250 -4160
rect 10160 -4790 10190 -4760
rect 10490 -4790 10520 -4760
rect 12040 -3580 12070 -3550
rect 11310 -4790 11340 -4760
rect 13100 -3700 13130 -3670
rect 12980 -3820 13010 -3790
rect 12250 -4060 12280 -4030
rect 13100 -4060 13130 -4030
rect 12160 -4670 12190 -4640
rect 11430 -4910 11460 -4880
rect 12250 -4550 12280 -4520
rect 12370 -4550 12400 -4520
rect 13920 -3460 13950 -3430
rect 14040 -4060 14070 -4030
rect 13190 -4670 13220 -4640
rect 13310 -4550 13340 -4520
rect 14980 -3700 15010 -3670
rect 14860 -3940 14890 -3910
rect 14130 -4430 14160 -4400
rect 14980 -4430 15010 -4400
rect 14250 -4550 14280 -4520
rect 14130 -4790 14160 -4760
rect 15800 -3460 15830 -3430
rect 15920 -4430 15950 -4400
rect 15070 -4550 15100 -4520
rect 15190 -4550 15220 -4520
rect 16860 -3700 16890 -3670
rect 17680 -3460 17710 -3430
rect 16950 -3700 16980 -3670
rect 16740 -3940 16770 -3910
rect 18740 -3700 18770 -3670
rect 19560 -3460 19590 -3430
rect 18830 -3700 18860 -3670
rect 18620 -3820 18650 -3790
rect 17890 -4060 17920 -4030
rect 18740 -4060 18770 -4030
rect 16010 -4430 16040 -4400
rect 16860 -4430 16890 -4400
rect 16130 -4550 16160 -4520
rect 16010 -4790 16040 -4760
rect 17800 -4430 17830 -4400
rect 17070 -4550 17100 -4520
rect 17890 -4550 17920 -4520
rect 18010 -4550 18040 -4520
rect 19680 -4060 19710 -4030
rect 18950 -4550 18980 -4520
rect 20500 -3460 20530 -3430
rect 20710 -3460 20740 -3430
rect 21440 -3580 21470 -3550
rect 21650 -3460 21680 -3430
rect 22380 -3460 22410 -3430
rect 21560 -3580 21590 -3550
rect 19770 -4910 19800 -4880
rect 19890 -4910 19920 -4880
rect 20620 -5030 20650 -5000
rect 20830 -5030 20860 -5000
rect 21560 -5030 21590 -5000
rect 21770 -5030 21800 -5000
rect 23320 -3460 23350 -3430
rect 24270 -4300 24410 -4160
rect 22710 -5030 22740 -5000
rect -1940 -6490 -1910 -6350
rect -1940 -6650 -1910 -6510
rect -6310 -7940 -6280 -7910
rect -6110 -7940 -6080 -7910
rect -5910 -7940 -5880 -7910
rect -5710 -7940 -5680 -7910
rect -5510 -7940 -5480 -7910
rect -5310 -7940 -5280 -7910
rect -5110 -7940 -5080 -7910
rect -4710 -7940 -4680 -7910
rect -4510 -7940 -4480 -7910
rect -4310 -7940 -4280 -7910
rect -4110 -7940 -4080 -7910
rect -3910 -7940 -3880 -7910
rect -3710 -7940 -3680 -7910
rect -3510 -7940 -3480 -7910
rect -6310 -8060 -6280 -8030
rect -6310 -8180 -6280 -8150
rect -6310 -8300 -6280 -8270
rect -6310 -8420 -6280 -8390
rect -6310 -8540 -6280 -8510
rect -6310 -8660 -6280 -8630
rect -6310 -8910 -6280 -8880
rect -6310 -9030 -6280 -9000
rect -6310 -9150 -6280 -9120
rect -6310 -9270 -6280 -9240
rect -6310 -9390 -6280 -9360
rect -6310 -9510 -6280 -9480
rect -1850 -6490 -1820 -6350
rect -1850 -6650 -1820 -6510
rect -910 -6490 -880 -6350
rect -910 -6650 -880 -6510
rect 970 -6490 1000 -6350
rect 970 -6650 1000 -6510
rect 2850 -6490 2880 -6350
rect 2850 -6650 2880 -6510
rect 4730 -6490 4760 -6350
rect 4730 -6650 4760 -6510
rect 6610 -6490 6640 -6350
rect 6610 -6650 6640 -6510
rect 9430 -6490 9460 -6350
rect 9430 -6650 9460 -6510
rect 11220 -6490 11250 -6350
rect 11220 -6650 11250 -6510
rect 14040 -6490 14070 -6350
rect 14040 -6650 14070 -6510
rect 15920 -6490 15950 -6350
rect 15920 -6650 15950 -6510
rect 17800 -6490 17830 -6350
rect 17800 -6650 17830 -6510
rect 19680 -6490 19710 -6350
rect 19680 -6650 19710 -6510
rect 21560 -6490 21590 -6350
rect 21560 -6650 21590 -6510
rect 22500 -6490 22530 -6350
rect 22500 -6650 22530 -6510
rect 22590 -6490 22620 -6350
rect 22590 -6650 22620 -6510
rect -2060 -8000 -2030 -7970
rect -2670 -9570 -2640 -9540
rect -6310 -9630 -6280 -9600
rect -6110 -9630 -6080 -9600
rect -5910 -9630 -5880 -9600
rect -5710 -9630 -5680 -9600
rect -5510 -9630 -5480 -9600
rect -5310 -9630 -5280 -9600
rect -5110 -9630 -5080 -9600
rect -4710 -9630 -4680 -9600
rect -4510 -9630 -4480 -9600
rect -4310 -9630 -4280 -9600
rect -4110 -9630 -4080 -9600
rect -3910 -9630 -3880 -9600
rect -3710 -9630 -3680 -9600
rect -3510 -9630 -3480 -9600
rect -1120 -8000 -1090 -7970
rect -910 -8000 -880 -7970
rect -180 -8000 -150 -7970
rect 30 -8000 60 -7970
rect 760 -8120 790 -8090
rect 880 -8120 910 -8090
rect -910 -9450 -880 -9420
rect -1730 -9570 -1700 -9540
rect -1000 -9570 -970 -9540
rect -790 -9450 -760 -9420
rect -60 -9570 -30 -9540
rect 150 -9570 180 -9540
rect 1700 -8480 1730 -8450
rect 970 -8970 1000 -8940
rect 2640 -8480 2670 -8450
rect 2760 -8480 2790 -8450
rect 3580 -8480 3610 -8450
rect 2850 -8600 2880 -8570
rect 4640 -8240 4670 -8210
rect 4520 -8480 4550 -8450
rect 3790 -8600 3820 -8570
rect 4640 -8600 4670 -8570
rect 1910 -8970 1940 -8940
rect 2760 -8970 2790 -8940
rect 2030 -9210 2060 -9180
rect 1820 -9330 1850 -9300
rect 1090 -9570 1120 -9540
rect 1910 -9330 1940 -9300
rect 3910 -9090 3940 -9060
rect 3700 -9330 3730 -9300
rect 2970 -9570 3000 -9540
rect 3790 -9330 3820 -9300
rect 5460 -8480 5490 -8450
rect 5580 -8480 5610 -8450
rect 4730 -8600 4760 -8570
rect 4850 -9570 4880 -9540
rect 6520 -8240 6550 -8210
rect 6400 -8480 6430 -8450
rect 5670 -8600 5700 -8570
rect 6520 -8600 6550 -8570
rect 5790 -9090 5820 -9060
rect 5670 -9330 5700 -9300
rect 7340 -8480 7370 -8450
rect 7460 -8360 7490 -8330
rect 6610 -8970 6640 -8940
rect 6730 -9570 6760 -9540
rect 8280 -8480 8310 -8450
rect 8400 -8480 8430 -8450
rect 9220 -8120 9250 -8090
rect 8490 -8360 8520 -8330
rect 7550 -8970 7580 -8940
rect 8400 -8970 8430 -8940
rect 7670 -9210 7700 -9180
rect 7550 -9330 7580 -9300
rect 9340 -8240 9370 -8210
rect 8610 -9450 8640 -9420
rect 10160 -8240 10190 -8210
rect 10490 -8240 10520 -8210
rect 9430 -8840 9460 -8700
rect 9550 -8360 9580 -8330
rect 11100 -8360 11130 -8330
rect 10280 -8840 10310 -8700
rect 10370 -8840 10400 -8700
rect 11220 -8840 11250 -8700
rect 11430 -8120 11460 -8090
rect 11310 -8240 11340 -8210
rect 12160 -8360 12190 -8330
rect 12040 -9450 12070 -9420
rect 12250 -8480 12280 -8450
rect 12370 -8480 12400 -8450
rect 12250 -8970 12280 -8940
rect 13100 -8970 13130 -8940
rect 13190 -8360 13220 -8330
rect 12980 -9210 13010 -9180
rect 13100 -9330 13130 -9300
rect 13310 -8480 13340 -8450
rect 14130 -8240 14160 -8210
rect 14250 -8480 14280 -8450
rect 14040 -8970 14070 -8940
rect 14130 -8600 14160 -8570
rect 13920 -9570 13950 -9540
rect 14980 -8600 15010 -8570
rect 15070 -8480 15100 -8450
rect 14860 -9090 14890 -9060
rect 14980 -9330 15010 -9300
rect 15190 -8480 15220 -8450
rect 16010 -8240 16040 -8210
rect 16130 -8480 16160 -8450
rect 15920 -8600 15950 -8570
rect 16010 -8600 16040 -8570
rect 15800 -9570 15830 -9540
rect 17070 -8480 17100 -8450
rect 16860 -8600 16890 -8570
rect 17890 -8480 17920 -8450
rect 18010 -8480 18040 -8450
rect 17800 -8600 17830 -8570
rect 17890 -8970 17920 -8940
rect 16740 -9090 16770 -9060
rect 16860 -9330 16890 -9300
rect 16950 -9330 16980 -9300
rect 17680 -9570 17710 -9540
rect 18950 -8480 18980 -8450
rect 18740 -8970 18770 -8940
rect 19680 -8970 19710 -8940
rect 19770 -8120 19800 -8090
rect 18620 -9210 18650 -9180
rect 18740 -9330 18770 -9300
rect 18830 -9330 18860 -9300
rect 19560 -9570 19590 -9540
rect 20620 -8000 20650 -7970
rect 20830 -8000 20860 -7970
rect 21560 -8000 21590 -7970
rect 21770 -8000 21800 -7970
rect 19890 -8120 19920 -8090
rect 21440 -9450 21470 -9420
rect 20500 -9570 20530 -9540
rect 20710 -9570 20740 -9540
rect 21560 -9450 21590 -9420
rect 21650 -9570 21680 -9540
rect 22380 -9570 22410 -9540
rect 23440 -6490 23470 -6350
rect 23440 -6650 23470 -6510
rect 22710 -8000 22740 -7970
rect 24270 -8840 24410 -8700
rect 23320 -9570 23350 -9540
rect -2790 -12770 -2760 -12630
rect -2790 -12930 -2760 -12790
rect -1940 -12770 -1910 -12630
rect -1940 -12930 -1910 -12790
rect -1000 -12770 -970 -12630
rect -1000 -12930 -970 -12790
rect 880 -12770 910 -12630
rect 880 -12930 910 -12790
rect 1820 -12770 1850 -12630
rect 1820 -12930 1850 -12790
rect 3700 -12770 3730 -12630
rect 3700 -12930 3730 -12790
rect 5580 -12770 5610 -12630
rect 5580 -12930 5610 -12790
rect 7460 -12770 7490 -12630
rect 7460 -12930 7490 -12790
rect 10280 -12770 10310 -12630
rect 10280 -12930 10310 -12790
rect 10370 -12770 10400 -12630
rect 10370 -12930 10400 -12790
rect 13190 -12770 13220 -12630
rect 13190 -12930 13220 -12790
rect 15070 -12770 15100 -12630
rect 15070 -12930 15100 -12790
rect 16950 -12770 16980 -12630
rect 16950 -12930 16980 -12790
rect 18830 -12770 18860 -12630
rect 18830 -12930 18860 -12790
rect 19770 -12770 19800 -12630
rect 19770 -12930 19800 -12790
rect 21650 -12770 21680 -12630
rect 21650 -12930 21680 -12790
rect 22590 -12770 22620 -12630
rect 22590 -12930 22620 -12790
rect 23440 -12770 23470 -12630
rect 23440 -12930 23470 -12790
rect -6310 -15960 -6280 -15930
rect -6110 -15960 -6080 -15930
rect -5910 -15960 -5880 -15930
rect -5710 -15960 -5680 -15930
rect -5510 -15960 -5480 -15930
rect -5310 -15960 -5280 -15930
rect -5110 -15960 -5080 -15930
rect -4710 -15960 -4680 -15930
rect -4510 -15960 -4480 -15930
rect -4310 -15960 -4280 -15930
rect -4110 -15960 -4080 -15930
rect -3910 -15960 -3880 -15930
rect -3710 -15960 -3680 -15930
rect -3510 -15960 -3480 -15930
rect -6310 -16080 -6280 -16050
rect -6310 -16200 -6280 -16170
rect -6310 -16320 -6280 -16290
rect -6310 -16440 -6280 -16410
rect -6310 -16560 -6280 -16530
rect -6310 -16680 -6280 -16650
rect -6310 -16930 -6280 -16900
rect -6310 -17050 -6280 -17020
rect -6310 -17170 -6280 -17140
rect -6310 -17290 -6280 -17260
rect -6310 -17410 -6280 -17380
rect -6310 -17530 -6280 -17500
rect -2670 -16020 -2640 -15990
rect -2060 -17590 -2030 -17560
rect -6310 -17650 -6280 -17620
rect -6110 -17650 -6080 -17620
rect -5910 -17650 -5880 -17620
rect -5710 -17650 -5680 -17620
rect -5510 -17650 -5480 -17620
rect -5310 -17650 -5280 -17620
rect -5110 -17650 -5080 -17620
rect -4710 -17650 -4680 -17620
rect -4510 -17650 -4480 -17620
rect -4310 -17650 -4280 -17620
rect -4110 -17650 -4080 -17620
rect -3910 -17650 -3880 -17620
rect -3710 -17650 -3680 -17620
rect -3510 -17650 -3480 -17620
rect -2790 -19050 -2760 -18910
rect -2790 -19210 -2760 -19070
rect -1730 -16020 -1700 -15990
rect -1000 -16020 -970 -15990
rect -910 -16140 -880 -16110
rect -60 -16020 -30 -15990
rect 150 -16020 180 -15990
rect -790 -16140 -760 -16110
rect 760 -17470 790 -17440
rect -1120 -17590 -1090 -17560
rect -910 -17590 -880 -17560
rect -180 -17590 -150 -17560
rect 30 -17590 60 -17560
rect 1090 -16020 1120 -15990
rect 1820 -16260 1850 -16230
rect 1910 -16260 1940 -16230
rect 2030 -16380 2060 -16350
rect 880 -17470 910 -17440
rect 970 -16620 1000 -16590
rect 1910 -16620 1940 -16590
rect 1700 -17110 1730 -17080
rect 2970 -16020 3000 -15990
rect 3700 -16260 3730 -16230
rect 3790 -16260 3820 -16230
rect 3910 -16500 3940 -16470
rect 2760 -16620 2790 -16590
rect 2850 -16990 2880 -16960
rect 2640 -17110 2670 -17080
rect 2760 -17110 2790 -17080
rect 3790 -16990 3820 -16960
rect 3580 -17110 3610 -17080
rect 4850 -16020 4880 -15990
rect 4640 -16990 4670 -16960
rect 4730 -16990 4760 -16960
rect 4520 -17110 4550 -17080
rect 4640 -17350 4670 -17320
rect 5460 -17110 5490 -17080
rect 5670 -16260 5700 -16230
rect 5790 -16500 5820 -16470
rect 5580 -17110 5610 -17080
rect 5670 -16990 5700 -16960
rect 6730 -16020 6760 -15990
rect 6520 -16990 6550 -16960
rect 6610 -16620 6640 -16590
rect 6400 -17110 6430 -17080
rect 6520 -17350 6550 -17320
rect 7340 -17110 7370 -17080
rect 7550 -16260 7580 -16230
rect 7670 -16380 7700 -16350
rect 7460 -17230 7490 -17200
rect 7550 -16620 7580 -16590
rect 8400 -16620 8430 -16590
rect 8280 -17110 8310 -17080
rect 8400 -17110 8430 -17080
rect 8610 -16140 8640 -16110
rect 8490 -17230 8520 -17200
rect 9340 -17350 9370 -17320
rect 9220 -17470 9250 -17440
rect 9430 -16860 9460 -16720
rect 10280 -16860 10310 -16720
rect 10370 -16860 10400 -16720
rect 9550 -17230 9580 -17200
rect 11100 -17230 11130 -17200
rect 11220 -16860 11250 -16720
rect 10160 -17350 10190 -17320
rect 10490 -17350 10520 -17320
rect 12040 -16140 12070 -16110
rect 11310 -17350 11340 -17320
rect 13100 -16260 13130 -16230
rect 12980 -16380 13010 -16350
rect 12250 -16620 12280 -16590
rect 13100 -16620 13130 -16590
rect 12160 -17230 12190 -17200
rect 11430 -17470 11460 -17440
rect 12250 -17110 12280 -17080
rect 12370 -17110 12400 -17080
rect 13920 -16020 13950 -15990
rect 14040 -16620 14070 -16590
rect 13190 -17230 13220 -17200
rect 13310 -17110 13340 -17080
rect 14980 -16260 15010 -16230
rect 14860 -16500 14890 -16470
rect 14130 -16990 14160 -16960
rect 14980 -16990 15010 -16960
rect 14250 -17110 14280 -17080
rect 14130 -17350 14160 -17320
rect 15800 -16020 15830 -15990
rect 15920 -16990 15950 -16960
rect 15070 -17110 15100 -17080
rect 15190 -17110 15220 -17080
rect 16860 -16260 16890 -16230
rect 17680 -16020 17710 -15990
rect 16950 -16260 16980 -16230
rect 16740 -16500 16770 -16470
rect 18740 -16260 18770 -16230
rect 19560 -16020 19590 -15990
rect 18830 -16260 18860 -16230
rect 18620 -16380 18650 -16350
rect 17890 -16620 17920 -16590
rect 18740 -16620 18770 -16590
rect 16010 -16990 16040 -16960
rect 16860 -16990 16890 -16960
rect 16130 -17110 16160 -17080
rect 16010 -17350 16040 -17320
rect 17800 -16990 17830 -16960
rect 17070 -17110 17100 -17080
rect 17890 -17110 17920 -17080
rect 18010 -17110 18040 -17080
rect 19680 -16620 19710 -16590
rect 18950 -17110 18980 -17080
rect 20500 -16020 20530 -15990
rect 20710 -16020 20740 -15990
rect 21440 -16140 21470 -16110
rect 21650 -16020 21680 -15990
rect 22380 -16020 22410 -15990
rect 21560 -16140 21590 -16110
rect 19770 -17470 19800 -17440
rect 19890 -17470 19920 -17440
rect 20620 -17590 20650 -17560
rect 20830 -17590 20860 -17560
rect 21560 -17590 21590 -17560
rect 21770 -17590 21800 -17560
rect 23320 -16020 23350 -15990
rect 24270 -16860 24410 -16720
rect 22710 -17590 22740 -17560
rect -1940 -19050 -1910 -18910
rect -1940 -19210 -1910 -19070
rect -6310 -20500 -6280 -20470
rect -6110 -20500 -6080 -20470
rect -5910 -20500 -5880 -20470
rect -5710 -20500 -5680 -20470
rect -5510 -20500 -5480 -20470
rect -5310 -20500 -5280 -20470
rect -5110 -20500 -5080 -20470
rect -4710 -20500 -4680 -20470
rect -4510 -20500 -4480 -20470
rect -4310 -20500 -4280 -20470
rect -4110 -20500 -4080 -20470
rect -3910 -20500 -3880 -20470
rect -3710 -20500 -3680 -20470
rect -3510 -20500 -3480 -20470
rect -6310 -20620 -6280 -20590
rect -6310 -20740 -6280 -20710
rect -6310 -20860 -6280 -20830
rect -6310 -20980 -6280 -20950
rect -6310 -21100 -6280 -21070
rect -6310 -21220 -6280 -21190
rect -6310 -21470 -6280 -21440
rect -6310 -21590 -6280 -21560
rect -6310 -21710 -6280 -21680
rect -6310 -21830 -6280 -21800
rect -6310 -21950 -6280 -21920
rect -6310 -22070 -6280 -22040
rect -1850 -19050 -1820 -18910
rect -1850 -19210 -1820 -19070
rect -910 -19050 -880 -18910
rect -910 -19210 -880 -19070
rect 970 -19050 1000 -18910
rect 970 -19210 1000 -19070
rect 2850 -19050 2880 -18910
rect 2850 -19210 2880 -19070
rect 4730 -19050 4760 -18910
rect 4730 -19210 4760 -19070
rect 6610 -19050 6640 -18910
rect 6610 -19210 6640 -19070
rect 9430 -19050 9460 -18910
rect 9430 -19210 9460 -19070
rect 11220 -19050 11250 -18910
rect 11220 -19210 11250 -19070
rect 14040 -19050 14070 -18910
rect 14040 -19210 14070 -19070
rect 15920 -19050 15950 -18910
rect 15920 -19210 15950 -19070
rect 17800 -19050 17830 -18910
rect 17800 -19210 17830 -19070
rect 19680 -19050 19710 -18910
rect 19680 -19210 19710 -19070
rect 21560 -19050 21590 -18910
rect 21560 -19210 21590 -19070
rect 22500 -19050 22530 -18910
rect 22500 -19210 22530 -19070
rect 22590 -19050 22620 -18910
rect 22590 -19210 22620 -19070
rect -2060 -20560 -2030 -20530
rect -2670 -22130 -2640 -22100
rect -6310 -22190 -6280 -22160
rect -6110 -22190 -6080 -22160
rect -5910 -22190 -5880 -22160
rect -5710 -22190 -5680 -22160
rect -5510 -22190 -5480 -22160
rect -5310 -22190 -5280 -22160
rect -5110 -22190 -5080 -22160
rect -4710 -22190 -4680 -22160
rect -4510 -22190 -4480 -22160
rect -4310 -22190 -4280 -22160
rect -4110 -22190 -4080 -22160
rect -3910 -22190 -3880 -22160
rect -3710 -22190 -3680 -22160
rect -3510 -22190 -3480 -22160
rect -1120 -20560 -1090 -20530
rect -910 -20560 -880 -20530
rect -180 -20560 -150 -20530
rect 30 -20560 60 -20530
rect 760 -20680 790 -20650
rect 880 -20680 910 -20650
rect -910 -22010 -880 -21980
rect -1730 -22130 -1700 -22100
rect -1000 -22130 -970 -22100
rect -790 -22010 -760 -21980
rect -60 -22130 -30 -22100
rect 150 -22130 180 -22100
rect 1700 -21040 1730 -21010
rect 970 -21530 1000 -21500
rect 2640 -21040 2670 -21010
rect 2760 -21040 2790 -21010
rect 3580 -21040 3610 -21010
rect 2850 -21160 2880 -21130
rect 4640 -20800 4670 -20770
rect 4520 -21040 4550 -21010
rect 3790 -21160 3820 -21130
rect 4640 -21160 4670 -21130
rect 1910 -21530 1940 -21500
rect 2760 -21530 2790 -21500
rect 2030 -21770 2060 -21740
rect 1820 -21890 1850 -21860
rect 1090 -22130 1120 -22100
rect 1910 -21890 1940 -21860
rect 3910 -21650 3940 -21620
rect 3700 -21890 3730 -21860
rect 2970 -22130 3000 -22100
rect 3790 -21890 3820 -21860
rect 5460 -21040 5490 -21010
rect 5580 -21040 5610 -21010
rect 4730 -21160 4760 -21130
rect 4850 -22130 4880 -22100
rect 6520 -20800 6550 -20770
rect 6400 -21040 6430 -21010
rect 5670 -21160 5700 -21130
rect 6520 -21160 6550 -21130
rect 5790 -21650 5820 -21620
rect 5670 -21890 5700 -21860
rect 7340 -21040 7370 -21010
rect 7460 -20920 7490 -20890
rect 6610 -21530 6640 -21500
rect 6730 -22130 6760 -22100
rect 8280 -21040 8310 -21010
rect 8400 -21040 8430 -21010
rect 9220 -20680 9250 -20650
rect 8490 -20920 8520 -20890
rect 7550 -21530 7580 -21500
rect 8400 -21530 8430 -21500
rect 7670 -21770 7700 -21740
rect 7550 -21890 7580 -21860
rect 9340 -20800 9370 -20770
rect 8610 -22010 8640 -21980
rect 10160 -20800 10190 -20770
rect 10490 -20800 10520 -20770
rect 9430 -21400 9460 -21260
rect 9550 -20920 9580 -20890
rect 11100 -20920 11130 -20890
rect 10280 -21400 10310 -21260
rect 10370 -21400 10400 -21260
rect 11220 -21400 11250 -21260
rect 11430 -20680 11460 -20650
rect 11310 -20800 11340 -20770
rect 12160 -20920 12190 -20890
rect 12040 -22010 12070 -21980
rect 12250 -21040 12280 -21010
rect 12370 -21040 12400 -21010
rect 12250 -21530 12280 -21500
rect 13100 -21530 13130 -21500
rect 13190 -20920 13220 -20890
rect 12980 -21770 13010 -21740
rect 13100 -21890 13130 -21860
rect 13310 -21040 13340 -21010
rect 14130 -20800 14160 -20770
rect 14250 -21040 14280 -21010
rect 14040 -21530 14070 -21500
rect 14130 -21160 14160 -21130
rect 13920 -22130 13950 -22100
rect 14980 -21160 15010 -21130
rect 15070 -21040 15100 -21010
rect 14860 -21650 14890 -21620
rect 14980 -21890 15010 -21860
rect 15190 -21040 15220 -21010
rect 16010 -20800 16040 -20770
rect 16130 -21040 16160 -21010
rect 15920 -21160 15950 -21130
rect 16010 -21160 16040 -21130
rect 15800 -22130 15830 -22100
rect 17070 -21040 17100 -21010
rect 16860 -21160 16890 -21130
rect 17890 -21040 17920 -21010
rect 18010 -21040 18040 -21010
rect 17800 -21160 17830 -21130
rect 17890 -21530 17920 -21500
rect 16740 -21650 16770 -21620
rect 16860 -21890 16890 -21860
rect 16950 -21890 16980 -21860
rect 17680 -22130 17710 -22100
rect 18950 -21040 18980 -21010
rect 18740 -21530 18770 -21500
rect 19680 -21530 19710 -21500
rect 19770 -20680 19800 -20650
rect 18620 -21770 18650 -21740
rect 18740 -21890 18770 -21860
rect 18830 -21890 18860 -21860
rect 19560 -22130 19590 -22100
rect 20620 -20560 20650 -20530
rect 20830 -20560 20860 -20530
rect 21560 -20560 21590 -20530
rect 21770 -20560 21800 -20530
rect 19890 -20680 19920 -20650
rect 21440 -22010 21470 -21980
rect 20500 -22130 20530 -22100
rect 20710 -22130 20740 -22100
rect 21560 -22010 21590 -21980
rect 21650 -22130 21680 -22100
rect 22380 -22130 22410 -22100
rect 23440 -19050 23470 -18910
rect 23440 -19210 23470 -19070
rect 22710 -20560 22740 -20530
rect 24270 -21400 24410 -21260
rect 23320 -22130 23350 -22100
rect -2790 -25330 -2760 -25190
rect -1940 -25330 -1910 -25190
rect -1000 -25330 -970 -25190
rect 880 -25330 910 -25190
rect 1820 -25330 1850 -25190
rect 3700 -25330 3730 -25190
rect 5580 -25330 5610 -25190
rect 7460 -25330 7490 -25190
rect 10280 -25330 10310 -25190
rect 10370 -25330 10400 -25190
rect 13190 -25330 13220 -25190
rect 15070 -25330 15100 -25190
rect 16950 -25330 16980 -25190
rect 18830 -25330 18860 -25190
rect 19770 -25330 19800 -25190
rect 21650 -25330 21680 -25190
rect 22590 -25330 22620 -25190
rect 23440 -25330 23470 -25190
<< metal2 >>
rect -3420 -230 24420 -220
rect -3420 -370 -3410 -230
rect -3270 -370 -2790 -230
rect -2760 -370 -1940 -230
rect -1910 -370 -1000 -230
rect -970 -370 880 -230
rect 910 -370 1820 -230
rect 1850 -370 3700 -230
rect 3730 -370 5580 -230
rect 5610 -370 7460 -230
rect 7490 -370 10280 -230
rect 10310 -370 10370 -230
rect 10400 -370 13190 -230
rect 13220 -370 15070 -230
rect 15100 -370 16950 -230
rect 16980 -370 18830 -230
rect 18860 -370 19770 -230
rect 19800 -370 21650 -230
rect 21680 -370 22590 -230
rect 22620 -370 23440 -230
rect 23470 -370 23950 -230
rect 24090 -370 24420 -230
rect -3420 -380 24420 -370
rect -6320 -3370 -6270 -3360
rect -6120 -3370 -6070 -3360
rect -5920 -3370 -5870 -3360
rect -5720 -3370 -5670 -3360
rect -5520 -3370 -5470 -3360
rect -5320 -3370 -5270 -3360
rect -5120 -3370 -5070 -3360
rect -4720 -3370 -4670 -3360
rect -4520 -3370 -4470 -3360
rect -4320 -3370 -4270 -3360
rect -4120 -3370 -4070 -3360
rect -3920 -3370 -3870 -3360
rect -3720 -3370 -3670 -3360
rect -3520 -3370 -3470 -3360
rect -6320 -3400 -6310 -3370
rect -6280 -3400 -6110 -3370
rect -6080 -3400 -5910 -3370
rect -5880 -3400 -5710 -3370
rect -5680 -3400 -5510 -3370
rect -5480 -3400 -5310 -3370
rect -5280 -3400 -5110 -3370
rect -5080 -3400 -4710 -3370
rect -4680 -3400 -4510 -3370
rect -4480 -3400 -4310 -3370
rect -4280 -3400 -4110 -3370
rect -4080 -3400 -3910 -3370
rect -3880 -3400 -3710 -3370
rect -3680 -3400 -3510 -3370
rect -3480 -3400 23620 -3370
rect -6320 -3410 -6270 -3400
rect -6120 -3410 -6070 -3400
rect -5920 -3410 -5870 -3400
rect -5720 -3410 -5670 -3400
rect -5520 -3410 -5470 -3400
rect -5320 -3410 -5270 -3400
rect -5120 -3410 -5070 -3400
rect -4720 -3410 -4670 -3400
rect -4520 -3410 -4470 -3400
rect -4320 -3410 -4270 -3400
rect -4120 -3410 -4070 -3400
rect -3920 -3410 -3870 -3400
rect -3720 -3410 -3670 -3400
rect -3520 -3410 -3470 -3400
rect -6220 -3430 -6170 -3420
rect -6310 -3460 -6210 -3430
rect -6180 -3460 -2670 -3430
rect -2640 -3460 -1730 -3430
rect -1700 -3460 -1000 -3430
rect -970 -3460 -60 -3430
rect -30 -3460 150 -3430
rect 180 -3460 1090 -3430
rect 1120 -3460 2970 -3430
rect 3000 -3460 4850 -3430
rect 4880 -3460 6730 -3430
rect 6760 -3460 13920 -3430
rect 13950 -3460 15800 -3430
rect 15830 -3460 17680 -3430
rect 17710 -3460 19560 -3430
rect 19590 -3460 20500 -3430
rect 20530 -3460 20710 -3430
rect 20740 -3460 21650 -3430
rect 21680 -3460 22380 -3430
rect 22410 -3460 23320 -3430
rect 23350 -3460 23620 -3430
rect -6220 -3470 -6170 -3460
rect -6320 -3490 -6270 -3480
rect -6320 -3520 -6310 -3490
rect -6280 -3520 23620 -3490
rect -6320 -3530 -6270 -3520
rect -6020 -3550 -5970 -3540
rect -6310 -3580 -6010 -3550
rect -5980 -3580 -910 -3550
rect -880 -3580 -790 -3550
rect -760 -3580 8610 -3550
rect 8640 -3580 12040 -3550
rect 12070 -3580 21440 -3550
rect 21470 -3580 21560 -3550
rect 21590 -3580 23620 -3550
rect -6020 -3590 -5970 -3580
rect -6320 -3610 -6270 -3600
rect -6320 -3640 -6310 -3610
rect -6280 -3640 23620 -3610
rect -6320 -3650 -6270 -3640
rect -5820 -3670 -5770 -3660
rect -6310 -3700 -5810 -3670
rect -5780 -3700 1820 -3670
rect 1850 -3700 1910 -3670
rect 1940 -3700 3700 -3670
rect 3730 -3700 3790 -3670
rect 3820 -3700 5670 -3670
rect 5700 -3700 7550 -3670
rect 7580 -3700 13100 -3670
rect 13130 -3700 14980 -3670
rect 15010 -3700 16860 -3670
rect 16890 -3700 16950 -3670
rect 16980 -3700 18740 -3670
rect 18770 -3700 18830 -3670
rect 18860 -3700 23620 -3670
rect -5820 -3710 -5770 -3700
rect -6320 -3730 -6270 -3720
rect -6320 -3760 -6310 -3730
rect -6280 -3760 23620 -3730
rect -6320 -3770 -6270 -3760
rect -5620 -3790 -5570 -3780
rect -6310 -3820 -5610 -3790
rect -5580 -3820 2030 -3790
rect 2060 -3820 7670 -3790
rect 7700 -3820 12980 -3790
rect 13010 -3820 18620 -3790
rect 18650 -3820 23620 -3790
rect -5620 -3830 -5570 -3820
rect -6320 -3850 -6270 -3840
rect -6320 -3880 -6310 -3850
rect -6280 -3880 23620 -3850
rect -6320 -3890 -6270 -3880
rect -5420 -3910 -5370 -3900
rect -6310 -3940 -5410 -3910
rect -5380 -3940 3910 -3910
rect 3940 -3940 5790 -3910
rect 5820 -3940 14860 -3910
rect 14890 -3940 16740 -3910
rect 16770 -3940 23620 -3910
rect -5420 -3950 -5370 -3940
rect -6320 -3970 -6270 -3960
rect -6320 -4000 -6310 -3970
rect -6280 -4000 23620 -3970
rect -6320 -4010 -6270 -4000
rect -5220 -4030 -5170 -4020
rect -6310 -4060 -5210 -4030
rect -5180 -4060 970 -4030
rect 1000 -4060 1910 -4030
rect 1940 -4060 2760 -4030
rect 2790 -4060 6610 -4030
rect 6640 -4060 7550 -4030
rect 7580 -4060 8400 -4030
rect 8430 -4060 12250 -4030
rect 12280 -4060 13100 -4030
rect 13130 -4060 14040 -4030
rect 14070 -4060 17890 -4030
rect 17920 -4060 18740 -4030
rect 18770 -4060 19680 -4030
rect 19710 -4060 23620 -4030
rect -5220 -4070 -5170 -4060
rect -6320 -4090 -6270 -4080
rect -6320 -4120 -6310 -4090
rect -6280 -4120 23620 -4090
rect -6320 -4130 -6270 -4120
rect -6310 -4160 23620 -4150
rect -6310 -4300 -5000 -4160
rect -4790 -4300 9430 -4160
rect 9460 -4300 10280 -4160
rect 10310 -4300 10370 -4160
rect 10400 -4300 11220 -4160
rect 11250 -4300 23620 -4160
rect -6310 -4310 23620 -4300
rect 24260 -4160 24420 -4150
rect 24260 -4300 24270 -4160
rect 24410 -4300 24420 -4160
rect 24260 -4310 24420 -4300
rect -6320 -4340 -6270 -4330
rect -6320 -4370 -6310 -4340
rect -6280 -4370 23620 -4340
rect -6320 -4380 -6270 -4370
rect -4620 -4400 -4570 -4390
rect -6310 -4430 -4610 -4400
rect -4580 -4430 2850 -4400
rect 2880 -4430 3790 -4400
rect 3820 -4430 4640 -4400
rect 4670 -4430 4730 -4400
rect 4760 -4430 5670 -4400
rect 5700 -4430 6520 -4400
rect 6550 -4430 14130 -4400
rect 14160 -4430 14980 -4400
rect 15010 -4430 15920 -4400
rect 15950 -4430 16010 -4400
rect 16040 -4430 16860 -4400
rect 16890 -4430 17800 -4400
rect 17830 -4430 23620 -4400
rect -4620 -4440 -4570 -4430
rect -6320 -4460 -6270 -4450
rect -6320 -4490 -6310 -4460
rect -6280 -4490 23620 -4460
rect -6320 -4500 -6270 -4490
rect -4420 -4520 -4370 -4510
rect -6310 -4550 -4410 -4520
rect -4380 -4550 1700 -4520
rect 1730 -4550 2640 -4520
rect 2670 -4550 2760 -4520
rect 2790 -4550 3580 -4520
rect 3610 -4550 4520 -4520
rect 4550 -4550 5460 -4520
rect 5490 -4550 5580 -4520
rect 5610 -4550 6400 -4520
rect 6430 -4550 7340 -4520
rect 7370 -4550 8280 -4520
rect 8310 -4550 8400 -4520
rect 8430 -4550 12250 -4520
rect 12280 -4550 12370 -4520
rect 12400 -4550 13310 -4520
rect 13340 -4550 14250 -4520
rect 14280 -4550 15070 -4520
rect 15100 -4550 15190 -4520
rect 15220 -4550 16130 -4520
rect 16160 -4550 17070 -4520
rect 17100 -4550 17890 -4520
rect 17920 -4550 18010 -4520
rect 18040 -4550 18950 -4520
rect 18980 -4550 23620 -4520
rect -4420 -4560 -4370 -4550
rect -6320 -4580 -6270 -4570
rect -6320 -4610 -6310 -4580
rect -6280 -4610 23620 -4580
rect -6320 -4620 -6270 -4610
rect -4220 -4640 -4170 -4630
rect -6310 -4670 -4210 -4640
rect -4180 -4670 7460 -4640
rect 7490 -4670 8490 -4640
rect 8520 -4670 9550 -4640
rect 9580 -4670 11100 -4640
rect 11130 -4670 12160 -4640
rect 12190 -4670 13190 -4640
rect 13220 -4670 23620 -4640
rect -4220 -4680 -4170 -4670
rect -6320 -4700 -6270 -4690
rect -6320 -4730 -6310 -4700
rect -6280 -4730 23620 -4700
rect -6320 -4740 -6270 -4730
rect -4020 -4760 -3970 -4750
rect -6310 -4790 -4010 -4760
rect -3980 -4790 4640 -4760
rect 4670 -4790 6520 -4760
rect 6550 -4790 9340 -4760
rect 9370 -4790 10160 -4760
rect 10190 -4790 10490 -4760
rect 10520 -4790 11310 -4760
rect 11340 -4790 14130 -4760
rect 14160 -4790 16010 -4760
rect 16040 -4790 23620 -4760
rect -4020 -4800 -3970 -4790
rect -6320 -4820 -6270 -4810
rect -6320 -4850 -6310 -4820
rect -6280 -4850 23620 -4820
rect -6320 -4860 -6270 -4850
rect -3820 -4880 -3770 -4870
rect -6310 -4910 -3810 -4880
rect -3780 -4910 760 -4880
rect 790 -4910 880 -4880
rect 910 -4910 9220 -4880
rect 9250 -4910 11430 -4880
rect 11460 -4910 19770 -4880
rect 19800 -4910 19890 -4880
rect 19920 -4910 23620 -4880
rect -3820 -4920 -3770 -4910
rect -6320 -4940 -6270 -4930
rect -6320 -4970 -6310 -4940
rect -6280 -4970 23620 -4940
rect -6320 -4980 -6270 -4970
rect -3620 -5000 -3570 -4990
rect -6310 -5030 -3610 -5000
rect -3580 -5030 -2060 -5000
rect -2030 -5030 -1120 -5000
rect -1090 -5030 -910 -5000
rect -880 -5030 -180 -5000
rect -150 -5030 30 -5000
rect 60 -5030 20620 -5000
rect 20650 -5030 20830 -5000
rect 20860 -5030 21560 -5000
rect 21590 -5030 21770 -5000
rect 21800 -5030 22710 -5000
rect 22740 -5030 23620 -5000
rect -3620 -5040 -3570 -5030
rect -6320 -5060 -6270 -5050
rect -6120 -5060 -6070 -5050
rect -5920 -5060 -5870 -5050
rect -5720 -5060 -5670 -5050
rect -5520 -5060 -5470 -5050
rect -5320 -5060 -5270 -5050
rect -5120 -5060 -5070 -5050
rect -4720 -5060 -4670 -5050
rect -4520 -5060 -4470 -5050
rect -4320 -5060 -4270 -5050
rect -4120 -5060 -4070 -5050
rect -3920 -5060 -3870 -5050
rect -3720 -5060 -3670 -5050
rect -3520 -5060 -3470 -5050
rect -6320 -5090 -6310 -5060
rect -6280 -5090 -6110 -5060
rect -6080 -5090 -5910 -5060
rect -5880 -5090 -5710 -5060
rect -5680 -5090 -5510 -5060
rect -5480 -5090 -5310 -5060
rect -5280 -5090 -5110 -5060
rect -5080 -5090 -4710 -5060
rect -4680 -5090 -4510 -5060
rect -4480 -5090 -4310 -5060
rect -4280 -5090 -4110 -5060
rect -4080 -5090 -3910 -5060
rect -3880 -5090 -3710 -5060
rect -3680 -5090 -3510 -5060
rect -3480 -5090 23620 -5060
rect -6320 -5100 -6270 -5090
rect -6120 -5100 -6070 -5090
rect -5920 -5100 -5870 -5090
rect -5720 -5100 -5670 -5090
rect -5520 -5100 -5470 -5090
rect -5320 -5100 -5270 -5090
rect -5120 -5100 -5070 -5090
rect -4720 -5100 -4670 -5090
rect -4520 -5100 -4470 -5090
rect -4320 -5100 -4270 -5090
rect -4120 -5100 -4070 -5090
rect -3920 -5100 -3870 -5090
rect -3720 -5100 -3670 -5090
rect -3520 -5100 -3470 -5090
rect -3100 -6350 24420 -6340
rect -3100 -6490 -3090 -6350
rect -2950 -6490 -2790 -6350
rect -2760 -6490 -1940 -6350
rect -1910 -6490 -1850 -6350
rect -1820 -6490 -910 -6350
rect -880 -6490 970 -6350
rect 1000 -6490 2850 -6350
rect 2880 -6490 4730 -6350
rect 4760 -6490 6610 -6350
rect 6640 -6490 9430 -6350
rect 9460 -6490 11220 -6350
rect 11250 -6490 14040 -6350
rect 14070 -6490 15920 -6350
rect 15950 -6490 17800 -6350
rect 17830 -6490 19680 -6350
rect 19710 -6490 21560 -6350
rect 21590 -6490 22500 -6350
rect 22530 -6490 22590 -6350
rect 22620 -6490 23440 -6350
rect 23470 -6490 23630 -6350
rect 23770 -6490 24420 -6350
rect -3100 -6510 24420 -6490
rect -3100 -6650 -3090 -6510
rect -2950 -6650 -2790 -6510
rect -2760 -6650 -1940 -6510
rect -1910 -6650 -1850 -6510
rect -1820 -6650 -910 -6510
rect -880 -6650 970 -6510
rect 1000 -6650 2850 -6510
rect 2880 -6650 4730 -6510
rect 4760 -6650 6610 -6510
rect 6640 -6650 9430 -6510
rect 9460 -6650 11220 -6510
rect 11250 -6650 14040 -6510
rect 14070 -6650 15920 -6510
rect 15950 -6650 17800 -6510
rect 17830 -6650 19680 -6510
rect 19710 -6650 21560 -6510
rect 21590 -6650 22500 -6510
rect 22530 -6650 22590 -6510
rect 22620 -6650 23440 -6510
rect 23470 -6650 23630 -6510
rect 23770 -6650 24420 -6510
rect -3100 -6660 24420 -6650
rect -6320 -7910 -6270 -7900
rect -6120 -7910 -6070 -7900
rect -5920 -7910 -5870 -7900
rect -5720 -7910 -5670 -7900
rect -5520 -7910 -5470 -7900
rect -5320 -7910 -5270 -7900
rect -5120 -7910 -5070 -7900
rect -4720 -7910 -4670 -7900
rect -4520 -7910 -4470 -7900
rect -4320 -7910 -4270 -7900
rect -4120 -7910 -4070 -7900
rect -3920 -7910 -3870 -7900
rect -3720 -7910 -3670 -7900
rect -3520 -7910 -3470 -7900
rect -6320 -7940 -6310 -7910
rect -6280 -7940 -6110 -7910
rect -6080 -7940 -5910 -7910
rect -5880 -7940 -5710 -7910
rect -5680 -7940 -5510 -7910
rect -5480 -7940 -5310 -7910
rect -5280 -7940 -5110 -7910
rect -5080 -7940 -4710 -7910
rect -4680 -7940 -4510 -7910
rect -4480 -7940 -4310 -7910
rect -4280 -7940 -4110 -7910
rect -4080 -7940 -3910 -7910
rect -3880 -7940 -3710 -7910
rect -3680 -7940 -3510 -7910
rect -3480 -7940 23620 -7910
rect -6320 -7950 -6270 -7940
rect -6120 -7950 -6070 -7940
rect -5920 -7950 -5870 -7940
rect -5720 -7950 -5670 -7940
rect -5520 -7950 -5470 -7940
rect -5320 -7950 -5270 -7940
rect -5120 -7950 -5070 -7940
rect -4720 -7950 -4670 -7940
rect -4520 -7950 -4470 -7940
rect -4320 -7950 -4270 -7940
rect -4120 -7950 -4070 -7940
rect -3920 -7950 -3870 -7940
rect -3720 -7950 -3670 -7940
rect -3520 -7950 -3470 -7940
rect -3620 -7970 -3570 -7960
rect -6310 -8000 -3610 -7970
rect -3580 -8000 -2060 -7970
rect -2030 -8000 -1120 -7970
rect -1090 -8000 -910 -7970
rect -880 -8000 -180 -7970
rect -150 -8000 30 -7970
rect 60 -8000 20620 -7970
rect 20650 -8000 20830 -7970
rect 20860 -8000 21560 -7970
rect 21590 -8000 21770 -7970
rect 21800 -8000 22710 -7970
rect 22740 -8000 23620 -7970
rect -3620 -8010 -3570 -8000
rect -6320 -8030 -6270 -8020
rect -6320 -8060 -6310 -8030
rect -6280 -8060 23620 -8030
rect -6320 -8070 -6270 -8060
rect -3820 -8090 -3770 -8080
rect -6310 -8120 -3810 -8090
rect -3780 -8120 760 -8090
rect 790 -8120 880 -8090
rect 910 -8120 9220 -8090
rect 9250 -8120 11430 -8090
rect 11460 -8120 19770 -8090
rect 19800 -8120 19890 -8090
rect 19920 -8120 23620 -8090
rect -3820 -8130 -3770 -8120
rect -6320 -8150 -6270 -8140
rect -6320 -8180 -6310 -8150
rect -6280 -8180 23620 -8150
rect -6320 -8190 -6270 -8180
rect -4020 -8210 -3970 -8200
rect -6310 -8240 -4010 -8210
rect -3980 -8240 4640 -8210
rect 4670 -8240 6520 -8210
rect 6550 -8240 9340 -8210
rect 9370 -8240 10160 -8210
rect 10190 -8240 10490 -8210
rect 10520 -8240 11310 -8210
rect 11340 -8240 14130 -8210
rect 14160 -8240 16010 -8210
rect 16040 -8240 23620 -8210
rect -4020 -8250 -3970 -8240
rect -6320 -8270 -6270 -8260
rect -6320 -8300 -6310 -8270
rect -6280 -8300 23620 -8270
rect -6320 -8310 -6270 -8300
rect -4220 -8330 -4170 -8320
rect -6310 -8360 -4210 -8330
rect -4180 -8360 7460 -8330
rect 7490 -8360 8490 -8330
rect 8520 -8360 9550 -8330
rect 9580 -8360 11100 -8330
rect 11130 -8360 12160 -8330
rect 12190 -8360 13190 -8330
rect 13220 -8360 23620 -8330
rect -4220 -8370 -4170 -8360
rect -6320 -8390 -6270 -8380
rect -6320 -8420 -6310 -8390
rect -6280 -8420 23620 -8390
rect -6320 -8430 -6270 -8420
rect -4420 -8450 -4370 -8440
rect -6310 -8480 -4410 -8450
rect -4380 -8480 1700 -8450
rect 1730 -8480 2640 -8450
rect 2670 -8480 2760 -8450
rect 2790 -8480 3580 -8450
rect 3610 -8480 4520 -8450
rect 4550 -8480 5460 -8450
rect 5490 -8480 5580 -8450
rect 5610 -8480 6400 -8450
rect 6430 -8480 7340 -8450
rect 7370 -8480 8280 -8450
rect 8310 -8480 8400 -8450
rect 8430 -8480 12250 -8450
rect 12280 -8480 12370 -8450
rect 12400 -8480 13310 -8450
rect 13340 -8480 14250 -8450
rect 14280 -8480 15070 -8450
rect 15100 -8480 15190 -8450
rect 15220 -8480 16130 -8450
rect 16160 -8480 17070 -8450
rect 17100 -8480 17890 -8450
rect 17920 -8480 18010 -8450
rect 18040 -8480 18950 -8450
rect 18980 -8480 23620 -8450
rect -4420 -8490 -4370 -8480
rect -6320 -8510 -6270 -8500
rect -6320 -8540 -6310 -8510
rect -6280 -8540 23620 -8510
rect -6320 -8550 -6270 -8540
rect -4620 -8570 -4570 -8560
rect -6310 -8600 -4610 -8570
rect -4580 -8600 2850 -8570
rect 2880 -8600 3790 -8570
rect 3820 -8600 4640 -8570
rect 4670 -8600 4730 -8570
rect 4760 -8600 5670 -8570
rect 5700 -8600 6520 -8570
rect 6550 -8600 14130 -8570
rect 14160 -8600 14980 -8570
rect 15010 -8600 15920 -8570
rect 15950 -8600 16010 -8570
rect 16040 -8600 16860 -8570
rect 16890 -8600 17800 -8570
rect 17830 -8600 23620 -8570
rect -4620 -8610 -4570 -8600
rect -6320 -8630 -6270 -8620
rect -6320 -8660 -6310 -8630
rect -6280 -8660 23620 -8630
rect -6320 -8670 -6270 -8660
rect -6310 -8700 23620 -8690
rect -6310 -8840 -5000 -8700
rect -4790 -8840 9430 -8700
rect 9460 -8840 10280 -8700
rect 10310 -8840 10370 -8700
rect 10400 -8840 11220 -8700
rect 11250 -8840 23620 -8700
rect -6310 -8850 23620 -8840
rect 24260 -8700 24420 -8690
rect 24260 -8840 24270 -8700
rect 24410 -8840 24420 -8700
rect 24260 -8850 24420 -8840
rect -6320 -8880 -6270 -8870
rect -6320 -8910 -6310 -8880
rect -6280 -8910 23620 -8880
rect -6320 -8920 -6270 -8910
rect -5220 -8940 -5170 -8930
rect -6310 -8970 -5210 -8940
rect -5180 -8970 970 -8940
rect 1000 -8970 1910 -8940
rect 1940 -8970 2760 -8940
rect 2790 -8970 6610 -8940
rect 6640 -8970 7550 -8940
rect 7580 -8970 8400 -8940
rect 8430 -8970 12250 -8940
rect 12280 -8970 13100 -8940
rect 13130 -8970 14040 -8940
rect 14070 -8970 17890 -8940
rect 17920 -8970 18740 -8940
rect 18770 -8970 19680 -8940
rect 19710 -8970 23620 -8940
rect -5220 -8980 -5170 -8970
rect -6320 -9000 -6270 -8990
rect -6320 -9030 -6310 -9000
rect -6280 -9030 23620 -9000
rect -6320 -9040 -6270 -9030
rect -5420 -9060 -5370 -9050
rect -6310 -9090 -5410 -9060
rect -5380 -9090 3910 -9060
rect 3940 -9090 5790 -9060
rect 5820 -9090 14860 -9060
rect 14890 -9090 16740 -9060
rect 16770 -9090 23620 -9060
rect -5420 -9100 -5370 -9090
rect -6320 -9120 -6270 -9110
rect -6320 -9150 -6310 -9120
rect -6280 -9150 23620 -9120
rect -6320 -9160 -6270 -9150
rect -5620 -9180 -5570 -9170
rect -6310 -9210 -5610 -9180
rect -5580 -9210 2030 -9180
rect 2060 -9210 7670 -9180
rect 7700 -9210 12980 -9180
rect 13010 -9210 18620 -9180
rect 18650 -9210 23620 -9180
rect -5620 -9220 -5570 -9210
rect -6320 -9240 -6270 -9230
rect -6320 -9270 -6310 -9240
rect -6280 -9270 23620 -9240
rect -6320 -9280 -6270 -9270
rect -5820 -9300 -5770 -9290
rect -6310 -9330 -5810 -9300
rect -5780 -9330 1820 -9300
rect 1850 -9330 1910 -9300
rect 1940 -9330 3700 -9300
rect 3730 -9330 3790 -9300
rect 3820 -9330 5670 -9300
rect 5700 -9330 7550 -9300
rect 7580 -9330 13100 -9300
rect 13130 -9330 14980 -9300
rect 15010 -9330 16860 -9300
rect 16890 -9330 16950 -9300
rect 16980 -9330 18740 -9300
rect 18770 -9330 18830 -9300
rect 18860 -9330 23620 -9300
rect -5820 -9340 -5770 -9330
rect -6320 -9360 -6270 -9350
rect -6320 -9390 -6310 -9360
rect -6280 -9390 23620 -9360
rect -6320 -9400 -6270 -9390
rect -6020 -9420 -5970 -9410
rect -6310 -9450 -6010 -9420
rect -5980 -9450 -910 -9420
rect -880 -9450 -790 -9420
rect -760 -9450 8610 -9420
rect 8640 -9450 12040 -9420
rect 12070 -9450 21440 -9420
rect 21470 -9450 21560 -9420
rect 21590 -9450 23620 -9420
rect -6020 -9460 -5970 -9450
rect -6320 -9480 -6270 -9470
rect -6320 -9510 -6310 -9480
rect -6280 -9510 23620 -9480
rect -6320 -9520 -6270 -9510
rect -6220 -9540 -6170 -9530
rect -6310 -9570 -6210 -9540
rect -6180 -9570 -2670 -9540
rect -2640 -9570 -1730 -9540
rect -1700 -9570 -1000 -9540
rect -970 -9570 -60 -9540
rect -30 -9570 150 -9540
rect 180 -9570 1090 -9540
rect 1120 -9570 2970 -9540
rect 3000 -9570 4850 -9540
rect 4880 -9570 6730 -9540
rect 6760 -9570 13920 -9540
rect 13950 -9570 15800 -9540
rect 15830 -9570 17680 -9540
rect 17710 -9570 19560 -9540
rect 19590 -9570 20500 -9540
rect 20530 -9570 20710 -9540
rect 20740 -9570 21650 -9540
rect 21680 -9570 22380 -9540
rect 22410 -9570 23320 -9540
rect 23350 -9570 23620 -9540
rect -6220 -9580 -6170 -9570
rect -6320 -9600 -6270 -9590
rect -6120 -9600 -6070 -9590
rect -5920 -9600 -5870 -9590
rect -5720 -9600 -5670 -9590
rect -5520 -9600 -5470 -9590
rect -5320 -9600 -5270 -9590
rect -5120 -9600 -5070 -9590
rect -4720 -9600 -4670 -9590
rect -4520 -9600 -4470 -9590
rect -4320 -9600 -4270 -9590
rect -4120 -9600 -4070 -9590
rect -3920 -9600 -3870 -9590
rect -3720 -9600 -3670 -9590
rect -3520 -9600 -3470 -9590
rect -6320 -9630 -6310 -9600
rect -6280 -9630 -6110 -9600
rect -6080 -9630 -5910 -9600
rect -5880 -9630 -5710 -9600
rect -5680 -9630 -5510 -9600
rect -5480 -9630 -5310 -9600
rect -5280 -9630 -5110 -9600
rect -5080 -9630 -4710 -9600
rect -4680 -9630 -4510 -9600
rect -4480 -9630 -4310 -9600
rect -4280 -9630 -4110 -9600
rect -4080 -9630 -3910 -9600
rect -3880 -9630 -3710 -9600
rect -3680 -9630 -3510 -9600
rect -3480 -9630 23620 -9600
rect -6320 -9640 -6270 -9630
rect -6120 -9640 -6070 -9630
rect -5920 -9640 -5870 -9630
rect -5720 -9640 -5670 -9630
rect -5520 -9640 -5470 -9630
rect -5320 -9640 -5270 -9630
rect -5120 -9640 -5070 -9630
rect -4720 -9640 -4670 -9630
rect -4520 -9640 -4470 -9630
rect -4320 -9640 -4270 -9630
rect -4120 -9640 -4070 -9630
rect -3920 -9640 -3870 -9630
rect -3720 -9640 -3670 -9630
rect -3520 -9640 -3470 -9630
rect -3420 -12630 24420 -12620
rect -3420 -12770 -3410 -12630
rect -3270 -12770 -2790 -12630
rect -2760 -12770 -1940 -12630
rect -1910 -12770 -1000 -12630
rect -970 -12770 880 -12630
rect 910 -12770 1820 -12630
rect 1850 -12770 3700 -12630
rect 3730 -12770 5580 -12630
rect 5610 -12770 7460 -12630
rect 7490 -12770 10280 -12630
rect 10310 -12770 10370 -12630
rect 10400 -12770 13190 -12630
rect 13220 -12770 15070 -12630
rect 15100 -12770 16950 -12630
rect 16980 -12770 18830 -12630
rect 18860 -12770 19770 -12630
rect 19800 -12770 21650 -12630
rect 21680 -12770 22590 -12630
rect 22620 -12770 23440 -12630
rect 23470 -12770 23950 -12630
rect 24090 -12770 24420 -12630
rect -3420 -12790 24420 -12770
rect -3420 -12930 -3410 -12790
rect -3270 -12930 -2790 -12790
rect -2760 -12930 -1940 -12790
rect -1910 -12930 -1000 -12790
rect -970 -12930 880 -12790
rect 910 -12930 1820 -12790
rect 1850 -12930 3700 -12790
rect 3730 -12930 5580 -12790
rect 5610 -12930 7460 -12790
rect 7490 -12930 10280 -12790
rect 10310 -12930 10370 -12790
rect 10400 -12930 13190 -12790
rect 13220 -12930 15070 -12790
rect 15100 -12930 16950 -12790
rect 16980 -12930 18830 -12790
rect 18860 -12930 19770 -12790
rect 19800 -12930 21650 -12790
rect 21680 -12930 22590 -12790
rect 22620 -12930 23440 -12790
rect 23470 -12930 23950 -12790
rect 24090 -12930 24420 -12790
rect -3420 -12940 24420 -12930
rect -6320 -15930 -6270 -15920
rect -6120 -15930 -6070 -15920
rect -5920 -15930 -5870 -15920
rect -5720 -15930 -5670 -15920
rect -5520 -15930 -5470 -15920
rect -5320 -15930 -5270 -15920
rect -5120 -15930 -5070 -15920
rect -4720 -15930 -4670 -15920
rect -4520 -15930 -4470 -15920
rect -4320 -15930 -4270 -15920
rect -4120 -15930 -4070 -15920
rect -3920 -15930 -3870 -15920
rect -3720 -15930 -3670 -15920
rect -3520 -15930 -3470 -15920
rect -6320 -15960 -6310 -15930
rect -6280 -15960 -6110 -15930
rect -6080 -15960 -5910 -15930
rect -5880 -15960 -5710 -15930
rect -5680 -15960 -5510 -15930
rect -5480 -15960 -5310 -15930
rect -5280 -15960 -5110 -15930
rect -5080 -15960 -4710 -15930
rect -4680 -15960 -4510 -15930
rect -4480 -15960 -4310 -15930
rect -4280 -15960 -4110 -15930
rect -4080 -15960 -3910 -15930
rect -3880 -15960 -3710 -15930
rect -3680 -15960 -3510 -15930
rect -3480 -15960 23620 -15930
rect -6320 -15970 -6270 -15960
rect -6120 -15970 -6070 -15960
rect -5920 -15970 -5870 -15960
rect -5720 -15970 -5670 -15960
rect -5520 -15970 -5470 -15960
rect -5320 -15970 -5270 -15960
rect -5120 -15970 -5070 -15960
rect -4720 -15970 -4670 -15960
rect -4520 -15970 -4470 -15960
rect -4320 -15970 -4270 -15960
rect -4120 -15970 -4070 -15960
rect -3920 -15970 -3870 -15960
rect -3720 -15970 -3670 -15960
rect -3520 -15970 -3470 -15960
rect -6220 -15990 -6170 -15980
rect -6310 -16020 -6210 -15990
rect -6180 -16020 -2670 -15990
rect -2640 -16020 -1730 -15990
rect -1700 -16020 -1000 -15990
rect -970 -16020 -60 -15990
rect -30 -16020 150 -15990
rect 180 -16020 1090 -15990
rect 1120 -16020 2970 -15990
rect 3000 -16020 4850 -15990
rect 4880 -16020 6730 -15990
rect 6760 -16020 13920 -15990
rect 13950 -16020 15800 -15990
rect 15830 -16020 17680 -15990
rect 17710 -16020 19560 -15990
rect 19590 -16020 20500 -15990
rect 20530 -16020 20710 -15990
rect 20740 -16020 21650 -15990
rect 21680 -16020 22380 -15990
rect 22410 -16020 23320 -15990
rect 23350 -16020 23620 -15990
rect -6220 -16030 -6170 -16020
rect -6320 -16050 -6270 -16040
rect -6320 -16080 -6310 -16050
rect -6280 -16080 23620 -16050
rect -6320 -16090 -6270 -16080
rect -6020 -16110 -5970 -16100
rect -6310 -16140 -6010 -16110
rect -5980 -16140 -910 -16110
rect -880 -16140 -790 -16110
rect -760 -16140 8610 -16110
rect 8640 -16140 12040 -16110
rect 12070 -16140 21440 -16110
rect 21470 -16140 21560 -16110
rect 21590 -16140 23620 -16110
rect -6020 -16150 -5970 -16140
rect -6320 -16170 -6270 -16160
rect -6320 -16200 -6310 -16170
rect -6280 -16200 23620 -16170
rect -6320 -16210 -6270 -16200
rect -5820 -16230 -5770 -16220
rect -6310 -16260 -5810 -16230
rect -5780 -16260 1820 -16230
rect 1850 -16260 1910 -16230
rect 1940 -16260 3700 -16230
rect 3730 -16260 3790 -16230
rect 3820 -16260 5670 -16230
rect 5700 -16260 7550 -16230
rect 7580 -16260 13100 -16230
rect 13130 -16260 14980 -16230
rect 15010 -16260 16860 -16230
rect 16890 -16260 16950 -16230
rect 16980 -16260 18740 -16230
rect 18770 -16260 18830 -16230
rect 18860 -16260 23620 -16230
rect -5820 -16270 -5770 -16260
rect -6320 -16290 -6270 -16280
rect -6320 -16320 -6310 -16290
rect -6280 -16320 23620 -16290
rect -6320 -16330 -6270 -16320
rect -5620 -16350 -5570 -16340
rect -6310 -16380 -5610 -16350
rect -5580 -16380 2030 -16350
rect 2060 -16380 7670 -16350
rect 7700 -16380 12980 -16350
rect 13010 -16380 18620 -16350
rect 18650 -16380 23620 -16350
rect -5620 -16390 -5570 -16380
rect -6320 -16410 -6270 -16400
rect -6320 -16440 -6310 -16410
rect -6280 -16440 23620 -16410
rect -6320 -16450 -6270 -16440
rect -5420 -16470 -5370 -16460
rect -6310 -16500 -5410 -16470
rect -5380 -16500 3910 -16470
rect 3940 -16500 5790 -16470
rect 5820 -16500 14860 -16470
rect 14890 -16500 16740 -16470
rect 16770 -16500 23620 -16470
rect -5420 -16510 -5370 -16500
rect -6320 -16530 -6270 -16520
rect -6320 -16560 -6310 -16530
rect -6280 -16560 23620 -16530
rect -6320 -16570 -6270 -16560
rect -5220 -16590 -5170 -16580
rect -6310 -16620 -5210 -16590
rect -5180 -16620 970 -16590
rect 1000 -16620 1910 -16590
rect 1940 -16620 2760 -16590
rect 2790 -16620 6610 -16590
rect 6640 -16620 7550 -16590
rect 7580 -16620 8400 -16590
rect 8430 -16620 12250 -16590
rect 12280 -16620 13100 -16590
rect 13130 -16620 14040 -16590
rect 14070 -16620 17890 -16590
rect 17920 -16620 18740 -16590
rect 18770 -16620 19680 -16590
rect 19710 -16620 23620 -16590
rect -5220 -16630 -5170 -16620
rect -6320 -16650 -6270 -16640
rect -6320 -16680 -6310 -16650
rect -6280 -16680 23620 -16650
rect -6320 -16690 -6270 -16680
rect -6310 -16720 23620 -16710
rect -6310 -16860 -5000 -16720
rect -4790 -16860 9430 -16720
rect 9460 -16860 10280 -16720
rect 10310 -16860 10370 -16720
rect 10400 -16860 11220 -16720
rect 11250 -16860 23620 -16720
rect -6310 -16870 23620 -16860
rect 24260 -16720 24420 -16710
rect 24260 -16860 24270 -16720
rect 24410 -16860 24420 -16720
rect 24260 -16870 24420 -16860
rect -6320 -16900 -6270 -16890
rect -6320 -16930 -6310 -16900
rect -6280 -16930 23620 -16900
rect -6320 -16940 -6270 -16930
rect -4620 -16960 -4570 -16950
rect -6310 -16990 -4610 -16960
rect -4580 -16990 2850 -16960
rect 2880 -16990 3790 -16960
rect 3820 -16990 4640 -16960
rect 4670 -16990 4730 -16960
rect 4760 -16990 5670 -16960
rect 5700 -16990 6520 -16960
rect 6550 -16990 14130 -16960
rect 14160 -16990 14980 -16960
rect 15010 -16990 15920 -16960
rect 15950 -16990 16010 -16960
rect 16040 -16990 16860 -16960
rect 16890 -16990 17800 -16960
rect 17830 -16990 23620 -16960
rect -4620 -17000 -4570 -16990
rect -6320 -17020 -6270 -17010
rect -6320 -17050 -6310 -17020
rect -6280 -17050 23620 -17020
rect -6320 -17060 -6270 -17050
rect -4420 -17080 -4370 -17070
rect -6310 -17110 -4410 -17080
rect -4380 -17110 1700 -17080
rect 1730 -17110 2640 -17080
rect 2670 -17110 2760 -17080
rect 2790 -17110 3580 -17080
rect 3610 -17110 4520 -17080
rect 4550 -17110 5460 -17080
rect 5490 -17110 5580 -17080
rect 5610 -17110 6400 -17080
rect 6430 -17110 7340 -17080
rect 7370 -17110 8280 -17080
rect 8310 -17110 8400 -17080
rect 8430 -17110 12250 -17080
rect 12280 -17110 12370 -17080
rect 12400 -17110 13310 -17080
rect 13340 -17110 14250 -17080
rect 14280 -17110 15070 -17080
rect 15100 -17110 15190 -17080
rect 15220 -17110 16130 -17080
rect 16160 -17110 17070 -17080
rect 17100 -17110 17890 -17080
rect 17920 -17110 18010 -17080
rect 18040 -17110 18950 -17080
rect 18980 -17110 23620 -17080
rect -4420 -17120 -4370 -17110
rect -6320 -17140 -6270 -17130
rect -6320 -17170 -6310 -17140
rect -6280 -17170 23620 -17140
rect -6320 -17180 -6270 -17170
rect -4220 -17200 -4170 -17190
rect -6310 -17230 -4210 -17200
rect -4180 -17230 7460 -17200
rect 7490 -17230 8490 -17200
rect 8520 -17230 9550 -17200
rect 9580 -17230 11100 -17200
rect 11130 -17230 12160 -17200
rect 12190 -17230 13190 -17200
rect 13220 -17230 23620 -17200
rect -4220 -17240 -4170 -17230
rect -6320 -17260 -6270 -17250
rect -6320 -17290 -6310 -17260
rect -6280 -17290 23620 -17260
rect -6320 -17300 -6270 -17290
rect -4020 -17320 -3970 -17310
rect -6310 -17350 -4010 -17320
rect -3980 -17350 4640 -17320
rect 4670 -17350 6520 -17320
rect 6550 -17350 9340 -17320
rect 9370 -17350 10160 -17320
rect 10190 -17350 10490 -17320
rect 10520 -17350 11310 -17320
rect 11340 -17350 14130 -17320
rect 14160 -17350 16010 -17320
rect 16040 -17350 23620 -17320
rect -4020 -17360 -3970 -17350
rect -6320 -17380 -6270 -17370
rect -6320 -17410 -6310 -17380
rect -6280 -17410 23620 -17380
rect -6320 -17420 -6270 -17410
rect -3820 -17440 -3770 -17430
rect -6310 -17470 -3810 -17440
rect -3780 -17470 760 -17440
rect 790 -17470 880 -17440
rect 910 -17470 9220 -17440
rect 9250 -17470 11430 -17440
rect 11460 -17470 19770 -17440
rect 19800 -17470 19890 -17440
rect 19920 -17470 23620 -17440
rect -3820 -17480 -3770 -17470
rect -6320 -17500 -6270 -17490
rect -6320 -17530 -6310 -17500
rect -6280 -17530 23620 -17500
rect -6320 -17540 -6270 -17530
rect -3620 -17560 -3570 -17550
rect -6310 -17590 -3610 -17560
rect -3580 -17590 -2060 -17560
rect -2030 -17590 -1120 -17560
rect -1090 -17590 -910 -17560
rect -880 -17590 -180 -17560
rect -150 -17590 30 -17560
rect 60 -17590 20620 -17560
rect 20650 -17590 20830 -17560
rect 20860 -17590 21560 -17560
rect 21590 -17590 21770 -17560
rect 21800 -17590 22710 -17560
rect 22740 -17590 23620 -17560
rect -3620 -17600 -3570 -17590
rect -6320 -17620 -6270 -17610
rect -6120 -17620 -6070 -17610
rect -5920 -17620 -5870 -17610
rect -5720 -17620 -5670 -17610
rect -5520 -17620 -5470 -17610
rect -5320 -17620 -5270 -17610
rect -5120 -17620 -5070 -17610
rect -4720 -17620 -4670 -17610
rect -4520 -17620 -4470 -17610
rect -4320 -17620 -4270 -17610
rect -4120 -17620 -4070 -17610
rect -3920 -17620 -3870 -17610
rect -3720 -17620 -3670 -17610
rect -3520 -17620 -3470 -17610
rect -6320 -17650 -6310 -17620
rect -6280 -17650 -6110 -17620
rect -6080 -17650 -5910 -17620
rect -5880 -17650 -5710 -17620
rect -5680 -17650 -5510 -17620
rect -5480 -17650 -5310 -17620
rect -5280 -17650 -5110 -17620
rect -5080 -17650 -4710 -17620
rect -4680 -17650 -4510 -17620
rect -4480 -17650 -4310 -17620
rect -4280 -17650 -4110 -17620
rect -4080 -17650 -3910 -17620
rect -3880 -17650 -3710 -17620
rect -3680 -17650 -3510 -17620
rect -3480 -17650 23620 -17620
rect -6320 -17660 -6270 -17650
rect -6120 -17660 -6070 -17650
rect -5920 -17660 -5870 -17650
rect -5720 -17660 -5670 -17650
rect -5520 -17660 -5470 -17650
rect -5320 -17660 -5270 -17650
rect -5120 -17660 -5070 -17650
rect -4720 -17660 -4670 -17650
rect -4520 -17660 -4470 -17650
rect -4320 -17660 -4270 -17650
rect -4120 -17660 -4070 -17650
rect -3920 -17660 -3870 -17650
rect -3720 -17660 -3670 -17650
rect -3520 -17660 -3470 -17650
rect -3100 -18910 24420 -18900
rect -3100 -19050 -3090 -18910
rect -2950 -19050 -2790 -18910
rect -2760 -19050 -1940 -18910
rect -1910 -19050 -1850 -18910
rect -1820 -19050 -910 -18910
rect -880 -19050 970 -18910
rect 1000 -19050 2850 -18910
rect 2880 -19050 4730 -18910
rect 4760 -19050 6610 -18910
rect 6640 -19050 9430 -18910
rect 9460 -19050 11220 -18910
rect 11250 -19050 14040 -18910
rect 14070 -19050 15920 -18910
rect 15950 -19050 17800 -18910
rect 17830 -19050 19680 -18910
rect 19710 -19050 21560 -18910
rect 21590 -19050 22500 -18910
rect 22530 -19050 22590 -18910
rect 22620 -19050 23440 -18910
rect 23470 -19050 23630 -18910
rect 23770 -19050 24420 -18910
rect -3100 -19070 24420 -19050
rect -3100 -19210 -3090 -19070
rect -2950 -19210 -2790 -19070
rect -2760 -19210 -1940 -19070
rect -1910 -19210 -1850 -19070
rect -1820 -19210 -910 -19070
rect -880 -19210 970 -19070
rect 1000 -19210 2850 -19070
rect 2880 -19210 4730 -19070
rect 4760 -19210 6610 -19070
rect 6640 -19210 9430 -19070
rect 9460 -19210 11220 -19070
rect 11250 -19210 14040 -19070
rect 14070 -19210 15920 -19070
rect 15950 -19210 17800 -19070
rect 17830 -19210 19680 -19070
rect 19710 -19210 21560 -19070
rect 21590 -19210 22500 -19070
rect 22530 -19210 22590 -19070
rect 22620 -19210 23440 -19070
rect 23470 -19210 23630 -19070
rect 23770 -19210 24420 -19070
rect -3100 -19220 24420 -19210
rect -6320 -20470 -6270 -20460
rect -6120 -20470 -6070 -20460
rect -5920 -20470 -5870 -20460
rect -5720 -20470 -5670 -20460
rect -5520 -20470 -5470 -20460
rect -5320 -20470 -5270 -20460
rect -5120 -20470 -5070 -20460
rect -4720 -20470 -4670 -20460
rect -4520 -20470 -4470 -20460
rect -4320 -20470 -4270 -20460
rect -4120 -20470 -4070 -20460
rect -3920 -20470 -3870 -20460
rect -3720 -20470 -3670 -20460
rect -3520 -20470 -3470 -20460
rect -6320 -20500 -6310 -20470
rect -6280 -20500 -6110 -20470
rect -6080 -20500 -5910 -20470
rect -5880 -20500 -5710 -20470
rect -5680 -20500 -5510 -20470
rect -5480 -20500 -5310 -20470
rect -5280 -20500 -5110 -20470
rect -5080 -20500 -4710 -20470
rect -4680 -20500 -4510 -20470
rect -4480 -20500 -4310 -20470
rect -4280 -20500 -4110 -20470
rect -4080 -20500 -3910 -20470
rect -3880 -20500 -3710 -20470
rect -3680 -20500 -3510 -20470
rect -3480 -20500 23620 -20470
rect -6320 -20510 -6270 -20500
rect -6120 -20510 -6070 -20500
rect -5920 -20510 -5870 -20500
rect -5720 -20510 -5670 -20500
rect -5520 -20510 -5470 -20500
rect -5320 -20510 -5270 -20500
rect -5120 -20510 -5070 -20500
rect -4720 -20510 -4670 -20500
rect -4520 -20510 -4470 -20500
rect -4320 -20510 -4270 -20500
rect -4120 -20510 -4070 -20500
rect -3920 -20510 -3870 -20500
rect -3720 -20510 -3670 -20500
rect -3520 -20510 -3470 -20500
rect -3620 -20530 -3570 -20520
rect -6310 -20560 -3610 -20530
rect -3580 -20560 -2060 -20530
rect -2030 -20560 -1120 -20530
rect -1090 -20560 -910 -20530
rect -880 -20560 -180 -20530
rect -150 -20560 30 -20530
rect 60 -20560 20620 -20530
rect 20650 -20560 20830 -20530
rect 20860 -20560 21560 -20530
rect 21590 -20560 21770 -20530
rect 21800 -20560 22710 -20530
rect 22740 -20560 23620 -20530
rect -3620 -20570 -3570 -20560
rect -6320 -20590 -6270 -20580
rect -6320 -20620 -6310 -20590
rect -6280 -20620 23620 -20590
rect -6320 -20630 -6270 -20620
rect -3820 -20650 -3770 -20640
rect -6310 -20680 -3810 -20650
rect -3780 -20680 760 -20650
rect 790 -20680 880 -20650
rect 910 -20680 9220 -20650
rect 9250 -20680 11430 -20650
rect 11460 -20680 19770 -20650
rect 19800 -20680 19890 -20650
rect 19920 -20680 23620 -20650
rect -3820 -20690 -3770 -20680
rect -6320 -20710 -6270 -20700
rect -6320 -20740 -6310 -20710
rect -6280 -20740 23620 -20710
rect -6320 -20750 -6270 -20740
rect -4020 -20770 -3970 -20760
rect -6310 -20800 -4010 -20770
rect -3980 -20800 4640 -20770
rect 4670 -20800 6520 -20770
rect 6550 -20800 9340 -20770
rect 9370 -20800 10160 -20770
rect 10190 -20800 10490 -20770
rect 10520 -20800 11310 -20770
rect 11340 -20800 14130 -20770
rect 14160 -20800 16010 -20770
rect 16040 -20800 23620 -20770
rect -4020 -20810 -3970 -20800
rect -6320 -20830 -6270 -20820
rect -6320 -20860 -6310 -20830
rect -6280 -20860 23620 -20830
rect -6320 -20870 -6270 -20860
rect -4220 -20890 -4170 -20880
rect -6310 -20920 -4210 -20890
rect -4180 -20920 7460 -20890
rect 7490 -20920 8490 -20890
rect 8520 -20920 9550 -20890
rect 9580 -20920 11100 -20890
rect 11130 -20920 12160 -20890
rect 12190 -20920 13190 -20890
rect 13220 -20920 23620 -20890
rect -4220 -20930 -4170 -20920
rect -6320 -20950 -6270 -20940
rect -6320 -20980 -6310 -20950
rect -6280 -20980 23620 -20950
rect -6320 -20990 -6270 -20980
rect -4420 -21010 -4370 -21000
rect -6310 -21040 -4410 -21010
rect -4380 -21040 1700 -21010
rect 1730 -21040 2640 -21010
rect 2670 -21040 2760 -21010
rect 2790 -21040 3580 -21010
rect 3610 -21040 4520 -21010
rect 4550 -21040 5460 -21010
rect 5490 -21040 5580 -21010
rect 5610 -21040 6400 -21010
rect 6430 -21040 7340 -21010
rect 7370 -21040 8280 -21010
rect 8310 -21040 8400 -21010
rect 8430 -21040 12250 -21010
rect 12280 -21040 12370 -21010
rect 12400 -21040 13310 -21010
rect 13340 -21040 14250 -21010
rect 14280 -21040 15070 -21010
rect 15100 -21040 15190 -21010
rect 15220 -21040 16130 -21010
rect 16160 -21040 17070 -21010
rect 17100 -21040 17890 -21010
rect 17920 -21040 18010 -21010
rect 18040 -21040 18950 -21010
rect 18980 -21040 23620 -21010
rect -4420 -21050 -4370 -21040
rect -6320 -21070 -6270 -21060
rect -6320 -21100 -6310 -21070
rect -6280 -21100 23620 -21070
rect -6320 -21110 -6270 -21100
rect -4620 -21130 -4570 -21120
rect -6310 -21160 -4610 -21130
rect -4580 -21160 2850 -21130
rect 2880 -21160 3790 -21130
rect 3820 -21160 4640 -21130
rect 4670 -21160 4730 -21130
rect 4760 -21160 5670 -21130
rect 5700 -21160 6520 -21130
rect 6550 -21160 14130 -21130
rect 14160 -21160 14980 -21130
rect 15010 -21160 15920 -21130
rect 15950 -21160 16010 -21130
rect 16040 -21160 16860 -21130
rect 16890 -21160 17800 -21130
rect 17830 -21160 23620 -21130
rect -4620 -21170 -4570 -21160
rect -6320 -21190 -6270 -21180
rect -6320 -21220 -6310 -21190
rect -6280 -21220 23620 -21190
rect -6320 -21230 -6270 -21220
rect -6310 -21260 23620 -21250
rect -6310 -21400 -5000 -21260
rect -4790 -21400 9430 -21260
rect 9460 -21400 10280 -21260
rect 10310 -21400 10370 -21260
rect 10400 -21400 11220 -21260
rect 11250 -21400 23620 -21260
rect -6310 -21410 23620 -21400
rect 24260 -21260 24420 -21250
rect 24260 -21400 24270 -21260
rect 24410 -21400 24420 -21260
rect 24260 -21410 24420 -21400
rect -6320 -21440 -6270 -21430
rect -6320 -21470 -6310 -21440
rect -6280 -21470 23620 -21440
rect -6320 -21480 -6270 -21470
rect -5220 -21500 -5170 -21490
rect -6310 -21530 -5210 -21500
rect -5180 -21530 970 -21500
rect 1000 -21530 1910 -21500
rect 1940 -21530 2760 -21500
rect 2790 -21530 6610 -21500
rect 6640 -21530 7550 -21500
rect 7580 -21530 8400 -21500
rect 8430 -21530 12250 -21500
rect 12280 -21530 13100 -21500
rect 13130 -21530 14040 -21500
rect 14070 -21530 17890 -21500
rect 17920 -21530 18740 -21500
rect 18770 -21530 19680 -21500
rect 19710 -21530 23620 -21500
rect -5220 -21540 -5170 -21530
rect -6320 -21560 -6270 -21550
rect -6320 -21590 -6310 -21560
rect -6280 -21590 23620 -21560
rect -6320 -21600 -6270 -21590
rect -5420 -21620 -5370 -21610
rect -6310 -21650 -5410 -21620
rect -5380 -21650 3910 -21620
rect 3940 -21650 5790 -21620
rect 5820 -21650 14860 -21620
rect 14890 -21650 16740 -21620
rect 16770 -21650 23620 -21620
rect -5420 -21660 -5370 -21650
rect -6320 -21680 -6270 -21670
rect -6320 -21710 -6310 -21680
rect -6280 -21710 23620 -21680
rect -6320 -21720 -6270 -21710
rect -5620 -21740 -5570 -21730
rect -6310 -21770 -5610 -21740
rect -5580 -21770 2030 -21740
rect 2060 -21770 7670 -21740
rect 7700 -21770 12980 -21740
rect 13010 -21770 18620 -21740
rect 18650 -21770 23620 -21740
rect -5620 -21780 -5570 -21770
rect -6320 -21800 -6270 -21790
rect -6320 -21830 -6310 -21800
rect -6280 -21830 23620 -21800
rect -6320 -21840 -6270 -21830
rect -5820 -21860 -5770 -21850
rect -6310 -21890 -5810 -21860
rect -5780 -21890 1820 -21860
rect 1850 -21890 1910 -21860
rect 1940 -21890 3700 -21860
rect 3730 -21890 3790 -21860
rect 3820 -21890 5670 -21860
rect 5700 -21890 7550 -21860
rect 7580 -21890 13100 -21860
rect 13130 -21890 14980 -21860
rect 15010 -21890 16860 -21860
rect 16890 -21890 16950 -21860
rect 16980 -21890 18740 -21860
rect 18770 -21890 18830 -21860
rect 18860 -21890 23620 -21860
rect -5820 -21900 -5770 -21890
rect -6320 -21920 -6270 -21910
rect -6320 -21950 -6310 -21920
rect -6280 -21950 23620 -21920
rect -6320 -21960 -6270 -21950
rect -6020 -21980 -5970 -21970
rect -6310 -22010 -6010 -21980
rect -5980 -22010 -910 -21980
rect -880 -22010 -790 -21980
rect -760 -22010 8610 -21980
rect 8640 -22010 12040 -21980
rect 12070 -22010 21440 -21980
rect 21470 -22010 21560 -21980
rect 21590 -22010 23620 -21980
rect -6020 -22020 -5970 -22010
rect -6320 -22040 -6270 -22030
rect -6320 -22070 -6310 -22040
rect -6280 -22070 23620 -22040
rect -6320 -22080 -6270 -22070
rect -6220 -22100 -6170 -22090
rect -6310 -22130 -6210 -22100
rect -6180 -22130 -2670 -22100
rect -2640 -22130 -1730 -22100
rect -1700 -22130 -1000 -22100
rect -970 -22130 -60 -22100
rect -30 -22130 150 -22100
rect 180 -22130 1090 -22100
rect 1120 -22130 2970 -22100
rect 3000 -22130 4850 -22100
rect 4880 -22130 6730 -22100
rect 6760 -22130 13920 -22100
rect 13950 -22130 15800 -22100
rect 15830 -22130 17680 -22100
rect 17710 -22130 19560 -22100
rect 19590 -22130 20500 -22100
rect 20530 -22130 20710 -22100
rect 20740 -22130 21650 -22100
rect 21680 -22130 22380 -22100
rect 22410 -22130 23320 -22100
rect 23350 -22130 23620 -22100
rect -6220 -22140 -6170 -22130
rect -6320 -22160 -6270 -22150
rect -6120 -22160 -6070 -22150
rect -5920 -22160 -5870 -22150
rect -5720 -22160 -5670 -22150
rect -5520 -22160 -5470 -22150
rect -5320 -22160 -5270 -22150
rect -5120 -22160 -5070 -22150
rect -4720 -22160 -4670 -22150
rect -4520 -22160 -4470 -22150
rect -4320 -22160 -4270 -22150
rect -4120 -22160 -4070 -22150
rect -3920 -22160 -3870 -22150
rect -3720 -22160 -3670 -22150
rect -3520 -22160 -3470 -22150
rect -6320 -22190 -6310 -22160
rect -6280 -22190 -6110 -22160
rect -6080 -22190 -5910 -22160
rect -5880 -22190 -5710 -22160
rect -5680 -22190 -5510 -22160
rect -5480 -22190 -5310 -22160
rect -5280 -22190 -5110 -22160
rect -5080 -22190 -4710 -22160
rect -4680 -22190 -4510 -22160
rect -4480 -22190 -4310 -22160
rect -4280 -22190 -4110 -22160
rect -4080 -22190 -3910 -22160
rect -3880 -22190 -3710 -22160
rect -3680 -22190 -3510 -22160
rect -3480 -22190 23620 -22160
rect -6320 -22200 -6270 -22190
rect -6120 -22200 -6070 -22190
rect -5920 -22200 -5870 -22190
rect -5720 -22200 -5670 -22190
rect -5520 -22200 -5470 -22190
rect -5320 -22200 -5270 -22190
rect -5120 -22200 -5070 -22190
rect -4720 -22200 -4670 -22190
rect -4520 -22200 -4470 -22190
rect -4320 -22200 -4270 -22190
rect -4120 -22200 -4070 -22190
rect -3920 -22200 -3870 -22190
rect -3720 -22200 -3670 -22190
rect -3520 -22200 -3470 -22190
rect -3420 -25190 24420 -25180
rect -3420 -25330 -3410 -25190
rect -3270 -25330 -2790 -25190
rect -2760 -25330 -1940 -25190
rect -1910 -25330 -1000 -25190
rect -970 -25330 880 -25190
rect 910 -25330 1820 -25190
rect 1850 -25330 3700 -25190
rect 3730 -25330 5580 -25190
rect 5610 -25330 7460 -25190
rect 7490 -25330 10280 -25190
rect 10310 -25330 10370 -25190
rect 10400 -25330 13190 -25190
rect 13220 -25330 15070 -25190
rect 15100 -25330 16950 -25190
rect 16980 -25330 18830 -25190
rect 18860 -25330 19770 -25190
rect 19800 -25330 21650 -25190
rect 21680 -25330 22590 -25190
rect 22620 -25330 23440 -25190
rect 23470 -25330 23950 -25190
rect 24090 -25330 24420 -25190
rect -3420 -25340 24420 -25330
<< via2 >>
rect -3410 -370 -3270 -230
rect 23950 -370 24090 -230
rect -6310 -3400 -6280 -3370
rect -6110 -3400 -6080 -3370
rect -5910 -3400 -5880 -3370
rect -5710 -3400 -5680 -3370
rect -5510 -3400 -5480 -3370
rect -5310 -3400 -5280 -3370
rect -5110 -3400 -5080 -3370
rect -4710 -3400 -4680 -3370
rect -4510 -3400 -4480 -3370
rect -4310 -3400 -4280 -3370
rect -4110 -3400 -4080 -3370
rect -3910 -3400 -3880 -3370
rect -3710 -3400 -3680 -3370
rect -3510 -3400 -3480 -3370
rect -6210 -3460 -6180 -3430
rect -6310 -3520 -6280 -3490
rect -6010 -3580 -5980 -3550
rect -6310 -3640 -6280 -3610
rect -5810 -3700 -5780 -3670
rect -6310 -3760 -6280 -3730
rect -5610 -3820 -5580 -3790
rect -6310 -3880 -6280 -3850
rect -5410 -3940 -5380 -3910
rect -6310 -4000 -6280 -3970
rect -5210 -4060 -5180 -4030
rect -6310 -4120 -6280 -4090
rect -5000 -4300 -4790 -4160
rect 24270 -4300 24410 -4160
rect -6310 -4370 -6280 -4340
rect -4610 -4430 -4580 -4400
rect -6310 -4490 -6280 -4460
rect -4410 -4550 -4380 -4520
rect -6310 -4610 -6280 -4580
rect -4210 -4670 -4180 -4640
rect -6310 -4730 -6280 -4700
rect -4010 -4790 -3980 -4760
rect -6310 -4850 -6280 -4820
rect -3810 -4910 -3780 -4880
rect -6310 -4970 -6280 -4940
rect -3610 -5030 -3580 -5000
rect -6310 -5090 -6280 -5060
rect -6110 -5090 -6080 -5060
rect -5910 -5090 -5880 -5060
rect -5710 -5090 -5680 -5060
rect -5510 -5090 -5480 -5060
rect -5310 -5090 -5280 -5060
rect -5110 -5090 -5080 -5060
rect -4710 -5090 -4680 -5060
rect -4510 -5090 -4480 -5060
rect -4310 -5090 -4280 -5060
rect -4110 -5090 -4080 -5060
rect -3910 -5090 -3880 -5060
rect -3710 -5090 -3680 -5060
rect -3510 -5090 -3480 -5060
rect -3090 -6490 -2950 -6350
rect 23630 -6490 23770 -6350
rect -3090 -6650 -2950 -6510
rect 23630 -6650 23770 -6510
rect -6310 -7940 -6280 -7910
rect -6110 -7940 -6080 -7910
rect -5910 -7940 -5880 -7910
rect -5710 -7940 -5680 -7910
rect -5510 -7940 -5480 -7910
rect -5310 -7940 -5280 -7910
rect -5110 -7940 -5080 -7910
rect -4710 -7940 -4680 -7910
rect -4510 -7940 -4480 -7910
rect -4310 -7940 -4280 -7910
rect -4110 -7940 -4080 -7910
rect -3910 -7940 -3880 -7910
rect -3710 -7940 -3680 -7910
rect -3510 -7940 -3480 -7910
rect -3610 -8000 -3580 -7970
rect -6310 -8060 -6280 -8030
rect -3810 -8120 -3780 -8090
rect -6310 -8180 -6280 -8150
rect -4010 -8240 -3980 -8210
rect -6310 -8300 -6280 -8270
rect -4210 -8360 -4180 -8330
rect -6310 -8420 -6280 -8390
rect -4410 -8480 -4380 -8450
rect -6310 -8540 -6280 -8510
rect -4610 -8600 -4580 -8570
rect -6310 -8660 -6280 -8630
rect -5000 -8840 -4790 -8700
rect 24270 -8840 24410 -8700
rect -6310 -8910 -6280 -8880
rect -5210 -8970 -5180 -8940
rect -6310 -9030 -6280 -9000
rect -5410 -9090 -5380 -9060
rect -6310 -9150 -6280 -9120
rect -5610 -9210 -5580 -9180
rect -6310 -9270 -6280 -9240
rect -5810 -9330 -5780 -9300
rect -6310 -9390 -6280 -9360
rect -6010 -9450 -5980 -9420
rect -6310 -9510 -6280 -9480
rect -6210 -9570 -6180 -9540
rect -6310 -9630 -6280 -9600
rect -6110 -9630 -6080 -9600
rect -5910 -9630 -5880 -9600
rect -5710 -9630 -5680 -9600
rect -5510 -9630 -5480 -9600
rect -5310 -9630 -5280 -9600
rect -5110 -9630 -5080 -9600
rect -4710 -9630 -4680 -9600
rect -4510 -9630 -4480 -9600
rect -4310 -9630 -4280 -9600
rect -4110 -9630 -4080 -9600
rect -3910 -9630 -3880 -9600
rect -3710 -9630 -3680 -9600
rect -3510 -9630 -3480 -9600
rect -3410 -12770 -3270 -12630
rect 23950 -12770 24090 -12630
rect -3410 -12930 -3270 -12790
rect 23950 -12930 24090 -12790
rect -6310 -15960 -6280 -15930
rect -6110 -15960 -6080 -15930
rect -5910 -15960 -5880 -15930
rect -5710 -15960 -5680 -15930
rect -5510 -15960 -5480 -15930
rect -5310 -15960 -5280 -15930
rect -5110 -15960 -5080 -15930
rect -4710 -15960 -4680 -15930
rect -4510 -15960 -4480 -15930
rect -4310 -15960 -4280 -15930
rect -4110 -15960 -4080 -15930
rect -3910 -15960 -3880 -15930
rect -3710 -15960 -3680 -15930
rect -3510 -15960 -3480 -15930
rect -6210 -16020 -6180 -15990
rect -6310 -16080 -6280 -16050
rect -6010 -16140 -5980 -16110
rect -6310 -16200 -6280 -16170
rect -5810 -16260 -5780 -16230
rect -6310 -16320 -6280 -16290
rect -5610 -16380 -5580 -16350
rect -6310 -16440 -6280 -16410
rect -5410 -16500 -5380 -16470
rect -6310 -16560 -6280 -16530
rect -5210 -16620 -5180 -16590
rect -6310 -16680 -6280 -16650
rect -5000 -16860 -4790 -16720
rect 24270 -16860 24410 -16720
rect -6310 -16930 -6280 -16900
rect -4610 -16990 -4580 -16960
rect -6310 -17050 -6280 -17020
rect -4410 -17110 -4380 -17080
rect -6310 -17170 -6280 -17140
rect -4210 -17230 -4180 -17200
rect -6310 -17290 -6280 -17260
rect -4010 -17350 -3980 -17320
rect -6310 -17410 -6280 -17380
rect -3810 -17470 -3780 -17440
rect -6310 -17530 -6280 -17500
rect -3610 -17590 -3580 -17560
rect -6310 -17650 -6280 -17620
rect -6110 -17650 -6080 -17620
rect -5910 -17650 -5880 -17620
rect -5710 -17650 -5680 -17620
rect -5510 -17650 -5480 -17620
rect -5310 -17650 -5280 -17620
rect -5110 -17650 -5080 -17620
rect -4710 -17650 -4680 -17620
rect -4510 -17650 -4480 -17620
rect -4310 -17650 -4280 -17620
rect -4110 -17650 -4080 -17620
rect -3910 -17650 -3880 -17620
rect -3710 -17650 -3680 -17620
rect -3510 -17650 -3480 -17620
rect -3090 -19050 -2950 -18910
rect 23630 -19050 23770 -18910
rect -3090 -19210 -2950 -19070
rect 23630 -19210 23770 -19070
rect -6310 -20500 -6280 -20470
rect -6110 -20500 -6080 -20470
rect -5910 -20500 -5880 -20470
rect -5710 -20500 -5680 -20470
rect -5510 -20500 -5480 -20470
rect -5310 -20500 -5280 -20470
rect -5110 -20500 -5080 -20470
rect -4710 -20500 -4680 -20470
rect -4510 -20500 -4480 -20470
rect -4310 -20500 -4280 -20470
rect -4110 -20500 -4080 -20470
rect -3910 -20500 -3880 -20470
rect -3710 -20500 -3680 -20470
rect -3510 -20500 -3480 -20470
rect -3610 -20560 -3580 -20530
rect -6310 -20620 -6280 -20590
rect -3810 -20680 -3780 -20650
rect -6310 -20740 -6280 -20710
rect -4010 -20800 -3980 -20770
rect -6310 -20860 -6280 -20830
rect -4210 -20920 -4180 -20890
rect -6310 -20980 -6280 -20950
rect -4410 -21040 -4380 -21010
rect -6310 -21100 -6280 -21070
rect -4610 -21160 -4580 -21130
rect -6310 -21220 -6280 -21190
rect -5000 -21400 -4790 -21260
rect 24270 -21400 24410 -21260
rect -6310 -21470 -6280 -21440
rect -5210 -21530 -5180 -21500
rect -6310 -21590 -6280 -21560
rect -5410 -21650 -5380 -21620
rect -6310 -21710 -6280 -21680
rect -5610 -21770 -5580 -21740
rect -6310 -21830 -6280 -21800
rect -5810 -21890 -5780 -21860
rect -6310 -21950 -6280 -21920
rect -6010 -22010 -5980 -21980
rect -6310 -22070 -6280 -22040
rect -6210 -22130 -6180 -22100
rect -6310 -22190 -6280 -22160
rect -6110 -22190 -6080 -22160
rect -5910 -22190 -5880 -22160
rect -5710 -22190 -5680 -22160
rect -5510 -22190 -5480 -22160
rect -5310 -22190 -5280 -22160
rect -5110 -22190 -5080 -22160
rect -4710 -22190 -4680 -22160
rect -4510 -22190 -4480 -22160
rect -4310 -22190 -4280 -22160
rect -4110 -22190 -4080 -22160
rect -3910 -22190 -3880 -22160
rect -3710 -22190 -3680 -22160
rect -3510 -22190 -3480 -22160
rect -3410 -25330 -3270 -25190
rect 23950 -25330 24090 -25190
<< metal3 >>
rect -6310 -3360 -6280 -220
rect -6320 -3370 -6270 -3360
rect -6320 -3400 -6310 -3370
rect -6280 -3400 -6270 -3370
rect -6320 -3410 -6270 -3400
rect -6310 -3480 -6280 -3410
rect -6210 -3420 -6180 -190
rect -6110 -3360 -6080 -220
rect -6120 -3370 -6070 -3360
rect -6120 -3400 -6110 -3370
rect -6080 -3400 -6070 -3370
rect -6120 -3410 -6070 -3400
rect -6220 -3430 -6170 -3420
rect -6220 -3460 -6210 -3430
rect -6180 -3460 -6170 -3430
rect -6220 -3470 -6170 -3460
rect -6320 -3490 -6270 -3480
rect -6320 -3520 -6310 -3490
rect -6280 -3520 -6270 -3490
rect -6320 -3530 -6270 -3520
rect -6310 -3600 -6280 -3530
rect -6320 -3610 -6270 -3600
rect -6320 -3640 -6310 -3610
rect -6280 -3640 -6270 -3610
rect -6320 -3650 -6270 -3640
rect -6310 -3720 -6280 -3650
rect -6320 -3730 -6270 -3720
rect -6320 -3760 -6310 -3730
rect -6280 -3760 -6270 -3730
rect -6320 -3770 -6270 -3760
rect -6310 -3840 -6280 -3770
rect -6320 -3850 -6270 -3840
rect -6320 -3880 -6310 -3850
rect -6280 -3880 -6270 -3850
rect -6320 -3890 -6270 -3880
rect -6310 -3960 -6280 -3890
rect -6320 -3970 -6270 -3960
rect -6320 -4000 -6310 -3970
rect -6280 -4000 -6270 -3970
rect -6320 -4010 -6270 -4000
rect -6310 -4080 -6280 -4010
rect -6320 -4090 -6270 -4080
rect -6320 -4120 -6310 -4090
rect -6280 -4120 -6270 -4090
rect -6320 -4130 -6270 -4120
rect -6310 -4330 -6280 -4130
rect -6320 -4340 -6270 -4330
rect -6320 -4370 -6310 -4340
rect -6280 -4370 -6270 -4340
rect -6320 -4380 -6270 -4370
rect -6310 -4450 -6280 -4380
rect -6320 -4460 -6270 -4450
rect -6320 -4490 -6310 -4460
rect -6280 -4490 -6270 -4460
rect -6320 -4500 -6270 -4490
rect -6310 -4570 -6280 -4500
rect -6320 -4580 -6270 -4570
rect -6320 -4610 -6310 -4580
rect -6280 -4610 -6270 -4580
rect -6320 -4620 -6270 -4610
rect -6310 -4690 -6280 -4620
rect -6320 -4700 -6270 -4690
rect -6320 -4730 -6310 -4700
rect -6280 -4730 -6270 -4700
rect -6320 -4740 -6270 -4730
rect -6310 -4810 -6280 -4740
rect -6320 -4820 -6270 -4810
rect -6320 -4850 -6310 -4820
rect -6280 -4850 -6270 -4820
rect -6320 -4860 -6270 -4850
rect -6310 -4930 -6280 -4860
rect -6320 -4940 -6270 -4930
rect -6320 -4970 -6310 -4940
rect -6280 -4970 -6270 -4940
rect -6320 -4980 -6270 -4970
rect -6310 -5050 -6280 -4980
rect -6320 -5060 -6270 -5050
rect -6320 -5090 -6310 -5060
rect -6280 -5090 -6270 -5060
rect -6320 -5100 -6270 -5090
rect -6310 -7900 -6280 -5100
rect -6320 -7910 -6270 -7900
rect -6320 -7940 -6310 -7910
rect -6280 -7940 -6270 -7910
rect -6320 -7950 -6270 -7940
rect -6310 -8020 -6280 -7950
rect -6320 -8030 -6270 -8020
rect -6320 -8060 -6310 -8030
rect -6280 -8060 -6270 -8030
rect -6320 -8070 -6270 -8060
rect -6310 -8140 -6280 -8070
rect -6320 -8150 -6270 -8140
rect -6320 -8180 -6310 -8150
rect -6280 -8180 -6270 -8150
rect -6320 -8190 -6270 -8180
rect -6310 -8260 -6280 -8190
rect -6320 -8270 -6270 -8260
rect -6320 -8300 -6310 -8270
rect -6280 -8300 -6270 -8270
rect -6320 -8310 -6270 -8300
rect -6310 -8380 -6280 -8310
rect -6320 -8390 -6270 -8380
rect -6320 -8420 -6310 -8390
rect -6280 -8420 -6270 -8390
rect -6320 -8430 -6270 -8420
rect -6310 -8500 -6280 -8430
rect -6320 -8510 -6270 -8500
rect -6320 -8540 -6310 -8510
rect -6280 -8540 -6270 -8510
rect -6320 -8550 -6270 -8540
rect -6310 -8620 -6280 -8550
rect -6320 -8630 -6270 -8620
rect -6320 -8660 -6310 -8630
rect -6280 -8660 -6270 -8630
rect -6320 -8670 -6270 -8660
rect -6310 -8870 -6280 -8670
rect -6320 -8880 -6270 -8870
rect -6320 -8910 -6310 -8880
rect -6280 -8910 -6270 -8880
rect -6320 -8920 -6270 -8910
rect -6310 -8990 -6280 -8920
rect -6320 -9000 -6270 -8990
rect -6320 -9030 -6310 -9000
rect -6280 -9030 -6270 -9000
rect -6320 -9040 -6270 -9030
rect -6310 -9110 -6280 -9040
rect -6320 -9120 -6270 -9110
rect -6320 -9150 -6310 -9120
rect -6280 -9150 -6270 -9120
rect -6320 -9160 -6270 -9150
rect -6310 -9230 -6280 -9160
rect -6320 -9240 -6270 -9230
rect -6320 -9270 -6310 -9240
rect -6280 -9270 -6270 -9240
rect -6320 -9280 -6270 -9270
rect -6310 -9350 -6280 -9280
rect -6320 -9360 -6270 -9350
rect -6320 -9390 -6310 -9360
rect -6280 -9390 -6270 -9360
rect -6320 -9400 -6270 -9390
rect -6310 -9470 -6280 -9400
rect -6320 -9480 -6270 -9470
rect -6320 -9510 -6310 -9480
rect -6280 -9510 -6270 -9480
rect -6320 -9520 -6270 -9510
rect -6310 -9590 -6280 -9520
rect -6210 -9530 -6180 -3470
rect -6110 -5050 -6080 -3410
rect -6010 -3540 -5980 -190
rect -5910 -3360 -5880 -220
rect -5920 -3370 -5870 -3360
rect -5920 -3400 -5910 -3370
rect -5880 -3400 -5870 -3370
rect -5920 -3410 -5870 -3400
rect -6020 -3550 -5970 -3540
rect -6020 -3580 -6010 -3550
rect -5980 -3580 -5970 -3550
rect -6020 -3590 -5970 -3580
rect -6120 -5060 -6070 -5050
rect -6120 -5090 -6110 -5060
rect -6080 -5090 -6070 -5060
rect -6120 -5100 -6070 -5090
rect -6110 -7900 -6080 -5100
rect -6120 -7910 -6070 -7900
rect -6120 -7940 -6110 -7910
rect -6080 -7940 -6070 -7910
rect -6120 -7950 -6070 -7940
rect -6220 -9540 -6170 -9530
rect -6220 -9570 -6210 -9540
rect -6180 -9570 -6170 -9540
rect -6220 -9580 -6170 -9570
rect -6320 -9600 -6270 -9590
rect -6320 -9630 -6310 -9600
rect -6280 -9630 -6270 -9600
rect -6320 -9640 -6270 -9630
rect -6310 -15920 -6280 -9640
rect -6320 -15930 -6270 -15920
rect -6320 -15960 -6310 -15930
rect -6280 -15960 -6270 -15930
rect -6320 -15970 -6270 -15960
rect -6310 -16040 -6280 -15970
rect -6210 -15980 -6180 -9580
rect -6110 -9590 -6080 -7950
rect -6010 -9410 -5980 -3590
rect -5910 -5050 -5880 -3410
rect -5810 -3660 -5780 -190
rect -5710 -3360 -5680 -220
rect -5720 -3370 -5670 -3360
rect -5720 -3400 -5710 -3370
rect -5680 -3400 -5670 -3370
rect -5720 -3410 -5670 -3400
rect -5820 -3670 -5770 -3660
rect -5820 -3700 -5810 -3670
rect -5780 -3700 -5770 -3670
rect -5820 -3710 -5770 -3700
rect -5920 -5060 -5870 -5050
rect -5920 -5090 -5910 -5060
rect -5880 -5090 -5870 -5060
rect -5920 -5100 -5870 -5090
rect -5910 -7900 -5880 -5100
rect -5920 -7910 -5870 -7900
rect -5920 -7940 -5910 -7910
rect -5880 -7940 -5870 -7910
rect -5920 -7950 -5870 -7940
rect -6020 -9420 -5970 -9410
rect -6020 -9450 -6010 -9420
rect -5980 -9450 -5970 -9420
rect -6020 -9460 -5970 -9450
rect -6120 -9600 -6070 -9590
rect -6120 -9630 -6110 -9600
rect -6080 -9630 -6070 -9600
rect -6120 -9640 -6070 -9630
rect -6110 -15920 -6080 -9640
rect -6120 -15930 -6070 -15920
rect -6120 -15960 -6110 -15930
rect -6080 -15960 -6070 -15930
rect -6120 -15970 -6070 -15960
rect -6220 -15990 -6170 -15980
rect -6220 -16020 -6210 -15990
rect -6180 -16020 -6170 -15990
rect -6220 -16030 -6170 -16020
rect -6320 -16050 -6270 -16040
rect -6320 -16080 -6310 -16050
rect -6280 -16080 -6270 -16050
rect -6320 -16090 -6270 -16080
rect -6310 -16160 -6280 -16090
rect -6320 -16170 -6270 -16160
rect -6320 -16200 -6310 -16170
rect -6280 -16200 -6270 -16170
rect -6320 -16210 -6270 -16200
rect -6310 -16280 -6280 -16210
rect -6320 -16290 -6270 -16280
rect -6320 -16320 -6310 -16290
rect -6280 -16320 -6270 -16290
rect -6320 -16330 -6270 -16320
rect -6310 -16400 -6280 -16330
rect -6320 -16410 -6270 -16400
rect -6320 -16440 -6310 -16410
rect -6280 -16440 -6270 -16410
rect -6320 -16450 -6270 -16440
rect -6310 -16520 -6280 -16450
rect -6320 -16530 -6270 -16520
rect -6320 -16560 -6310 -16530
rect -6280 -16560 -6270 -16530
rect -6320 -16570 -6270 -16560
rect -6310 -16640 -6280 -16570
rect -6320 -16650 -6270 -16640
rect -6320 -16680 -6310 -16650
rect -6280 -16680 -6270 -16650
rect -6320 -16690 -6270 -16680
rect -6310 -16890 -6280 -16690
rect -6320 -16900 -6270 -16890
rect -6320 -16930 -6310 -16900
rect -6280 -16930 -6270 -16900
rect -6320 -16940 -6270 -16930
rect -6310 -17010 -6280 -16940
rect -6320 -17020 -6270 -17010
rect -6320 -17050 -6310 -17020
rect -6280 -17050 -6270 -17020
rect -6320 -17060 -6270 -17050
rect -6310 -17130 -6280 -17060
rect -6320 -17140 -6270 -17130
rect -6320 -17170 -6310 -17140
rect -6280 -17170 -6270 -17140
rect -6320 -17180 -6270 -17170
rect -6310 -17250 -6280 -17180
rect -6320 -17260 -6270 -17250
rect -6320 -17290 -6310 -17260
rect -6280 -17290 -6270 -17260
rect -6320 -17300 -6270 -17290
rect -6310 -17370 -6280 -17300
rect -6320 -17380 -6270 -17370
rect -6320 -17410 -6310 -17380
rect -6280 -17410 -6270 -17380
rect -6320 -17420 -6270 -17410
rect -6310 -17490 -6280 -17420
rect -6320 -17500 -6270 -17490
rect -6320 -17530 -6310 -17500
rect -6280 -17530 -6270 -17500
rect -6320 -17540 -6270 -17530
rect -6310 -17610 -6280 -17540
rect -6320 -17620 -6270 -17610
rect -6320 -17650 -6310 -17620
rect -6280 -17650 -6270 -17620
rect -6320 -17660 -6270 -17650
rect -6310 -20460 -6280 -17660
rect -6320 -20470 -6270 -20460
rect -6320 -20500 -6310 -20470
rect -6280 -20500 -6270 -20470
rect -6320 -20510 -6270 -20500
rect -6310 -20580 -6280 -20510
rect -6320 -20590 -6270 -20580
rect -6320 -20620 -6310 -20590
rect -6280 -20620 -6270 -20590
rect -6320 -20630 -6270 -20620
rect -6310 -20700 -6280 -20630
rect -6320 -20710 -6270 -20700
rect -6320 -20740 -6310 -20710
rect -6280 -20740 -6270 -20710
rect -6320 -20750 -6270 -20740
rect -6310 -20820 -6280 -20750
rect -6320 -20830 -6270 -20820
rect -6320 -20860 -6310 -20830
rect -6280 -20860 -6270 -20830
rect -6320 -20870 -6270 -20860
rect -6310 -20940 -6280 -20870
rect -6320 -20950 -6270 -20940
rect -6320 -20980 -6310 -20950
rect -6280 -20980 -6270 -20950
rect -6320 -20990 -6270 -20980
rect -6310 -21060 -6280 -20990
rect -6320 -21070 -6270 -21060
rect -6320 -21100 -6310 -21070
rect -6280 -21100 -6270 -21070
rect -6320 -21110 -6270 -21100
rect -6310 -21180 -6280 -21110
rect -6320 -21190 -6270 -21180
rect -6320 -21220 -6310 -21190
rect -6280 -21220 -6270 -21190
rect -6320 -21230 -6270 -21220
rect -6310 -21430 -6280 -21230
rect -6320 -21440 -6270 -21430
rect -6320 -21470 -6310 -21440
rect -6280 -21470 -6270 -21440
rect -6320 -21480 -6270 -21470
rect -6310 -21550 -6280 -21480
rect -6320 -21560 -6270 -21550
rect -6320 -21590 -6310 -21560
rect -6280 -21590 -6270 -21560
rect -6320 -21600 -6270 -21590
rect -6310 -21670 -6280 -21600
rect -6320 -21680 -6270 -21670
rect -6320 -21710 -6310 -21680
rect -6280 -21710 -6270 -21680
rect -6320 -21720 -6270 -21710
rect -6310 -21790 -6280 -21720
rect -6320 -21800 -6270 -21790
rect -6320 -21830 -6310 -21800
rect -6280 -21830 -6270 -21800
rect -6320 -21840 -6270 -21830
rect -6310 -21910 -6280 -21840
rect -6320 -21920 -6270 -21910
rect -6320 -21950 -6310 -21920
rect -6280 -21950 -6270 -21920
rect -6320 -21960 -6270 -21950
rect -6310 -22030 -6280 -21960
rect -6320 -22040 -6270 -22030
rect -6320 -22070 -6310 -22040
rect -6280 -22070 -6270 -22040
rect -6320 -22080 -6270 -22070
rect -6310 -22150 -6280 -22080
rect -6210 -22090 -6180 -16030
rect -6110 -17610 -6080 -15970
rect -6010 -16100 -5980 -9460
rect -5910 -9590 -5880 -7950
rect -5810 -9290 -5780 -3710
rect -5710 -5050 -5680 -3410
rect -5610 -3780 -5580 -190
rect -5510 -3360 -5480 -220
rect -5520 -3370 -5470 -3360
rect -5520 -3400 -5510 -3370
rect -5480 -3400 -5470 -3370
rect -5520 -3410 -5470 -3400
rect -5620 -3790 -5570 -3780
rect -5620 -3820 -5610 -3790
rect -5580 -3820 -5570 -3790
rect -5620 -3830 -5570 -3820
rect -5720 -5060 -5670 -5050
rect -5720 -5090 -5710 -5060
rect -5680 -5090 -5670 -5060
rect -5720 -5100 -5670 -5090
rect -5710 -7900 -5680 -5100
rect -5720 -7910 -5670 -7900
rect -5720 -7940 -5710 -7910
rect -5680 -7940 -5670 -7910
rect -5720 -7950 -5670 -7940
rect -5820 -9300 -5770 -9290
rect -5820 -9330 -5810 -9300
rect -5780 -9330 -5770 -9300
rect -5820 -9340 -5770 -9330
rect -5920 -9600 -5870 -9590
rect -5920 -9630 -5910 -9600
rect -5880 -9630 -5870 -9600
rect -5920 -9640 -5870 -9630
rect -5910 -15920 -5880 -9640
rect -5920 -15930 -5870 -15920
rect -5920 -15960 -5910 -15930
rect -5880 -15960 -5870 -15930
rect -5920 -15970 -5870 -15960
rect -6020 -16110 -5970 -16100
rect -6020 -16140 -6010 -16110
rect -5980 -16140 -5970 -16110
rect -6020 -16150 -5970 -16140
rect -6120 -17620 -6070 -17610
rect -6120 -17650 -6110 -17620
rect -6080 -17650 -6070 -17620
rect -6120 -17660 -6070 -17650
rect -6110 -20460 -6080 -17660
rect -6120 -20470 -6070 -20460
rect -6120 -20500 -6110 -20470
rect -6080 -20500 -6070 -20470
rect -6120 -20510 -6070 -20500
rect -6220 -22100 -6170 -22090
rect -6220 -22130 -6210 -22100
rect -6180 -22130 -6170 -22100
rect -6220 -22140 -6170 -22130
rect -6320 -22160 -6270 -22150
rect -6320 -22190 -6310 -22160
rect -6280 -22190 -6270 -22160
rect -6320 -22200 -6270 -22190
rect -6310 -28520 -6280 -22200
rect -6210 -28520 -6180 -22140
rect -6110 -22150 -6080 -20510
rect -6010 -21970 -5980 -16150
rect -5910 -17610 -5880 -15970
rect -5810 -16220 -5780 -9340
rect -5710 -9590 -5680 -7950
rect -5610 -9170 -5580 -3830
rect -5510 -5050 -5480 -3410
rect -5410 -3900 -5380 -190
rect -5310 -3360 -5280 -220
rect -5320 -3370 -5270 -3360
rect -5320 -3400 -5310 -3370
rect -5280 -3400 -5270 -3370
rect -5320 -3410 -5270 -3400
rect -5420 -3910 -5370 -3900
rect -5420 -3940 -5410 -3910
rect -5380 -3940 -5370 -3910
rect -5420 -3950 -5370 -3940
rect -5520 -5060 -5470 -5050
rect -5520 -5090 -5510 -5060
rect -5480 -5090 -5470 -5060
rect -5520 -5100 -5470 -5090
rect -5510 -7900 -5480 -5100
rect -5520 -7910 -5470 -7900
rect -5520 -7940 -5510 -7910
rect -5480 -7940 -5470 -7910
rect -5520 -7950 -5470 -7940
rect -5620 -9180 -5570 -9170
rect -5620 -9210 -5610 -9180
rect -5580 -9210 -5570 -9180
rect -5620 -9220 -5570 -9210
rect -5720 -9600 -5670 -9590
rect -5720 -9630 -5710 -9600
rect -5680 -9630 -5670 -9600
rect -5720 -9640 -5670 -9630
rect -5710 -15920 -5680 -9640
rect -5720 -15930 -5670 -15920
rect -5720 -15960 -5710 -15930
rect -5680 -15960 -5670 -15930
rect -5720 -15970 -5670 -15960
rect -5820 -16230 -5770 -16220
rect -5820 -16260 -5810 -16230
rect -5780 -16260 -5770 -16230
rect -5820 -16270 -5770 -16260
rect -5920 -17620 -5870 -17610
rect -5920 -17650 -5910 -17620
rect -5880 -17650 -5870 -17620
rect -5920 -17660 -5870 -17650
rect -5910 -20460 -5880 -17660
rect -5920 -20470 -5870 -20460
rect -5920 -20500 -5910 -20470
rect -5880 -20500 -5870 -20470
rect -5920 -20510 -5870 -20500
rect -6020 -21980 -5970 -21970
rect -6020 -22010 -6010 -21980
rect -5980 -22010 -5970 -21980
rect -6020 -22020 -5970 -22010
rect -6120 -22160 -6070 -22150
rect -6120 -22190 -6110 -22160
rect -6080 -22190 -6070 -22160
rect -6120 -22200 -6070 -22190
rect -6110 -28520 -6080 -22200
rect -6010 -28520 -5980 -22020
rect -5910 -22150 -5880 -20510
rect -5810 -21850 -5780 -16270
rect -5710 -17610 -5680 -15970
rect -5610 -16340 -5580 -9220
rect -5510 -9590 -5480 -7950
rect -5410 -9050 -5380 -3950
rect -5310 -5050 -5280 -3410
rect -5210 -4020 -5180 -190
rect -5110 -3360 -5080 -220
rect -5120 -3370 -5070 -3360
rect -5120 -3400 -5110 -3370
rect -5080 -3400 -5070 -3370
rect -5120 -3410 -5070 -3400
rect -5220 -4030 -5170 -4020
rect -5220 -4060 -5210 -4030
rect -5180 -4060 -5170 -4030
rect -5220 -4070 -5170 -4060
rect -5320 -5060 -5270 -5050
rect -5320 -5090 -5310 -5060
rect -5280 -5090 -5270 -5060
rect -5320 -5100 -5270 -5090
rect -5310 -7900 -5280 -5100
rect -5320 -7910 -5270 -7900
rect -5320 -7940 -5310 -7910
rect -5280 -7940 -5270 -7910
rect -5320 -7950 -5270 -7940
rect -5420 -9060 -5370 -9050
rect -5420 -9090 -5410 -9060
rect -5380 -9090 -5370 -9060
rect -5420 -9100 -5370 -9090
rect -5520 -9600 -5470 -9590
rect -5520 -9630 -5510 -9600
rect -5480 -9630 -5470 -9600
rect -5520 -9640 -5470 -9630
rect -5510 -15920 -5480 -9640
rect -5520 -15930 -5470 -15920
rect -5520 -15960 -5510 -15930
rect -5480 -15960 -5470 -15930
rect -5520 -15970 -5470 -15960
rect -5620 -16350 -5570 -16340
rect -5620 -16380 -5610 -16350
rect -5580 -16380 -5570 -16350
rect -5620 -16390 -5570 -16380
rect -5720 -17620 -5670 -17610
rect -5720 -17650 -5710 -17620
rect -5680 -17650 -5670 -17620
rect -5720 -17660 -5670 -17650
rect -5710 -20460 -5680 -17660
rect -5720 -20470 -5670 -20460
rect -5720 -20500 -5710 -20470
rect -5680 -20500 -5670 -20470
rect -5720 -20510 -5670 -20500
rect -5820 -21860 -5770 -21850
rect -5820 -21890 -5810 -21860
rect -5780 -21890 -5770 -21860
rect -5820 -21900 -5770 -21890
rect -5920 -22160 -5870 -22150
rect -5920 -22190 -5910 -22160
rect -5880 -22190 -5870 -22160
rect -5920 -22200 -5870 -22190
rect -5910 -28520 -5880 -22200
rect -5810 -28520 -5780 -21900
rect -5710 -22150 -5680 -20510
rect -5610 -21730 -5580 -16390
rect -5510 -17610 -5480 -15970
rect -5410 -16460 -5380 -9100
rect -5310 -9590 -5280 -7950
rect -5210 -8930 -5180 -4070
rect -5110 -5050 -5080 -3410
rect -5010 -4160 -4780 -190
rect -4710 -3360 -4680 -220
rect -4720 -3370 -4670 -3360
rect -4720 -3400 -4710 -3370
rect -4680 -3400 -4670 -3370
rect -4720 -3410 -4670 -3400
rect -5010 -4300 -5000 -4160
rect -4790 -4300 -4780 -4160
rect -5120 -5060 -5070 -5050
rect -5120 -5090 -5110 -5060
rect -5080 -5090 -5070 -5060
rect -5120 -5100 -5070 -5090
rect -5110 -7900 -5080 -5100
rect -5120 -7910 -5070 -7900
rect -5120 -7940 -5110 -7910
rect -5080 -7940 -5070 -7910
rect -5120 -7950 -5070 -7940
rect -5220 -8940 -5170 -8930
rect -5220 -8970 -5210 -8940
rect -5180 -8970 -5170 -8940
rect -5220 -8980 -5170 -8970
rect -5320 -9600 -5270 -9590
rect -5320 -9630 -5310 -9600
rect -5280 -9630 -5270 -9600
rect -5320 -9640 -5270 -9630
rect -5310 -15920 -5280 -9640
rect -5320 -15930 -5270 -15920
rect -5320 -15960 -5310 -15930
rect -5280 -15960 -5270 -15930
rect -5320 -15970 -5270 -15960
rect -5420 -16470 -5370 -16460
rect -5420 -16500 -5410 -16470
rect -5380 -16500 -5370 -16470
rect -5420 -16510 -5370 -16500
rect -5520 -17620 -5470 -17610
rect -5520 -17650 -5510 -17620
rect -5480 -17650 -5470 -17620
rect -5520 -17660 -5470 -17650
rect -5510 -20460 -5480 -17660
rect -5520 -20470 -5470 -20460
rect -5520 -20500 -5510 -20470
rect -5480 -20500 -5470 -20470
rect -5520 -20510 -5470 -20500
rect -5620 -21740 -5570 -21730
rect -5620 -21770 -5610 -21740
rect -5580 -21770 -5570 -21740
rect -5620 -21780 -5570 -21770
rect -5720 -22160 -5670 -22150
rect -5720 -22190 -5710 -22160
rect -5680 -22190 -5670 -22160
rect -5720 -22200 -5670 -22190
rect -5710 -28520 -5680 -22200
rect -5610 -28520 -5580 -21780
rect -5510 -22150 -5480 -20510
rect -5410 -21610 -5380 -16510
rect -5310 -17610 -5280 -15970
rect -5210 -16580 -5180 -8980
rect -5110 -9590 -5080 -7950
rect -5010 -8700 -4780 -4300
rect -4710 -5050 -4680 -3410
rect -4610 -4390 -4580 -190
rect -4510 -3360 -4480 -220
rect -4520 -3370 -4470 -3360
rect -4520 -3400 -4510 -3370
rect -4480 -3400 -4470 -3370
rect -4520 -3410 -4470 -3400
rect -4620 -4400 -4570 -4390
rect -4620 -4430 -4610 -4400
rect -4580 -4430 -4570 -4400
rect -4620 -4440 -4570 -4430
rect -4720 -5060 -4670 -5050
rect -4720 -5090 -4710 -5060
rect -4680 -5090 -4670 -5060
rect -4720 -5100 -4670 -5090
rect -4710 -7900 -4680 -5100
rect -4720 -7910 -4670 -7900
rect -4720 -7940 -4710 -7910
rect -4680 -7940 -4670 -7910
rect -4720 -7950 -4670 -7940
rect -5010 -8840 -5000 -8700
rect -4790 -8840 -4780 -8700
rect -5120 -9600 -5070 -9590
rect -5120 -9630 -5110 -9600
rect -5080 -9630 -5070 -9600
rect -5120 -9640 -5070 -9630
rect -5110 -15920 -5080 -9640
rect -5120 -15930 -5070 -15920
rect -5120 -15960 -5110 -15930
rect -5080 -15960 -5070 -15930
rect -5120 -15970 -5070 -15960
rect -5220 -16590 -5170 -16580
rect -5220 -16620 -5210 -16590
rect -5180 -16620 -5170 -16590
rect -5220 -16630 -5170 -16620
rect -5320 -17620 -5270 -17610
rect -5320 -17650 -5310 -17620
rect -5280 -17650 -5270 -17620
rect -5320 -17660 -5270 -17650
rect -5310 -20460 -5280 -17660
rect -5320 -20470 -5270 -20460
rect -5320 -20500 -5310 -20470
rect -5280 -20500 -5270 -20470
rect -5320 -20510 -5270 -20500
rect -5420 -21620 -5370 -21610
rect -5420 -21650 -5410 -21620
rect -5380 -21650 -5370 -21620
rect -5420 -21660 -5370 -21650
rect -5520 -22160 -5470 -22150
rect -5520 -22190 -5510 -22160
rect -5480 -22190 -5470 -22160
rect -5520 -22200 -5470 -22190
rect -5510 -28520 -5480 -22200
rect -5410 -28520 -5380 -21660
rect -5310 -22150 -5280 -20510
rect -5210 -21490 -5180 -16630
rect -5110 -17610 -5080 -15970
rect -5010 -16720 -4780 -8840
rect -4710 -9590 -4680 -7950
rect -4610 -8560 -4580 -4440
rect -4510 -5050 -4480 -3410
rect -4410 -4510 -4380 -190
rect -4310 -3360 -4280 -220
rect -4320 -3370 -4270 -3360
rect -4320 -3400 -4310 -3370
rect -4280 -3400 -4270 -3370
rect -4320 -3410 -4270 -3400
rect -4420 -4520 -4370 -4510
rect -4420 -4550 -4410 -4520
rect -4380 -4550 -4370 -4520
rect -4420 -4560 -4370 -4550
rect -4520 -5060 -4470 -5050
rect -4520 -5090 -4510 -5060
rect -4480 -5090 -4470 -5060
rect -4520 -5100 -4470 -5090
rect -4510 -7900 -4480 -5100
rect -4520 -7910 -4470 -7900
rect -4520 -7940 -4510 -7910
rect -4480 -7940 -4470 -7910
rect -4520 -7950 -4470 -7940
rect -4620 -8570 -4570 -8560
rect -4620 -8600 -4610 -8570
rect -4580 -8600 -4570 -8570
rect -4620 -8610 -4570 -8600
rect -4720 -9600 -4670 -9590
rect -4720 -9630 -4710 -9600
rect -4680 -9630 -4670 -9600
rect -4720 -9640 -4670 -9630
rect -4710 -15920 -4680 -9640
rect -4720 -15930 -4670 -15920
rect -4720 -15960 -4710 -15930
rect -4680 -15960 -4670 -15930
rect -4720 -15970 -4670 -15960
rect -5010 -16860 -5000 -16720
rect -4790 -16860 -4780 -16720
rect -5120 -17620 -5070 -17610
rect -5120 -17650 -5110 -17620
rect -5080 -17650 -5070 -17620
rect -5120 -17660 -5070 -17650
rect -5110 -20460 -5080 -17660
rect -5120 -20470 -5070 -20460
rect -5120 -20500 -5110 -20470
rect -5080 -20500 -5070 -20470
rect -5120 -20510 -5070 -20500
rect -5220 -21500 -5170 -21490
rect -5220 -21530 -5210 -21500
rect -5180 -21530 -5170 -21500
rect -5220 -21540 -5170 -21530
rect -5320 -22160 -5270 -22150
rect -5320 -22190 -5310 -22160
rect -5280 -22190 -5270 -22160
rect -5320 -22200 -5270 -22190
rect -5310 -28520 -5280 -22200
rect -5210 -28520 -5180 -21540
rect -5110 -22150 -5080 -20510
rect -5010 -21260 -4780 -16860
rect -4710 -17610 -4680 -15970
rect -4610 -16950 -4580 -8610
rect -4510 -9590 -4480 -7950
rect -4410 -8440 -4380 -4560
rect -4310 -5050 -4280 -3410
rect -4210 -4630 -4180 -190
rect -4110 -3360 -4080 -220
rect -4120 -3370 -4070 -3360
rect -4120 -3400 -4110 -3370
rect -4080 -3400 -4070 -3370
rect -4120 -3410 -4070 -3400
rect -4220 -4640 -4170 -4630
rect -4220 -4670 -4210 -4640
rect -4180 -4670 -4170 -4640
rect -4220 -4680 -4170 -4670
rect -4320 -5060 -4270 -5050
rect -4320 -5090 -4310 -5060
rect -4280 -5090 -4270 -5060
rect -4320 -5100 -4270 -5090
rect -4310 -7900 -4280 -5100
rect -4320 -7910 -4270 -7900
rect -4320 -7940 -4310 -7910
rect -4280 -7940 -4270 -7910
rect -4320 -7950 -4270 -7940
rect -4420 -8450 -4370 -8440
rect -4420 -8480 -4410 -8450
rect -4380 -8480 -4370 -8450
rect -4420 -8490 -4370 -8480
rect -4520 -9600 -4470 -9590
rect -4520 -9630 -4510 -9600
rect -4480 -9630 -4470 -9600
rect -4520 -9640 -4470 -9630
rect -4510 -15920 -4480 -9640
rect -4520 -15930 -4470 -15920
rect -4520 -15960 -4510 -15930
rect -4480 -15960 -4470 -15930
rect -4520 -15970 -4470 -15960
rect -4620 -16960 -4570 -16950
rect -4620 -16990 -4610 -16960
rect -4580 -16990 -4570 -16960
rect -4620 -17000 -4570 -16990
rect -4720 -17620 -4670 -17610
rect -4720 -17650 -4710 -17620
rect -4680 -17650 -4670 -17620
rect -4720 -17660 -4670 -17650
rect -4710 -20460 -4680 -17660
rect -4720 -20470 -4670 -20460
rect -4720 -20500 -4710 -20470
rect -4680 -20500 -4670 -20470
rect -4720 -20510 -4670 -20500
rect -5010 -21400 -5000 -21260
rect -4790 -21400 -4780 -21260
rect -5120 -22160 -5070 -22150
rect -5120 -22190 -5110 -22160
rect -5080 -22190 -5070 -22160
rect -5120 -22200 -5070 -22190
rect -5110 -28520 -5080 -22200
rect -5010 -26910 -4780 -21400
rect -4710 -22150 -4680 -20510
rect -4610 -21120 -4580 -17000
rect -4510 -17610 -4480 -15970
rect -4410 -17070 -4380 -8490
rect -4310 -9590 -4280 -7950
rect -4210 -8320 -4180 -4680
rect -4110 -5050 -4080 -3410
rect -4010 -4750 -3980 -190
rect -3910 -3360 -3880 -220
rect -3920 -3370 -3870 -3360
rect -3920 -3400 -3910 -3370
rect -3880 -3400 -3870 -3370
rect -3920 -3410 -3870 -3400
rect -4020 -4760 -3970 -4750
rect -4020 -4790 -4010 -4760
rect -3980 -4790 -3970 -4760
rect -4020 -4800 -3970 -4790
rect -4120 -5060 -4070 -5050
rect -4120 -5090 -4110 -5060
rect -4080 -5090 -4070 -5060
rect -4120 -5100 -4070 -5090
rect -4110 -7900 -4080 -5100
rect -4120 -7910 -4070 -7900
rect -4120 -7940 -4110 -7910
rect -4080 -7940 -4070 -7910
rect -4120 -7950 -4070 -7940
rect -4220 -8330 -4170 -8320
rect -4220 -8360 -4210 -8330
rect -4180 -8360 -4170 -8330
rect -4220 -8370 -4170 -8360
rect -4320 -9600 -4270 -9590
rect -4320 -9630 -4310 -9600
rect -4280 -9630 -4270 -9600
rect -4320 -9640 -4270 -9630
rect -4310 -15920 -4280 -9640
rect -4320 -15930 -4270 -15920
rect -4320 -15960 -4310 -15930
rect -4280 -15960 -4270 -15930
rect -4320 -15970 -4270 -15960
rect -4420 -17080 -4370 -17070
rect -4420 -17110 -4410 -17080
rect -4380 -17110 -4370 -17080
rect -4420 -17120 -4370 -17110
rect -4520 -17620 -4470 -17610
rect -4520 -17650 -4510 -17620
rect -4480 -17650 -4470 -17620
rect -4520 -17660 -4470 -17650
rect -4510 -20460 -4480 -17660
rect -4520 -20470 -4470 -20460
rect -4520 -20500 -4510 -20470
rect -4480 -20500 -4470 -20470
rect -4520 -20510 -4470 -20500
rect -4620 -21130 -4570 -21120
rect -4620 -21160 -4610 -21130
rect -4580 -21160 -4570 -21130
rect -4620 -21170 -4570 -21160
rect -4720 -22160 -4670 -22150
rect -4720 -22190 -4710 -22160
rect -4680 -22190 -4670 -22160
rect -4720 -22200 -4670 -22190
rect -5010 -27050 -5000 -26910
rect -4790 -27050 -4780 -26910
rect -5010 -28520 -4780 -27050
rect -4710 -28520 -4680 -22200
rect -4610 -28520 -4580 -21170
rect -4510 -22150 -4480 -20510
rect -4410 -21000 -4380 -17120
rect -4310 -17610 -4280 -15970
rect -4210 -17190 -4180 -8370
rect -4110 -9590 -4080 -7950
rect -4010 -8200 -3980 -4800
rect -3910 -5050 -3880 -3410
rect -3810 -4870 -3780 -190
rect -3710 -3360 -3680 -220
rect -3720 -3370 -3670 -3360
rect -3720 -3400 -3710 -3370
rect -3680 -3400 -3670 -3370
rect -3720 -3410 -3670 -3400
rect -3820 -4880 -3770 -4870
rect -3820 -4910 -3810 -4880
rect -3780 -4910 -3770 -4880
rect -3820 -4920 -3770 -4910
rect -3920 -5060 -3870 -5050
rect -3920 -5090 -3910 -5060
rect -3880 -5090 -3870 -5060
rect -3920 -5100 -3870 -5090
rect -3910 -7900 -3880 -5100
rect -3920 -7910 -3870 -7900
rect -3920 -7940 -3910 -7910
rect -3880 -7940 -3870 -7910
rect -3920 -7950 -3870 -7940
rect -4020 -8210 -3970 -8200
rect -4020 -8240 -4010 -8210
rect -3980 -8240 -3970 -8210
rect -4020 -8250 -3970 -8240
rect -4120 -9600 -4070 -9590
rect -4120 -9630 -4110 -9600
rect -4080 -9630 -4070 -9600
rect -4120 -9640 -4070 -9630
rect -4110 -15920 -4080 -9640
rect -4120 -15930 -4070 -15920
rect -4120 -15960 -4110 -15930
rect -4080 -15960 -4070 -15930
rect -4120 -15970 -4070 -15960
rect -4220 -17200 -4170 -17190
rect -4220 -17230 -4210 -17200
rect -4180 -17230 -4170 -17200
rect -4220 -17240 -4170 -17230
rect -4320 -17620 -4270 -17610
rect -4320 -17650 -4310 -17620
rect -4280 -17650 -4270 -17620
rect -4320 -17660 -4270 -17650
rect -4310 -20460 -4280 -17660
rect -4320 -20470 -4270 -20460
rect -4320 -20500 -4310 -20470
rect -4280 -20500 -4270 -20470
rect -4320 -20510 -4270 -20500
rect -4420 -21010 -4370 -21000
rect -4420 -21040 -4410 -21010
rect -4380 -21040 -4370 -21010
rect -4420 -21050 -4370 -21040
rect -4520 -22160 -4470 -22150
rect -4520 -22190 -4510 -22160
rect -4480 -22190 -4470 -22160
rect -4520 -22200 -4470 -22190
rect -4510 -28520 -4480 -22200
rect -4410 -28520 -4380 -21050
rect -4310 -22150 -4280 -20510
rect -4210 -20880 -4180 -17240
rect -4110 -17610 -4080 -15970
rect -4010 -17310 -3980 -8250
rect -3910 -9590 -3880 -7950
rect -3810 -8080 -3780 -4920
rect -3710 -5050 -3680 -3410
rect -3610 -4990 -3580 -190
rect -3510 -3360 -3480 -220
rect -3420 -230 -3260 -220
rect -3420 -370 -3410 -230
rect -3270 -370 -3260 -230
rect -3520 -3370 -3470 -3360
rect -3520 -3400 -3510 -3370
rect -3480 -3400 -3470 -3370
rect -3520 -3410 -3470 -3400
rect -3620 -5000 -3570 -4990
rect -3620 -5030 -3610 -5000
rect -3580 -5030 -3570 -5000
rect -3620 -5040 -3570 -5030
rect -3720 -5060 -3670 -5050
rect -3720 -5090 -3710 -5060
rect -3680 -5090 -3670 -5060
rect -3720 -5100 -3670 -5090
rect -3710 -7900 -3680 -5100
rect -3720 -7910 -3670 -7900
rect -3720 -7940 -3710 -7910
rect -3680 -7940 -3670 -7910
rect -3720 -7950 -3670 -7940
rect -3820 -8090 -3770 -8080
rect -3820 -8120 -3810 -8090
rect -3780 -8120 -3770 -8090
rect -3820 -8130 -3770 -8120
rect -3920 -9600 -3870 -9590
rect -3920 -9630 -3910 -9600
rect -3880 -9630 -3870 -9600
rect -3920 -9640 -3870 -9630
rect -3910 -15920 -3880 -9640
rect -3920 -15930 -3870 -15920
rect -3920 -15960 -3910 -15930
rect -3880 -15960 -3870 -15930
rect -3920 -15970 -3870 -15960
rect -4020 -17320 -3970 -17310
rect -4020 -17350 -4010 -17320
rect -3980 -17350 -3970 -17320
rect -4020 -17360 -3970 -17350
rect -4120 -17620 -4070 -17610
rect -4120 -17650 -4110 -17620
rect -4080 -17650 -4070 -17620
rect -4120 -17660 -4070 -17650
rect -4110 -20460 -4080 -17660
rect -4120 -20470 -4070 -20460
rect -4120 -20500 -4110 -20470
rect -4080 -20500 -4070 -20470
rect -4120 -20510 -4070 -20500
rect -4220 -20890 -4170 -20880
rect -4220 -20920 -4210 -20890
rect -4180 -20920 -4170 -20890
rect -4220 -20930 -4170 -20920
rect -4320 -22160 -4270 -22150
rect -4320 -22190 -4310 -22160
rect -4280 -22190 -4270 -22160
rect -4320 -22200 -4270 -22190
rect -4310 -28520 -4280 -22200
rect -4210 -26700 -4180 -20930
rect -4110 -22150 -4080 -20510
rect -4010 -20760 -3980 -17360
rect -3910 -17610 -3880 -15970
rect -3810 -17430 -3780 -8130
rect -3710 -9590 -3680 -7950
rect -3610 -7960 -3580 -5040
rect -3510 -5050 -3480 -3410
rect -3520 -5060 -3470 -5050
rect -3520 -5090 -3510 -5060
rect -3480 -5090 -3470 -5060
rect -3520 -5100 -3470 -5090
rect -3510 -7900 -3480 -5100
rect -3520 -7910 -3470 -7900
rect -3520 -7940 -3510 -7910
rect -3480 -7940 -3470 -7910
rect -3520 -7950 -3470 -7940
rect -3620 -7970 -3570 -7960
rect -3620 -8000 -3610 -7970
rect -3580 -8000 -3570 -7970
rect -3620 -8010 -3570 -8000
rect -3720 -9600 -3670 -9590
rect -3720 -9630 -3710 -9600
rect -3680 -9630 -3670 -9600
rect -3720 -9640 -3670 -9630
rect -3710 -15920 -3680 -9640
rect -3720 -15930 -3670 -15920
rect -3720 -15960 -3710 -15930
rect -3680 -15960 -3670 -15930
rect -3720 -15970 -3670 -15960
rect -3820 -17440 -3770 -17430
rect -3820 -17470 -3810 -17440
rect -3780 -17470 -3770 -17440
rect -3820 -17480 -3770 -17470
rect -3920 -17620 -3870 -17610
rect -3920 -17650 -3910 -17620
rect -3880 -17650 -3870 -17620
rect -3920 -17660 -3870 -17650
rect -3910 -20460 -3880 -17660
rect -3920 -20470 -3870 -20460
rect -3920 -20500 -3910 -20470
rect -3880 -20500 -3870 -20470
rect -3920 -20510 -3870 -20500
rect -4020 -20770 -3970 -20760
rect -4020 -20800 -4010 -20770
rect -3980 -20800 -3970 -20770
rect -4020 -20810 -3970 -20800
rect -4120 -22160 -4070 -22150
rect -4120 -22190 -4110 -22160
rect -4080 -22190 -4070 -22160
rect -4120 -22200 -4070 -22190
rect -4230 -26710 -4160 -26700
rect -4230 -26850 -4220 -26710
rect -4170 -26850 -4160 -26710
rect -4230 -26860 -4160 -26850
rect -4210 -28520 -4180 -26860
rect -4110 -28520 -4080 -22200
rect -4010 -27100 -3980 -20810
rect -3910 -22150 -3880 -20510
rect -3810 -20640 -3780 -17480
rect -3710 -17610 -3680 -15970
rect -3610 -17550 -3580 -8010
rect -3510 -9590 -3480 -7950
rect -3520 -9600 -3470 -9590
rect -3520 -9630 -3510 -9600
rect -3480 -9630 -3470 -9600
rect -3520 -9640 -3470 -9630
rect -3510 -15920 -3480 -9640
rect -3420 -12630 -3260 -370
rect -3420 -12770 -3410 -12630
rect -3270 -12770 -3260 -12630
rect -3420 -12790 -3260 -12770
rect -3420 -12930 -3410 -12790
rect -3270 -12930 -3260 -12790
rect -3520 -15930 -3470 -15920
rect -3520 -15960 -3510 -15930
rect -3480 -15960 -3470 -15930
rect -3520 -15970 -3470 -15960
rect -3620 -17560 -3570 -17550
rect -3620 -17590 -3610 -17560
rect -3580 -17590 -3570 -17560
rect -3620 -17600 -3570 -17590
rect -3720 -17620 -3670 -17610
rect -3720 -17650 -3710 -17620
rect -3680 -17650 -3670 -17620
rect -3720 -17660 -3670 -17650
rect -3710 -20460 -3680 -17660
rect -3720 -20470 -3670 -20460
rect -3720 -20500 -3710 -20470
rect -3680 -20500 -3670 -20470
rect -3720 -20510 -3670 -20500
rect -3820 -20650 -3770 -20640
rect -3820 -20680 -3810 -20650
rect -3780 -20680 -3770 -20650
rect -3820 -20690 -3770 -20680
rect -3920 -22160 -3870 -22150
rect -3920 -22190 -3910 -22160
rect -3880 -22190 -3870 -22160
rect -3920 -22200 -3870 -22190
rect -4030 -27110 -3960 -27100
rect -4030 -27250 -4020 -27110
rect -3970 -27250 -3960 -27110
rect -4030 -27260 -3960 -27250
rect -4010 -28520 -3980 -27260
rect -3910 -28520 -3880 -22200
rect -3810 -28520 -3780 -20690
rect -3710 -22150 -3680 -20510
rect -3610 -20520 -3580 -17600
rect -3510 -17610 -3480 -15970
rect -3520 -17620 -3470 -17610
rect -3520 -17650 -3510 -17620
rect -3480 -17650 -3470 -17620
rect -3520 -17660 -3470 -17650
rect -3510 -20460 -3480 -17660
rect -3520 -20470 -3470 -20460
rect -3520 -20500 -3510 -20470
rect -3480 -20500 -3470 -20470
rect -3520 -20510 -3470 -20500
rect -3620 -20530 -3570 -20520
rect -3620 -20560 -3610 -20530
rect -3580 -20560 -3570 -20530
rect -3620 -20570 -3570 -20560
rect -3720 -22160 -3670 -22150
rect -3720 -22190 -3710 -22160
rect -3680 -22190 -3670 -22160
rect -3720 -22200 -3670 -22190
rect -3710 -28520 -3680 -22200
rect -3610 -28520 -3580 -20570
rect -3510 -22150 -3480 -20510
rect -3520 -22160 -3470 -22150
rect -3520 -22190 -3510 -22160
rect -3480 -22190 -3470 -22160
rect -3520 -22200 -3470 -22190
rect -3510 -28300 -3480 -22200
rect -3420 -25190 -3260 -12930
rect -3420 -25330 -3410 -25190
rect -3270 -25330 -3260 -25190
rect -3420 -25340 -3260 -25330
rect -3100 -6350 -2940 -220
rect -3100 -6490 -3090 -6350
rect -2950 -6490 -2940 -6350
rect -3100 -6510 -2940 -6490
rect -3100 -6650 -3090 -6510
rect -2950 -6650 -2940 -6510
rect -3100 -18910 -2940 -6650
rect -3100 -19050 -3090 -18910
rect -2950 -19050 -2940 -18910
rect -3100 -19070 -2940 -19050
rect -3100 -19210 -3090 -19070
rect -2950 -19210 -2940 -19070
rect -3100 -25340 -2940 -19210
rect 23620 -6350 23780 -190
rect 23620 -6490 23630 -6350
rect 23770 -6490 23780 -6350
rect 23620 -6510 23780 -6490
rect 23620 -6650 23630 -6510
rect 23770 -6650 23780 -6510
rect 23620 -18910 23780 -6650
rect 23620 -19050 23630 -18910
rect 23770 -19050 23780 -18910
rect 23620 -19070 23780 -19050
rect 23620 -19210 23630 -19070
rect 23770 -19210 23780 -19070
rect 23620 -25340 23780 -19210
rect 23940 -230 24100 -190
rect 23940 -370 23950 -230
rect 24090 -370 24100 -230
rect 23940 -12630 24100 -370
rect 23940 -12770 23950 -12630
rect 24090 -12770 24100 -12630
rect 23940 -12790 24100 -12770
rect 23940 -12930 23950 -12790
rect 24090 -12930 24100 -12790
rect 23940 -25190 24100 -12930
rect 23940 -25330 23950 -25190
rect 24090 -25330 24100 -25190
rect 23940 -25340 24100 -25330
rect 24260 -3440 24420 -190
rect 24260 -3570 24270 -3440
rect 24410 -3570 24420 -3440
rect 24260 -3680 24420 -3570
rect 24260 -3810 24270 -3680
rect 24410 -3810 24420 -3680
rect 24260 -3920 24420 -3810
rect 24260 -4050 24270 -3920
rect 24410 -4050 24420 -3920
rect 24260 -4160 24420 -4050
rect 24260 -4300 24270 -4160
rect 24410 -4300 24420 -4160
rect 24260 -4410 24420 -4300
rect 24260 -4540 24270 -4410
rect 24410 -4540 24420 -4410
rect 24260 -4650 24420 -4540
rect 24260 -4780 24270 -4650
rect 24410 -4780 24420 -4650
rect 24260 -4890 24420 -4780
rect 24260 -5020 24270 -4890
rect 24410 -5020 24420 -4890
rect 24260 -7980 24420 -5020
rect 24260 -8110 24270 -7980
rect 24410 -8110 24420 -7980
rect 24260 -8220 24420 -8110
rect 24260 -8350 24270 -8220
rect 24410 -8350 24420 -8220
rect 24260 -8460 24420 -8350
rect 24260 -8590 24270 -8460
rect 24410 -8590 24420 -8460
rect 24260 -8700 24420 -8590
rect 24260 -8840 24270 -8700
rect 24410 -8840 24420 -8700
rect 24260 -8950 24420 -8840
rect 24260 -9080 24270 -8950
rect 24410 -9080 24420 -8950
rect 24260 -9190 24420 -9080
rect 24260 -9320 24270 -9190
rect 24410 -9320 24420 -9190
rect 24260 -9430 24420 -9320
rect 24260 -9560 24270 -9430
rect 24410 -9560 24420 -9430
rect 24260 -16000 24420 -9560
rect 24260 -16130 24270 -16000
rect 24410 -16130 24420 -16000
rect 24260 -16240 24420 -16130
rect 24260 -16370 24270 -16240
rect 24410 -16370 24420 -16240
rect 24260 -16480 24420 -16370
rect 24260 -16610 24270 -16480
rect 24410 -16610 24420 -16480
rect 24260 -16720 24420 -16610
rect 24260 -16860 24270 -16720
rect 24410 -16860 24420 -16720
rect 24260 -16970 24420 -16860
rect 24260 -17100 24270 -16970
rect 24410 -17100 24420 -16970
rect 24260 -17210 24420 -17100
rect 24260 -17340 24270 -17210
rect 24410 -17340 24420 -17210
rect 24260 -17450 24420 -17340
rect 24260 -17580 24270 -17450
rect 24410 -17580 24420 -17450
rect 24260 -20540 24420 -17580
rect 24260 -20670 24270 -20540
rect 24410 -20670 24420 -20540
rect 24260 -20780 24420 -20670
rect 24260 -20910 24270 -20780
rect 24410 -20910 24420 -20780
rect 24260 -21020 24420 -20910
rect 24260 -21150 24270 -21020
rect 24410 -21150 24420 -21020
rect 24260 -21260 24420 -21150
rect 24260 -21400 24270 -21260
rect 24410 -21400 24420 -21260
rect 24260 -21510 24420 -21400
rect 24260 -21640 24270 -21510
rect 24410 -21640 24420 -21510
rect 24260 -21750 24420 -21640
rect 24260 -21880 24270 -21750
rect 24410 -21880 24420 -21750
rect 24260 -21990 24420 -21880
rect 24260 -22120 24270 -21990
rect 24410 -22120 24420 -21990
rect 24260 -25510 24420 -22120
rect 24260 -25650 24270 -25510
rect 24410 -25650 24420 -25510
rect -2380 -26900 -1340 -25820
rect -1290 -26900 -250 -25820
rect -200 -26900 840 -25820
rect 890 -26900 1930 -25820
rect 1980 -26900 3020 -25820
rect 3070 -26900 4110 -25820
rect 4160 -26900 5200 -25820
rect 5250 -26900 6290 -25820
rect 6340 -26900 7380 -25820
rect 7430 -26900 8470 -25820
rect 8520 -26900 9560 -25820
rect 9610 -26900 10650 -25820
rect 10700 -26900 11740 -25820
rect 11790 -26900 12830 -25820
rect 12880 -26900 13920 -25820
rect 13970 -26900 15010 -25820
rect 15060 -26900 16100 -25820
rect 16150 -26900 17190 -25820
rect 17240 -26900 18280 -25820
rect 18330 -26900 19370 -25820
rect 19420 -26900 20460 -25820
rect 20510 -26900 21550 -25820
rect 21600 -26900 22640 -25820
rect 22690 -26900 23730 -25820
rect -2380 -26920 23730 -26900
rect -2380 -27040 -2360 -26920
rect -1360 -27040 -1270 -26920
rect -270 -27040 -180 -26920
rect 820 -27040 910 -26920
rect 1910 -27040 2000 -26920
rect 3000 -27040 3090 -26920
rect 4090 -27040 4180 -26920
rect 5180 -27040 5270 -26920
rect 6270 -27040 6360 -26920
rect 7360 -27040 7450 -26920
rect 8450 -27040 8540 -26920
rect 9540 -27040 9630 -26920
rect 10630 -27040 10720 -26920
rect 11720 -27040 11810 -26920
rect 12810 -27040 12900 -26920
rect 13900 -27040 13990 -26920
rect 14990 -27040 15080 -26920
rect 16080 -27040 16170 -26920
rect 17170 -27040 17260 -26920
rect 18260 -27040 18350 -26920
rect 19350 -27040 19440 -26920
rect 20440 -27040 20530 -26920
rect 21530 -27040 21620 -26920
rect 22620 -27040 22710 -26920
rect 23710 -27040 23730 -26920
rect -2380 -27060 23730 -27040
rect -2380 -28140 -1340 -27060
rect -1290 -28140 -250 -27060
rect -200 -28140 840 -27060
rect 890 -28140 1930 -27060
rect 1980 -28140 3020 -27060
rect 3070 -28140 4110 -27060
rect 4160 -28140 5200 -27060
rect 5250 -28140 6290 -27060
rect 6340 -28140 7380 -27060
rect 7430 -28140 8470 -27060
rect 8520 -28140 9560 -27060
rect 9610 -28140 10650 -27060
rect 10700 -28140 11740 -27060
rect 11790 -28140 12830 -27060
rect 12880 -28140 13920 -27060
rect 13970 -28140 15010 -27060
rect 15060 -28140 16100 -27060
rect 16150 -28140 17190 -27060
rect 17240 -28140 18280 -27060
rect 18330 -28140 19370 -27060
rect 19420 -28140 20460 -27060
rect 20510 -28140 21550 -27060
rect 21600 -28140 22640 -27060
rect 22690 -28140 23730 -27060
rect -3530 -28310 -3460 -28300
rect -3530 -28450 -3520 -28310
rect -3470 -28450 -3460 -28310
rect -3530 -28460 -3460 -28450
rect 24260 -28310 24420 -25650
rect 24260 -28450 24270 -28310
rect 24410 -28450 24420 -28310
rect 24260 -28460 24420 -28450
rect -3510 -28520 -3480 -28460
<< via3 >>
rect -5000 -27050 -4790 -26910
rect -4220 -26850 -4170 -26710
rect -4020 -27250 -3970 -27110
rect 24270 -3570 24410 -3440
rect 24270 -3810 24410 -3680
rect 24270 -4050 24410 -3920
rect 24270 -4300 24410 -4160
rect 24270 -4540 24410 -4410
rect 24270 -4780 24410 -4650
rect 24270 -5020 24410 -4890
rect 24270 -8110 24410 -7980
rect 24270 -8350 24410 -8220
rect 24270 -8590 24410 -8460
rect 24270 -8840 24410 -8700
rect 24270 -9080 24410 -8950
rect 24270 -9320 24410 -9190
rect 24270 -9560 24410 -9430
rect 24270 -16130 24410 -16000
rect 24270 -16370 24410 -16240
rect 24270 -16610 24410 -16480
rect 24270 -16860 24410 -16720
rect 24270 -17100 24410 -16970
rect 24270 -17340 24410 -17210
rect 24270 -17580 24410 -17450
rect 24270 -20670 24410 -20540
rect 24270 -20910 24410 -20780
rect 24270 -21150 24410 -21020
rect 24270 -21400 24410 -21260
rect 24270 -21640 24410 -21510
rect 24270 -21880 24410 -21750
rect 24270 -22120 24410 -21990
rect 24270 -25650 24410 -25510
rect -2360 -27040 -1360 -26920
rect -1270 -27040 -270 -26920
rect -180 -27040 820 -26920
rect 910 -27040 1910 -26920
rect 2000 -27040 3000 -26920
rect 3090 -27040 4090 -26920
rect 4180 -27040 5180 -26920
rect 5270 -27040 6270 -26920
rect 6360 -27040 7360 -26920
rect 7450 -27040 8450 -26920
rect 8540 -27040 9540 -26920
rect 9630 -27040 10630 -26920
rect 10720 -27040 11720 -26920
rect 11810 -27040 12810 -26920
rect 12900 -27040 13900 -26920
rect 13990 -27040 14990 -26920
rect 15080 -27040 16080 -26920
rect 16170 -27040 17170 -26920
rect 17260 -27040 18260 -26920
rect 18350 -27040 19350 -26920
rect 19440 -27040 20440 -26920
rect 20530 -27040 21530 -26920
rect 21620 -27040 22620 -26920
rect 22710 -27040 23710 -26920
rect -3520 -28450 -3470 -28310
rect 24270 -28450 24410 -28310
<< mimcap >>
rect -2360 -25850 -1360 -25840
rect -2360 -26830 -2350 -25850
rect -1370 -26830 -1360 -25850
rect -2360 -26840 -1360 -26830
rect -1270 -25850 -270 -25840
rect -1270 -26830 -1260 -25850
rect -280 -26830 -270 -25850
rect -1270 -26840 -270 -26830
rect -180 -25850 820 -25840
rect -180 -26830 -170 -25850
rect 810 -26830 820 -25850
rect -180 -26840 820 -26830
rect 910 -25850 1910 -25840
rect 910 -26830 920 -25850
rect 1900 -26830 1910 -25850
rect 910 -26840 1910 -26830
rect 2000 -25850 3000 -25840
rect 2000 -26830 2010 -25850
rect 2990 -26830 3000 -25850
rect 2000 -26840 3000 -26830
rect 3090 -25850 4090 -25840
rect 3090 -26830 3100 -25850
rect 4080 -26830 4090 -25850
rect 3090 -26840 4090 -26830
rect 4180 -25850 5180 -25840
rect 4180 -26830 4190 -25850
rect 5170 -26830 5180 -25850
rect 4180 -26840 5180 -26830
rect 5270 -25850 6270 -25840
rect 5270 -26830 5280 -25850
rect 6260 -26830 6270 -25850
rect 5270 -26840 6270 -26830
rect 6360 -25850 7360 -25840
rect 6360 -26830 6370 -25850
rect 7350 -26830 7360 -25850
rect 6360 -26840 7360 -26830
rect 7450 -25850 8450 -25840
rect 7450 -26830 7460 -25850
rect 8440 -26830 8450 -25850
rect 7450 -26840 8450 -26830
rect 8540 -25850 9540 -25840
rect 8540 -26830 8550 -25850
rect 9530 -26830 9540 -25850
rect 8540 -26840 9540 -26830
rect 9630 -25850 10630 -25840
rect 9630 -26830 9640 -25850
rect 10620 -26830 10630 -25850
rect 9630 -26840 10630 -26830
rect 10720 -25850 11720 -25840
rect 10720 -26830 10730 -25850
rect 11710 -26830 11720 -25850
rect 10720 -26840 11720 -26830
rect 11810 -25850 12810 -25840
rect 11810 -26830 11820 -25850
rect 12800 -26830 12810 -25850
rect 11810 -26840 12810 -26830
rect 12900 -25850 13900 -25840
rect 12900 -26830 12910 -25850
rect 13890 -26830 13900 -25850
rect 12900 -26840 13900 -26830
rect 13990 -25850 14990 -25840
rect 13990 -26830 14000 -25850
rect 14980 -26830 14990 -25850
rect 13990 -26840 14990 -26830
rect 15080 -25850 16080 -25840
rect 15080 -26830 15090 -25850
rect 16070 -26830 16080 -25850
rect 15080 -26840 16080 -26830
rect 16170 -25850 17170 -25840
rect 16170 -26830 16180 -25850
rect 17160 -26830 17170 -25850
rect 16170 -26840 17170 -26830
rect 17260 -25850 18260 -25840
rect 17260 -26830 17270 -25850
rect 18250 -26830 18260 -25850
rect 17260 -26840 18260 -26830
rect 18350 -25850 19350 -25840
rect 18350 -26830 18360 -25850
rect 19340 -26830 19350 -25850
rect 18350 -26840 19350 -26830
rect 19440 -25850 20440 -25840
rect 19440 -26830 19450 -25850
rect 20430 -26830 20440 -25850
rect 19440 -26840 20440 -26830
rect 20530 -25850 21530 -25840
rect 20530 -26830 20540 -25850
rect 21520 -26830 21530 -25850
rect 20530 -26840 21530 -26830
rect 21620 -25850 22620 -25840
rect 21620 -26830 21630 -25850
rect 22610 -26830 22620 -25850
rect 21620 -26840 22620 -26830
rect 22710 -25850 23710 -25840
rect 22710 -26830 22720 -25850
rect 23700 -26830 23710 -25850
rect 22710 -26840 23710 -26830
rect -2360 -27130 -1360 -27120
rect -2360 -28110 -2350 -27130
rect -1370 -28110 -1360 -27130
rect -2360 -28120 -1360 -28110
rect -1270 -27130 -270 -27120
rect -1270 -28110 -1260 -27130
rect -280 -28110 -270 -27130
rect -1270 -28120 -270 -28110
rect -180 -27130 820 -27120
rect -180 -28110 -170 -27130
rect 810 -28110 820 -27130
rect -180 -28120 820 -28110
rect 910 -27130 1910 -27120
rect 910 -28110 920 -27130
rect 1900 -28110 1910 -27130
rect 910 -28120 1910 -28110
rect 2000 -27130 3000 -27120
rect 2000 -28110 2010 -27130
rect 2990 -28110 3000 -27130
rect 2000 -28120 3000 -28110
rect 3090 -27130 4090 -27120
rect 3090 -28110 3100 -27130
rect 4080 -28110 4090 -27130
rect 3090 -28120 4090 -28110
rect 4180 -27130 5180 -27120
rect 4180 -28110 4190 -27130
rect 5170 -28110 5180 -27130
rect 4180 -28120 5180 -28110
rect 5270 -27130 6270 -27120
rect 5270 -28110 5280 -27130
rect 6260 -28110 6270 -27130
rect 5270 -28120 6270 -28110
rect 6360 -27130 7360 -27120
rect 6360 -28110 6370 -27130
rect 7350 -28110 7360 -27130
rect 6360 -28120 7360 -28110
rect 7450 -27130 8450 -27120
rect 7450 -28110 7460 -27130
rect 8440 -28110 8450 -27130
rect 7450 -28120 8450 -28110
rect 8540 -27130 9540 -27120
rect 8540 -28110 8550 -27130
rect 9530 -28110 9540 -27130
rect 8540 -28120 9540 -28110
rect 9630 -27130 10630 -27120
rect 9630 -28110 9640 -27130
rect 10620 -28110 10630 -27130
rect 9630 -28120 10630 -28110
rect 10720 -27130 11720 -27120
rect 10720 -28110 10730 -27130
rect 11710 -28110 11720 -27130
rect 10720 -28120 11720 -28110
rect 11810 -27130 12810 -27120
rect 11810 -28110 11820 -27130
rect 12800 -28110 12810 -27130
rect 11810 -28120 12810 -28110
rect 12900 -27130 13900 -27120
rect 12900 -28110 12910 -27130
rect 13890 -28110 13900 -27130
rect 12900 -28120 13900 -28110
rect 13990 -27130 14990 -27120
rect 13990 -28110 14000 -27130
rect 14980 -28110 14990 -27130
rect 13990 -28120 14990 -28110
rect 15080 -27130 16080 -27120
rect 15080 -28110 15090 -27130
rect 16070 -28110 16080 -27130
rect 15080 -28120 16080 -28110
rect 16170 -27130 17170 -27120
rect 16170 -28110 16180 -27130
rect 17160 -28110 17170 -27130
rect 16170 -28120 17170 -28110
rect 17260 -27130 18260 -27120
rect 17260 -28110 17270 -27130
rect 18250 -28110 18260 -27130
rect 17260 -28120 18260 -28110
rect 18350 -27130 19350 -27120
rect 18350 -28110 18360 -27130
rect 19340 -28110 19350 -27130
rect 18350 -28120 19350 -28110
rect 19440 -27130 20440 -27120
rect 19440 -28110 19450 -27130
rect 20430 -28110 20440 -27130
rect 19440 -28120 20440 -28110
rect 20530 -27130 21530 -27120
rect 20530 -28110 20540 -27130
rect 21520 -28110 21530 -27130
rect 20530 -28120 21530 -28110
rect 21620 -27130 22620 -27120
rect 21620 -28110 21630 -27130
rect 22610 -28110 22620 -27130
rect 21620 -28120 22620 -28110
rect 22710 -27130 23710 -27120
rect 22710 -28110 22720 -27130
rect 23700 -28110 23710 -27130
rect 22710 -28120 23710 -28110
<< mimcapcontact >>
rect -2350 -26830 -1370 -25850
rect -1260 -26830 -280 -25850
rect -170 -26830 810 -25850
rect 920 -26830 1900 -25850
rect 2010 -26830 2990 -25850
rect 3100 -26830 4080 -25850
rect 4190 -26830 5170 -25850
rect 5280 -26830 6260 -25850
rect 6370 -26830 7350 -25850
rect 7460 -26830 8440 -25850
rect 8550 -26830 9530 -25850
rect 9640 -26830 10620 -25850
rect 10730 -26830 11710 -25850
rect 11820 -26830 12800 -25850
rect 12910 -26830 13890 -25850
rect 14000 -26830 14980 -25850
rect 15090 -26830 16070 -25850
rect 16180 -26830 17160 -25850
rect 17270 -26830 18250 -25850
rect 18360 -26830 19340 -25850
rect 19450 -26830 20430 -25850
rect 20540 -26830 21520 -25850
rect 21630 -26830 22610 -25850
rect 22720 -26830 23700 -25850
rect -2350 -28110 -1370 -27130
rect -1260 -28110 -280 -27130
rect -170 -28110 810 -27130
rect 920 -28110 1900 -27130
rect 2010 -28110 2990 -27130
rect 3100 -28110 4080 -27130
rect 4190 -28110 5170 -27130
rect 5280 -28110 6260 -27130
rect 6370 -28110 7350 -27130
rect 7460 -28110 8440 -27130
rect 8550 -28110 9530 -27130
rect 9640 -28110 10620 -27130
rect 10730 -28110 11710 -27130
rect 11820 -28110 12800 -27130
rect 12910 -28110 13890 -27130
rect 14000 -28110 14980 -27130
rect 15090 -28110 16070 -27130
rect 16180 -28110 17160 -27130
rect 17270 -28110 18250 -27130
rect 18360 -28110 19340 -27130
rect 19450 -28110 20430 -27130
rect 20540 -28110 21520 -27130
rect 21630 -28110 22610 -27130
rect 22720 -28110 23700 -27130
<< metal4 >>
rect -3510 -3440 24420 -3430
rect -3510 -3570 24270 -3440
rect 24410 -3570 24420 -3440
rect -3510 -3580 24420 -3570
rect -3510 -3680 24420 -3670
rect -3510 -3810 24270 -3680
rect 24410 -3810 24420 -3680
rect -3510 -3820 24420 -3810
rect -3510 -3920 24420 -3910
rect -3510 -4050 24270 -3920
rect 24410 -4050 24420 -3920
rect -3510 -4060 24420 -4050
rect -3510 -4160 24420 -4150
rect -3510 -4300 24270 -4160
rect 24410 -4300 24420 -4160
rect -3510 -4310 24420 -4300
rect -3510 -4410 24420 -4400
rect -3510 -4540 24270 -4410
rect 24410 -4540 24420 -4410
rect -3510 -4550 24420 -4540
rect -3510 -4650 24420 -4640
rect -3510 -4780 24270 -4650
rect 24410 -4780 24420 -4650
rect -3510 -4790 24420 -4780
rect -3510 -4890 24420 -4880
rect -3510 -5020 24270 -4890
rect 24410 -5020 24420 -4890
rect -3510 -5030 24420 -5020
rect -3510 -7980 24420 -7970
rect -3510 -8110 24270 -7980
rect 24410 -8110 24420 -7980
rect -3510 -8120 24420 -8110
rect -3510 -8220 24420 -8210
rect -3510 -8350 24270 -8220
rect 24410 -8350 24420 -8220
rect -3510 -8360 24420 -8350
rect -3510 -8460 24420 -8450
rect -3510 -8590 24270 -8460
rect 24410 -8590 24420 -8460
rect -3510 -8600 24420 -8590
rect -3510 -8700 24420 -8690
rect -3510 -8840 24270 -8700
rect 24410 -8840 24420 -8700
rect -3510 -8850 24420 -8840
rect -3510 -8950 24420 -8940
rect -3510 -9080 24270 -8950
rect 24410 -9080 24420 -8950
rect -3510 -9090 24420 -9080
rect -3510 -9190 24420 -9180
rect -3510 -9320 24270 -9190
rect 24410 -9320 24420 -9190
rect -3510 -9330 24420 -9320
rect -3510 -9430 24420 -9420
rect -3510 -9560 24270 -9430
rect 24410 -9560 24420 -9430
rect -3510 -9570 24420 -9560
rect -3510 -16000 24420 -15990
rect -3510 -16130 24270 -16000
rect 24410 -16130 24420 -16000
rect -3510 -16140 24420 -16130
rect -3510 -16240 24420 -16230
rect -3510 -16370 24270 -16240
rect 24410 -16370 24420 -16240
rect -3510 -16380 24420 -16370
rect -3510 -16480 24420 -16470
rect -3510 -16610 24270 -16480
rect 24410 -16610 24420 -16480
rect -3510 -16620 24420 -16610
rect -3510 -16720 24420 -16710
rect -3510 -16860 24270 -16720
rect 24410 -16860 24420 -16720
rect -3510 -16870 24420 -16860
rect -3510 -16970 24420 -16960
rect -3510 -17100 24270 -16970
rect 24410 -17100 24420 -16970
rect -3510 -17110 24420 -17100
rect -3510 -17210 24420 -17200
rect -3510 -17340 24270 -17210
rect 24410 -17340 24420 -17210
rect -3510 -17350 24420 -17340
rect -3510 -17450 24420 -17440
rect -3510 -17580 24270 -17450
rect 24410 -17580 24420 -17450
rect -3510 -17590 24420 -17580
rect -3510 -20540 24420 -20530
rect -3510 -20670 24270 -20540
rect 24410 -20670 24420 -20540
rect -3510 -20680 24420 -20670
rect -3510 -20780 24420 -20770
rect -3510 -20910 24270 -20780
rect 24410 -20910 24420 -20780
rect -3510 -20920 24420 -20910
rect -3510 -21020 24420 -21010
rect -3510 -21150 24270 -21020
rect 24410 -21150 24420 -21020
rect -3510 -21160 24420 -21150
rect -3510 -21260 24420 -21250
rect -3510 -21400 24270 -21260
rect 24410 -21400 24420 -21260
rect -3510 -21410 24420 -21400
rect -3510 -21510 24420 -21500
rect -3510 -21640 24270 -21510
rect 24410 -21640 24420 -21510
rect -3510 -21650 24420 -21640
rect -3510 -21750 24420 -21740
rect -3510 -21880 24270 -21750
rect 24410 -21880 24420 -21750
rect -3510 -21890 24420 -21880
rect -3510 -21990 24420 -21980
rect -3510 -22120 24270 -21990
rect 24410 -22120 24420 -21990
rect -3510 -22130 24420 -22120
rect -6210 -25510 24420 -25500
rect -6210 -25650 24270 -25510
rect 24410 -25650 24420 -25510
rect -6210 -25660 24420 -25650
rect -2380 -25850 23730 -25820
rect -2380 -26700 -2350 -25850
rect -4230 -26710 -2350 -26700
rect -4230 -26850 -4220 -26710
rect -4170 -26830 -2350 -26710
rect -1370 -25980 -1260 -25850
rect -1370 -26830 -1340 -25980
rect -4170 -26850 -1340 -26830
rect -4230 -26860 -1340 -26850
rect -1290 -26830 -1260 -25980
rect -280 -25980 -170 -25850
rect -280 -26830 -250 -25980
rect -1290 -26860 -250 -26830
rect -200 -26830 -170 -25980
rect 810 -25980 920 -25850
rect 810 -26830 840 -25980
rect -200 -26860 840 -26830
rect 890 -26830 920 -25980
rect 1900 -25980 2010 -25850
rect 1900 -26830 1930 -25980
rect 890 -26860 1930 -26830
rect 1980 -26830 2010 -25980
rect 2990 -25980 3100 -25850
rect 2990 -26830 3020 -25980
rect 1980 -26860 3020 -26830
rect 3070 -26830 3100 -25980
rect 4080 -25980 4190 -25850
rect 4080 -26830 4110 -25980
rect 3070 -26860 4110 -26830
rect 4160 -26830 4190 -25980
rect 5170 -25980 5280 -25850
rect 5170 -26830 5200 -25980
rect 4160 -26860 5200 -26830
rect 5250 -26830 5280 -25980
rect 6260 -25980 6370 -25850
rect 6260 -26830 6290 -25980
rect 5250 -26860 6290 -26830
rect 6340 -26830 6370 -25980
rect 7350 -25980 7460 -25850
rect 7350 -26830 7380 -25980
rect 6340 -26860 7380 -26830
rect 7430 -26830 7460 -25980
rect 8440 -25980 8550 -25850
rect 8440 -26830 8470 -25980
rect 7430 -26860 8470 -26830
rect 8520 -26830 8550 -25980
rect 9530 -25980 9640 -25850
rect 9530 -26830 9560 -25980
rect 8520 -26860 9560 -26830
rect 9610 -26830 9640 -25980
rect 10620 -25980 10730 -25850
rect 10620 -26830 10650 -25980
rect 9610 -26860 10650 -26830
rect 10700 -26830 10730 -25980
rect 11710 -25980 11820 -25850
rect 11710 -26830 11740 -25980
rect 10700 -26860 11740 -26830
rect 11790 -26830 11820 -25980
rect 12800 -25980 12910 -25850
rect 12800 -26830 12830 -25980
rect 11790 -26860 12830 -26830
rect 12880 -26830 12910 -25980
rect 13890 -25980 14000 -25850
rect 13890 -26830 13920 -25980
rect 12880 -26860 13920 -26830
rect 13970 -26830 14000 -25980
rect 14980 -25980 15090 -25850
rect 14980 -26830 15010 -25980
rect 13970 -26860 15010 -26830
rect 15060 -26830 15090 -25980
rect 16070 -25980 16180 -25850
rect 16070 -26830 16100 -25980
rect 15060 -26860 16100 -26830
rect 16150 -26830 16180 -25980
rect 17160 -25980 17270 -25850
rect 17160 -26830 17190 -25980
rect 16150 -26860 17190 -26830
rect 17240 -26830 17270 -25980
rect 18250 -25980 18360 -25850
rect 18250 -26830 18280 -25980
rect 17240 -26860 18280 -26830
rect 18330 -26830 18360 -25980
rect 19340 -25980 19450 -25850
rect 19340 -26830 19370 -25980
rect 18330 -26860 19370 -26830
rect 19420 -26830 19450 -25980
rect 20430 -25980 20540 -25850
rect 20430 -26830 20460 -25980
rect 19420 -26860 20460 -26830
rect 20510 -26830 20540 -25980
rect 21520 -25980 21630 -25850
rect 21520 -26830 21550 -25980
rect 20510 -26860 21550 -26830
rect 21600 -26830 21630 -25980
rect 22610 -25980 22720 -25850
rect 22610 -26830 22640 -25980
rect 21600 -26860 22640 -26830
rect 22690 -26830 22720 -25980
rect 23700 -26830 23730 -25850
rect 22690 -26860 23730 -26830
rect -5010 -26910 23730 -26900
rect -5010 -27050 -5000 -26910
rect -4790 -26920 23730 -26910
rect -4790 -27040 -2360 -26920
rect -1360 -27040 -1270 -26920
rect -270 -27040 -180 -26920
rect 820 -27040 910 -26920
rect 1910 -27040 2000 -26920
rect 3000 -27040 3090 -26920
rect 4090 -27040 4180 -26920
rect 5180 -27040 5270 -26920
rect 6270 -27040 6360 -26920
rect 7360 -27040 7450 -26920
rect 8450 -27040 8540 -26920
rect 9540 -27040 9630 -26920
rect 10630 -27040 10720 -26920
rect 11720 -27040 11810 -26920
rect 12810 -27040 12900 -26920
rect 13900 -27040 13990 -26920
rect 14990 -27040 15080 -26920
rect 16080 -27040 16170 -26920
rect 17170 -27040 17260 -26920
rect 18260 -27040 18350 -26920
rect 19350 -27040 19440 -26920
rect 20440 -27040 20530 -26920
rect 21530 -27040 21620 -26920
rect 22620 -27040 22710 -26920
rect 23710 -27040 23730 -26920
rect -4790 -27050 23730 -27040
rect -5010 -27060 23730 -27050
rect -4030 -27110 -1340 -27100
rect -4030 -27250 -4020 -27110
rect -3970 -27130 -1340 -27110
rect -3970 -27250 -2350 -27130
rect -4030 -27260 -2350 -27250
rect -2380 -28110 -2350 -27260
rect -1370 -27980 -1340 -27130
rect -1290 -27130 -250 -27100
rect -1290 -27980 -1260 -27130
rect -1370 -28110 -1260 -27980
rect -280 -27980 -250 -27130
rect -200 -27130 840 -27100
rect -200 -27980 -170 -27130
rect -280 -28110 -170 -27980
rect 810 -27980 840 -27130
rect 890 -27130 1930 -27100
rect 890 -27980 920 -27130
rect 810 -28110 920 -27980
rect 1900 -27980 1930 -27130
rect 1980 -27130 3020 -27100
rect 1980 -27980 2010 -27130
rect 1900 -28110 2010 -27980
rect 2990 -27980 3020 -27130
rect 3070 -27130 4110 -27100
rect 3070 -27980 3100 -27130
rect 2990 -28110 3100 -27980
rect 4080 -27980 4110 -27130
rect 4160 -27130 5200 -27100
rect 4160 -27980 4190 -27130
rect 4080 -28110 4190 -27980
rect 5170 -27980 5200 -27130
rect 5250 -27130 6290 -27100
rect 5250 -27980 5280 -27130
rect 5170 -28110 5280 -27980
rect 6260 -27980 6290 -27130
rect 6340 -27130 7380 -27100
rect 6340 -27980 6370 -27130
rect 6260 -28110 6370 -27980
rect 7350 -27980 7380 -27130
rect 7430 -27130 8470 -27100
rect 7430 -27980 7460 -27130
rect 7350 -28110 7460 -27980
rect 8440 -27980 8470 -27130
rect 8520 -27130 9560 -27100
rect 8520 -27980 8550 -27130
rect 8440 -28110 8550 -27980
rect 9530 -27980 9560 -27130
rect 9610 -27130 10650 -27100
rect 9610 -27980 9640 -27130
rect 9530 -28110 9640 -27980
rect 10620 -27980 10650 -27130
rect 10700 -27130 11740 -27100
rect 10700 -27980 10730 -27130
rect 10620 -28110 10730 -27980
rect 11710 -27980 11740 -27130
rect 11790 -27130 12830 -27100
rect 11790 -27980 11820 -27130
rect 11710 -28110 11820 -27980
rect 12800 -27980 12830 -27130
rect 12880 -27130 13920 -27100
rect 12880 -27980 12910 -27130
rect 12800 -28110 12910 -27980
rect 13890 -27980 13920 -27130
rect 13970 -27130 15010 -27100
rect 13970 -27980 14000 -27130
rect 13890 -28110 14000 -27980
rect 14980 -27980 15010 -27130
rect 15060 -27130 16100 -27100
rect 15060 -27980 15090 -27130
rect 14980 -28110 15090 -27980
rect 16070 -27980 16100 -27130
rect 16150 -27130 17190 -27100
rect 16150 -27980 16180 -27130
rect 16070 -28110 16180 -27980
rect 17160 -27980 17190 -27130
rect 17240 -27130 18280 -27100
rect 17240 -27980 17270 -27130
rect 17160 -28110 17270 -27980
rect 18250 -27980 18280 -27130
rect 18330 -27130 19370 -27100
rect 18330 -27980 18360 -27130
rect 18250 -28110 18360 -27980
rect 19340 -27980 19370 -27130
rect 19420 -27130 20460 -27100
rect 19420 -27980 19450 -27130
rect 19340 -28110 19450 -27980
rect 20430 -27980 20460 -27130
rect 20510 -27130 21550 -27100
rect 20510 -27980 20540 -27130
rect 20430 -28110 20540 -27980
rect 21520 -27980 21550 -27130
rect 21600 -27130 22640 -27100
rect 21600 -27980 21630 -27130
rect 21520 -28110 21630 -27980
rect 22610 -27980 22640 -27130
rect 22690 -27130 23730 -27100
rect 22690 -27980 22720 -27130
rect 22610 -28110 22720 -27980
rect 23700 -28110 23730 -27130
rect -2380 -28140 23730 -28110
rect -6310 -28310 24420 -28300
rect -6310 -28450 -3520 -28310
rect -3470 -28450 24270 -28310
rect 24410 -28450 24420 -28310
rect -6310 -28460 24420 -28450
<< metal5 >>
rect -6210 -28520 -5980 -220
rect -5810 -28520 -5580 -220
rect -5410 -28520 -5180 -220
rect -5010 -28520 -4780 -220
rect -4610 -28520 -4380 -220
rect -4210 -28520 -3980 -220
rect -3810 -28520 -3580 -220
use p8_1  p8_1_35
timestamp 1634440961
transform 1 0 -2820 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_27
timestamp 1634440922
transform 1 0 -1880 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_34
timestamp 1634440961
transform 1 0 -940 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_28
timestamp 1634440922
transform 1 0 0 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_29
timestamp 1634440922
transform 1 0 940 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_32
timestamp 1634440961
transform 1 0 1880 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_26
timestamp 1634440922
transform 1 0 2820 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_33
timestamp 1634440961
transform 1 0 3760 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_30
timestamp 1634440961
transform 1 0 5640 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_24
timestamp 1634440922
transform 1 0 4700 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_31
timestamp 1634440961
transform 1 0 7520 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_25
timestamp 1634440922
transform 1 0 6580 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_29
timestamp 1634440961
transform 1 0 8460 0 -1 -22200
box 0 0 940 2970
use p4_2  p4_2_4
timestamp 1634665005
transform 1 0 9400 0 -1 -22200
box 0 0 940 2970
use p4_2  p4_2_5
timestamp 1634665005
transform -1 0 11280 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_26
timestamp 1634440961
transform -1 0 12220 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_27
timestamp 1634440961
transform -1 0 13160 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_23
timestamp 1634440922
transform -1 0 14100 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_28
timestamp 1634440961
transform -1 0 15040 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_21
timestamp 1634440922
transform -1 0 15980 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_24
timestamp 1634440961
transform -1 0 16920 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_22
timestamp 1634440922
transform -1 0 17860 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_25
timestamp 1634440961
transform -1 0 18800 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_19
timestamp 1634440922
transform -1 0 19740 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_20
timestamp 1634440922
transform -1 0 20680 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_23
timestamp 1634440961
transform -1 0 21620 0 -1 -22200
box 0 0 940 2970
use p8_1  p8_1_22
timestamp 1634440961
transform -1 0 23500 0 -1 -22200
box 0 0 940 2970
use p1_8  p1_8_18
timestamp 1634440922
transform -1 0 22560 0 -1 -22200
box 0 0 940 2970
use n8_1  n8_1_48
timestamp 1634429522
transform 1 0 -2820 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_49
timestamp 1634429522
transform 1 0 -2820 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_36
timestamp 1634337365
transform 1 0 -1880 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_39
timestamp 1634337365
transform 1 0 -1880 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_37
timestamp 1634337365
transform 1 0 -940 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_46
timestamp 1634429522
transform 1 0 0 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_40
timestamp 1634337365
transform 1 0 -940 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_47
timestamp 1634429522
transform 1 0 0 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_38
timestamp 1634337365
transform 1 0 940 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_41
timestamp 1634337365
transform 1 0 940 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_42
timestamp 1634429522
transform 1 0 1880 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_44
timestamp 1634429522
transform 1 0 1880 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_34
timestamp 1634337365
transform 1 0 2820 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_43
timestamp 1634429522
transform 1 0 3760 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_35
timestamp 1634337365
transform 1 0 2820 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_45
timestamp 1634429522
transform 1 0 3760 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_30
timestamp 1634337365
transform 1 0 4700 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_38
timestamp 1634429522
transform 1 0 5640 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_32
timestamp 1634337365
transform 1 0 4700 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_40
timestamp 1634429522
transform 1 0 5640 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_31
timestamp 1634337365
transform 1 0 6580 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_39
timestamp 1634429522
transform 1 0 7520 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_33
timestamp 1634337365
transform 1 0 6580 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_41
timestamp 1634429522
transform 1 0 7520 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_36
timestamp 1634429522
transform 1 0 8460 0 1 -18890
box 0 0 940 1230
use n4_2  n4_2_4
timestamp 1634664854
transform 1 0 9400 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_37
timestamp 1634429522
transform 1 0 8460 0 -1 -19230
box 0 0 940 1230
use n4_2  n4_2_6
timestamp 1634664854
transform 1 0 9400 0 -1 -19230
box 0 0 940 1230
use n4_2  n4_2_5
timestamp 1634664854
transform -1 0 11280 0 1 -18890
box 0 0 940 1230
use n4_2  n4_2_7
timestamp 1634664854
transform -1 0 11280 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_30
timestamp 1634429522
transform -1 0 12220 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_31
timestamp 1634429522
transform -1 0 13160 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_28
timestamp 1634337365
transform -1 0 14100 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_33
timestamp 1634429522
transform -1 0 12220 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_34
timestamp 1634429522
transform -1 0 13160 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_29
timestamp 1634337365
transform -1 0 14100 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_32
timestamp 1634429522
transform -1 0 15040 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_35
timestamp 1634429522
transform -1 0 15040 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_24
timestamp 1634337365
transform -1 0 15980 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_26
timestamp 1634429522
transform -1 0 16920 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_25
timestamp 1634337365
transform -1 0 17860 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_26
timestamp 1634337365
transform -1 0 15980 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_28
timestamp 1634429522
transform -1 0 16920 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_27
timestamp 1634337365
transform -1 0 17860 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_27
timestamp 1634429522
transform -1 0 18800 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_29
timestamp 1634429522
transform -1 0 18800 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_20
timestamp 1634337365
transform -1 0 19740 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_24
timestamp 1634429522
transform -1 0 20680 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_21
timestamp 1634337365
transform -1 0 21620 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_22
timestamp 1634337365
transform -1 0 19740 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_25
timestamp 1634429522
transform -1 0 20680 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_23
timestamp 1634337365
transform -1 0 21620 0 -1 -19230
box 0 0 940 1230
use n1_8  n1_8_18
timestamp 1634337365
transform -1 0 22560 0 1 -18890
box 0 0 940 1230
use n8_1  n8_1_22
timestamp 1634429522
transform -1 0 23500 0 1 -18890
box 0 0 940 1230
use n1_8  n1_8_19
timestamp 1634337365
transform -1 0 22560 0 -1 -19230
box 0 0 940 1230
use n8_1  n8_1_23
timestamp 1634429522
transform -1 0 23500 0 -1 -19230
box 0 0 940 1230
use p8_1  p8_1_49
timestamp 1634440961
transform 1 0 -2820 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_39
timestamp 1634440922
transform 1 0 -1880 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_48
timestamp 1634440961
transform 1 0 -940 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_40
timestamp 1634440922
transform 1 0 0 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_41
timestamp 1634440922
transform 1 0 940 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_46
timestamp 1634440961
transform 1 0 1880 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_38
timestamp 1634440922
transform 1 0 2820 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_47
timestamp 1634440961
transform 1 0 3760 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_36
timestamp 1634440922
transform 1 0 4700 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_44
timestamp 1634440961
transform 1 0 5640 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_37
timestamp 1634440922
transform 1 0 6580 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_45
timestamp 1634440961
transform 1 0 7520 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_43
timestamp 1634440961
transform 1 0 8460 0 1 -15920
box 0 0 940 2970
use p4_2  p4_2_6
timestamp 1634665005
transform 1 0 9400 0 1 -15920
box 0 0 940 2970
use p4_2  p4_2_7
timestamp 1634665005
transform -1 0 11280 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_40
timestamp 1634440961
transform -1 0 12220 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_41
timestamp 1634440961
transform -1 0 13160 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_35
timestamp 1634440922
transform -1 0 14100 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_42
timestamp 1634440961
transform -1 0 15040 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_33
timestamp 1634440922
transform -1 0 15980 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_38
timestamp 1634440961
transform -1 0 16920 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_34
timestamp 1634440922
transform -1 0 17860 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_39
timestamp 1634440961
transform -1 0 18800 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_31
timestamp 1634440922
transform -1 0 19740 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_32
timestamp 1634440922
transform -1 0 20680 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_37
timestamp 1634440961
transform -1 0 21620 0 1 -15920
box 0 0 940 2970
use p1_8  p1_8_30
timestamp 1634440922
transform -1 0 22560 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_36
timestamp 1634440961
transform -1 0 23500 0 1 -15920
box 0 0 940 2970
use p8_1  p8_1_21
timestamp 1634440961
transform 1 0 -2820 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_16
timestamp 1634440922
transform 1 0 -1880 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_20
timestamp 1634440961
transform 1 0 -940 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_17
timestamp 1634440922
transform 1 0 0 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_14
timestamp 1634440922
transform 1 0 940 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_18
timestamp 1634440961
transform 1 0 1880 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_15
timestamp 1634440922
transform 1 0 2820 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_19
timestamp 1634440961
transform 1 0 3760 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_12
timestamp 1634440922
transform 1 0 4700 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_17
timestamp 1634440961
transform 1 0 5640 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_13
timestamp 1634440922
transform 1 0 6580 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_15
timestamp 1634440961
transform 1 0 7520 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_16
timestamp 1634440961
transform 1 0 8460 0 -1 -9640
box 0 0 940 2970
use p4_2  p4_2_2
timestamp 1634665005
transform 1 0 9400 0 -1 -9640
box 0 0 940 2970
use p4_2  p4_2_3
timestamp 1634665005
transform -1 0 11280 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_13
timestamp 1634440961
transform -1 0 12220 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_14
timestamp 1634440961
transform -1 0 13160 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_11
timestamp 1634440922
transform -1 0 14100 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_11
timestamp 1634440961
transform -1 0 15040 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_9
timestamp 1634440922
transform -1 0 15980 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_12
timestamp 1634440961
transform -1 0 16920 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_10
timestamp 1634440922
transform -1 0 17860 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_9
timestamp 1634440961
transform -1 0 18800 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_7
timestamp 1634440922
transform -1 0 19740 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_8
timestamp 1634440922
transform -1 0 20680 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_10
timestamp 1634440961
transform -1 0 21620 0 -1 -9640
box 0 0 940 2970
use p1_8  p1_8_6
timestamp 1634440922
transform -1 0 22560 0 -1 -9640
box 0 0 940 2970
use p8_1  p8_1_6
timestamp 1634440961
transform -1 0 23500 0 -1 -9640
box 0 0 940 2970
use n8_1  n8_1_21
timestamp 1634429522
transform 1 0 -2820 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_16
timestamp 1634337365
transform 1 0 -1880 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_17
timestamp 1634337365
transform 1 0 -940 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_20
timestamp 1634429522
transform 1 0 0 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_18
timestamp 1634429522
transform 1 0 1880 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_15
timestamp 1634337365
transform 1 0 940 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_14
timestamp 1634337365
transform 1 0 2820 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_19
timestamp 1634429522
transform 1 0 3760 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_12
timestamp 1634337365
transform 1 0 4700 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_17
timestamp 1634429522
transform 1 0 5640 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_13
timestamp 1634337365
transform 1 0 6580 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_15
timestamp 1634429522
transform 1 0 8460 0 -1 -6670
box 0 0 940 1230
use n4_2  n4_2_2
timestamp 1634664854
transform 1 0 9400 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_16
timestamp 1634429522
transform 1 0 7520 0 -1 -6670
box 0 0 940 1230
use n4_2  n4_2_3
timestamp 1634664854
transform -1 0 11280 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_13
timestamp 1634429522
transform -1 0 12220 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_14
timestamp 1634429522
transform -1 0 13160 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_11
timestamp 1634337365
transform -1 0 14100 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_12
timestamp 1634429522
transform -1 0 15040 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_9
timestamp 1634337365
transform -1 0 15980 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_11
timestamp 1634429522
transform -1 0 16920 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_10
timestamp 1634337365
transform -1 0 17860 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_9
timestamp 1634429522
transform -1 0 18800 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_7
timestamp 1634337365
transform -1 0 19740 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_10
timestamp 1634429522
transform -1 0 20680 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_8
timestamp 1634337365
transform -1 0 21620 0 -1 -6670
box 0 0 940 1230
use n1_8  n1_8_6
timestamp 1634337365
transform -1 0 22560 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_6
timestamp 1634429522
transform -1 0 23500 0 -1 -6670
box 0 0 940 1230
use n8_1  n8_1_8
timestamp 1634429522
transform 1 0 -2820 0 1 -6330
box 0 0 940 1230
use n1_8  na4_1
timestamp 1634337365
transform 1 0 -1880 0 1 -6330
box 0 0 940 1230
use p1_8  pa1_1
timestamp 1634440922
transform 1 0 -1880 0 1 -3360
box 0 0 940 2970
use p8_1  p8_1_7
timestamp 1634440961
transform 1 0 -2820 0 1 -3360
box 0 0 940 2970
use n1_8  nb4_1
timestamp 1634337365
transform 1 0 -940 0 1 -6330
box 0 0 940 1230
use n8_1  nb3_1
timestamp 1634429522
transform 1 0 0 0 1 -6330
box 0 0 940 1230
use n1_8  ne4_1
timestamp 1634337365
transform 1 0 940 0 1 -6330
box 0 0 940 1230
use n8_1  ne3_1
timestamp 1634429522
transform 1 0 1880 0 1 -6330
box 0 0 940 1230
use p8_1  pa2_1
timestamp 1634440961
transform 1 0 -940 0 1 -3360
box 0 0 940 2970
use p1_8  pb1_1
timestamp 1634440922
transform 1 0 0 0 1 -3360
box 0 0 940 2970
use p1_8  pc1_1
timestamp 1634440922
transform 1 0 940 0 1 -3360
box 0 0 940 2970
use p8_1  pc2_1
timestamp 1634440961
transform 1 0 1880 0 1 -3360
box 0 0 940 2970
use n1_8  nf4_1
timestamp 1634337365
transform 1 0 2820 0 1 -6330
box 0 0 940 1230
use n8_1  nf3_1
timestamp 1634429522
transform 1 0 3760 0 1 -6330
box 0 0 940 1230
use n1_8  nf4_2
timestamp 1634337365
transform 1 0 4700 0 1 -6330
box 0 0 940 1230
use n8_1  nf3_2
timestamp 1634429522
transform 1 0 5640 0 1 -6330
box 0 0 940 1230
use p1_8  pd1_1
timestamp 1634440922
transform 1 0 2820 0 1 -3360
box 0 0 940 2970
use p8_1  pd2_1
timestamp 1634440961
transform 1 0 3760 0 1 -3360
box 0 0 940 2970
use p1_8  pe1_1
timestamp 1634440922
transform 1 0 4700 0 1 -3360
box 0 0 940 2970
use p8_1  pd2_2
timestamp 1634440961
transform 1 0 5640 0 1 -3360
box 0 0 940 2970
use n1_8  ne4_2
timestamp 1634337365
transform 1 0 6580 0 1 -6330
box 0 0 940 1230
use n8_1  ne3_2
timestamp 1634429522
transform 1 0 7520 0 1 -6330
box 0 0 940 1230
use n8_1  nf2_1
timestamp 1634429522
transform 1 0 8460 0 1 -6330
box 0 0 940 1230
use n4_2  n4_2_0
timestamp 1634664854
transform 1 0 9400 0 1 -6330
box 0 0 940 1230
use p1_8  pf1_1
timestamp 1634440922
transform 1 0 6580 0 1 -3360
box 0 0 940 2970
use p8_1  pc2_2
timestamp 1634440961
transform 1 0 7520 0 1 -3360
box 0 0 940 2970
use p8_1  pf2_1
timestamp 1634440961
transform 1 0 8460 0 1 -3360
box 0 0 940 2970
use p4_2  p4_2_0
timestamp 1634665005
transform 1 0 9400 0 1 -3360
box 0 0 940 2970
use n4_2  n4_2_1
timestamp 1634664854
transform -1 0 11280 0 1 -6330
box 0 0 940 1230
use n8_1  n8_1_5
timestamp 1634429522
transform -1 0 12220 0 1 -6330
box 0 0 940 1230
use n8_1  n8_1_4
timestamp 1634429522
transform -1 0 13160 0 1 -6330
box 0 0 940 1230
use n1_8  n1_8_5
timestamp 1634337365
transform -1 0 14100 0 1 -6330
box 0 0 940 1230
use p4_2  p4_2_1
timestamp 1634665005
transform -1 0 11280 0 1 -3360
box 0 0 940 2970
use p8_1  p8_1_5
timestamp 1634440961
transform -1 0 12220 0 1 -3360
box 0 0 940 2970
use p8_1  p8_1_4
timestamp 1634440961
transform -1 0 13160 0 1 -3360
box 0 0 940 2970
use p1_8  p1_8_5
timestamp 1634440922
transform -1 0 14100 0 1 -3360
box 0 0 940 2970
use n8_1  n8_1_3
timestamp 1634429522
transform -1 0 15040 0 1 -6330
box 0 0 940 1230
use n1_8  n1_8_4
timestamp 1634337365
transform -1 0 15980 0 1 -6330
box 0 0 940 1230
use n8_1  n8_1_2
timestamp 1634429522
transform -1 0 16920 0 1 -6330
box 0 0 940 1230
use n1_8  n1_8_3
timestamp 1634337365
transform -1 0 17860 0 1 -6330
box 0 0 940 1230
use p8_1  p8_1_3
timestamp 1634440961
transform -1 0 15040 0 1 -3360
box 0 0 940 2970
use p1_8  p1_8_4
timestamp 1634440922
transform -1 0 15980 0 1 -3360
box 0 0 940 2970
use p8_1  p8_1_2
timestamp 1634440961
transform -1 0 16920 0 1 -3360
box 0 0 940 2970
use p1_8  p1_8_3
timestamp 1634440922
transform -1 0 17860 0 1 -3360
box 0 0 940 2970
use n8_1  n8_1_1
timestamp 1634429522
transform -1 0 18800 0 1 -6330
box 0 0 940 1230
use n1_8  n1_8_2
timestamp 1634337365
transform -1 0 19740 0 1 -6330
box 0 0 940 1230
use n8_1  n8_1_0
timestamp 1634429522
transform -1 0 20680 0 1 -6330
box 0 0 940 1230
use n1_8  n1_8_0
timestamp 1634337365
transform -1 0 21620 0 1 -6330
box 0 0 940 1230
use p8_1  p8_1_1
timestamp 1634440961
transform -1 0 18800 0 1 -3360
box 0 0 940 2970
use p1_8  p1_8_2
timestamp 1634440922
transform -1 0 19740 0 1 -3360
box 0 0 940 2970
use p1_8  p1_8_1
timestamp 1634440922
transform -1 0 20680 0 1 -3360
box 0 0 940 2970
use p8_1  p8_1_0
timestamp 1634440961
transform -1 0 21620 0 1 -3360
box 0 0 940 2970
use n1_8  n1_8_1
timestamp 1634337365
transform -1 0 22560 0 1 -6330
box 0 0 940 1230
use n8_1  n8_1_7
timestamp 1634429522
transform -1 0 23500 0 1 -6330
box 0 0 940 1230
use p1_8  p1_8_0
timestamp 1634440922
transform -1 0 22560 0 1 -3360
box 0 0 940 2970
use p8_1  p8_1_8
timestamp 1634440961
transform -1 0 23500 0 1 -3360
box 0 0 940 2970
<< labels >>
rlabel metal3 23940 -220 24100 -190 1 vdda
port 5 n
rlabel metal3 24260 -220 24420 -190 1 gnda
port 6 n
rlabel metal3 23620 -220 23780 -190 1 vssa
port 7 n
rlabel metal3 -3610 -220 -3580 -190 1 n1
rlabel metal3 -3810 -220 -3780 -190 1 n2
rlabel metal3 -4010 -220 -3980 -190 1 c
rlabel metal3 -4210 -220 -4180 -190 1 b
rlabel metal3 -4410 -220 -4380 -190 1 a
rlabel metal3 -4610 -220 -4580 -190 1 xp
rlabel metal3 -5010 -220 -4780 -190 1 out
port 3 n
rlabel metal3 -5610 -220 -5580 -190 1 inm
port 1 n
rlabel metal3 -5410 -220 -5380 -190 1 inp
port 2 n
rlabel metal3 -5210 -220 -5180 -190 1 xm
rlabel metal3 -5810 -220 -5780 -190 1 x
rlabel metal3 -6210 -220 -6180 -190 1 p1
rlabel metal3 -6010 -220 -5980 -190 1 ib
port 4 n
rlabel metal2 -6310 -3820 -6300 -3790 3 inm
<< end >>
