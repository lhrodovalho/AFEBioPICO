magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< error_p >>
rect -472 4240 4552 4312
rect -472 4160 -400 4240
rect -386 4200 4466 4226
rect -386 3240 -360 4200
rect -320 4134 4400 4160
rect -320 3352 -248 4134
rect 4374 3352 4400 4134
rect -320 3280 4400 3352
rect 4440 3240 4466 4200
rect 4480 3280 4552 4240
rect 8008 4240 13032 4312
rect 8008 4160 8080 4240
rect 8094 4200 12946 4226
rect -386 3214 4466 3240
rect 8094 3240 8120 4200
rect 8160 4134 12880 4160
rect 8160 3352 8232 4134
rect 12854 3352 12880 4134
rect 8160 3280 12880 3352
rect 12920 3240 12946 4200
rect 12960 3280 13032 4240
rect 8094 3214 12946 3240
rect -472 2960 4552 3032
rect -472 2880 -400 2960
rect -386 2920 4466 2946
rect -386 1960 -360 2920
rect -320 2854 4400 2880
rect -320 2072 -248 2854
rect 4374 2072 4400 2854
rect -320 2000 4400 2072
rect 4440 1960 4466 2920
rect 4480 2000 4552 2960
rect 8008 2960 13032 3032
rect 8008 2880 8080 2960
rect 8094 2920 12946 2946
rect -386 1934 4466 1960
rect 8094 1960 8120 2920
rect 8160 2854 12880 2880
rect 8160 2072 8232 2854
rect 12854 2072 12880 2854
rect 8160 2000 12880 2072
rect 12920 1960 12946 2920
rect 12960 2000 13032 2960
rect 8094 1934 12946 1960
rect -472 1680 4552 1752
rect -472 1600 -400 1680
rect -386 1640 4466 1666
rect -386 680 -360 1640
rect -320 1574 4400 1600
rect -320 792 -248 1574
rect 4374 792 4400 1574
rect -320 720 4400 792
rect 4440 680 4466 1640
rect 4480 720 4552 1680
rect 8008 1680 13032 1752
rect 8008 1600 8080 1680
rect 8094 1640 12946 1666
rect -386 654 4466 680
rect 8094 680 8120 1640
rect 8160 1574 12880 1600
rect 8160 792 8232 1574
rect 12854 792 12880 1574
rect 8160 720 12880 792
rect 12920 680 12946 1640
rect 12960 720 13032 1680
rect 8094 654 12946 680
rect -472 400 4552 472
rect -472 320 -400 400
rect -386 360 4466 386
rect -386 -600 -360 360
rect -320 294 4400 320
rect -320 -488 -248 294
rect 4374 -488 4400 294
rect -320 -560 4400 -488
rect 4440 -600 4466 360
rect 4480 -560 4552 400
rect 8008 400 13032 472
rect 8008 320 8080 400
rect 8094 360 12946 386
rect -386 -626 4466 -600
rect 8094 -600 8120 360
rect 8160 294 12880 320
rect 8160 -488 8232 294
rect 12854 -488 12880 294
rect 8160 -560 12880 -488
rect 12920 -600 12946 360
rect 12960 -560 13032 400
rect 8094 -626 12946 -600
<< nwell >>
rect -360 3240 4440 4200
rect -360 1960 4440 2920
rect -360 680 4440 1640
rect -360 -600 4440 360
rect 8120 3240 12920 4200
rect 8120 1960 12920 2920
rect 8120 680 12920 1640
rect 8120 -600 12920 360
<< pwell >>
rect -506 4214 4586 4346
rect -506 3226 -374 4214
rect 4454 3226 4586 4214
rect -506 2934 4586 3226
rect -506 1946 -374 2934
rect 4454 1946 4586 2934
rect -506 1654 4586 1946
rect -506 666 -374 1654
rect 4454 666 4586 1654
rect -506 374 4586 666
rect -506 -614 -374 374
rect 4454 -614 4586 374
rect -506 -746 4586 -614
rect 7974 4214 13066 4346
rect 7974 3226 8106 4214
rect 12934 3226 13066 4214
rect 7974 2934 13066 3226
rect 7974 1946 8106 2934
rect 12934 1946 13066 2934
rect 7974 1654 13066 1946
rect 7974 666 8106 1654
rect 12934 666 13066 1654
rect 7974 374 13066 666
rect 7974 -614 8106 374
rect 12934 -614 13066 374
rect 7974 -746 13066 -614
<< mvpmos >>
rect 40 3916 4040 4000
rect 40 3596 4040 3680
rect 8520 3916 12520 4000
rect 8520 3596 12520 3680
rect 40 2480 4040 2564
rect 40 2160 4040 2244
rect 8520 2480 12520 2564
rect 8520 2160 12520 2244
rect 40 1356 4040 1440
rect 40 1036 4040 1120
rect 8520 1356 12520 1440
rect 8520 1036 12520 1120
rect 40 -80 4040 4
rect 40 -400 4040 -316
rect 8520 -80 12520 4
rect 8520 -400 12520 -316
<< mvpdiff >>
rect -160 3977 40 4000
rect -160 3943 -137 3977
rect -103 3943 40 3977
rect -160 3916 40 3943
rect 4040 3977 4240 4000
rect 4040 3943 4183 3977
rect 4217 3943 4240 3977
rect 4040 3916 4240 3943
rect -160 3657 40 3680
rect -160 3623 -137 3657
rect -103 3623 40 3657
rect -160 3596 40 3623
rect 4040 3657 4240 3680
rect 4040 3623 4183 3657
rect 4217 3623 4240 3657
rect 4040 3596 4240 3623
rect 8320 3977 8520 4000
rect 8320 3943 8343 3977
rect 8377 3943 8520 3977
rect 8320 3916 8520 3943
rect 12520 3977 12720 4000
rect 12520 3943 12663 3977
rect 12697 3943 12720 3977
rect 12520 3916 12720 3943
rect 8320 3657 8520 3680
rect 8320 3623 8343 3657
rect 8377 3623 8520 3657
rect 8320 3596 8520 3623
rect 12520 3657 12720 3680
rect 12520 3623 12663 3657
rect 12697 3623 12720 3657
rect 12520 3596 12720 3623
rect -160 2537 40 2564
rect -160 2503 -137 2537
rect -103 2503 40 2537
rect -160 2480 40 2503
rect 4040 2537 4240 2564
rect 4040 2503 4183 2537
rect 4217 2503 4240 2537
rect 4040 2480 4240 2503
rect -160 2217 40 2244
rect -160 2183 -137 2217
rect -103 2183 40 2217
rect -160 2160 40 2183
rect 4040 2217 4240 2244
rect 4040 2183 4183 2217
rect 4217 2183 4240 2217
rect 4040 2160 4240 2183
rect 8320 2537 8520 2564
rect 8320 2503 8343 2537
rect 8377 2503 8520 2537
rect 8320 2480 8520 2503
rect 12520 2537 12720 2564
rect 12520 2503 12663 2537
rect 12697 2503 12720 2537
rect 12520 2480 12720 2503
rect 8320 2217 8520 2244
rect 8320 2183 8343 2217
rect 8377 2183 8520 2217
rect 8320 2160 8520 2183
rect 12520 2217 12720 2244
rect 12520 2183 12663 2217
rect 12697 2183 12720 2217
rect 12520 2160 12720 2183
rect -160 1417 40 1440
rect -160 1383 -137 1417
rect -103 1383 40 1417
rect -160 1356 40 1383
rect 4040 1417 4240 1440
rect 4040 1383 4183 1417
rect 4217 1383 4240 1417
rect 4040 1356 4240 1383
rect -160 1097 40 1120
rect -160 1063 -137 1097
rect -103 1063 40 1097
rect -160 1036 40 1063
rect 4040 1097 4240 1120
rect 4040 1063 4183 1097
rect 4217 1063 4240 1097
rect 4040 1036 4240 1063
rect 8320 1417 8520 1440
rect 8320 1383 8343 1417
rect 8377 1383 8520 1417
rect 8320 1356 8520 1383
rect 12520 1417 12720 1440
rect 12520 1383 12663 1417
rect 12697 1383 12720 1417
rect 12520 1356 12720 1383
rect 8320 1097 8520 1120
rect 8320 1063 8343 1097
rect 8377 1063 8520 1097
rect 8320 1036 8520 1063
rect 12520 1097 12720 1120
rect 12520 1063 12663 1097
rect 12697 1063 12720 1097
rect 12520 1036 12720 1063
rect -160 -23 40 4
rect -160 -57 -137 -23
rect -103 -57 40 -23
rect -160 -80 40 -57
rect 4040 -23 4240 4
rect 4040 -57 4183 -23
rect 4217 -57 4240 -23
rect 4040 -80 4240 -57
rect -160 -343 40 -316
rect -160 -377 -137 -343
rect -103 -377 40 -343
rect -160 -400 40 -377
rect 4040 -343 4240 -316
rect 4040 -377 4183 -343
rect 4217 -377 4240 -343
rect 4040 -400 4240 -377
rect 8320 -23 8520 4
rect 8320 -57 8343 -23
rect 8377 -57 8520 -23
rect 8320 -80 8520 -57
rect 12520 -23 12720 4
rect 12520 -57 12663 -23
rect 12697 -57 12720 -23
rect 12520 -80 12720 -57
rect 8320 -343 8520 -316
rect 8320 -377 8343 -343
rect 8377 -377 8520 -343
rect 8320 -400 8520 -377
rect 12520 -343 12720 -316
rect 12520 -377 12663 -343
rect 12697 -377 12720 -343
rect 12520 -400 12720 -377
<< mvpdiffc >>
rect -137 3943 -103 3977
rect 4183 3943 4217 3977
rect -137 3623 -103 3657
rect 4183 3623 4217 3657
rect 8343 3943 8377 3977
rect 12663 3943 12697 3977
rect 8343 3623 8377 3657
rect 12663 3623 12697 3657
rect -137 2503 -103 2537
rect 4183 2503 4217 2537
rect -137 2183 -103 2217
rect 4183 2183 4217 2217
rect 8343 2503 8377 2537
rect 12663 2503 12697 2537
rect 8343 2183 8377 2217
rect 12663 2183 12697 2217
rect -137 1383 -103 1417
rect 4183 1383 4217 1417
rect -137 1063 -103 1097
rect 4183 1063 4217 1097
rect 8343 1383 8377 1417
rect 12663 1383 12697 1417
rect 8343 1063 8377 1097
rect 12663 1063 12697 1097
rect -137 -57 -103 -23
rect 4183 -57 4217 -23
rect -137 -377 -103 -343
rect 4183 -377 4217 -343
rect 8343 -57 8377 -23
rect 12663 -57 12697 -23
rect 8343 -377 8377 -343
rect 12663 -377 12697 -343
<< psubdiff >>
rect -480 4297 4560 4320
rect -480 4263 -357 4297
rect -323 4263 -289 4297
rect -255 4263 -221 4297
rect -187 4263 -153 4297
rect -119 4263 -85 4297
rect -51 4263 -17 4297
rect 17 4263 51 4297
rect 85 4263 119 4297
rect 153 4263 187 4297
rect 221 4263 255 4297
rect 289 4263 323 4297
rect 357 4263 391 4297
rect 425 4263 459 4297
rect 493 4263 527 4297
rect 561 4263 595 4297
rect 629 4263 663 4297
rect 697 4263 731 4297
rect 765 4263 799 4297
rect 833 4263 867 4297
rect 901 4263 935 4297
rect 969 4263 1003 4297
rect 1037 4263 1071 4297
rect 1105 4263 1139 4297
rect 1173 4263 1207 4297
rect 1241 4263 1275 4297
rect 1309 4263 1343 4297
rect 1377 4263 1411 4297
rect 1445 4263 1479 4297
rect 1513 4263 1547 4297
rect 1581 4263 1615 4297
rect 1649 4263 1683 4297
rect 1717 4263 1751 4297
rect 1785 4263 1819 4297
rect 1853 4263 1887 4297
rect 1921 4263 1955 4297
rect 1989 4263 2023 4297
rect 2057 4263 2091 4297
rect 2125 4263 2159 4297
rect 2193 4263 2227 4297
rect 2261 4263 2295 4297
rect 2329 4263 2363 4297
rect 2397 4263 2431 4297
rect 2465 4263 2499 4297
rect 2533 4263 2567 4297
rect 2601 4263 2635 4297
rect 2669 4263 2703 4297
rect 2737 4263 2771 4297
rect 2805 4263 2839 4297
rect 2873 4263 2907 4297
rect 2941 4263 2975 4297
rect 3009 4263 3043 4297
rect 3077 4263 3111 4297
rect 3145 4263 3179 4297
rect 3213 4263 3247 4297
rect 3281 4263 3315 4297
rect 3349 4263 3383 4297
rect 3417 4263 3451 4297
rect 3485 4263 3519 4297
rect 3553 4263 3587 4297
rect 3621 4263 3655 4297
rect 3689 4263 3723 4297
rect 3757 4263 3791 4297
rect 3825 4263 3859 4297
rect 3893 4263 3927 4297
rect 3961 4263 3995 4297
rect 4029 4263 4063 4297
rect 4097 4263 4131 4297
rect 4165 4263 4199 4297
rect 4233 4263 4267 4297
rect 4301 4263 4335 4297
rect 4369 4263 4403 4297
rect 4437 4263 4560 4297
rect -480 4240 4560 4263
rect -480 4199 -400 4240
rect -480 4165 -457 4199
rect -423 4165 -400 4199
rect -480 4131 -400 4165
rect 4480 4199 4560 4240
rect 4480 4165 4503 4199
rect 4537 4165 4560 4199
rect -480 4097 -457 4131
rect -423 4097 -400 4131
rect -480 4063 -400 4097
rect -480 4029 -457 4063
rect -423 4029 -400 4063
rect -480 3995 -400 4029
rect -480 3961 -457 3995
rect -423 3961 -400 3995
rect -480 3927 -400 3961
rect -480 3893 -457 3927
rect -423 3893 -400 3927
rect -480 3859 -400 3893
rect -480 3825 -457 3859
rect -423 3825 -400 3859
rect -480 3791 -400 3825
rect -480 3757 -457 3791
rect -423 3757 -400 3791
rect -480 3723 -400 3757
rect -480 3689 -457 3723
rect -423 3689 -400 3723
rect -480 3655 -400 3689
rect -480 3621 -457 3655
rect -423 3621 -400 3655
rect -480 3587 -400 3621
rect -480 3553 -457 3587
rect -423 3553 -400 3587
rect -480 3519 -400 3553
rect -480 3485 -457 3519
rect -423 3485 -400 3519
rect -480 3451 -400 3485
rect -480 3417 -457 3451
rect -423 3417 -400 3451
rect -480 3383 -400 3417
rect -480 3349 -457 3383
rect -423 3349 -400 3383
rect -480 3315 -400 3349
rect -480 3281 -457 3315
rect -423 3281 -400 3315
rect -480 3200 -400 3281
rect 4480 4131 4560 4165
rect 4480 4097 4503 4131
rect 4537 4097 4560 4131
rect 4480 4063 4560 4097
rect 4480 4029 4503 4063
rect 4537 4029 4560 4063
rect 4480 3995 4560 4029
rect 4480 3961 4503 3995
rect 4537 3961 4560 3995
rect 4480 3927 4560 3961
rect 4480 3893 4503 3927
rect 4537 3893 4560 3927
rect 4480 3859 4560 3893
rect 4480 3825 4503 3859
rect 4537 3825 4560 3859
rect 4480 3791 4560 3825
rect 4480 3757 4503 3791
rect 4537 3757 4560 3791
rect 4480 3723 4560 3757
rect 4480 3689 4503 3723
rect 4537 3689 4560 3723
rect 4480 3655 4560 3689
rect 4480 3621 4503 3655
rect 4537 3621 4560 3655
rect 4480 3587 4560 3621
rect 4480 3553 4503 3587
rect 4537 3553 4560 3587
rect 4480 3519 4560 3553
rect 4480 3485 4503 3519
rect 4537 3485 4560 3519
rect 4480 3451 4560 3485
rect 4480 3417 4503 3451
rect 4537 3417 4560 3451
rect 4480 3383 4560 3417
rect 4480 3349 4503 3383
rect 4537 3349 4560 3383
rect 4480 3315 4560 3349
rect 4480 3281 4503 3315
rect 4537 3281 4560 3315
rect 4480 3200 4560 3281
rect -480 3177 4560 3200
rect -480 3143 -357 3177
rect -323 3143 -289 3177
rect -255 3143 -221 3177
rect -187 3143 -153 3177
rect -119 3143 -85 3177
rect -51 3143 -17 3177
rect 17 3143 51 3177
rect 85 3143 119 3177
rect 153 3143 187 3177
rect 221 3143 255 3177
rect 289 3143 323 3177
rect 357 3143 391 3177
rect 425 3143 459 3177
rect 493 3143 527 3177
rect 561 3143 595 3177
rect 629 3143 663 3177
rect 697 3143 731 3177
rect 765 3143 799 3177
rect 833 3143 867 3177
rect 901 3143 935 3177
rect 969 3143 1003 3177
rect 1037 3143 1071 3177
rect 1105 3143 1139 3177
rect 1173 3143 1207 3177
rect 1241 3143 1275 3177
rect 1309 3143 1343 3177
rect 1377 3143 1411 3177
rect 1445 3143 1479 3177
rect 1513 3143 1547 3177
rect 1581 3143 1615 3177
rect 1649 3143 1683 3177
rect 1717 3143 1751 3177
rect 1785 3143 1819 3177
rect 1853 3143 1887 3177
rect 1921 3143 1955 3177
rect 1989 3143 2023 3177
rect 2057 3143 2091 3177
rect 2125 3143 2159 3177
rect 2193 3143 2227 3177
rect 2261 3143 2295 3177
rect 2329 3143 2363 3177
rect 2397 3143 2431 3177
rect 2465 3143 2499 3177
rect 2533 3143 2567 3177
rect 2601 3143 2635 3177
rect 2669 3143 2703 3177
rect 2737 3143 2771 3177
rect 2805 3143 2839 3177
rect 2873 3143 2907 3177
rect 2941 3143 2975 3177
rect 3009 3143 3043 3177
rect 3077 3143 3111 3177
rect 3145 3143 3179 3177
rect 3213 3143 3247 3177
rect 3281 3143 3315 3177
rect 3349 3143 3383 3177
rect 3417 3143 3451 3177
rect 3485 3143 3519 3177
rect 3553 3143 3587 3177
rect 3621 3143 3655 3177
rect 3689 3143 3723 3177
rect 3757 3143 3791 3177
rect 3825 3143 3859 3177
rect 3893 3143 3927 3177
rect 3961 3143 3995 3177
rect 4029 3143 4063 3177
rect 4097 3143 4131 3177
rect 4165 3143 4199 3177
rect 4233 3143 4267 3177
rect 4301 3143 4335 3177
rect 4369 3143 4403 3177
rect 4437 3143 4560 3177
rect -480 3120 4560 3143
rect 8000 4297 13040 4320
rect 8000 4263 8123 4297
rect 8157 4263 8191 4297
rect 8225 4263 8259 4297
rect 8293 4263 8327 4297
rect 8361 4263 8395 4297
rect 8429 4263 8463 4297
rect 8497 4263 8531 4297
rect 8565 4263 8599 4297
rect 8633 4263 8667 4297
rect 8701 4263 8735 4297
rect 8769 4263 8803 4297
rect 8837 4263 8871 4297
rect 8905 4263 8939 4297
rect 8973 4263 9007 4297
rect 9041 4263 9075 4297
rect 9109 4263 9143 4297
rect 9177 4263 9211 4297
rect 9245 4263 9279 4297
rect 9313 4263 9347 4297
rect 9381 4263 9415 4297
rect 9449 4263 9483 4297
rect 9517 4263 9551 4297
rect 9585 4263 9619 4297
rect 9653 4263 9687 4297
rect 9721 4263 9755 4297
rect 9789 4263 9823 4297
rect 9857 4263 9891 4297
rect 9925 4263 9959 4297
rect 9993 4263 10027 4297
rect 10061 4263 10095 4297
rect 10129 4263 10163 4297
rect 10197 4263 10231 4297
rect 10265 4263 10299 4297
rect 10333 4263 10367 4297
rect 10401 4263 10435 4297
rect 10469 4263 10503 4297
rect 10537 4263 10571 4297
rect 10605 4263 10639 4297
rect 10673 4263 10707 4297
rect 10741 4263 10775 4297
rect 10809 4263 10843 4297
rect 10877 4263 10911 4297
rect 10945 4263 10979 4297
rect 11013 4263 11047 4297
rect 11081 4263 11115 4297
rect 11149 4263 11183 4297
rect 11217 4263 11251 4297
rect 11285 4263 11319 4297
rect 11353 4263 11387 4297
rect 11421 4263 11455 4297
rect 11489 4263 11523 4297
rect 11557 4263 11591 4297
rect 11625 4263 11659 4297
rect 11693 4263 11727 4297
rect 11761 4263 11795 4297
rect 11829 4263 11863 4297
rect 11897 4263 11931 4297
rect 11965 4263 11999 4297
rect 12033 4263 12067 4297
rect 12101 4263 12135 4297
rect 12169 4263 12203 4297
rect 12237 4263 12271 4297
rect 12305 4263 12339 4297
rect 12373 4263 12407 4297
rect 12441 4263 12475 4297
rect 12509 4263 12543 4297
rect 12577 4263 12611 4297
rect 12645 4263 12679 4297
rect 12713 4263 12747 4297
rect 12781 4263 12815 4297
rect 12849 4263 12883 4297
rect 12917 4263 13040 4297
rect 8000 4240 13040 4263
rect 8000 4199 8080 4240
rect 8000 4165 8023 4199
rect 8057 4165 8080 4199
rect 8000 4131 8080 4165
rect 12960 4199 13040 4240
rect 12960 4165 12983 4199
rect 13017 4165 13040 4199
rect 8000 4097 8023 4131
rect 8057 4097 8080 4131
rect 8000 4063 8080 4097
rect 8000 4029 8023 4063
rect 8057 4029 8080 4063
rect 8000 3995 8080 4029
rect 8000 3961 8023 3995
rect 8057 3961 8080 3995
rect 8000 3927 8080 3961
rect 8000 3893 8023 3927
rect 8057 3893 8080 3927
rect 8000 3859 8080 3893
rect 8000 3825 8023 3859
rect 8057 3825 8080 3859
rect 8000 3791 8080 3825
rect 8000 3757 8023 3791
rect 8057 3757 8080 3791
rect 8000 3723 8080 3757
rect 8000 3689 8023 3723
rect 8057 3689 8080 3723
rect 8000 3655 8080 3689
rect 8000 3621 8023 3655
rect 8057 3621 8080 3655
rect 8000 3587 8080 3621
rect 8000 3553 8023 3587
rect 8057 3553 8080 3587
rect 8000 3519 8080 3553
rect 8000 3485 8023 3519
rect 8057 3485 8080 3519
rect 8000 3451 8080 3485
rect 8000 3417 8023 3451
rect 8057 3417 8080 3451
rect 8000 3383 8080 3417
rect 8000 3349 8023 3383
rect 8057 3349 8080 3383
rect 8000 3315 8080 3349
rect 8000 3281 8023 3315
rect 8057 3281 8080 3315
rect 8000 3200 8080 3281
rect 12960 4131 13040 4165
rect 12960 4097 12983 4131
rect 13017 4097 13040 4131
rect 12960 4063 13040 4097
rect 12960 4029 12983 4063
rect 13017 4029 13040 4063
rect 12960 3995 13040 4029
rect 12960 3961 12983 3995
rect 13017 3961 13040 3995
rect 12960 3927 13040 3961
rect 12960 3893 12983 3927
rect 13017 3893 13040 3927
rect 12960 3859 13040 3893
rect 12960 3825 12983 3859
rect 13017 3825 13040 3859
rect 12960 3791 13040 3825
rect 12960 3757 12983 3791
rect 13017 3757 13040 3791
rect 12960 3723 13040 3757
rect 12960 3689 12983 3723
rect 13017 3689 13040 3723
rect 12960 3655 13040 3689
rect 12960 3621 12983 3655
rect 13017 3621 13040 3655
rect 12960 3587 13040 3621
rect 12960 3553 12983 3587
rect 13017 3553 13040 3587
rect 12960 3519 13040 3553
rect 12960 3485 12983 3519
rect 13017 3485 13040 3519
rect 12960 3451 13040 3485
rect 12960 3417 12983 3451
rect 13017 3417 13040 3451
rect 12960 3383 13040 3417
rect 12960 3349 12983 3383
rect 13017 3349 13040 3383
rect 12960 3315 13040 3349
rect 12960 3281 12983 3315
rect 13017 3281 13040 3315
rect 12960 3200 13040 3281
rect 8000 3177 13040 3200
rect 8000 3143 8123 3177
rect 8157 3143 8191 3177
rect 8225 3143 8259 3177
rect 8293 3143 8327 3177
rect 8361 3143 8395 3177
rect 8429 3143 8463 3177
rect 8497 3143 8531 3177
rect 8565 3143 8599 3177
rect 8633 3143 8667 3177
rect 8701 3143 8735 3177
rect 8769 3143 8803 3177
rect 8837 3143 8871 3177
rect 8905 3143 8939 3177
rect 8973 3143 9007 3177
rect 9041 3143 9075 3177
rect 9109 3143 9143 3177
rect 9177 3143 9211 3177
rect 9245 3143 9279 3177
rect 9313 3143 9347 3177
rect 9381 3143 9415 3177
rect 9449 3143 9483 3177
rect 9517 3143 9551 3177
rect 9585 3143 9619 3177
rect 9653 3143 9687 3177
rect 9721 3143 9755 3177
rect 9789 3143 9823 3177
rect 9857 3143 9891 3177
rect 9925 3143 9959 3177
rect 9993 3143 10027 3177
rect 10061 3143 10095 3177
rect 10129 3143 10163 3177
rect 10197 3143 10231 3177
rect 10265 3143 10299 3177
rect 10333 3143 10367 3177
rect 10401 3143 10435 3177
rect 10469 3143 10503 3177
rect 10537 3143 10571 3177
rect 10605 3143 10639 3177
rect 10673 3143 10707 3177
rect 10741 3143 10775 3177
rect 10809 3143 10843 3177
rect 10877 3143 10911 3177
rect 10945 3143 10979 3177
rect 11013 3143 11047 3177
rect 11081 3143 11115 3177
rect 11149 3143 11183 3177
rect 11217 3143 11251 3177
rect 11285 3143 11319 3177
rect 11353 3143 11387 3177
rect 11421 3143 11455 3177
rect 11489 3143 11523 3177
rect 11557 3143 11591 3177
rect 11625 3143 11659 3177
rect 11693 3143 11727 3177
rect 11761 3143 11795 3177
rect 11829 3143 11863 3177
rect 11897 3143 11931 3177
rect 11965 3143 11999 3177
rect 12033 3143 12067 3177
rect 12101 3143 12135 3177
rect 12169 3143 12203 3177
rect 12237 3143 12271 3177
rect 12305 3143 12339 3177
rect 12373 3143 12407 3177
rect 12441 3143 12475 3177
rect 12509 3143 12543 3177
rect 12577 3143 12611 3177
rect 12645 3143 12679 3177
rect 12713 3143 12747 3177
rect 12781 3143 12815 3177
rect 12849 3143 12883 3177
rect 12917 3143 13040 3177
rect 8000 3120 13040 3143
rect -480 3017 4560 3040
rect -480 2983 -357 3017
rect -323 2983 -289 3017
rect -255 2983 -221 3017
rect -187 2983 -153 3017
rect -119 2983 -85 3017
rect -51 2983 -17 3017
rect 17 2983 51 3017
rect 85 2983 119 3017
rect 153 2983 187 3017
rect 221 2983 255 3017
rect 289 2983 323 3017
rect 357 2983 391 3017
rect 425 2983 459 3017
rect 493 2983 527 3017
rect 561 2983 595 3017
rect 629 2983 663 3017
rect 697 2983 731 3017
rect 765 2983 799 3017
rect 833 2983 867 3017
rect 901 2983 935 3017
rect 969 2983 1003 3017
rect 1037 2983 1071 3017
rect 1105 2983 1139 3017
rect 1173 2983 1207 3017
rect 1241 2983 1275 3017
rect 1309 2983 1343 3017
rect 1377 2983 1411 3017
rect 1445 2983 1479 3017
rect 1513 2983 1547 3017
rect 1581 2983 1615 3017
rect 1649 2983 1683 3017
rect 1717 2983 1751 3017
rect 1785 2983 1819 3017
rect 1853 2983 1887 3017
rect 1921 2983 1955 3017
rect 1989 2983 2023 3017
rect 2057 2983 2091 3017
rect 2125 2983 2159 3017
rect 2193 2983 2227 3017
rect 2261 2983 2295 3017
rect 2329 2983 2363 3017
rect 2397 2983 2431 3017
rect 2465 2983 2499 3017
rect 2533 2983 2567 3017
rect 2601 2983 2635 3017
rect 2669 2983 2703 3017
rect 2737 2983 2771 3017
rect 2805 2983 2839 3017
rect 2873 2983 2907 3017
rect 2941 2983 2975 3017
rect 3009 2983 3043 3017
rect 3077 2983 3111 3017
rect 3145 2983 3179 3017
rect 3213 2983 3247 3017
rect 3281 2983 3315 3017
rect 3349 2983 3383 3017
rect 3417 2983 3451 3017
rect 3485 2983 3519 3017
rect 3553 2983 3587 3017
rect 3621 2983 3655 3017
rect 3689 2983 3723 3017
rect 3757 2983 3791 3017
rect 3825 2983 3859 3017
rect 3893 2983 3927 3017
rect 3961 2983 3995 3017
rect 4029 2983 4063 3017
rect 4097 2983 4131 3017
rect 4165 2983 4199 3017
rect 4233 2983 4267 3017
rect 4301 2983 4335 3017
rect 4369 2983 4403 3017
rect 4437 2983 4560 3017
rect -480 2960 4560 2983
rect -480 2879 -400 2960
rect -480 2845 -457 2879
rect -423 2845 -400 2879
rect -480 2811 -400 2845
rect -480 2777 -457 2811
rect -423 2777 -400 2811
rect -480 2743 -400 2777
rect -480 2709 -457 2743
rect -423 2709 -400 2743
rect -480 2675 -400 2709
rect -480 2641 -457 2675
rect -423 2641 -400 2675
rect -480 2607 -400 2641
rect -480 2573 -457 2607
rect -423 2573 -400 2607
rect -480 2539 -400 2573
rect -480 2505 -457 2539
rect -423 2505 -400 2539
rect -480 2471 -400 2505
rect -480 2437 -457 2471
rect -423 2437 -400 2471
rect -480 2403 -400 2437
rect -480 2369 -457 2403
rect -423 2369 -400 2403
rect -480 2335 -400 2369
rect -480 2301 -457 2335
rect -423 2301 -400 2335
rect -480 2267 -400 2301
rect -480 2233 -457 2267
rect -423 2233 -400 2267
rect -480 2199 -400 2233
rect -480 2165 -457 2199
rect -423 2165 -400 2199
rect -480 2131 -400 2165
rect -480 2097 -457 2131
rect -423 2097 -400 2131
rect -480 2063 -400 2097
rect -480 2029 -457 2063
rect -423 2029 -400 2063
rect -480 1995 -400 2029
rect 4480 2879 4560 2960
rect 4480 2845 4503 2879
rect 4537 2845 4560 2879
rect 4480 2811 4560 2845
rect 4480 2777 4503 2811
rect 4537 2777 4560 2811
rect 4480 2743 4560 2777
rect 4480 2709 4503 2743
rect 4537 2709 4560 2743
rect 4480 2675 4560 2709
rect 4480 2641 4503 2675
rect 4537 2641 4560 2675
rect 4480 2607 4560 2641
rect 4480 2573 4503 2607
rect 4537 2573 4560 2607
rect 4480 2539 4560 2573
rect 4480 2505 4503 2539
rect 4537 2505 4560 2539
rect 4480 2471 4560 2505
rect 4480 2437 4503 2471
rect 4537 2437 4560 2471
rect 4480 2403 4560 2437
rect 4480 2369 4503 2403
rect 4537 2369 4560 2403
rect 4480 2335 4560 2369
rect 4480 2301 4503 2335
rect 4537 2301 4560 2335
rect 4480 2267 4560 2301
rect 4480 2233 4503 2267
rect 4537 2233 4560 2267
rect 4480 2199 4560 2233
rect 4480 2165 4503 2199
rect 4537 2165 4560 2199
rect 4480 2131 4560 2165
rect 4480 2097 4503 2131
rect 4537 2097 4560 2131
rect 4480 2063 4560 2097
rect 4480 2029 4503 2063
rect 4537 2029 4560 2063
rect -480 1961 -457 1995
rect -423 1961 -400 1995
rect -480 1920 -400 1961
rect 4480 1995 4560 2029
rect 4480 1961 4503 1995
rect 4537 1961 4560 1995
rect 4480 1920 4560 1961
rect -480 1897 4560 1920
rect -480 1863 -357 1897
rect -323 1863 -289 1897
rect -255 1863 -221 1897
rect -187 1863 -153 1897
rect -119 1863 -85 1897
rect -51 1863 -17 1897
rect 17 1863 51 1897
rect 85 1863 119 1897
rect 153 1863 187 1897
rect 221 1863 255 1897
rect 289 1863 323 1897
rect 357 1863 391 1897
rect 425 1863 459 1897
rect 493 1863 527 1897
rect 561 1863 595 1897
rect 629 1863 663 1897
rect 697 1863 731 1897
rect 765 1863 799 1897
rect 833 1863 867 1897
rect 901 1863 935 1897
rect 969 1863 1003 1897
rect 1037 1863 1071 1897
rect 1105 1863 1139 1897
rect 1173 1863 1207 1897
rect 1241 1863 1275 1897
rect 1309 1863 1343 1897
rect 1377 1863 1411 1897
rect 1445 1863 1479 1897
rect 1513 1863 1547 1897
rect 1581 1863 1615 1897
rect 1649 1863 1683 1897
rect 1717 1863 1751 1897
rect 1785 1863 1819 1897
rect 1853 1863 1887 1897
rect 1921 1863 1955 1897
rect 1989 1863 2023 1897
rect 2057 1863 2091 1897
rect 2125 1863 2159 1897
rect 2193 1863 2227 1897
rect 2261 1863 2295 1897
rect 2329 1863 2363 1897
rect 2397 1863 2431 1897
rect 2465 1863 2499 1897
rect 2533 1863 2567 1897
rect 2601 1863 2635 1897
rect 2669 1863 2703 1897
rect 2737 1863 2771 1897
rect 2805 1863 2839 1897
rect 2873 1863 2907 1897
rect 2941 1863 2975 1897
rect 3009 1863 3043 1897
rect 3077 1863 3111 1897
rect 3145 1863 3179 1897
rect 3213 1863 3247 1897
rect 3281 1863 3315 1897
rect 3349 1863 3383 1897
rect 3417 1863 3451 1897
rect 3485 1863 3519 1897
rect 3553 1863 3587 1897
rect 3621 1863 3655 1897
rect 3689 1863 3723 1897
rect 3757 1863 3791 1897
rect 3825 1863 3859 1897
rect 3893 1863 3927 1897
rect 3961 1863 3995 1897
rect 4029 1863 4063 1897
rect 4097 1863 4131 1897
rect 4165 1863 4199 1897
rect 4233 1863 4267 1897
rect 4301 1863 4335 1897
rect 4369 1863 4403 1897
rect 4437 1863 4560 1897
rect -480 1840 4560 1863
rect 8000 3017 13040 3040
rect 8000 2983 8123 3017
rect 8157 2983 8191 3017
rect 8225 2983 8259 3017
rect 8293 2983 8327 3017
rect 8361 2983 8395 3017
rect 8429 2983 8463 3017
rect 8497 2983 8531 3017
rect 8565 2983 8599 3017
rect 8633 2983 8667 3017
rect 8701 2983 8735 3017
rect 8769 2983 8803 3017
rect 8837 2983 8871 3017
rect 8905 2983 8939 3017
rect 8973 2983 9007 3017
rect 9041 2983 9075 3017
rect 9109 2983 9143 3017
rect 9177 2983 9211 3017
rect 9245 2983 9279 3017
rect 9313 2983 9347 3017
rect 9381 2983 9415 3017
rect 9449 2983 9483 3017
rect 9517 2983 9551 3017
rect 9585 2983 9619 3017
rect 9653 2983 9687 3017
rect 9721 2983 9755 3017
rect 9789 2983 9823 3017
rect 9857 2983 9891 3017
rect 9925 2983 9959 3017
rect 9993 2983 10027 3017
rect 10061 2983 10095 3017
rect 10129 2983 10163 3017
rect 10197 2983 10231 3017
rect 10265 2983 10299 3017
rect 10333 2983 10367 3017
rect 10401 2983 10435 3017
rect 10469 2983 10503 3017
rect 10537 2983 10571 3017
rect 10605 2983 10639 3017
rect 10673 2983 10707 3017
rect 10741 2983 10775 3017
rect 10809 2983 10843 3017
rect 10877 2983 10911 3017
rect 10945 2983 10979 3017
rect 11013 2983 11047 3017
rect 11081 2983 11115 3017
rect 11149 2983 11183 3017
rect 11217 2983 11251 3017
rect 11285 2983 11319 3017
rect 11353 2983 11387 3017
rect 11421 2983 11455 3017
rect 11489 2983 11523 3017
rect 11557 2983 11591 3017
rect 11625 2983 11659 3017
rect 11693 2983 11727 3017
rect 11761 2983 11795 3017
rect 11829 2983 11863 3017
rect 11897 2983 11931 3017
rect 11965 2983 11999 3017
rect 12033 2983 12067 3017
rect 12101 2983 12135 3017
rect 12169 2983 12203 3017
rect 12237 2983 12271 3017
rect 12305 2983 12339 3017
rect 12373 2983 12407 3017
rect 12441 2983 12475 3017
rect 12509 2983 12543 3017
rect 12577 2983 12611 3017
rect 12645 2983 12679 3017
rect 12713 2983 12747 3017
rect 12781 2983 12815 3017
rect 12849 2983 12883 3017
rect 12917 2983 13040 3017
rect 8000 2960 13040 2983
rect 8000 2879 8080 2960
rect 8000 2845 8023 2879
rect 8057 2845 8080 2879
rect 8000 2811 8080 2845
rect 8000 2777 8023 2811
rect 8057 2777 8080 2811
rect 8000 2743 8080 2777
rect 8000 2709 8023 2743
rect 8057 2709 8080 2743
rect 8000 2675 8080 2709
rect 8000 2641 8023 2675
rect 8057 2641 8080 2675
rect 8000 2607 8080 2641
rect 8000 2573 8023 2607
rect 8057 2573 8080 2607
rect 8000 2539 8080 2573
rect 8000 2505 8023 2539
rect 8057 2505 8080 2539
rect 8000 2471 8080 2505
rect 8000 2437 8023 2471
rect 8057 2437 8080 2471
rect 8000 2403 8080 2437
rect 8000 2369 8023 2403
rect 8057 2369 8080 2403
rect 8000 2335 8080 2369
rect 8000 2301 8023 2335
rect 8057 2301 8080 2335
rect 8000 2267 8080 2301
rect 8000 2233 8023 2267
rect 8057 2233 8080 2267
rect 8000 2199 8080 2233
rect 8000 2165 8023 2199
rect 8057 2165 8080 2199
rect 8000 2131 8080 2165
rect 8000 2097 8023 2131
rect 8057 2097 8080 2131
rect 8000 2063 8080 2097
rect 8000 2029 8023 2063
rect 8057 2029 8080 2063
rect 8000 1995 8080 2029
rect 12960 2879 13040 2960
rect 12960 2845 12983 2879
rect 13017 2845 13040 2879
rect 12960 2811 13040 2845
rect 12960 2777 12983 2811
rect 13017 2777 13040 2811
rect 12960 2743 13040 2777
rect 12960 2709 12983 2743
rect 13017 2709 13040 2743
rect 12960 2675 13040 2709
rect 12960 2641 12983 2675
rect 13017 2641 13040 2675
rect 12960 2607 13040 2641
rect 12960 2573 12983 2607
rect 13017 2573 13040 2607
rect 12960 2539 13040 2573
rect 12960 2505 12983 2539
rect 13017 2505 13040 2539
rect 12960 2471 13040 2505
rect 12960 2437 12983 2471
rect 13017 2437 13040 2471
rect 12960 2403 13040 2437
rect 12960 2369 12983 2403
rect 13017 2369 13040 2403
rect 12960 2335 13040 2369
rect 12960 2301 12983 2335
rect 13017 2301 13040 2335
rect 12960 2267 13040 2301
rect 12960 2233 12983 2267
rect 13017 2233 13040 2267
rect 12960 2199 13040 2233
rect 12960 2165 12983 2199
rect 13017 2165 13040 2199
rect 12960 2131 13040 2165
rect 12960 2097 12983 2131
rect 13017 2097 13040 2131
rect 12960 2063 13040 2097
rect 12960 2029 12983 2063
rect 13017 2029 13040 2063
rect 8000 1961 8023 1995
rect 8057 1961 8080 1995
rect 8000 1920 8080 1961
rect 12960 1995 13040 2029
rect 12960 1961 12983 1995
rect 13017 1961 13040 1995
rect 12960 1920 13040 1961
rect 8000 1897 13040 1920
rect 8000 1863 8123 1897
rect 8157 1863 8191 1897
rect 8225 1863 8259 1897
rect 8293 1863 8327 1897
rect 8361 1863 8395 1897
rect 8429 1863 8463 1897
rect 8497 1863 8531 1897
rect 8565 1863 8599 1897
rect 8633 1863 8667 1897
rect 8701 1863 8735 1897
rect 8769 1863 8803 1897
rect 8837 1863 8871 1897
rect 8905 1863 8939 1897
rect 8973 1863 9007 1897
rect 9041 1863 9075 1897
rect 9109 1863 9143 1897
rect 9177 1863 9211 1897
rect 9245 1863 9279 1897
rect 9313 1863 9347 1897
rect 9381 1863 9415 1897
rect 9449 1863 9483 1897
rect 9517 1863 9551 1897
rect 9585 1863 9619 1897
rect 9653 1863 9687 1897
rect 9721 1863 9755 1897
rect 9789 1863 9823 1897
rect 9857 1863 9891 1897
rect 9925 1863 9959 1897
rect 9993 1863 10027 1897
rect 10061 1863 10095 1897
rect 10129 1863 10163 1897
rect 10197 1863 10231 1897
rect 10265 1863 10299 1897
rect 10333 1863 10367 1897
rect 10401 1863 10435 1897
rect 10469 1863 10503 1897
rect 10537 1863 10571 1897
rect 10605 1863 10639 1897
rect 10673 1863 10707 1897
rect 10741 1863 10775 1897
rect 10809 1863 10843 1897
rect 10877 1863 10911 1897
rect 10945 1863 10979 1897
rect 11013 1863 11047 1897
rect 11081 1863 11115 1897
rect 11149 1863 11183 1897
rect 11217 1863 11251 1897
rect 11285 1863 11319 1897
rect 11353 1863 11387 1897
rect 11421 1863 11455 1897
rect 11489 1863 11523 1897
rect 11557 1863 11591 1897
rect 11625 1863 11659 1897
rect 11693 1863 11727 1897
rect 11761 1863 11795 1897
rect 11829 1863 11863 1897
rect 11897 1863 11931 1897
rect 11965 1863 11999 1897
rect 12033 1863 12067 1897
rect 12101 1863 12135 1897
rect 12169 1863 12203 1897
rect 12237 1863 12271 1897
rect 12305 1863 12339 1897
rect 12373 1863 12407 1897
rect 12441 1863 12475 1897
rect 12509 1863 12543 1897
rect 12577 1863 12611 1897
rect 12645 1863 12679 1897
rect 12713 1863 12747 1897
rect 12781 1863 12815 1897
rect 12849 1863 12883 1897
rect 12917 1863 13040 1897
rect 8000 1840 13040 1863
rect -480 1737 4560 1760
rect -480 1703 -357 1737
rect -323 1703 -289 1737
rect -255 1703 -221 1737
rect -187 1703 -153 1737
rect -119 1703 -85 1737
rect -51 1703 -17 1737
rect 17 1703 51 1737
rect 85 1703 119 1737
rect 153 1703 187 1737
rect 221 1703 255 1737
rect 289 1703 323 1737
rect 357 1703 391 1737
rect 425 1703 459 1737
rect 493 1703 527 1737
rect 561 1703 595 1737
rect 629 1703 663 1737
rect 697 1703 731 1737
rect 765 1703 799 1737
rect 833 1703 867 1737
rect 901 1703 935 1737
rect 969 1703 1003 1737
rect 1037 1703 1071 1737
rect 1105 1703 1139 1737
rect 1173 1703 1207 1737
rect 1241 1703 1275 1737
rect 1309 1703 1343 1737
rect 1377 1703 1411 1737
rect 1445 1703 1479 1737
rect 1513 1703 1547 1737
rect 1581 1703 1615 1737
rect 1649 1703 1683 1737
rect 1717 1703 1751 1737
rect 1785 1703 1819 1737
rect 1853 1703 1887 1737
rect 1921 1703 1955 1737
rect 1989 1703 2023 1737
rect 2057 1703 2091 1737
rect 2125 1703 2159 1737
rect 2193 1703 2227 1737
rect 2261 1703 2295 1737
rect 2329 1703 2363 1737
rect 2397 1703 2431 1737
rect 2465 1703 2499 1737
rect 2533 1703 2567 1737
rect 2601 1703 2635 1737
rect 2669 1703 2703 1737
rect 2737 1703 2771 1737
rect 2805 1703 2839 1737
rect 2873 1703 2907 1737
rect 2941 1703 2975 1737
rect 3009 1703 3043 1737
rect 3077 1703 3111 1737
rect 3145 1703 3179 1737
rect 3213 1703 3247 1737
rect 3281 1703 3315 1737
rect 3349 1703 3383 1737
rect 3417 1703 3451 1737
rect 3485 1703 3519 1737
rect 3553 1703 3587 1737
rect 3621 1703 3655 1737
rect 3689 1703 3723 1737
rect 3757 1703 3791 1737
rect 3825 1703 3859 1737
rect 3893 1703 3927 1737
rect 3961 1703 3995 1737
rect 4029 1703 4063 1737
rect 4097 1703 4131 1737
rect 4165 1703 4199 1737
rect 4233 1703 4267 1737
rect 4301 1703 4335 1737
rect 4369 1703 4403 1737
rect 4437 1703 4560 1737
rect -480 1680 4560 1703
rect -480 1639 -400 1680
rect -480 1605 -457 1639
rect -423 1605 -400 1639
rect -480 1571 -400 1605
rect 4480 1639 4560 1680
rect 4480 1605 4503 1639
rect 4537 1605 4560 1639
rect -480 1537 -457 1571
rect -423 1537 -400 1571
rect -480 1503 -400 1537
rect -480 1469 -457 1503
rect -423 1469 -400 1503
rect -480 1435 -400 1469
rect -480 1401 -457 1435
rect -423 1401 -400 1435
rect -480 1367 -400 1401
rect -480 1333 -457 1367
rect -423 1333 -400 1367
rect -480 1299 -400 1333
rect -480 1265 -457 1299
rect -423 1265 -400 1299
rect -480 1231 -400 1265
rect -480 1197 -457 1231
rect -423 1197 -400 1231
rect -480 1163 -400 1197
rect -480 1129 -457 1163
rect -423 1129 -400 1163
rect -480 1095 -400 1129
rect -480 1061 -457 1095
rect -423 1061 -400 1095
rect -480 1027 -400 1061
rect -480 993 -457 1027
rect -423 993 -400 1027
rect -480 959 -400 993
rect -480 925 -457 959
rect -423 925 -400 959
rect -480 891 -400 925
rect -480 857 -457 891
rect -423 857 -400 891
rect -480 823 -400 857
rect -480 789 -457 823
rect -423 789 -400 823
rect -480 755 -400 789
rect -480 721 -457 755
rect -423 721 -400 755
rect -480 640 -400 721
rect 4480 1571 4560 1605
rect 4480 1537 4503 1571
rect 4537 1537 4560 1571
rect 4480 1503 4560 1537
rect 4480 1469 4503 1503
rect 4537 1469 4560 1503
rect 4480 1435 4560 1469
rect 4480 1401 4503 1435
rect 4537 1401 4560 1435
rect 4480 1367 4560 1401
rect 4480 1333 4503 1367
rect 4537 1333 4560 1367
rect 4480 1299 4560 1333
rect 4480 1265 4503 1299
rect 4537 1265 4560 1299
rect 4480 1231 4560 1265
rect 4480 1197 4503 1231
rect 4537 1197 4560 1231
rect 4480 1163 4560 1197
rect 4480 1129 4503 1163
rect 4537 1129 4560 1163
rect 4480 1095 4560 1129
rect 4480 1061 4503 1095
rect 4537 1061 4560 1095
rect 4480 1027 4560 1061
rect 4480 993 4503 1027
rect 4537 993 4560 1027
rect 4480 959 4560 993
rect 4480 925 4503 959
rect 4537 925 4560 959
rect 4480 891 4560 925
rect 4480 857 4503 891
rect 4537 857 4560 891
rect 4480 823 4560 857
rect 4480 789 4503 823
rect 4537 789 4560 823
rect 4480 755 4560 789
rect 4480 721 4503 755
rect 4537 721 4560 755
rect 4480 640 4560 721
rect -480 617 4560 640
rect -480 583 -357 617
rect -323 583 -289 617
rect -255 583 -221 617
rect -187 583 -153 617
rect -119 583 -85 617
rect -51 583 -17 617
rect 17 583 51 617
rect 85 583 119 617
rect 153 583 187 617
rect 221 583 255 617
rect 289 583 323 617
rect 357 583 391 617
rect 425 583 459 617
rect 493 583 527 617
rect 561 583 595 617
rect 629 583 663 617
rect 697 583 731 617
rect 765 583 799 617
rect 833 583 867 617
rect 901 583 935 617
rect 969 583 1003 617
rect 1037 583 1071 617
rect 1105 583 1139 617
rect 1173 583 1207 617
rect 1241 583 1275 617
rect 1309 583 1343 617
rect 1377 583 1411 617
rect 1445 583 1479 617
rect 1513 583 1547 617
rect 1581 583 1615 617
rect 1649 583 1683 617
rect 1717 583 1751 617
rect 1785 583 1819 617
rect 1853 583 1887 617
rect 1921 583 1955 617
rect 1989 583 2023 617
rect 2057 583 2091 617
rect 2125 583 2159 617
rect 2193 583 2227 617
rect 2261 583 2295 617
rect 2329 583 2363 617
rect 2397 583 2431 617
rect 2465 583 2499 617
rect 2533 583 2567 617
rect 2601 583 2635 617
rect 2669 583 2703 617
rect 2737 583 2771 617
rect 2805 583 2839 617
rect 2873 583 2907 617
rect 2941 583 2975 617
rect 3009 583 3043 617
rect 3077 583 3111 617
rect 3145 583 3179 617
rect 3213 583 3247 617
rect 3281 583 3315 617
rect 3349 583 3383 617
rect 3417 583 3451 617
rect 3485 583 3519 617
rect 3553 583 3587 617
rect 3621 583 3655 617
rect 3689 583 3723 617
rect 3757 583 3791 617
rect 3825 583 3859 617
rect 3893 583 3927 617
rect 3961 583 3995 617
rect 4029 583 4063 617
rect 4097 583 4131 617
rect 4165 583 4199 617
rect 4233 583 4267 617
rect 4301 583 4335 617
rect 4369 583 4403 617
rect 4437 583 4560 617
rect -480 560 4560 583
rect 8000 1737 13040 1760
rect 8000 1703 8123 1737
rect 8157 1703 8191 1737
rect 8225 1703 8259 1737
rect 8293 1703 8327 1737
rect 8361 1703 8395 1737
rect 8429 1703 8463 1737
rect 8497 1703 8531 1737
rect 8565 1703 8599 1737
rect 8633 1703 8667 1737
rect 8701 1703 8735 1737
rect 8769 1703 8803 1737
rect 8837 1703 8871 1737
rect 8905 1703 8939 1737
rect 8973 1703 9007 1737
rect 9041 1703 9075 1737
rect 9109 1703 9143 1737
rect 9177 1703 9211 1737
rect 9245 1703 9279 1737
rect 9313 1703 9347 1737
rect 9381 1703 9415 1737
rect 9449 1703 9483 1737
rect 9517 1703 9551 1737
rect 9585 1703 9619 1737
rect 9653 1703 9687 1737
rect 9721 1703 9755 1737
rect 9789 1703 9823 1737
rect 9857 1703 9891 1737
rect 9925 1703 9959 1737
rect 9993 1703 10027 1737
rect 10061 1703 10095 1737
rect 10129 1703 10163 1737
rect 10197 1703 10231 1737
rect 10265 1703 10299 1737
rect 10333 1703 10367 1737
rect 10401 1703 10435 1737
rect 10469 1703 10503 1737
rect 10537 1703 10571 1737
rect 10605 1703 10639 1737
rect 10673 1703 10707 1737
rect 10741 1703 10775 1737
rect 10809 1703 10843 1737
rect 10877 1703 10911 1737
rect 10945 1703 10979 1737
rect 11013 1703 11047 1737
rect 11081 1703 11115 1737
rect 11149 1703 11183 1737
rect 11217 1703 11251 1737
rect 11285 1703 11319 1737
rect 11353 1703 11387 1737
rect 11421 1703 11455 1737
rect 11489 1703 11523 1737
rect 11557 1703 11591 1737
rect 11625 1703 11659 1737
rect 11693 1703 11727 1737
rect 11761 1703 11795 1737
rect 11829 1703 11863 1737
rect 11897 1703 11931 1737
rect 11965 1703 11999 1737
rect 12033 1703 12067 1737
rect 12101 1703 12135 1737
rect 12169 1703 12203 1737
rect 12237 1703 12271 1737
rect 12305 1703 12339 1737
rect 12373 1703 12407 1737
rect 12441 1703 12475 1737
rect 12509 1703 12543 1737
rect 12577 1703 12611 1737
rect 12645 1703 12679 1737
rect 12713 1703 12747 1737
rect 12781 1703 12815 1737
rect 12849 1703 12883 1737
rect 12917 1703 13040 1737
rect 8000 1680 13040 1703
rect 8000 1639 8080 1680
rect 8000 1605 8023 1639
rect 8057 1605 8080 1639
rect 8000 1571 8080 1605
rect 12960 1639 13040 1680
rect 12960 1605 12983 1639
rect 13017 1605 13040 1639
rect 8000 1537 8023 1571
rect 8057 1537 8080 1571
rect 8000 1503 8080 1537
rect 8000 1469 8023 1503
rect 8057 1469 8080 1503
rect 8000 1435 8080 1469
rect 8000 1401 8023 1435
rect 8057 1401 8080 1435
rect 8000 1367 8080 1401
rect 8000 1333 8023 1367
rect 8057 1333 8080 1367
rect 8000 1299 8080 1333
rect 8000 1265 8023 1299
rect 8057 1265 8080 1299
rect 8000 1231 8080 1265
rect 8000 1197 8023 1231
rect 8057 1197 8080 1231
rect 8000 1163 8080 1197
rect 8000 1129 8023 1163
rect 8057 1129 8080 1163
rect 8000 1095 8080 1129
rect 8000 1061 8023 1095
rect 8057 1061 8080 1095
rect 8000 1027 8080 1061
rect 8000 993 8023 1027
rect 8057 993 8080 1027
rect 8000 959 8080 993
rect 8000 925 8023 959
rect 8057 925 8080 959
rect 8000 891 8080 925
rect 8000 857 8023 891
rect 8057 857 8080 891
rect 8000 823 8080 857
rect 8000 789 8023 823
rect 8057 789 8080 823
rect 8000 755 8080 789
rect 8000 721 8023 755
rect 8057 721 8080 755
rect 8000 640 8080 721
rect 12960 1571 13040 1605
rect 12960 1537 12983 1571
rect 13017 1537 13040 1571
rect 12960 1503 13040 1537
rect 12960 1469 12983 1503
rect 13017 1469 13040 1503
rect 12960 1435 13040 1469
rect 12960 1401 12983 1435
rect 13017 1401 13040 1435
rect 12960 1367 13040 1401
rect 12960 1333 12983 1367
rect 13017 1333 13040 1367
rect 12960 1299 13040 1333
rect 12960 1265 12983 1299
rect 13017 1265 13040 1299
rect 12960 1231 13040 1265
rect 12960 1197 12983 1231
rect 13017 1197 13040 1231
rect 12960 1163 13040 1197
rect 12960 1129 12983 1163
rect 13017 1129 13040 1163
rect 12960 1095 13040 1129
rect 12960 1061 12983 1095
rect 13017 1061 13040 1095
rect 12960 1027 13040 1061
rect 12960 993 12983 1027
rect 13017 993 13040 1027
rect 12960 959 13040 993
rect 12960 925 12983 959
rect 13017 925 13040 959
rect 12960 891 13040 925
rect 12960 857 12983 891
rect 13017 857 13040 891
rect 12960 823 13040 857
rect 12960 789 12983 823
rect 13017 789 13040 823
rect 12960 755 13040 789
rect 12960 721 12983 755
rect 13017 721 13040 755
rect 12960 640 13040 721
rect 8000 617 13040 640
rect 8000 583 8123 617
rect 8157 583 8191 617
rect 8225 583 8259 617
rect 8293 583 8327 617
rect 8361 583 8395 617
rect 8429 583 8463 617
rect 8497 583 8531 617
rect 8565 583 8599 617
rect 8633 583 8667 617
rect 8701 583 8735 617
rect 8769 583 8803 617
rect 8837 583 8871 617
rect 8905 583 8939 617
rect 8973 583 9007 617
rect 9041 583 9075 617
rect 9109 583 9143 617
rect 9177 583 9211 617
rect 9245 583 9279 617
rect 9313 583 9347 617
rect 9381 583 9415 617
rect 9449 583 9483 617
rect 9517 583 9551 617
rect 9585 583 9619 617
rect 9653 583 9687 617
rect 9721 583 9755 617
rect 9789 583 9823 617
rect 9857 583 9891 617
rect 9925 583 9959 617
rect 9993 583 10027 617
rect 10061 583 10095 617
rect 10129 583 10163 617
rect 10197 583 10231 617
rect 10265 583 10299 617
rect 10333 583 10367 617
rect 10401 583 10435 617
rect 10469 583 10503 617
rect 10537 583 10571 617
rect 10605 583 10639 617
rect 10673 583 10707 617
rect 10741 583 10775 617
rect 10809 583 10843 617
rect 10877 583 10911 617
rect 10945 583 10979 617
rect 11013 583 11047 617
rect 11081 583 11115 617
rect 11149 583 11183 617
rect 11217 583 11251 617
rect 11285 583 11319 617
rect 11353 583 11387 617
rect 11421 583 11455 617
rect 11489 583 11523 617
rect 11557 583 11591 617
rect 11625 583 11659 617
rect 11693 583 11727 617
rect 11761 583 11795 617
rect 11829 583 11863 617
rect 11897 583 11931 617
rect 11965 583 11999 617
rect 12033 583 12067 617
rect 12101 583 12135 617
rect 12169 583 12203 617
rect 12237 583 12271 617
rect 12305 583 12339 617
rect 12373 583 12407 617
rect 12441 583 12475 617
rect 12509 583 12543 617
rect 12577 583 12611 617
rect 12645 583 12679 617
rect 12713 583 12747 617
rect 12781 583 12815 617
rect 12849 583 12883 617
rect 12917 583 13040 617
rect 8000 560 13040 583
rect -480 457 4560 480
rect -480 423 -357 457
rect -323 423 -289 457
rect -255 423 -221 457
rect -187 423 -153 457
rect -119 423 -85 457
rect -51 423 -17 457
rect 17 423 51 457
rect 85 423 119 457
rect 153 423 187 457
rect 221 423 255 457
rect 289 423 323 457
rect 357 423 391 457
rect 425 423 459 457
rect 493 423 527 457
rect 561 423 595 457
rect 629 423 663 457
rect 697 423 731 457
rect 765 423 799 457
rect 833 423 867 457
rect 901 423 935 457
rect 969 423 1003 457
rect 1037 423 1071 457
rect 1105 423 1139 457
rect 1173 423 1207 457
rect 1241 423 1275 457
rect 1309 423 1343 457
rect 1377 423 1411 457
rect 1445 423 1479 457
rect 1513 423 1547 457
rect 1581 423 1615 457
rect 1649 423 1683 457
rect 1717 423 1751 457
rect 1785 423 1819 457
rect 1853 423 1887 457
rect 1921 423 1955 457
rect 1989 423 2023 457
rect 2057 423 2091 457
rect 2125 423 2159 457
rect 2193 423 2227 457
rect 2261 423 2295 457
rect 2329 423 2363 457
rect 2397 423 2431 457
rect 2465 423 2499 457
rect 2533 423 2567 457
rect 2601 423 2635 457
rect 2669 423 2703 457
rect 2737 423 2771 457
rect 2805 423 2839 457
rect 2873 423 2907 457
rect 2941 423 2975 457
rect 3009 423 3043 457
rect 3077 423 3111 457
rect 3145 423 3179 457
rect 3213 423 3247 457
rect 3281 423 3315 457
rect 3349 423 3383 457
rect 3417 423 3451 457
rect 3485 423 3519 457
rect 3553 423 3587 457
rect 3621 423 3655 457
rect 3689 423 3723 457
rect 3757 423 3791 457
rect 3825 423 3859 457
rect 3893 423 3927 457
rect 3961 423 3995 457
rect 4029 423 4063 457
rect 4097 423 4131 457
rect 4165 423 4199 457
rect 4233 423 4267 457
rect 4301 423 4335 457
rect 4369 423 4403 457
rect 4437 423 4560 457
rect -480 400 4560 423
rect -480 319 -400 400
rect -480 285 -457 319
rect -423 285 -400 319
rect -480 251 -400 285
rect -480 217 -457 251
rect -423 217 -400 251
rect -480 183 -400 217
rect -480 149 -457 183
rect -423 149 -400 183
rect -480 115 -400 149
rect -480 81 -457 115
rect -423 81 -400 115
rect -480 47 -400 81
rect -480 13 -457 47
rect -423 13 -400 47
rect -480 -21 -400 13
rect -480 -55 -457 -21
rect -423 -55 -400 -21
rect -480 -89 -400 -55
rect -480 -123 -457 -89
rect -423 -123 -400 -89
rect -480 -157 -400 -123
rect -480 -191 -457 -157
rect -423 -191 -400 -157
rect -480 -225 -400 -191
rect -480 -259 -457 -225
rect -423 -259 -400 -225
rect -480 -293 -400 -259
rect -480 -327 -457 -293
rect -423 -327 -400 -293
rect -480 -361 -400 -327
rect -480 -395 -457 -361
rect -423 -395 -400 -361
rect -480 -429 -400 -395
rect -480 -463 -457 -429
rect -423 -463 -400 -429
rect -480 -497 -400 -463
rect -480 -531 -457 -497
rect -423 -531 -400 -497
rect -480 -565 -400 -531
rect 4480 319 4560 400
rect 4480 285 4503 319
rect 4537 285 4560 319
rect 4480 251 4560 285
rect 4480 217 4503 251
rect 4537 217 4560 251
rect 4480 183 4560 217
rect 4480 149 4503 183
rect 4537 149 4560 183
rect 4480 115 4560 149
rect 4480 81 4503 115
rect 4537 81 4560 115
rect 4480 47 4560 81
rect 4480 13 4503 47
rect 4537 13 4560 47
rect 4480 -21 4560 13
rect 4480 -55 4503 -21
rect 4537 -55 4560 -21
rect 4480 -89 4560 -55
rect 4480 -123 4503 -89
rect 4537 -123 4560 -89
rect 4480 -157 4560 -123
rect 4480 -191 4503 -157
rect 4537 -191 4560 -157
rect 4480 -225 4560 -191
rect 4480 -259 4503 -225
rect 4537 -259 4560 -225
rect 4480 -293 4560 -259
rect 4480 -327 4503 -293
rect 4537 -327 4560 -293
rect 4480 -361 4560 -327
rect 4480 -395 4503 -361
rect 4537 -395 4560 -361
rect 4480 -429 4560 -395
rect 4480 -463 4503 -429
rect 4537 -463 4560 -429
rect 4480 -497 4560 -463
rect 4480 -531 4503 -497
rect 4537 -531 4560 -497
rect -480 -599 -457 -565
rect -423 -599 -400 -565
rect -480 -640 -400 -599
rect 4480 -565 4560 -531
rect 4480 -599 4503 -565
rect 4537 -599 4560 -565
rect 4480 -640 4560 -599
rect -480 -663 4560 -640
rect -480 -697 -357 -663
rect -323 -697 -289 -663
rect -255 -697 -221 -663
rect -187 -697 -153 -663
rect -119 -697 -85 -663
rect -51 -697 -17 -663
rect 17 -697 51 -663
rect 85 -697 119 -663
rect 153 -697 187 -663
rect 221 -697 255 -663
rect 289 -697 323 -663
rect 357 -697 391 -663
rect 425 -697 459 -663
rect 493 -697 527 -663
rect 561 -697 595 -663
rect 629 -697 663 -663
rect 697 -697 731 -663
rect 765 -697 799 -663
rect 833 -697 867 -663
rect 901 -697 935 -663
rect 969 -697 1003 -663
rect 1037 -697 1071 -663
rect 1105 -697 1139 -663
rect 1173 -697 1207 -663
rect 1241 -697 1275 -663
rect 1309 -697 1343 -663
rect 1377 -697 1411 -663
rect 1445 -697 1479 -663
rect 1513 -697 1547 -663
rect 1581 -697 1615 -663
rect 1649 -697 1683 -663
rect 1717 -697 1751 -663
rect 1785 -697 1819 -663
rect 1853 -697 1887 -663
rect 1921 -697 1955 -663
rect 1989 -697 2023 -663
rect 2057 -697 2091 -663
rect 2125 -697 2159 -663
rect 2193 -697 2227 -663
rect 2261 -697 2295 -663
rect 2329 -697 2363 -663
rect 2397 -697 2431 -663
rect 2465 -697 2499 -663
rect 2533 -697 2567 -663
rect 2601 -697 2635 -663
rect 2669 -697 2703 -663
rect 2737 -697 2771 -663
rect 2805 -697 2839 -663
rect 2873 -697 2907 -663
rect 2941 -697 2975 -663
rect 3009 -697 3043 -663
rect 3077 -697 3111 -663
rect 3145 -697 3179 -663
rect 3213 -697 3247 -663
rect 3281 -697 3315 -663
rect 3349 -697 3383 -663
rect 3417 -697 3451 -663
rect 3485 -697 3519 -663
rect 3553 -697 3587 -663
rect 3621 -697 3655 -663
rect 3689 -697 3723 -663
rect 3757 -697 3791 -663
rect 3825 -697 3859 -663
rect 3893 -697 3927 -663
rect 3961 -697 3995 -663
rect 4029 -697 4063 -663
rect 4097 -697 4131 -663
rect 4165 -697 4199 -663
rect 4233 -697 4267 -663
rect 4301 -697 4335 -663
rect 4369 -697 4403 -663
rect 4437 -697 4560 -663
rect -480 -720 4560 -697
rect 8000 457 13040 480
rect 8000 423 8123 457
rect 8157 423 8191 457
rect 8225 423 8259 457
rect 8293 423 8327 457
rect 8361 423 8395 457
rect 8429 423 8463 457
rect 8497 423 8531 457
rect 8565 423 8599 457
rect 8633 423 8667 457
rect 8701 423 8735 457
rect 8769 423 8803 457
rect 8837 423 8871 457
rect 8905 423 8939 457
rect 8973 423 9007 457
rect 9041 423 9075 457
rect 9109 423 9143 457
rect 9177 423 9211 457
rect 9245 423 9279 457
rect 9313 423 9347 457
rect 9381 423 9415 457
rect 9449 423 9483 457
rect 9517 423 9551 457
rect 9585 423 9619 457
rect 9653 423 9687 457
rect 9721 423 9755 457
rect 9789 423 9823 457
rect 9857 423 9891 457
rect 9925 423 9959 457
rect 9993 423 10027 457
rect 10061 423 10095 457
rect 10129 423 10163 457
rect 10197 423 10231 457
rect 10265 423 10299 457
rect 10333 423 10367 457
rect 10401 423 10435 457
rect 10469 423 10503 457
rect 10537 423 10571 457
rect 10605 423 10639 457
rect 10673 423 10707 457
rect 10741 423 10775 457
rect 10809 423 10843 457
rect 10877 423 10911 457
rect 10945 423 10979 457
rect 11013 423 11047 457
rect 11081 423 11115 457
rect 11149 423 11183 457
rect 11217 423 11251 457
rect 11285 423 11319 457
rect 11353 423 11387 457
rect 11421 423 11455 457
rect 11489 423 11523 457
rect 11557 423 11591 457
rect 11625 423 11659 457
rect 11693 423 11727 457
rect 11761 423 11795 457
rect 11829 423 11863 457
rect 11897 423 11931 457
rect 11965 423 11999 457
rect 12033 423 12067 457
rect 12101 423 12135 457
rect 12169 423 12203 457
rect 12237 423 12271 457
rect 12305 423 12339 457
rect 12373 423 12407 457
rect 12441 423 12475 457
rect 12509 423 12543 457
rect 12577 423 12611 457
rect 12645 423 12679 457
rect 12713 423 12747 457
rect 12781 423 12815 457
rect 12849 423 12883 457
rect 12917 423 13040 457
rect 8000 400 13040 423
rect 8000 319 8080 400
rect 8000 285 8023 319
rect 8057 285 8080 319
rect 8000 251 8080 285
rect 8000 217 8023 251
rect 8057 217 8080 251
rect 8000 183 8080 217
rect 8000 149 8023 183
rect 8057 149 8080 183
rect 8000 115 8080 149
rect 8000 81 8023 115
rect 8057 81 8080 115
rect 8000 47 8080 81
rect 8000 13 8023 47
rect 8057 13 8080 47
rect 8000 -21 8080 13
rect 8000 -55 8023 -21
rect 8057 -55 8080 -21
rect 8000 -89 8080 -55
rect 8000 -123 8023 -89
rect 8057 -123 8080 -89
rect 8000 -157 8080 -123
rect 8000 -191 8023 -157
rect 8057 -191 8080 -157
rect 8000 -225 8080 -191
rect 8000 -259 8023 -225
rect 8057 -259 8080 -225
rect 8000 -293 8080 -259
rect 8000 -327 8023 -293
rect 8057 -327 8080 -293
rect 8000 -361 8080 -327
rect 8000 -395 8023 -361
rect 8057 -395 8080 -361
rect 8000 -429 8080 -395
rect 8000 -463 8023 -429
rect 8057 -463 8080 -429
rect 8000 -497 8080 -463
rect 8000 -531 8023 -497
rect 8057 -531 8080 -497
rect 8000 -565 8080 -531
rect 12960 319 13040 400
rect 12960 285 12983 319
rect 13017 285 13040 319
rect 12960 251 13040 285
rect 12960 217 12983 251
rect 13017 217 13040 251
rect 12960 183 13040 217
rect 12960 149 12983 183
rect 13017 149 13040 183
rect 12960 115 13040 149
rect 12960 81 12983 115
rect 13017 81 13040 115
rect 12960 47 13040 81
rect 12960 13 12983 47
rect 13017 13 13040 47
rect 12960 -21 13040 13
rect 12960 -55 12983 -21
rect 13017 -55 13040 -21
rect 12960 -89 13040 -55
rect 12960 -123 12983 -89
rect 13017 -123 13040 -89
rect 12960 -157 13040 -123
rect 12960 -191 12983 -157
rect 13017 -191 13040 -157
rect 12960 -225 13040 -191
rect 12960 -259 12983 -225
rect 13017 -259 13040 -225
rect 12960 -293 13040 -259
rect 12960 -327 12983 -293
rect 13017 -327 13040 -293
rect 12960 -361 13040 -327
rect 12960 -395 12983 -361
rect 13017 -395 13040 -361
rect 12960 -429 13040 -395
rect 12960 -463 12983 -429
rect 13017 -463 13040 -429
rect 12960 -497 13040 -463
rect 12960 -531 12983 -497
rect 13017 -531 13040 -497
rect 8000 -599 8023 -565
rect 8057 -599 8080 -565
rect 8000 -640 8080 -599
rect 12960 -565 13040 -531
rect 12960 -599 12983 -565
rect 13017 -599 13040 -565
rect 12960 -640 13040 -599
rect 8000 -663 13040 -640
rect 8000 -697 8123 -663
rect 8157 -697 8191 -663
rect 8225 -697 8259 -663
rect 8293 -697 8327 -663
rect 8361 -697 8395 -663
rect 8429 -697 8463 -663
rect 8497 -697 8531 -663
rect 8565 -697 8599 -663
rect 8633 -697 8667 -663
rect 8701 -697 8735 -663
rect 8769 -697 8803 -663
rect 8837 -697 8871 -663
rect 8905 -697 8939 -663
rect 8973 -697 9007 -663
rect 9041 -697 9075 -663
rect 9109 -697 9143 -663
rect 9177 -697 9211 -663
rect 9245 -697 9279 -663
rect 9313 -697 9347 -663
rect 9381 -697 9415 -663
rect 9449 -697 9483 -663
rect 9517 -697 9551 -663
rect 9585 -697 9619 -663
rect 9653 -697 9687 -663
rect 9721 -697 9755 -663
rect 9789 -697 9823 -663
rect 9857 -697 9891 -663
rect 9925 -697 9959 -663
rect 9993 -697 10027 -663
rect 10061 -697 10095 -663
rect 10129 -697 10163 -663
rect 10197 -697 10231 -663
rect 10265 -697 10299 -663
rect 10333 -697 10367 -663
rect 10401 -697 10435 -663
rect 10469 -697 10503 -663
rect 10537 -697 10571 -663
rect 10605 -697 10639 -663
rect 10673 -697 10707 -663
rect 10741 -697 10775 -663
rect 10809 -697 10843 -663
rect 10877 -697 10911 -663
rect 10945 -697 10979 -663
rect 11013 -697 11047 -663
rect 11081 -697 11115 -663
rect 11149 -697 11183 -663
rect 11217 -697 11251 -663
rect 11285 -697 11319 -663
rect 11353 -697 11387 -663
rect 11421 -697 11455 -663
rect 11489 -697 11523 -663
rect 11557 -697 11591 -663
rect 11625 -697 11659 -663
rect 11693 -697 11727 -663
rect 11761 -697 11795 -663
rect 11829 -697 11863 -663
rect 11897 -697 11931 -663
rect 11965 -697 11999 -663
rect 12033 -697 12067 -663
rect 12101 -697 12135 -663
rect 12169 -697 12203 -663
rect 12237 -697 12271 -663
rect 12305 -697 12339 -663
rect 12373 -697 12407 -663
rect 12441 -697 12475 -663
rect 12509 -697 12543 -663
rect 12577 -697 12611 -663
rect 12645 -697 12679 -663
rect 12713 -697 12747 -663
rect 12781 -697 12815 -663
rect 12849 -697 12883 -663
rect 12917 -697 13040 -663
rect 8000 -720 13040 -697
<< mvnsubdiff >>
rect -320 4137 4400 4160
rect -320 4103 -187 4137
rect -153 4103 -119 4137
rect -85 4103 -51 4137
rect -17 4103 17 4137
rect 51 4103 85 4137
rect 119 4103 153 4137
rect 187 4103 221 4137
rect 255 4103 289 4137
rect 323 4103 357 4137
rect 391 4103 425 4137
rect 459 4103 493 4137
rect 527 4103 561 4137
rect 595 4103 629 4137
rect 663 4103 697 4137
rect 731 4103 765 4137
rect 799 4103 833 4137
rect 867 4103 901 4137
rect 935 4103 969 4137
rect 1003 4103 1037 4137
rect 1071 4103 1105 4137
rect 1139 4103 1173 4137
rect 1207 4103 1241 4137
rect 1275 4103 1309 4137
rect 1343 4103 1377 4137
rect 1411 4103 1445 4137
rect 1479 4103 1513 4137
rect 1547 4103 1581 4137
rect 1615 4103 1649 4137
rect 1683 4103 1717 4137
rect 1751 4103 1785 4137
rect 1819 4103 1853 4137
rect 1887 4103 1921 4137
rect 1955 4103 1989 4137
rect 2023 4103 2057 4137
rect 2091 4103 2125 4137
rect 2159 4103 2193 4137
rect 2227 4103 2261 4137
rect 2295 4103 2329 4137
rect 2363 4103 2397 4137
rect 2431 4103 2465 4137
rect 2499 4103 2533 4137
rect 2567 4103 2601 4137
rect 2635 4103 2669 4137
rect 2703 4103 2737 4137
rect 2771 4103 2805 4137
rect 2839 4103 2873 4137
rect 2907 4103 2941 4137
rect 2975 4103 3009 4137
rect 3043 4103 3077 4137
rect 3111 4103 3145 4137
rect 3179 4103 3213 4137
rect 3247 4103 3281 4137
rect 3315 4103 3349 4137
rect 3383 4103 3417 4137
rect 3451 4103 3485 4137
rect 3519 4103 3553 4137
rect 3587 4103 3621 4137
rect 3655 4103 3689 4137
rect 3723 4103 3757 4137
rect 3791 4103 3825 4137
rect 3859 4103 3893 4137
rect 3927 4103 3961 4137
rect 3995 4103 4029 4137
rect 4063 4103 4097 4137
rect 4131 4103 4165 4137
rect 4199 4103 4233 4137
rect 4267 4103 4400 4137
rect -320 4080 4400 4103
rect -320 4023 -240 4080
rect -320 3989 -297 4023
rect -263 3989 -240 4023
rect 4320 4023 4400 4080
rect -320 3955 -240 3989
rect -320 3921 -297 3955
rect -263 3921 -240 3955
rect -320 3887 -240 3921
rect 4320 3989 4343 4023
rect 4377 3989 4400 4023
rect 4320 3955 4400 3989
rect 4320 3921 4343 3955
rect 4377 3921 4400 3955
rect -320 3853 -297 3887
rect -263 3853 -240 3887
rect -320 3819 -240 3853
rect -320 3785 -297 3819
rect -263 3785 -240 3819
rect -320 3751 -240 3785
rect 4320 3887 4400 3921
rect 4320 3853 4343 3887
rect 4377 3853 4400 3887
rect 4320 3819 4400 3853
rect 4320 3785 4343 3819
rect 4377 3785 4400 3819
rect -320 3717 -297 3751
rect -263 3717 -240 3751
rect -320 3683 -240 3717
rect 4320 3751 4400 3785
rect 4320 3717 4343 3751
rect 4377 3717 4400 3751
rect -320 3649 -297 3683
rect -263 3649 -240 3683
rect 4320 3683 4400 3717
rect -320 3615 -240 3649
rect -320 3581 -297 3615
rect -263 3581 -240 3615
rect 4320 3649 4343 3683
rect 4377 3649 4400 3683
rect 4320 3615 4400 3649
rect -320 3547 -240 3581
rect -320 3513 -297 3547
rect -263 3513 -240 3547
rect -320 3479 -240 3513
rect -320 3445 -297 3479
rect -263 3445 -240 3479
rect -320 3411 -240 3445
rect 4320 3581 4343 3615
rect 4377 3581 4400 3615
rect 4320 3547 4400 3581
rect 4320 3513 4343 3547
rect 4377 3513 4400 3547
rect 4320 3479 4400 3513
rect 4320 3445 4343 3479
rect 4377 3445 4400 3479
rect -320 3377 -297 3411
rect -263 3377 -240 3411
rect -320 3360 -240 3377
rect 4320 3411 4400 3445
rect 4320 3377 4343 3411
rect 4377 3377 4400 3411
rect 4320 3360 4400 3377
rect -320 3337 4400 3360
rect -320 3303 -187 3337
rect -153 3303 -119 3337
rect -85 3303 -51 3337
rect -17 3303 17 3337
rect 51 3303 85 3337
rect 119 3303 153 3337
rect 187 3303 221 3337
rect 255 3303 289 3337
rect 323 3303 357 3337
rect 391 3303 425 3337
rect 459 3303 493 3337
rect 527 3303 561 3337
rect 595 3303 629 3337
rect 663 3303 697 3337
rect 731 3303 765 3337
rect 799 3303 833 3337
rect 867 3303 901 3337
rect 935 3303 969 3337
rect 1003 3303 1037 3337
rect 1071 3303 1105 3337
rect 1139 3303 1173 3337
rect 1207 3303 1241 3337
rect 1275 3303 1309 3337
rect 1343 3303 1377 3337
rect 1411 3303 1445 3337
rect 1479 3303 1513 3337
rect 1547 3303 1581 3337
rect 1615 3303 1649 3337
rect 1683 3303 1717 3337
rect 1751 3303 1785 3337
rect 1819 3303 1853 3337
rect 1887 3303 1921 3337
rect 1955 3303 1989 3337
rect 2023 3303 2057 3337
rect 2091 3303 2125 3337
rect 2159 3303 2193 3337
rect 2227 3303 2261 3337
rect 2295 3303 2329 3337
rect 2363 3303 2397 3337
rect 2431 3303 2465 3337
rect 2499 3303 2533 3337
rect 2567 3303 2601 3337
rect 2635 3303 2669 3337
rect 2703 3303 2737 3337
rect 2771 3303 2805 3337
rect 2839 3303 2873 3337
rect 2907 3303 2941 3337
rect 2975 3303 3009 3337
rect 3043 3303 3077 3337
rect 3111 3303 3145 3337
rect 3179 3303 3213 3337
rect 3247 3303 3281 3337
rect 3315 3303 3349 3337
rect 3383 3303 3417 3337
rect 3451 3303 3485 3337
rect 3519 3303 3553 3337
rect 3587 3303 3621 3337
rect 3655 3303 3689 3337
rect 3723 3303 3757 3337
rect 3791 3303 3825 3337
rect 3859 3303 3893 3337
rect 3927 3303 3961 3337
rect 3995 3303 4029 3337
rect 4063 3303 4097 3337
rect 4131 3303 4165 3337
rect 4199 3303 4233 3337
rect 4267 3303 4400 3337
rect -320 3280 4400 3303
rect 8160 4137 12880 4160
rect 8160 4103 8293 4137
rect 8327 4103 8361 4137
rect 8395 4103 8429 4137
rect 8463 4103 8497 4137
rect 8531 4103 8565 4137
rect 8599 4103 8633 4137
rect 8667 4103 8701 4137
rect 8735 4103 8769 4137
rect 8803 4103 8837 4137
rect 8871 4103 8905 4137
rect 8939 4103 8973 4137
rect 9007 4103 9041 4137
rect 9075 4103 9109 4137
rect 9143 4103 9177 4137
rect 9211 4103 9245 4137
rect 9279 4103 9313 4137
rect 9347 4103 9381 4137
rect 9415 4103 9449 4137
rect 9483 4103 9517 4137
rect 9551 4103 9585 4137
rect 9619 4103 9653 4137
rect 9687 4103 9721 4137
rect 9755 4103 9789 4137
rect 9823 4103 9857 4137
rect 9891 4103 9925 4137
rect 9959 4103 9993 4137
rect 10027 4103 10061 4137
rect 10095 4103 10129 4137
rect 10163 4103 10197 4137
rect 10231 4103 10265 4137
rect 10299 4103 10333 4137
rect 10367 4103 10401 4137
rect 10435 4103 10469 4137
rect 10503 4103 10537 4137
rect 10571 4103 10605 4137
rect 10639 4103 10673 4137
rect 10707 4103 10741 4137
rect 10775 4103 10809 4137
rect 10843 4103 10877 4137
rect 10911 4103 10945 4137
rect 10979 4103 11013 4137
rect 11047 4103 11081 4137
rect 11115 4103 11149 4137
rect 11183 4103 11217 4137
rect 11251 4103 11285 4137
rect 11319 4103 11353 4137
rect 11387 4103 11421 4137
rect 11455 4103 11489 4137
rect 11523 4103 11557 4137
rect 11591 4103 11625 4137
rect 11659 4103 11693 4137
rect 11727 4103 11761 4137
rect 11795 4103 11829 4137
rect 11863 4103 11897 4137
rect 11931 4103 11965 4137
rect 11999 4103 12033 4137
rect 12067 4103 12101 4137
rect 12135 4103 12169 4137
rect 12203 4103 12237 4137
rect 12271 4103 12305 4137
rect 12339 4103 12373 4137
rect 12407 4103 12441 4137
rect 12475 4103 12509 4137
rect 12543 4103 12577 4137
rect 12611 4103 12645 4137
rect 12679 4103 12713 4137
rect 12747 4103 12880 4137
rect 8160 4080 12880 4103
rect 8160 4023 8240 4080
rect 8160 3989 8183 4023
rect 8217 3989 8240 4023
rect 12800 4023 12880 4080
rect 8160 3955 8240 3989
rect 8160 3921 8183 3955
rect 8217 3921 8240 3955
rect 8160 3887 8240 3921
rect 12800 3989 12823 4023
rect 12857 3989 12880 4023
rect 12800 3955 12880 3989
rect 12800 3921 12823 3955
rect 12857 3921 12880 3955
rect 8160 3853 8183 3887
rect 8217 3853 8240 3887
rect 8160 3819 8240 3853
rect 8160 3785 8183 3819
rect 8217 3785 8240 3819
rect 8160 3751 8240 3785
rect 12800 3887 12880 3921
rect 12800 3853 12823 3887
rect 12857 3853 12880 3887
rect 12800 3819 12880 3853
rect 12800 3785 12823 3819
rect 12857 3785 12880 3819
rect 8160 3717 8183 3751
rect 8217 3717 8240 3751
rect 8160 3683 8240 3717
rect 12800 3751 12880 3785
rect 12800 3717 12823 3751
rect 12857 3717 12880 3751
rect 8160 3649 8183 3683
rect 8217 3649 8240 3683
rect 12800 3683 12880 3717
rect 8160 3615 8240 3649
rect 8160 3581 8183 3615
rect 8217 3581 8240 3615
rect 12800 3649 12823 3683
rect 12857 3649 12880 3683
rect 12800 3615 12880 3649
rect 8160 3547 8240 3581
rect 8160 3513 8183 3547
rect 8217 3513 8240 3547
rect 8160 3479 8240 3513
rect 8160 3445 8183 3479
rect 8217 3445 8240 3479
rect 8160 3411 8240 3445
rect 12800 3581 12823 3615
rect 12857 3581 12880 3615
rect 12800 3547 12880 3581
rect 12800 3513 12823 3547
rect 12857 3513 12880 3547
rect 12800 3479 12880 3513
rect 12800 3445 12823 3479
rect 12857 3445 12880 3479
rect 8160 3377 8183 3411
rect 8217 3377 8240 3411
rect 8160 3360 8240 3377
rect 12800 3411 12880 3445
rect 12800 3377 12823 3411
rect 12857 3377 12880 3411
rect 12800 3360 12880 3377
rect 8160 3337 12880 3360
rect 8160 3303 8293 3337
rect 8327 3303 8361 3337
rect 8395 3303 8429 3337
rect 8463 3303 8497 3337
rect 8531 3303 8565 3337
rect 8599 3303 8633 3337
rect 8667 3303 8701 3337
rect 8735 3303 8769 3337
rect 8803 3303 8837 3337
rect 8871 3303 8905 3337
rect 8939 3303 8973 3337
rect 9007 3303 9041 3337
rect 9075 3303 9109 3337
rect 9143 3303 9177 3337
rect 9211 3303 9245 3337
rect 9279 3303 9313 3337
rect 9347 3303 9381 3337
rect 9415 3303 9449 3337
rect 9483 3303 9517 3337
rect 9551 3303 9585 3337
rect 9619 3303 9653 3337
rect 9687 3303 9721 3337
rect 9755 3303 9789 3337
rect 9823 3303 9857 3337
rect 9891 3303 9925 3337
rect 9959 3303 9993 3337
rect 10027 3303 10061 3337
rect 10095 3303 10129 3337
rect 10163 3303 10197 3337
rect 10231 3303 10265 3337
rect 10299 3303 10333 3337
rect 10367 3303 10401 3337
rect 10435 3303 10469 3337
rect 10503 3303 10537 3337
rect 10571 3303 10605 3337
rect 10639 3303 10673 3337
rect 10707 3303 10741 3337
rect 10775 3303 10809 3337
rect 10843 3303 10877 3337
rect 10911 3303 10945 3337
rect 10979 3303 11013 3337
rect 11047 3303 11081 3337
rect 11115 3303 11149 3337
rect 11183 3303 11217 3337
rect 11251 3303 11285 3337
rect 11319 3303 11353 3337
rect 11387 3303 11421 3337
rect 11455 3303 11489 3337
rect 11523 3303 11557 3337
rect 11591 3303 11625 3337
rect 11659 3303 11693 3337
rect 11727 3303 11761 3337
rect 11795 3303 11829 3337
rect 11863 3303 11897 3337
rect 11931 3303 11965 3337
rect 11999 3303 12033 3337
rect 12067 3303 12101 3337
rect 12135 3303 12169 3337
rect 12203 3303 12237 3337
rect 12271 3303 12305 3337
rect 12339 3303 12373 3337
rect 12407 3303 12441 3337
rect 12475 3303 12509 3337
rect 12543 3303 12577 3337
rect 12611 3303 12645 3337
rect 12679 3303 12713 3337
rect 12747 3303 12880 3337
rect 8160 3280 12880 3303
rect -320 2857 4400 2880
rect -320 2823 -187 2857
rect -153 2823 -119 2857
rect -85 2823 -51 2857
rect -17 2823 17 2857
rect 51 2823 85 2857
rect 119 2823 153 2857
rect 187 2823 221 2857
rect 255 2823 289 2857
rect 323 2823 357 2857
rect 391 2823 425 2857
rect 459 2823 493 2857
rect 527 2823 561 2857
rect 595 2823 629 2857
rect 663 2823 697 2857
rect 731 2823 765 2857
rect 799 2823 833 2857
rect 867 2823 901 2857
rect 935 2823 969 2857
rect 1003 2823 1037 2857
rect 1071 2823 1105 2857
rect 1139 2823 1173 2857
rect 1207 2823 1241 2857
rect 1275 2823 1309 2857
rect 1343 2823 1377 2857
rect 1411 2823 1445 2857
rect 1479 2823 1513 2857
rect 1547 2823 1581 2857
rect 1615 2823 1649 2857
rect 1683 2823 1717 2857
rect 1751 2823 1785 2857
rect 1819 2823 1853 2857
rect 1887 2823 1921 2857
rect 1955 2823 1989 2857
rect 2023 2823 2057 2857
rect 2091 2823 2125 2857
rect 2159 2823 2193 2857
rect 2227 2823 2261 2857
rect 2295 2823 2329 2857
rect 2363 2823 2397 2857
rect 2431 2823 2465 2857
rect 2499 2823 2533 2857
rect 2567 2823 2601 2857
rect 2635 2823 2669 2857
rect 2703 2823 2737 2857
rect 2771 2823 2805 2857
rect 2839 2823 2873 2857
rect 2907 2823 2941 2857
rect 2975 2823 3009 2857
rect 3043 2823 3077 2857
rect 3111 2823 3145 2857
rect 3179 2823 3213 2857
rect 3247 2823 3281 2857
rect 3315 2823 3349 2857
rect 3383 2823 3417 2857
rect 3451 2823 3485 2857
rect 3519 2823 3553 2857
rect 3587 2823 3621 2857
rect 3655 2823 3689 2857
rect 3723 2823 3757 2857
rect 3791 2823 3825 2857
rect 3859 2823 3893 2857
rect 3927 2823 3961 2857
rect 3995 2823 4029 2857
rect 4063 2823 4097 2857
rect 4131 2823 4165 2857
rect 4199 2823 4233 2857
rect 4267 2823 4400 2857
rect -320 2800 4400 2823
rect -320 2783 -240 2800
rect -320 2749 -297 2783
rect -263 2749 -240 2783
rect -320 2715 -240 2749
rect 4320 2783 4400 2800
rect 4320 2749 4343 2783
rect 4377 2749 4400 2783
rect -320 2681 -297 2715
rect -263 2681 -240 2715
rect -320 2647 -240 2681
rect -320 2613 -297 2647
rect -263 2613 -240 2647
rect -320 2579 -240 2613
rect -320 2545 -297 2579
rect -263 2545 -240 2579
rect 4320 2715 4400 2749
rect 4320 2681 4343 2715
rect 4377 2681 4400 2715
rect 4320 2647 4400 2681
rect 4320 2613 4343 2647
rect 4377 2613 4400 2647
rect 4320 2579 4400 2613
rect -320 2511 -240 2545
rect -320 2477 -297 2511
rect -263 2477 -240 2511
rect 4320 2545 4343 2579
rect 4377 2545 4400 2579
rect 4320 2511 4400 2545
rect -320 2443 -240 2477
rect 4320 2477 4343 2511
rect 4377 2477 4400 2511
rect -320 2409 -297 2443
rect -263 2409 -240 2443
rect -320 2375 -240 2409
rect 4320 2443 4400 2477
rect 4320 2409 4343 2443
rect 4377 2409 4400 2443
rect -320 2341 -297 2375
rect -263 2341 -240 2375
rect -320 2307 -240 2341
rect -320 2273 -297 2307
rect -263 2273 -240 2307
rect -320 2239 -240 2273
rect 4320 2375 4400 2409
rect 4320 2341 4343 2375
rect 4377 2341 4400 2375
rect 4320 2307 4400 2341
rect 4320 2273 4343 2307
rect 4377 2273 4400 2307
rect -320 2205 -297 2239
rect -263 2205 -240 2239
rect -320 2171 -240 2205
rect -320 2137 -297 2171
rect -263 2137 -240 2171
rect 4320 2239 4400 2273
rect 4320 2205 4343 2239
rect 4377 2205 4400 2239
rect 4320 2171 4400 2205
rect -320 2080 -240 2137
rect 4320 2137 4343 2171
rect 4377 2137 4400 2171
rect 4320 2080 4400 2137
rect -320 2057 4400 2080
rect -320 2023 -187 2057
rect -153 2023 -119 2057
rect -85 2023 -51 2057
rect -17 2023 17 2057
rect 51 2023 85 2057
rect 119 2023 153 2057
rect 187 2023 221 2057
rect 255 2023 289 2057
rect 323 2023 357 2057
rect 391 2023 425 2057
rect 459 2023 493 2057
rect 527 2023 561 2057
rect 595 2023 629 2057
rect 663 2023 697 2057
rect 731 2023 765 2057
rect 799 2023 833 2057
rect 867 2023 901 2057
rect 935 2023 969 2057
rect 1003 2023 1037 2057
rect 1071 2023 1105 2057
rect 1139 2023 1173 2057
rect 1207 2023 1241 2057
rect 1275 2023 1309 2057
rect 1343 2023 1377 2057
rect 1411 2023 1445 2057
rect 1479 2023 1513 2057
rect 1547 2023 1581 2057
rect 1615 2023 1649 2057
rect 1683 2023 1717 2057
rect 1751 2023 1785 2057
rect 1819 2023 1853 2057
rect 1887 2023 1921 2057
rect 1955 2023 1989 2057
rect 2023 2023 2057 2057
rect 2091 2023 2125 2057
rect 2159 2023 2193 2057
rect 2227 2023 2261 2057
rect 2295 2023 2329 2057
rect 2363 2023 2397 2057
rect 2431 2023 2465 2057
rect 2499 2023 2533 2057
rect 2567 2023 2601 2057
rect 2635 2023 2669 2057
rect 2703 2023 2737 2057
rect 2771 2023 2805 2057
rect 2839 2023 2873 2057
rect 2907 2023 2941 2057
rect 2975 2023 3009 2057
rect 3043 2023 3077 2057
rect 3111 2023 3145 2057
rect 3179 2023 3213 2057
rect 3247 2023 3281 2057
rect 3315 2023 3349 2057
rect 3383 2023 3417 2057
rect 3451 2023 3485 2057
rect 3519 2023 3553 2057
rect 3587 2023 3621 2057
rect 3655 2023 3689 2057
rect 3723 2023 3757 2057
rect 3791 2023 3825 2057
rect 3859 2023 3893 2057
rect 3927 2023 3961 2057
rect 3995 2023 4029 2057
rect 4063 2023 4097 2057
rect 4131 2023 4165 2057
rect 4199 2023 4233 2057
rect 4267 2023 4400 2057
rect -320 2000 4400 2023
rect 8160 2857 12880 2880
rect 8160 2823 8293 2857
rect 8327 2823 8361 2857
rect 8395 2823 8429 2857
rect 8463 2823 8497 2857
rect 8531 2823 8565 2857
rect 8599 2823 8633 2857
rect 8667 2823 8701 2857
rect 8735 2823 8769 2857
rect 8803 2823 8837 2857
rect 8871 2823 8905 2857
rect 8939 2823 8973 2857
rect 9007 2823 9041 2857
rect 9075 2823 9109 2857
rect 9143 2823 9177 2857
rect 9211 2823 9245 2857
rect 9279 2823 9313 2857
rect 9347 2823 9381 2857
rect 9415 2823 9449 2857
rect 9483 2823 9517 2857
rect 9551 2823 9585 2857
rect 9619 2823 9653 2857
rect 9687 2823 9721 2857
rect 9755 2823 9789 2857
rect 9823 2823 9857 2857
rect 9891 2823 9925 2857
rect 9959 2823 9993 2857
rect 10027 2823 10061 2857
rect 10095 2823 10129 2857
rect 10163 2823 10197 2857
rect 10231 2823 10265 2857
rect 10299 2823 10333 2857
rect 10367 2823 10401 2857
rect 10435 2823 10469 2857
rect 10503 2823 10537 2857
rect 10571 2823 10605 2857
rect 10639 2823 10673 2857
rect 10707 2823 10741 2857
rect 10775 2823 10809 2857
rect 10843 2823 10877 2857
rect 10911 2823 10945 2857
rect 10979 2823 11013 2857
rect 11047 2823 11081 2857
rect 11115 2823 11149 2857
rect 11183 2823 11217 2857
rect 11251 2823 11285 2857
rect 11319 2823 11353 2857
rect 11387 2823 11421 2857
rect 11455 2823 11489 2857
rect 11523 2823 11557 2857
rect 11591 2823 11625 2857
rect 11659 2823 11693 2857
rect 11727 2823 11761 2857
rect 11795 2823 11829 2857
rect 11863 2823 11897 2857
rect 11931 2823 11965 2857
rect 11999 2823 12033 2857
rect 12067 2823 12101 2857
rect 12135 2823 12169 2857
rect 12203 2823 12237 2857
rect 12271 2823 12305 2857
rect 12339 2823 12373 2857
rect 12407 2823 12441 2857
rect 12475 2823 12509 2857
rect 12543 2823 12577 2857
rect 12611 2823 12645 2857
rect 12679 2823 12713 2857
rect 12747 2823 12880 2857
rect 8160 2800 12880 2823
rect 8160 2783 8240 2800
rect 8160 2749 8183 2783
rect 8217 2749 8240 2783
rect 8160 2715 8240 2749
rect 12800 2783 12880 2800
rect 12800 2749 12823 2783
rect 12857 2749 12880 2783
rect 8160 2681 8183 2715
rect 8217 2681 8240 2715
rect 8160 2647 8240 2681
rect 8160 2613 8183 2647
rect 8217 2613 8240 2647
rect 8160 2579 8240 2613
rect 8160 2545 8183 2579
rect 8217 2545 8240 2579
rect 12800 2715 12880 2749
rect 12800 2681 12823 2715
rect 12857 2681 12880 2715
rect 12800 2647 12880 2681
rect 12800 2613 12823 2647
rect 12857 2613 12880 2647
rect 12800 2579 12880 2613
rect 8160 2511 8240 2545
rect 8160 2477 8183 2511
rect 8217 2477 8240 2511
rect 12800 2545 12823 2579
rect 12857 2545 12880 2579
rect 12800 2511 12880 2545
rect 8160 2443 8240 2477
rect 12800 2477 12823 2511
rect 12857 2477 12880 2511
rect 8160 2409 8183 2443
rect 8217 2409 8240 2443
rect 8160 2375 8240 2409
rect 12800 2443 12880 2477
rect 12800 2409 12823 2443
rect 12857 2409 12880 2443
rect 8160 2341 8183 2375
rect 8217 2341 8240 2375
rect 8160 2307 8240 2341
rect 8160 2273 8183 2307
rect 8217 2273 8240 2307
rect 8160 2239 8240 2273
rect 12800 2375 12880 2409
rect 12800 2341 12823 2375
rect 12857 2341 12880 2375
rect 12800 2307 12880 2341
rect 12800 2273 12823 2307
rect 12857 2273 12880 2307
rect 8160 2205 8183 2239
rect 8217 2205 8240 2239
rect 8160 2171 8240 2205
rect 8160 2137 8183 2171
rect 8217 2137 8240 2171
rect 12800 2239 12880 2273
rect 12800 2205 12823 2239
rect 12857 2205 12880 2239
rect 12800 2171 12880 2205
rect 8160 2080 8240 2137
rect 12800 2137 12823 2171
rect 12857 2137 12880 2171
rect 12800 2080 12880 2137
rect 8160 2057 12880 2080
rect 8160 2023 8293 2057
rect 8327 2023 8361 2057
rect 8395 2023 8429 2057
rect 8463 2023 8497 2057
rect 8531 2023 8565 2057
rect 8599 2023 8633 2057
rect 8667 2023 8701 2057
rect 8735 2023 8769 2057
rect 8803 2023 8837 2057
rect 8871 2023 8905 2057
rect 8939 2023 8973 2057
rect 9007 2023 9041 2057
rect 9075 2023 9109 2057
rect 9143 2023 9177 2057
rect 9211 2023 9245 2057
rect 9279 2023 9313 2057
rect 9347 2023 9381 2057
rect 9415 2023 9449 2057
rect 9483 2023 9517 2057
rect 9551 2023 9585 2057
rect 9619 2023 9653 2057
rect 9687 2023 9721 2057
rect 9755 2023 9789 2057
rect 9823 2023 9857 2057
rect 9891 2023 9925 2057
rect 9959 2023 9993 2057
rect 10027 2023 10061 2057
rect 10095 2023 10129 2057
rect 10163 2023 10197 2057
rect 10231 2023 10265 2057
rect 10299 2023 10333 2057
rect 10367 2023 10401 2057
rect 10435 2023 10469 2057
rect 10503 2023 10537 2057
rect 10571 2023 10605 2057
rect 10639 2023 10673 2057
rect 10707 2023 10741 2057
rect 10775 2023 10809 2057
rect 10843 2023 10877 2057
rect 10911 2023 10945 2057
rect 10979 2023 11013 2057
rect 11047 2023 11081 2057
rect 11115 2023 11149 2057
rect 11183 2023 11217 2057
rect 11251 2023 11285 2057
rect 11319 2023 11353 2057
rect 11387 2023 11421 2057
rect 11455 2023 11489 2057
rect 11523 2023 11557 2057
rect 11591 2023 11625 2057
rect 11659 2023 11693 2057
rect 11727 2023 11761 2057
rect 11795 2023 11829 2057
rect 11863 2023 11897 2057
rect 11931 2023 11965 2057
rect 11999 2023 12033 2057
rect 12067 2023 12101 2057
rect 12135 2023 12169 2057
rect 12203 2023 12237 2057
rect 12271 2023 12305 2057
rect 12339 2023 12373 2057
rect 12407 2023 12441 2057
rect 12475 2023 12509 2057
rect 12543 2023 12577 2057
rect 12611 2023 12645 2057
rect 12679 2023 12713 2057
rect 12747 2023 12880 2057
rect 8160 2000 12880 2023
rect -320 1577 4400 1600
rect -320 1543 -187 1577
rect -153 1543 -119 1577
rect -85 1543 -51 1577
rect -17 1543 17 1577
rect 51 1543 85 1577
rect 119 1543 153 1577
rect 187 1543 221 1577
rect 255 1543 289 1577
rect 323 1543 357 1577
rect 391 1543 425 1577
rect 459 1543 493 1577
rect 527 1543 561 1577
rect 595 1543 629 1577
rect 663 1543 697 1577
rect 731 1543 765 1577
rect 799 1543 833 1577
rect 867 1543 901 1577
rect 935 1543 969 1577
rect 1003 1543 1037 1577
rect 1071 1543 1105 1577
rect 1139 1543 1173 1577
rect 1207 1543 1241 1577
rect 1275 1543 1309 1577
rect 1343 1543 1377 1577
rect 1411 1543 1445 1577
rect 1479 1543 1513 1577
rect 1547 1543 1581 1577
rect 1615 1543 1649 1577
rect 1683 1543 1717 1577
rect 1751 1543 1785 1577
rect 1819 1543 1853 1577
rect 1887 1543 1921 1577
rect 1955 1543 1989 1577
rect 2023 1543 2057 1577
rect 2091 1543 2125 1577
rect 2159 1543 2193 1577
rect 2227 1543 2261 1577
rect 2295 1543 2329 1577
rect 2363 1543 2397 1577
rect 2431 1543 2465 1577
rect 2499 1543 2533 1577
rect 2567 1543 2601 1577
rect 2635 1543 2669 1577
rect 2703 1543 2737 1577
rect 2771 1543 2805 1577
rect 2839 1543 2873 1577
rect 2907 1543 2941 1577
rect 2975 1543 3009 1577
rect 3043 1543 3077 1577
rect 3111 1543 3145 1577
rect 3179 1543 3213 1577
rect 3247 1543 3281 1577
rect 3315 1543 3349 1577
rect 3383 1543 3417 1577
rect 3451 1543 3485 1577
rect 3519 1543 3553 1577
rect 3587 1543 3621 1577
rect 3655 1543 3689 1577
rect 3723 1543 3757 1577
rect 3791 1543 3825 1577
rect 3859 1543 3893 1577
rect 3927 1543 3961 1577
rect 3995 1543 4029 1577
rect 4063 1543 4097 1577
rect 4131 1543 4165 1577
rect 4199 1543 4233 1577
rect 4267 1543 4400 1577
rect -320 1520 4400 1543
rect -320 1463 -240 1520
rect -320 1429 -297 1463
rect -263 1429 -240 1463
rect 4320 1463 4400 1520
rect -320 1395 -240 1429
rect -320 1361 -297 1395
rect -263 1361 -240 1395
rect -320 1327 -240 1361
rect 4320 1429 4343 1463
rect 4377 1429 4400 1463
rect 4320 1395 4400 1429
rect 4320 1361 4343 1395
rect 4377 1361 4400 1395
rect -320 1293 -297 1327
rect -263 1293 -240 1327
rect -320 1259 -240 1293
rect -320 1225 -297 1259
rect -263 1225 -240 1259
rect -320 1191 -240 1225
rect 4320 1327 4400 1361
rect 4320 1293 4343 1327
rect 4377 1293 4400 1327
rect 4320 1259 4400 1293
rect 4320 1225 4343 1259
rect 4377 1225 4400 1259
rect -320 1157 -297 1191
rect -263 1157 -240 1191
rect -320 1123 -240 1157
rect 4320 1191 4400 1225
rect 4320 1157 4343 1191
rect 4377 1157 4400 1191
rect -320 1089 -297 1123
rect -263 1089 -240 1123
rect 4320 1123 4400 1157
rect -320 1055 -240 1089
rect -320 1021 -297 1055
rect -263 1021 -240 1055
rect 4320 1089 4343 1123
rect 4377 1089 4400 1123
rect 4320 1055 4400 1089
rect -320 987 -240 1021
rect -320 953 -297 987
rect -263 953 -240 987
rect -320 919 -240 953
rect -320 885 -297 919
rect -263 885 -240 919
rect -320 851 -240 885
rect 4320 1021 4343 1055
rect 4377 1021 4400 1055
rect 4320 987 4400 1021
rect 4320 953 4343 987
rect 4377 953 4400 987
rect 4320 919 4400 953
rect 4320 885 4343 919
rect 4377 885 4400 919
rect -320 817 -297 851
rect -263 817 -240 851
rect -320 800 -240 817
rect 4320 851 4400 885
rect 4320 817 4343 851
rect 4377 817 4400 851
rect 4320 800 4400 817
rect -320 777 4400 800
rect -320 743 -187 777
rect -153 743 -119 777
rect -85 743 -51 777
rect -17 743 17 777
rect 51 743 85 777
rect 119 743 153 777
rect 187 743 221 777
rect 255 743 289 777
rect 323 743 357 777
rect 391 743 425 777
rect 459 743 493 777
rect 527 743 561 777
rect 595 743 629 777
rect 663 743 697 777
rect 731 743 765 777
rect 799 743 833 777
rect 867 743 901 777
rect 935 743 969 777
rect 1003 743 1037 777
rect 1071 743 1105 777
rect 1139 743 1173 777
rect 1207 743 1241 777
rect 1275 743 1309 777
rect 1343 743 1377 777
rect 1411 743 1445 777
rect 1479 743 1513 777
rect 1547 743 1581 777
rect 1615 743 1649 777
rect 1683 743 1717 777
rect 1751 743 1785 777
rect 1819 743 1853 777
rect 1887 743 1921 777
rect 1955 743 1989 777
rect 2023 743 2057 777
rect 2091 743 2125 777
rect 2159 743 2193 777
rect 2227 743 2261 777
rect 2295 743 2329 777
rect 2363 743 2397 777
rect 2431 743 2465 777
rect 2499 743 2533 777
rect 2567 743 2601 777
rect 2635 743 2669 777
rect 2703 743 2737 777
rect 2771 743 2805 777
rect 2839 743 2873 777
rect 2907 743 2941 777
rect 2975 743 3009 777
rect 3043 743 3077 777
rect 3111 743 3145 777
rect 3179 743 3213 777
rect 3247 743 3281 777
rect 3315 743 3349 777
rect 3383 743 3417 777
rect 3451 743 3485 777
rect 3519 743 3553 777
rect 3587 743 3621 777
rect 3655 743 3689 777
rect 3723 743 3757 777
rect 3791 743 3825 777
rect 3859 743 3893 777
rect 3927 743 3961 777
rect 3995 743 4029 777
rect 4063 743 4097 777
rect 4131 743 4165 777
rect 4199 743 4233 777
rect 4267 743 4400 777
rect -320 720 4400 743
rect 8160 1577 12880 1600
rect 8160 1543 8293 1577
rect 8327 1543 8361 1577
rect 8395 1543 8429 1577
rect 8463 1543 8497 1577
rect 8531 1543 8565 1577
rect 8599 1543 8633 1577
rect 8667 1543 8701 1577
rect 8735 1543 8769 1577
rect 8803 1543 8837 1577
rect 8871 1543 8905 1577
rect 8939 1543 8973 1577
rect 9007 1543 9041 1577
rect 9075 1543 9109 1577
rect 9143 1543 9177 1577
rect 9211 1543 9245 1577
rect 9279 1543 9313 1577
rect 9347 1543 9381 1577
rect 9415 1543 9449 1577
rect 9483 1543 9517 1577
rect 9551 1543 9585 1577
rect 9619 1543 9653 1577
rect 9687 1543 9721 1577
rect 9755 1543 9789 1577
rect 9823 1543 9857 1577
rect 9891 1543 9925 1577
rect 9959 1543 9993 1577
rect 10027 1543 10061 1577
rect 10095 1543 10129 1577
rect 10163 1543 10197 1577
rect 10231 1543 10265 1577
rect 10299 1543 10333 1577
rect 10367 1543 10401 1577
rect 10435 1543 10469 1577
rect 10503 1543 10537 1577
rect 10571 1543 10605 1577
rect 10639 1543 10673 1577
rect 10707 1543 10741 1577
rect 10775 1543 10809 1577
rect 10843 1543 10877 1577
rect 10911 1543 10945 1577
rect 10979 1543 11013 1577
rect 11047 1543 11081 1577
rect 11115 1543 11149 1577
rect 11183 1543 11217 1577
rect 11251 1543 11285 1577
rect 11319 1543 11353 1577
rect 11387 1543 11421 1577
rect 11455 1543 11489 1577
rect 11523 1543 11557 1577
rect 11591 1543 11625 1577
rect 11659 1543 11693 1577
rect 11727 1543 11761 1577
rect 11795 1543 11829 1577
rect 11863 1543 11897 1577
rect 11931 1543 11965 1577
rect 11999 1543 12033 1577
rect 12067 1543 12101 1577
rect 12135 1543 12169 1577
rect 12203 1543 12237 1577
rect 12271 1543 12305 1577
rect 12339 1543 12373 1577
rect 12407 1543 12441 1577
rect 12475 1543 12509 1577
rect 12543 1543 12577 1577
rect 12611 1543 12645 1577
rect 12679 1543 12713 1577
rect 12747 1543 12880 1577
rect 8160 1520 12880 1543
rect 8160 1463 8240 1520
rect 8160 1429 8183 1463
rect 8217 1429 8240 1463
rect 12800 1463 12880 1520
rect 8160 1395 8240 1429
rect 8160 1361 8183 1395
rect 8217 1361 8240 1395
rect 8160 1327 8240 1361
rect 12800 1429 12823 1463
rect 12857 1429 12880 1463
rect 12800 1395 12880 1429
rect 12800 1361 12823 1395
rect 12857 1361 12880 1395
rect 8160 1293 8183 1327
rect 8217 1293 8240 1327
rect 8160 1259 8240 1293
rect 8160 1225 8183 1259
rect 8217 1225 8240 1259
rect 8160 1191 8240 1225
rect 12800 1327 12880 1361
rect 12800 1293 12823 1327
rect 12857 1293 12880 1327
rect 12800 1259 12880 1293
rect 12800 1225 12823 1259
rect 12857 1225 12880 1259
rect 8160 1157 8183 1191
rect 8217 1157 8240 1191
rect 8160 1123 8240 1157
rect 12800 1191 12880 1225
rect 12800 1157 12823 1191
rect 12857 1157 12880 1191
rect 8160 1089 8183 1123
rect 8217 1089 8240 1123
rect 12800 1123 12880 1157
rect 8160 1055 8240 1089
rect 8160 1021 8183 1055
rect 8217 1021 8240 1055
rect 12800 1089 12823 1123
rect 12857 1089 12880 1123
rect 12800 1055 12880 1089
rect 8160 987 8240 1021
rect 8160 953 8183 987
rect 8217 953 8240 987
rect 8160 919 8240 953
rect 8160 885 8183 919
rect 8217 885 8240 919
rect 8160 851 8240 885
rect 12800 1021 12823 1055
rect 12857 1021 12880 1055
rect 12800 987 12880 1021
rect 12800 953 12823 987
rect 12857 953 12880 987
rect 12800 919 12880 953
rect 12800 885 12823 919
rect 12857 885 12880 919
rect 8160 817 8183 851
rect 8217 817 8240 851
rect 8160 800 8240 817
rect 12800 851 12880 885
rect 12800 817 12823 851
rect 12857 817 12880 851
rect 12800 800 12880 817
rect 8160 777 12880 800
rect 8160 743 8293 777
rect 8327 743 8361 777
rect 8395 743 8429 777
rect 8463 743 8497 777
rect 8531 743 8565 777
rect 8599 743 8633 777
rect 8667 743 8701 777
rect 8735 743 8769 777
rect 8803 743 8837 777
rect 8871 743 8905 777
rect 8939 743 8973 777
rect 9007 743 9041 777
rect 9075 743 9109 777
rect 9143 743 9177 777
rect 9211 743 9245 777
rect 9279 743 9313 777
rect 9347 743 9381 777
rect 9415 743 9449 777
rect 9483 743 9517 777
rect 9551 743 9585 777
rect 9619 743 9653 777
rect 9687 743 9721 777
rect 9755 743 9789 777
rect 9823 743 9857 777
rect 9891 743 9925 777
rect 9959 743 9993 777
rect 10027 743 10061 777
rect 10095 743 10129 777
rect 10163 743 10197 777
rect 10231 743 10265 777
rect 10299 743 10333 777
rect 10367 743 10401 777
rect 10435 743 10469 777
rect 10503 743 10537 777
rect 10571 743 10605 777
rect 10639 743 10673 777
rect 10707 743 10741 777
rect 10775 743 10809 777
rect 10843 743 10877 777
rect 10911 743 10945 777
rect 10979 743 11013 777
rect 11047 743 11081 777
rect 11115 743 11149 777
rect 11183 743 11217 777
rect 11251 743 11285 777
rect 11319 743 11353 777
rect 11387 743 11421 777
rect 11455 743 11489 777
rect 11523 743 11557 777
rect 11591 743 11625 777
rect 11659 743 11693 777
rect 11727 743 11761 777
rect 11795 743 11829 777
rect 11863 743 11897 777
rect 11931 743 11965 777
rect 11999 743 12033 777
rect 12067 743 12101 777
rect 12135 743 12169 777
rect 12203 743 12237 777
rect 12271 743 12305 777
rect 12339 743 12373 777
rect 12407 743 12441 777
rect 12475 743 12509 777
rect 12543 743 12577 777
rect 12611 743 12645 777
rect 12679 743 12713 777
rect 12747 743 12880 777
rect 8160 720 12880 743
rect -320 297 4400 320
rect -320 263 -187 297
rect -153 263 -119 297
rect -85 263 -51 297
rect -17 263 17 297
rect 51 263 85 297
rect 119 263 153 297
rect 187 263 221 297
rect 255 263 289 297
rect 323 263 357 297
rect 391 263 425 297
rect 459 263 493 297
rect 527 263 561 297
rect 595 263 629 297
rect 663 263 697 297
rect 731 263 765 297
rect 799 263 833 297
rect 867 263 901 297
rect 935 263 969 297
rect 1003 263 1037 297
rect 1071 263 1105 297
rect 1139 263 1173 297
rect 1207 263 1241 297
rect 1275 263 1309 297
rect 1343 263 1377 297
rect 1411 263 1445 297
rect 1479 263 1513 297
rect 1547 263 1581 297
rect 1615 263 1649 297
rect 1683 263 1717 297
rect 1751 263 1785 297
rect 1819 263 1853 297
rect 1887 263 1921 297
rect 1955 263 1989 297
rect 2023 263 2057 297
rect 2091 263 2125 297
rect 2159 263 2193 297
rect 2227 263 2261 297
rect 2295 263 2329 297
rect 2363 263 2397 297
rect 2431 263 2465 297
rect 2499 263 2533 297
rect 2567 263 2601 297
rect 2635 263 2669 297
rect 2703 263 2737 297
rect 2771 263 2805 297
rect 2839 263 2873 297
rect 2907 263 2941 297
rect 2975 263 3009 297
rect 3043 263 3077 297
rect 3111 263 3145 297
rect 3179 263 3213 297
rect 3247 263 3281 297
rect 3315 263 3349 297
rect 3383 263 3417 297
rect 3451 263 3485 297
rect 3519 263 3553 297
rect 3587 263 3621 297
rect 3655 263 3689 297
rect 3723 263 3757 297
rect 3791 263 3825 297
rect 3859 263 3893 297
rect 3927 263 3961 297
rect 3995 263 4029 297
rect 4063 263 4097 297
rect 4131 263 4165 297
rect 4199 263 4233 297
rect 4267 263 4400 297
rect -320 240 4400 263
rect -320 223 -240 240
rect -320 189 -297 223
rect -263 189 -240 223
rect -320 155 -240 189
rect 4320 223 4400 240
rect 4320 189 4343 223
rect 4377 189 4400 223
rect -320 121 -297 155
rect -263 121 -240 155
rect -320 87 -240 121
rect -320 53 -297 87
rect -263 53 -240 87
rect -320 19 -240 53
rect -320 -15 -297 19
rect -263 -15 -240 19
rect 4320 155 4400 189
rect 4320 121 4343 155
rect 4377 121 4400 155
rect 4320 87 4400 121
rect 4320 53 4343 87
rect 4377 53 4400 87
rect 4320 19 4400 53
rect -320 -49 -240 -15
rect -320 -83 -297 -49
rect -263 -83 -240 -49
rect 4320 -15 4343 19
rect 4377 -15 4400 19
rect 4320 -49 4400 -15
rect -320 -117 -240 -83
rect 4320 -83 4343 -49
rect 4377 -83 4400 -49
rect -320 -151 -297 -117
rect -263 -151 -240 -117
rect -320 -185 -240 -151
rect 4320 -117 4400 -83
rect 4320 -151 4343 -117
rect 4377 -151 4400 -117
rect -320 -219 -297 -185
rect -263 -219 -240 -185
rect -320 -253 -240 -219
rect -320 -287 -297 -253
rect -263 -287 -240 -253
rect -320 -321 -240 -287
rect 4320 -185 4400 -151
rect 4320 -219 4343 -185
rect 4377 -219 4400 -185
rect 4320 -253 4400 -219
rect 4320 -287 4343 -253
rect 4377 -287 4400 -253
rect -320 -355 -297 -321
rect -263 -355 -240 -321
rect -320 -389 -240 -355
rect -320 -423 -297 -389
rect -263 -423 -240 -389
rect 4320 -321 4400 -287
rect 4320 -355 4343 -321
rect 4377 -355 4400 -321
rect 4320 -389 4400 -355
rect -320 -480 -240 -423
rect 4320 -423 4343 -389
rect 4377 -423 4400 -389
rect 4320 -480 4400 -423
rect -320 -503 4400 -480
rect -320 -537 -187 -503
rect -153 -537 -119 -503
rect -85 -537 -51 -503
rect -17 -537 17 -503
rect 51 -537 85 -503
rect 119 -537 153 -503
rect 187 -537 221 -503
rect 255 -537 289 -503
rect 323 -537 357 -503
rect 391 -537 425 -503
rect 459 -537 493 -503
rect 527 -537 561 -503
rect 595 -537 629 -503
rect 663 -537 697 -503
rect 731 -537 765 -503
rect 799 -537 833 -503
rect 867 -537 901 -503
rect 935 -537 969 -503
rect 1003 -537 1037 -503
rect 1071 -537 1105 -503
rect 1139 -537 1173 -503
rect 1207 -537 1241 -503
rect 1275 -537 1309 -503
rect 1343 -537 1377 -503
rect 1411 -537 1445 -503
rect 1479 -537 1513 -503
rect 1547 -537 1581 -503
rect 1615 -537 1649 -503
rect 1683 -537 1717 -503
rect 1751 -537 1785 -503
rect 1819 -537 1853 -503
rect 1887 -537 1921 -503
rect 1955 -537 1989 -503
rect 2023 -537 2057 -503
rect 2091 -537 2125 -503
rect 2159 -537 2193 -503
rect 2227 -537 2261 -503
rect 2295 -537 2329 -503
rect 2363 -537 2397 -503
rect 2431 -537 2465 -503
rect 2499 -537 2533 -503
rect 2567 -537 2601 -503
rect 2635 -537 2669 -503
rect 2703 -537 2737 -503
rect 2771 -537 2805 -503
rect 2839 -537 2873 -503
rect 2907 -537 2941 -503
rect 2975 -537 3009 -503
rect 3043 -537 3077 -503
rect 3111 -537 3145 -503
rect 3179 -537 3213 -503
rect 3247 -537 3281 -503
rect 3315 -537 3349 -503
rect 3383 -537 3417 -503
rect 3451 -537 3485 -503
rect 3519 -537 3553 -503
rect 3587 -537 3621 -503
rect 3655 -537 3689 -503
rect 3723 -537 3757 -503
rect 3791 -537 3825 -503
rect 3859 -537 3893 -503
rect 3927 -537 3961 -503
rect 3995 -537 4029 -503
rect 4063 -537 4097 -503
rect 4131 -537 4165 -503
rect 4199 -537 4233 -503
rect 4267 -537 4400 -503
rect -320 -560 4400 -537
rect 8160 297 12880 320
rect 8160 263 8293 297
rect 8327 263 8361 297
rect 8395 263 8429 297
rect 8463 263 8497 297
rect 8531 263 8565 297
rect 8599 263 8633 297
rect 8667 263 8701 297
rect 8735 263 8769 297
rect 8803 263 8837 297
rect 8871 263 8905 297
rect 8939 263 8973 297
rect 9007 263 9041 297
rect 9075 263 9109 297
rect 9143 263 9177 297
rect 9211 263 9245 297
rect 9279 263 9313 297
rect 9347 263 9381 297
rect 9415 263 9449 297
rect 9483 263 9517 297
rect 9551 263 9585 297
rect 9619 263 9653 297
rect 9687 263 9721 297
rect 9755 263 9789 297
rect 9823 263 9857 297
rect 9891 263 9925 297
rect 9959 263 9993 297
rect 10027 263 10061 297
rect 10095 263 10129 297
rect 10163 263 10197 297
rect 10231 263 10265 297
rect 10299 263 10333 297
rect 10367 263 10401 297
rect 10435 263 10469 297
rect 10503 263 10537 297
rect 10571 263 10605 297
rect 10639 263 10673 297
rect 10707 263 10741 297
rect 10775 263 10809 297
rect 10843 263 10877 297
rect 10911 263 10945 297
rect 10979 263 11013 297
rect 11047 263 11081 297
rect 11115 263 11149 297
rect 11183 263 11217 297
rect 11251 263 11285 297
rect 11319 263 11353 297
rect 11387 263 11421 297
rect 11455 263 11489 297
rect 11523 263 11557 297
rect 11591 263 11625 297
rect 11659 263 11693 297
rect 11727 263 11761 297
rect 11795 263 11829 297
rect 11863 263 11897 297
rect 11931 263 11965 297
rect 11999 263 12033 297
rect 12067 263 12101 297
rect 12135 263 12169 297
rect 12203 263 12237 297
rect 12271 263 12305 297
rect 12339 263 12373 297
rect 12407 263 12441 297
rect 12475 263 12509 297
rect 12543 263 12577 297
rect 12611 263 12645 297
rect 12679 263 12713 297
rect 12747 263 12880 297
rect 8160 240 12880 263
rect 8160 223 8240 240
rect 8160 189 8183 223
rect 8217 189 8240 223
rect 8160 155 8240 189
rect 12800 223 12880 240
rect 12800 189 12823 223
rect 12857 189 12880 223
rect 8160 121 8183 155
rect 8217 121 8240 155
rect 8160 87 8240 121
rect 8160 53 8183 87
rect 8217 53 8240 87
rect 8160 19 8240 53
rect 8160 -15 8183 19
rect 8217 -15 8240 19
rect 12800 155 12880 189
rect 12800 121 12823 155
rect 12857 121 12880 155
rect 12800 87 12880 121
rect 12800 53 12823 87
rect 12857 53 12880 87
rect 12800 19 12880 53
rect 8160 -49 8240 -15
rect 8160 -83 8183 -49
rect 8217 -83 8240 -49
rect 12800 -15 12823 19
rect 12857 -15 12880 19
rect 12800 -49 12880 -15
rect 8160 -117 8240 -83
rect 12800 -83 12823 -49
rect 12857 -83 12880 -49
rect 8160 -151 8183 -117
rect 8217 -151 8240 -117
rect 8160 -185 8240 -151
rect 12800 -117 12880 -83
rect 12800 -151 12823 -117
rect 12857 -151 12880 -117
rect 8160 -219 8183 -185
rect 8217 -219 8240 -185
rect 8160 -253 8240 -219
rect 8160 -287 8183 -253
rect 8217 -287 8240 -253
rect 8160 -321 8240 -287
rect 12800 -185 12880 -151
rect 12800 -219 12823 -185
rect 12857 -219 12880 -185
rect 12800 -253 12880 -219
rect 12800 -287 12823 -253
rect 12857 -287 12880 -253
rect 8160 -355 8183 -321
rect 8217 -355 8240 -321
rect 8160 -389 8240 -355
rect 8160 -423 8183 -389
rect 8217 -423 8240 -389
rect 12800 -321 12880 -287
rect 12800 -355 12823 -321
rect 12857 -355 12880 -321
rect 12800 -389 12880 -355
rect 8160 -480 8240 -423
rect 12800 -423 12823 -389
rect 12857 -423 12880 -389
rect 12800 -480 12880 -423
rect 8160 -503 12880 -480
rect 8160 -537 8293 -503
rect 8327 -537 8361 -503
rect 8395 -537 8429 -503
rect 8463 -537 8497 -503
rect 8531 -537 8565 -503
rect 8599 -537 8633 -503
rect 8667 -537 8701 -503
rect 8735 -537 8769 -503
rect 8803 -537 8837 -503
rect 8871 -537 8905 -503
rect 8939 -537 8973 -503
rect 9007 -537 9041 -503
rect 9075 -537 9109 -503
rect 9143 -537 9177 -503
rect 9211 -537 9245 -503
rect 9279 -537 9313 -503
rect 9347 -537 9381 -503
rect 9415 -537 9449 -503
rect 9483 -537 9517 -503
rect 9551 -537 9585 -503
rect 9619 -537 9653 -503
rect 9687 -537 9721 -503
rect 9755 -537 9789 -503
rect 9823 -537 9857 -503
rect 9891 -537 9925 -503
rect 9959 -537 9993 -503
rect 10027 -537 10061 -503
rect 10095 -537 10129 -503
rect 10163 -537 10197 -503
rect 10231 -537 10265 -503
rect 10299 -537 10333 -503
rect 10367 -537 10401 -503
rect 10435 -537 10469 -503
rect 10503 -537 10537 -503
rect 10571 -537 10605 -503
rect 10639 -537 10673 -503
rect 10707 -537 10741 -503
rect 10775 -537 10809 -503
rect 10843 -537 10877 -503
rect 10911 -537 10945 -503
rect 10979 -537 11013 -503
rect 11047 -537 11081 -503
rect 11115 -537 11149 -503
rect 11183 -537 11217 -503
rect 11251 -537 11285 -503
rect 11319 -537 11353 -503
rect 11387 -537 11421 -503
rect 11455 -537 11489 -503
rect 11523 -537 11557 -503
rect 11591 -537 11625 -503
rect 11659 -537 11693 -503
rect 11727 -537 11761 -503
rect 11795 -537 11829 -503
rect 11863 -537 11897 -503
rect 11931 -537 11965 -503
rect 11999 -537 12033 -503
rect 12067 -537 12101 -503
rect 12135 -537 12169 -503
rect 12203 -537 12237 -503
rect 12271 -537 12305 -503
rect 12339 -537 12373 -503
rect 12407 -537 12441 -503
rect 12475 -537 12509 -503
rect 12543 -537 12577 -503
rect 12611 -537 12645 -503
rect 12679 -537 12713 -503
rect 12747 -537 12880 -503
rect 8160 -560 12880 -537
<< psubdiffcont >>
rect -357 4263 -323 4297
rect -289 4263 -255 4297
rect -221 4263 -187 4297
rect -153 4263 -119 4297
rect -85 4263 -51 4297
rect -17 4263 17 4297
rect 51 4263 85 4297
rect 119 4263 153 4297
rect 187 4263 221 4297
rect 255 4263 289 4297
rect 323 4263 357 4297
rect 391 4263 425 4297
rect 459 4263 493 4297
rect 527 4263 561 4297
rect 595 4263 629 4297
rect 663 4263 697 4297
rect 731 4263 765 4297
rect 799 4263 833 4297
rect 867 4263 901 4297
rect 935 4263 969 4297
rect 1003 4263 1037 4297
rect 1071 4263 1105 4297
rect 1139 4263 1173 4297
rect 1207 4263 1241 4297
rect 1275 4263 1309 4297
rect 1343 4263 1377 4297
rect 1411 4263 1445 4297
rect 1479 4263 1513 4297
rect 1547 4263 1581 4297
rect 1615 4263 1649 4297
rect 1683 4263 1717 4297
rect 1751 4263 1785 4297
rect 1819 4263 1853 4297
rect 1887 4263 1921 4297
rect 1955 4263 1989 4297
rect 2023 4263 2057 4297
rect 2091 4263 2125 4297
rect 2159 4263 2193 4297
rect 2227 4263 2261 4297
rect 2295 4263 2329 4297
rect 2363 4263 2397 4297
rect 2431 4263 2465 4297
rect 2499 4263 2533 4297
rect 2567 4263 2601 4297
rect 2635 4263 2669 4297
rect 2703 4263 2737 4297
rect 2771 4263 2805 4297
rect 2839 4263 2873 4297
rect 2907 4263 2941 4297
rect 2975 4263 3009 4297
rect 3043 4263 3077 4297
rect 3111 4263 3145 4297
rect 3179 4263 3213 4297
rect 3247 4263 3281 4297
rect 3315 4263 3349 4297
rect 3383 4263 3417 4297
rect 3451 4263 3485 4297
rect 3519 4263 3553 4297
rect 3587 4263 3621 4297
rect 3655 4263 3689 4297
rect 3723 4263 3757 4297
rect 3791 4263 3825 4297
rect 3859 4263 3893 4297
rect 3927 4263 3961 4297
rect 3995 4263 4029 4297
rect 4063 4263 4097 4297
rect 4131 4263 4165 4297
rect 4199 4263 4233 4297
rect 4267 4263 4301 4297
rect 4335 4263 4369 4297
rect 4403 4263 4437 4297
rect -457 4165 -423 4199
rect 4503 4165 4537 4199
rect -457 4097 -423 4131
rect -457 4029 -423 4063
rect -457 3961 -423 3995
rect -457 3893 -423 3927
rect -457 3825 -423 3859
rect -457 3757 -423 3791
rect -457 3689 -423 3723
rect -457 3621 -423 3655
rect -457 3553 -423 3587
rect -457 3485 -423 3519
rect -457 3417 -423 3451
rect -457 3349 -423 3383
rect -457 3281 -423 3315
rect 4503 4097 4537 4131
rect 4503 4029 4537 4063
rect 4503 3961 4537 3995
rect 4503 3893 4537 3927
rect 4503 3825 4537 3859
rect 4503 3757 4537 3791
rect 4503 3689 4537 3723
rect 4503 3621 4537 3655
rect 4503 3553 4537 3587
rect 4503 3485 4537 3519
rect 4503 3417 4537 3451
rect 4503 3349 4537 3383
rect 4503 3281 4537 3315
rect -357 3143 -323 3177
rect -289 3143 -255 3177
rect -221 3143 -187 3177
rect -153 3143 -119 3177
rect -85 3143 -51 3177
rect -17 3143 17 3177
rect 51 3143 85 3177
rect 119 3143 153 3177
rect 187 3143 221 3177
rect 255 3143 289 3177
rect 323 3143 357 3177
rect 391 3143 425 3177
rect 459 3143 493 3177
rect 527 3143 561 3177
rect 595 3143 629 3177
rect 663 3143 697 3177
rect 731 3143 765 3177
rect 799 3143 833 3177
rect 867 3143 901 3177
rect 935 3143 969 3177
rect 1003 3143 1037 3177
rect 1071 3143 1105 3177
rect 1139 3143 1173 3177
rect 1207 3143 1241 3177
rect 1275 3143 1309 3177
rect 1343 3143 1377 3177
rect 1411 3143 1445 3177
rect 1479 3143 1513 3177
rect 1547 3143 1581 3177
rect 1615 3143 1649 3177
rect 1683 3143 1717 3177
rect 1751 3143 1785 3177
rect 1819 3143 1853 3177
rect 1887 3143 1921 3177
rect 1955 3143 1989 3177
rect 2023 3143 2057 3177
rect 2091 3143 2125 3177
rect 2159 3143 2193 3177
rect 2227 3143 2261 3177
rect 2295 3143 2329 3177
rect 2363 3143 2397 3177
rect 2431 3143 2465 3177
rect 2499 3143 2533 3177
rect 2567 3143 2601 3177
rect 2635 3143 2669 3177
rect 2703 3143 2737 3177
rect 2771 3143 2805 3177
rect 2839 3143 2873 3177
rect 2907 3143 2941 3177
rect 2975 3143 3009 3177
rect 3043 3143 3077 3177
rect 3111 3143 3145 3177
rect 3179 3143 3213 3177
rect 3247 3143 3281 3177
rect 3315 3143 3349 3177
rect 3383 3143 3417 3177
rect 3451 3143 3485 3177
rect 3519 3143 3553 3177
rect 3587 3143 3621 3177
rect 3655 3143 3689 3177
rect 3723 3143 3757 3177
rect 3791 3143 3825 3177
rect 3859 3143 3893 3177
rect 3927 3143 3961 3177
rect 3995 3143 4029 3177
rect 4063 3143 4097 3177
rect 4131 3143 4165 3177
rect 4199 3143 4233 3177
rect 4267 3143 4301 3177
rect 4335 3143 4369 3177
rect 4403 3143 4437 3177
rect 8123 4263 8157 4297
rect 8191 4263 8225 4297
rect 8259 4263 8293 4297
rect 8327 4263 8361 4297
rect 8395 4263 8429 4297
rect 8463 4263 8497 4297
rect 8531 4263 8565 4297
rect 8599 4263 8633 4297
rect 8667 4263 8701 4297
rect 8735 4263 8769 4297
rect 8803 4263 8837 4297
rect 8871 4263 8905 4297
rect 8939 4263 8973 4297
rect 9007 4263 9041 4297
rect 9075 4263 9109 4297
rect 9143 4263 9177 4297
rect 9211 4263 9245 4297
rect 9279 4263 9313 4297
rect 9347 4263 9381 4297
rect 9415 4263 9449 4297
rect 9483 4263 9517 4297
rect 9551 4263 9585 4297
rect 9619 4263 9653 4297
rect 9687 4263 9721 4297
rect 9755 4263 9789 4297
rect 9823 4263 9857 4297
rect 9891 4263 9925 4297
rect 9959 4263 9993 4297
rect 10027 4263 10061 4297
rect 10095 4263 10129 4297
rect 10163 4263 10197 4297
rect 10231 4263 10265 4297
rect 10299 4263 10333 4297
rect 10367 4263 10401 4297
rect 10435 4263 10469 4297
rect 10503 4263 10537 4297
rect 10571 4263 10605 4297
rect 10639 4263 10673 4297
rect 10707 4263 10741 4297
rect 10775 4263 10809 4297
rect 10843 4263 10877 4297
rect 10911 4263 10945 4297
rect 10979 4263 11013 4297
rect 11047 4263 11081 4297
rect 11115 4263 11149 4297
rect 11183 4263 11217 4297
rect 11251 4263 11285 4297
rect 11319 4263 11353 4297
rect 11387 4263 11421 4297
rect 11455 4263 11489 4297
rect 11523 4263 11557 4297
rect 11591 4263 11625 4297
rect 11659 4263 11693 4297
rect 11727 4263 11761 4297
rect 11795 4263 11829 4297
rect 11863 4263 11897 4297
rect 11931 4263 11965 4297
rect 11999 4263 12033 4297
rect 12067 4263 12101 4297
rect 12135 4263 12169 4297
rect 12203 4263 12237 4297
rect 12271 4263 12305 4297
rect 12339 4263 12373 4297
rect 12407 4263 12441 4297
rect 12475 4263 12509 4297
rect 12543 4263 12577 4297
rect 12611 4263 12645 4297
rect 12679 4263 12713 4297
rect 12747 4263 12781 4297
rect 12815 4263 12849 4297
rect 12883 4263 12917 4297
rect 8023 4165 8057 4199
rect 12983 4165 13017 4199
rect 8023 4097 8057 4131
rect 8023 4029 8057 4063
rect 8023 3961 8057 3995
rect 8023 3893 8057 3927
rect 8023 3825 8057 3859
rect 8023 3757 8057 3791
rect 8023 3689 8057 3723
rect 8023 3621 8057 3655
rect 8023 3553 8057 3587
rect 8023 3485 8057 3519
rect 8023 3417 8057 3451
rect 8023 3349 8057 3383
rect 8023 3281 8057 3315
rect 12983 4097 13017 4131
rect 12983 4029 13017 4063
rect 12983 3961 13017 3995
rect 12983 3893 13017 3927
rect 12983 3825 13017 3859
rect 12983 3757 13017 3791
rect 12983 3689 13017 3723
rect 12983 3621 13017 3655
rect 12983 3553 13017 3587
rect 12983 3485 13017 3519
rect 12983 3417 13017 3451
rect 12983 3349 13017 3383
rect 12983 3281 13017 3315
rect 8123 3143 8157 3177
rect 8191 3143 8225 3177
rect 8259 3143 8293 3177
rect 8327 3143 8361 3177
rect 8395 3143 8429 3177
rect 8463 3143 8497 3177
rect 8531 3143 8565 3177
rect 8599 3143 8633 3177
rect 8667 3143 8701 3177
rect 8735 3143 8769 3177
rect 8803 3143 8837 3177
rect 8871 3143 8905 3177
rect 8939 3143 8973 3177
rect 9007 3143 9041 3177
rect 9075 3143 9109 3177
rect 9143 3143 9177 3177
rect 9211 3143 9245 3177
rect 9279 3143 9313 3177
rect 9347 3143 9381 3177
rect 9415 3143 9449 3177
rect 9483 3143 9517 3177
rect 9551 3143 9585 3177
rect 9619 3143 9653 3177
rect 9687 3143 9721 3177
rect 9755 3143 9789 3177
rect 9823 3143 9857 3177
rect 9891 3143 9925 3177
rect 9959 3143 9993 3177
rect 10027 3143 10061 3177
rect 10095 3143 10129 3177
rect 10163 3143 10197 3177
rect 10231 3143 10265 3177
rect 10299 3143 10333 3177
rect 10367 3143 10401 3177
rect 10435 3143 10469 3177
rect 10503 3143 10537 3177
rect 10571 3143 10605 3177
rect 10639 3143 10673 3177
rect 10707 3143 10741 3177
rect 10775 3143 10809 3177
rect 10843 3143 10877 3177
rect 10911 3143 10945 3177
rect 10979 3143 11013 3177
rect 11047 3143 11081 3177
rect 11115 3143 11149 3177
rect 11183 3143 11217 3177
rect 11251 3143 11285 3177
rect 11319 3143 11353 3177
rect 11387 3143 11421 3177
rect 11455 3143 11489 3177
rect 11523 3143 11557 3177
rect 11591 3143 11625 3177
rect 11659 3143 11693 3177
rect 11727 3143 11761 3177
rect 11795 3143 11829 3177
rect 11863 3143 11897 3177
rect 11931 3143 11965 3177
rect 11999 3143 12033 3177
rect 12067 3143 12101 3177
rect 12135 3143 12169 3177
rect 12203 3143 12237 3177
rect 12271 3143 12305 3177
rect 12339 3143 12373 3177
rect 12407 3143 12441 3177
rect 12475 3143 12509 3177
rect 12543 3143 12577 3177
rect 12611 3143 12645 3177
rect 12679 3143 12713 3177
rect 12747 3143 12781 3177
rect 12815 3143 12849 3177
rect 12883 3143 12917 3177
rect -357 2983 -323 3017
rect -289 2983 -255 3017
rect -221 2983 -187 3017
rect -153 2983 -119 3017
rect -85 2983 -51 3017
rect -17 2983 17 3017
rect 51 2983 85 3017
rect 119 2983 153 3017
rect 187 2983 221 3017
rect 255 2983 289 3017
rect 323 2983 357 3017
rect 391 2983 425 3017
rect 459 2983 493 3017
rect 527 2983 561 3017
rect 595 2983 629 3017
rect 663 2983 697 3017
rect 731 2983 765 3017
rect 799 2983 833 3017
rect 867 2983 901 3017
rect 935 2983 969 3017
rect 1003 2983 1037 3017
rect 1071 2983 1105 3017
rect 1139 2983 1173 3017
rect 1207 2983 1241 3017
rect 1275 2983 1309 3017
rect 1343 2983 1377 3017
rect 1411 2983 1445 3017
rect 1479 2983 1513 3017
rect 1547 2983 1581 3017
rect 1615 2983 1649 3017
rect 1683 2983 1717 3017
rect 1751 2983 1785 3017
rect 1819 2983 1853 3017
rect 1887 2983 1921 3017
rect 1955 2983 1989 3017
rect 2023 2983 2057 3017
rect 2091 2983 2125 3017
rect 2159 2983 2193 3017
rect 2227 2983 2261 3017
rect 2295 2983 2329 3017
rect 2363 2983 2397 3017
rect 2431 2983 2465 3017
rect 2499 2983 2533 3017
rect 2567 2983 2601 3017
rect 2635 2983 2669 3017
rect 2703 2983 2737 3017
rect 2771 2983 2805 3017
rect 2839 2983 2873 3017
rect 2907 2983 2941 3017
rect 2975 2983 3009 3017
rect 3043 2983 3077 3017
rect 3111 2983 3145 3017
rect 3179 2983 3213 3017
rect 3247 2983 3281 3017
rect 3315 2983 3349 3017
rect 3383 2983 3417 3017
rect 3451 2983 3485 3017
rect 3519 2983 3553 3017
rect 3587 2983 3621 3017
rect 3655 2983 3689 3017
rect 3723 2983 3757 3017
rect 3791 2983 3825 3017
rect 3859 2983 3893 3017
rect 3927 2983 3961 3017
rect 3995 2983 4029 3017
rect 4063 2983 4097 3017
rect 4131 2983 4165 3017
rect 4199 2983 4233 3017
rect 4267 2983 4301 3017
rect 4335 2983 4369 3017
rect 4403 2983 4437 3017
rect -457 2845 -423 2879
rect -457 2777 -423 2811
rect -457 2709 -423 2743
rect -457 2641 -423 2675
rect -457 2573 -423 2607
rect -457 2505 -423 2539
rect -457 2437 -423 2471
rect -457 2369 -423 2403
rect -457 2301 -423 2335
rect -457 2233 -423 2267
rect -457 2165 -423 2199
rect -457 2097 -423 2131
rect -457 2029 -423 2063
rect 4503 2845 4537 2879
rect 4503 2777 4537 2811
rect 4503 2709 4537 2743
rect 4503 2641 4537 2675
rect 4503 2573 4537 2607
rect 4503 2505 4537 2539
rect 4503 2437 4537 2471
rect 4503 2369 4537 2403
rect 4503 2301 4537 2335
rect 4503 2233 4537 2267
rect 4503 2165 4537 2199
rect 4503 2097 4537 2131
rect 4503 2029 4537 2063
rect -457 1961 -423 1995
rect 4503 1961 4537 1995
rect -357 1863 -323 1897
rect -289 1863 -255 1897
rect -221 1863 -187 1897
rect -153 1863 -119 1897
rect -85 1863 -51 1897
rect -17 1863 17 1897
rect 51 1863 85 1897
rect 119 1863 153 1897
rect 187 1863 221 1897
rect 255 1863 289 1897
rect 323 1863 357 1897
rect 391 1863 425 1897
rect 459 1863 493 1897
rect 527 1863 561 1897
rect 595 1863 629 1897
rect 663 1863 697 1897
rect 731 1863 765 1897
rect 799 1863 833 1897
rect 867 1863 901 1897
rect 935 1863 969 1897
rect 1003 1863 1037 1897
rect 1071 1863 1105 1897
rect 1139 1863 1173 1897
rect 1207 1863 1241 1897
rect 1275 1863 1309 1897
rect 1343 1863 1377 1897
rect 1411 1863 1445 1897
rect 1479 1863 1513 1897
rect 1547 1863 1581 1897
rect 1615 1863 1649 1897
rect 1683 1863 1717 1897
rect 1751 1863 1785 1897
rect 1819 1863 1853 1897
rect 1887 1863 1921 1897
rect 1955 1863 1989 1897
rect 2023 1863 2057 1897
rect 2091 1863 2125 1897
rect 2159 1863 2193 1897
rect 2227 1863 2261 1897
rect 2295 1863 2329 1897
rect 2363 1863 2397 1897
rect 2431 1863 2465 1897
rect 2499 1863 2533 1897
rect 2567 1863 2601 1897
rect 2635 1863 2669 1897
rect 2703 1863 2737 1897
rect 2771 1863 2805 1897
rect 2839 1863 2873 1897
rect 2907 1863 2941 1897
rect 2975 1863 3009 1897
rect 3043 1863 3077 1897
rect 3111 1863 3145 1897
rect 3179 1863 3213 1897
rect 3247 1863 3281 1897
rect 3315 1863 3349 1897
rect 3383 1863 3417 1897
rect 3451 1863 3485 1897
rect 3519 1863 3553 1897
rect 3587 1863 3621 1897
rect 3655 1863 3689 1897
rect 3723 1863 3757 1897
rect 3791 1863 3825 1897
rect 3859 1863 3893 1897
rect 3927 1863 3961 1897
rect 3995 1863 4029 1897
rect 4063 1863 4097 1897
rect 4131 1863 4165 1897
rect 4199 1863 4233 1897
rect 4267 1863 4301 1897
rect 4335 1863 4369 1897
rect 4403 1863 4437 1897
rect 8123 2983 8157 3017
rect 8191 2983 8225 3017
rect 8259 2983 8293 3017
rect 8327 2983 8361 3017
rect 8395 2983 8429 3017
rect 8463 2983 8497 3017
rect 8531 2983 8565 3017
rect 8599 2983 8633 3017
rect 8667 2983 8701 3017
rect 8735 2983 8769 3017
rect 8803 2983 8837 3017
rect 8871 2983 8905 3017
rect 8939 2983 8973 3017
rect 9007 2983 9041 3017
rect 9075 2983 9109 3017
rect 9143 2983 9177 3017
rect 9211 2983 9245 3017
rect 9279 2983 9313 3017
rect 9347 2983 9381 3017
rect 9415 2983 9449 3017
rect 9483 2983 9517 3017
rect 9551 2983 9585 3017
rect 9619 2983 9653 3017
rect 9687 2983 9721 3017
rect 9755 2983 9789 3017
rect 9823 2983 9857 3017
rect 9891 2983 9925 3017
rect 9959 2983 9993 3017
rect 10027 2983 10061 3017
rect 10095 2983 10129 3017
rect 10163 2983 10197 3017
rect 10231 2983 10265 3017
rect 10299 2983 10333 3017
rect 10367 2983 10401 3017
rect 10435 2983 10469 3017
rect 10503 2983 10537 3017
rect 10571 2983 10605 3017
rect 10639 2983 10673 3017
rect 10707 2983 10741 3017
rect 10775 2983 10809 3017
rect 10843 2983 10877 3017
rect 10911 2983 10945 3017
rect 10979 2983 11013 3017
rect 11047 2983 11081 3017
rect 11115 2983 11149 3017
rect 11183 2983 11217 3017
rect 11251 2983 11285 3017
rect 11319 2983 11353 3017
rect 11387 2983 11421 3017
rect 11455 2983 11489 3017
rect 11523 2983 11557 3017
rect 11591 2983 11625 3017
rect 11659 2983 11693 3017
rect 11727 2983 11761 3017
rect 11795 2983 11829 3017
rect 11863 2983 11897 3017
rect 11931 2983 11965 3017
rect 11999 2983 12033 3017
rect 12067 2983 12101 3017
rect 12135 2983 12169 3017
rect 12203 2983 12237 3017
rect 12271 2983 12305 3017
rect 12339 2983 12373 3017
rect 12407 2983 12441 3017
rect 12475 2983 12509 3017
rect 12543 2983 12577 3017
rect 12611 2983 12645 3017
rect 12679 2983 12713 3017
rect 12747 2983 12781 3017
rect 12815 2983 12849 3017
rect 12883 2983 12917 3017
rect 8023 2845 8057 2879
rect 8023 2777 8057 2811
rect 8023 2709 8057 2743
rect 8023 2641 8057 2675
rect 8023 2573 8057 2607
rect 8023 2505 8057 2539
rect 8023 2437 8057 2471
rect 8023 2369 8057 2403
rect 8023 2301 8057 2335
rect 8023 2233 8057 2267
rect 8023 2165 8057 2199
rect 8023 2097 8057 2131
rect 8023 2029 8057 2063
rect 12983 2845 13017 2879
rect 12983 2777 13017 2811
rect 12983 2709 13017 2743
rect 12983 2641 13017 2675
rect 12983 2573 13017 2607
rect 12983 2505 13017 2539
rect 12983 2437 13017 2471
rect 12983 2369 13017 2403
rect 12983 2301 13017 2335
rect 12983 2233 13017 2267
rect 12983 2165 13017 2199
rect 12983 2097 13017 2131
rect 12983 2029 13017 2063
rect 8023 1961 8057 1995
rect 12983 1961 13017 1995
rect 8123 1863 8157 1897
rect 8191 1863 8225 1897
rect 8259 1863 8293 1897
rect 8327 1863 8361 1897
rect 8395 1863 8429 1897
rect 8463 1863 8497 1897
rect 8531 1863 8565 1897
rect 8599 1863 8633 1897
rect 8667 1863 8701 1897
rect 8735 1863 8769 1897
rect 8803 1863 8837 1897
rect 8871 1863 8905 1897
rect 8939 1863 8973 1897
rect 9007 1863 9041 1897
rect 9075 1863 9109 1897
rect 9143 1863 9177 1897
rect 9211 1863 9245 1897
rect 9279 1863 9313 1897
rect 9347 1863 9381 1897
rect 9415 1863 9449 1897
rect 9483 1863 9517 1897
rect 9551 1863 9585 1897
rect 9619 1863 9653 1897
rect 9687 1863 9721 1897
rect 9755 1863 9789 1897
rect 9823 1863 9857 1897
rect 9891 1863 9925 1897
rect 9959 1863 9993 1897
rect 10027 1863 10061 1897
rect 10095 1863 10129 1897
rect 10163 1863 10197 1897
rect 10231 1863 10265 1897
rect 10299 1863 10333 1897
rect 10367 1863 10401 1897
rect 10435 1863 10469 1897
rect 10503 1863 10537 1897
rect 10571 1863 10605 1897
rect 10639 1863 10673 1897
rect 10707 1863 10741 1897
rect 10775 1863 10809 1897
rect 10843 1863 10877 1897
rect 10911 1863 10945 1897
rect 10979 1863 11013 1897
rect 11047 1863 11081 1897
rect 11115 1863 11149 1897
rect 11183 1863 11217 1897
rect 11251 1863 11285 1897
rect 11319 1863 11353 1897
rect 11387 1863 11421 1897
rect 11455 1863 11489 1897
rect 11523 1863 11557 1897
rect 11591 1863 11625 1897
rect 11659 1863 11693 1897
rect 11727 1863 11761 1897
rect 11795 1863 11829 1897
rect 11863 1863 11897 1897
rect 11931 1863 11965 1897
rect 11999 1863 12033 1897
rect 12067 1863 12101 1897
rect 12135 1863 12169 1897
rect 12203 1863 12237 1897
rect 12271 1863 12305 1897
rect 12339 1863 12373 1897
rect 12407 1863 12441 1897
rect 12475 1863 12509 1897
rect 12543 1863 12577 1897
rect 12611 1863 12645 1897
rect 12679 1863 12713 1897
rect 12747 1863 12781 1897
rect 12815 1863 12849 1897
rect 12883 1863 12917 1897
rect -357 1703 -323 1737
rect -289 1703 -255 1737
rect -221 1703 -187 1737
rect -153 1703 -119 1737
rect -85 1703 -51 1737
rect -17 1703 17 1737
rect 51 1703 85 1737
rect 119 1703 153 1737
rect 187 1703 221 1737
rect 255 1703 289 1737
rect 323 1703 357 1737
rect 391 1703 425 1737
rect 459 1703 493 1737
rect 527 1703 561 1737
rect 595 1703 629 1737
rect 663 1703 697 1737
rect 731 1703 765 1737
rect 799 1703 833 1737
rect 867 1703 901 1737
rect 935 1703 969 1737
rect 1003 1703 1037 1737
rect 1071 1703 1105 1737
rect 1139 1703 1173 1737
rect 1207 1703 1241 1737
rect 1275 1703 1309 1737
rect 1343 1703 1377 1737
rect 1411 1703 1445 1737
rect 1479 1703 1513 1737
rect 1547 1703 1581 1737
rect 1615 1703 1649 1737
rect 1683 1703 1717 1737
rect 1751 1703 1785 1737
rect 1819 1703 1853 1737
rect 1887 1703 1921 1737
rect 1955 1703 1989 1737
rect 2023 1703 2057 1737
rect 2091 1703 2125 1737
rect 2159 1703 2193 1737
rect 2227 1703 2261 1737
rect 2295 1703 2329 1737
rect 2363 1703 2397 1737
rect 2431 1703 2465 1737
rect 2499 1703 2533 1737
rect 2567 1703 2601 1737
rect 2635 1703 2669 1737
rect 2703 1703 2737 1737
rect 2771 1703 2805 1737
rect 2839 1703 2873 1737
rect 2907 1703 2941 1737
rect 2975 1703 3009 1737
rect 3043 1703 3077 1737
rect 3111 1703 3145 1737
rect 3179 1703 3213 1737
rect 3247 1703 3281 1737
rect 3315 1703 3349 1737
rect 3383 1703 3417 1737
rect 3451 1703 3485 1737
rect 3519 1703 3553 1737
rect 3587 1703 3621 1737
rect 3655 1703 3689 1737
rect 3723 1703 3757 1737
rect 3791 1703 3825 1737
rect 3859 1703 3893 1737
rect 3927 1703 3961 1737
rect 3995 1703 4029 1737
rect 4063 1703 4097 1737
rect 4131 1703 4165 1737
rect 4199 1703 4233 1737
rect 4267 1703 4301 1737
rect 4335 1703 4369 1737
rect 4403 1703 4437 1737
rect -457 1605 -423 1639
rect 4503 1605 4537 1639
rect -457 1537 -423 1571
rect -457 1469 -423 1503
rect -457 1401 -423 1435
rect -457 1333 -423 1367
rect -457 1265 -423 1299
rect -457 1197 -423 1231
rect -457 1129 -423 1163
rect -457 1061 -423 1095
rect -457 993 -423 1027
rect -457 925 -423 959
rect -457 857 -423 891
rect -457 789 -423 823
rect -457 721 -423 755
rect 4503 1537 4537 1571
rect 4503 1469 4537 1503
rect 4503 1401 4537 1435
rect 4503 1333 4537 1367
rect 4503 1265 4537 1299
rect 4503 1197 4537 1231
rect 4503 1129 4537 1163
rect 4503 1061 4537 1095
rect 4503 993 4537 1027
rect 4503 925 4537 959
rect 4503 857 4537 891
rect 4503 789 4537 823
rect 4503 721 4537 755
rect -357 583 -323 617
rect -289 583 -255 617
rect -221 583 -187 617
rect -153 583 -119 617
rect -85 583 -51 617
rect -17 583 17 617
rect 51 583 85 617
rect 119 583 153 617
rect 187 583 221 617
rect 255 583 289 617
rect 323 583 357 617
rect 391 583 425 617
rect 459 583 493 617
rect 527 583 561 617
rect 595 583 629 617
rect 663 583 697 617
rect 731 583 765 617
rect 799 583 833 617
rect 867 583 901 617
rect 935 583 969 617
rect 1003 583 1037 617
rect 1071 583 1105 617
rect 1139 583 1173 617
rect 1207 583 1241 617
rect 1275 583 1309 617
rect 1343 583 1377 617
rect 1411 583 1445 617
rect 1479 583 1513 617
rect 1547 583 1581 617
rect 1615 583 1649 617
rect 1683 583 1717 617
rect 1751 583 1785 617
rect 1819 583 1853 617
rect 1887 583 1921 617
rect 1955 583 1989 617
rect 2023 583 2057 617
rect 2091 583 2125 617
rect 2159 583 2193 617
rect 2227 583 2261 617
rect 2295 583 2329 617
rect 2363 583 2397 617
rect 2431 583 2465 617
rect 2499 583 2533 617
rect 2567 583 2601 617
rect 2635 583 2669 617
rect 2703 583 2737 617
rect 2771 583 2805 617
rect 2839 583 2873 617
rect 2907 583 2941 617
rect 2975 583 3009 617
rect 3043 583 3077 617
rect 3111 583 3145 617
rect 3179 583 3213 617
rect 3247 583 3281 617
rect 3315 583 3349 617
rect 3383 583 3417 617
rect 3451 583 3485 617
rect 3519 583 3553 617
rect 3587 583 3621 617
rect 3655 583 3689 617
rect 3723 583 3757 617
rect 3791 583 3825 617
rect 3859 583 3893 617
rect 3927 583 3961 617
rect 3995 583 4029 617
rect 4063 583 4097 617
rect 4131 583 4165 617
rect 4199 583 4233 617
rect 4267 583 4301 617
rect 4335 583 4369 617
rect 4403 583 4437 617
rect 8123 1703 8157 1737
rect 8191 1703 8225 1737
rect 8259 1703 8293 1737
rect 8327 1703 8361 1737
rect 8395 1703 8429 1737
rect 8463 1703 8497 1737
rect 8531 1703 8565 1737
rect 8599 1703 8633 1737
rect 8667 1703 8701 1737
rect 8735 1703 8769 1737
rect 8803 1703 8837 1737
rect 8871 1703 8905 1737
rect 8939 1703 8973 1737
rect 9007 1703 9041 1737
rect 9075 1703 9109 1737
rect 9143 1703 9177 1737
rect 9211 1703 9245 1737
rect 9279 1703 9313 1737
rect 9347 1703 9381 1737
rect 9415 1703 9449 1737
rect 9483 1703 9517 1737
rect 9551 1703 9585 1737
rect 9619 1703 9653 1737
rect 9687 1703 9721 1737
rect 9755 1703 9789 1737
rect 9823 1703 9857 1737
rect 9891 1703 9925 1737
rect 9959 1703 9993 1737
rect 10027 1703 10061 1737
rect 10095 1703 10129 1737
rect 10163 1703 10197 1737
rect 10231 1703 10265 1737
rect 10299 1703 10333 1737
rect 10367 1703 10401 1737
rect 10435 1703 10469 1737
rect 10503 1703 10537 1737
rect 10571 1703 10605 1737
rect 10639 1703 10673 1737
rect 10707 1703 10741 1737
rect 10775 1703 10809 1737
rect 10843 1703 10877 1737
rect 10911 1703 10945 1737
rect 10979 1703 11013 1737
rect 11047 1703 11081 1737
rect 11115 1703 11149 1737
rect 11183 1703 11217 1737
rect 11251 1703 11285 1737
rect 11319 1703 11353 1737
rect 11387 1703 11421 1737
rect 11455 1703 11489 1737
rect 11523 1703 11557 1737
rect 11591 1703 11625 1737
rect 11659 1703 11693 1737
rect 11727 1703 11761 1737
rect 11795 1703 11829 1737
rect 11863 1703 11897 1737
rect 11931 1703 11965 1737
rect 11999 1703 12033 1737
rect 12067 1703 12101 1737
rect 12135 1703 12169 1737
rect 12203 1703 12237 1737
rect 12271 1703 12305 1737
rect 12339 1703 12373 1737
rect 12407 1703 12441 1737
rect 12475 1703 12509 1737
rect 12543 1703 12577 1737
rect 12611 1703 12645 1737
rect 12679 1703 12713 1737
rect 12747 1703 12781 1737
rect 12815 1703 12849 1737
rect 12883 1703 12917 1737
rect 8023 1605 8057 1639
rect 12983 1605 13017 1639
rect 8023 1537 8057 1571
rect 8023 1469 8057 1503
rect 8023 1401 8057 1435
rect 8023 1333 8057 1367
rect 8023 1265 8057 1299
rect 8023 1197 8057 1231
rect 8023 1129 8057 1163
rect 8023 1061 8057 1095
rect 8023 993 8057 1027
rect 8023 925 8057 959
rect 8023 857 8057 891
rect 8023 789 8057 823
rect 8023 721 8057 755
rect 12983 1537 13017 1571
rect 12983 1469 13017 1503
rect 12983 1401 13017 1435
rect 12983 1333 13017 1367
rect 12983 1265 13017 1299
rect 12983 1197 13017 1231
rect 12983 1129 13017 1163
rect 12983 1061 13017 1095
rect 12983 993 13017 1027
rect 12983 925 13017 959
rect 12983 857 13017 891
rect 12983 789 13017 823
rect 12983 721 13017 755
rect 8123 583 8157 617
rect 8191 583 8225 617
rect 8259 583 8293 617
rect 8327 583 8361 617
rect 8395 583 8429 617
rect 8463 583 8497 617
rect 8531 583 8565 617
rect 8599 583 8633 617
rect 8667 583 8701 617
rect 8735 583 8769 617
rect 8803 583 8837 617
rect 8871 583 8905 617
rect 8939 583 8973 617
rect 9007 583 9041 617
rect 9075 583 9109 617
rect 9143 583 9177 617
rect 9211 583 9245 617
rect 9279 583 9313 617
rect 9347 583 9381 617
rect 9415 583 9449 617
rect 9483 583 9517 617
rect 9551 583 9585 617
rect 9619 583 9653 617
rect 9687 583 9721 617
rect 9755 583 9789 617
rect 9823 583 9857 617
rect 9891 583 9925 617
rect 9959 583 9993 617
rect 10027 583 10061 617
rect 10095 583 10129 617
rect 10163 583 10197 617
rect 10231 583 10265 617
rect 10299 583 10333 617
rect 10367 583 10401 617
rect 10435 583 10469 617
rect 10503 583 10537 617
rect 10571 583 10605 617
rect 10639 583 10673 617
rect 10707 583 10741 617
rect 10775 583 10809 617
rect 10843 583 10877 617
rect 10911 583 10945 617
rect 10979 583 11013 617
rect 11047 583 11081 617
rect 11115 583 11149 617
rect 11183 583 11217 617
rect 11251 583 11285 617
rect 11319 583 11353 617
rect 11387 583 11421 617
rect 11455 583 11489 617
rect 11523 583 11557 617
rect 11591 583 11625 617
rect 11659 583 11693 617
rect 11727 583 11761 617
rect 11795 583 11829 617
rect 11863 583 11897 617
rect 11931 583 11965 617
rect 11999 583 12033 617
rect 12067 583 12101 617
rect 12135 583 12169 617
rect 12203 583 12237 617
rect 12271 583 12305 617
rect 12339 583 12373 617
rect 12407 583 12441 617
rect 12475 583 12509 617
rect 12543 583 12577 617
rect 12611 583 12645 617
rect 12679 583 12713 617
rect 12747 583 12781 617
rect 12815 583 12849 617
rect 12883 583 12917 617
rect -357 423 -323 457
rect -289 423 -255 457
rect -221 423 -187 457
rect -153 423 -119 457
rect -85 423 -51 457
rect -17 423 17 457
rect 51 423 85 457
rect 119 423 153 457
rect 187 423 221 457
rect 255 423 289 457
rect 323 423 357 457
rect 391 423 425 457
rect 459 423 493 457
rect 527 423 561 457
rect 595 423 629 457
rect 663 423 697 457
rect 731 423 765 457
rect 799 423 833 457
rect 867 423 901 457
rect 935 423 969 457
rect 1003 423 1037 457
rect 1071 423 1105 457
rect 1139 423 1173 457
rect 1207 423 1241 457
rect 1275 423 1309 457
rect 1343 423 1377 457
rect 1411 423 1445 457
rect 1479 423 1513 457
rect 1547 423 1581 457
rect 1615 423 1649 457
rect 1683 423 1717 457
rect 1751 423 1785 457
rect 1819 423 1853 457
rect 1887 423 1921 457
rect 1955 423 1989 457
rect 2023 423 2057 457
rect 2091 423 2125 457
rect 2159 423 2193 457
rect 2227 423 2261 457
rect 2295 423 2329 457
rect 2363 423 2397 457
rect 2431 423 2465 457
rect 2499 423 2533 457
rect 2567 423 2601 457
rect 2635 423 2669 457
rect 2703 423 2737 457
rect 2771 423 2805 457
rect 2839 423 2873 457
rect 2907 423 2941 457
rect 2975 423 3009 457
rect 3043 423 3077 457
rect 3111 423 3145 457
rect 3179 423 3213 457
rect 3247 423 3281 457
rect 3315 423 3349 457
rect 3383 423 3417 457
rect 3451 423 3485 457
rect 3519 423 3553 457
rect 3587 423 3621 457
rect 3655 423 3689 457
rect 3723 423 3757 457
rect 3791 423 3825 457
rect 3859 423 3893 457
rect 3927 423 3961 457
rect 3995 423 4029 457
rect 4063 423 4097 457
rect 4131 423 4165 457
rect 4199 423 4233 457
rect 4267 423 4301 457
rect 4335 423 4369 457
rect 4403 423 4437 457
rect -457 285 -423 319
rect -457 217 -423 251
rect -457 149 -423 183
rect -457 81 -423 115
rect -457 13 -423 47
rect -457 -55 -423 -21
rect -457 -123 -423 -89
rect -457 -191 -423 -157
rect -457 -259 -423 -225
rect -457 -327 -423 -293
rect -457 -395 -423 -361
rect -457 -463 -423 -429
rect -457 -531 -423 -497
rect 4503 285 4537 319
rect 4503 217 4537 251
rect 4503 149 4537 183
rect 4503 81 4537 115
rect 4503 13 4537 47
rect 4503 -55 4537 -21
rect 4503 -123 4537 -89
rect 4503 -191 4537 -157
rect 4503 -259 4537 -225
rect 4503 -327 4537 -293
rect 4503 -395 4537 -361
rect 4503 -463 4537 -429
rect 4503 -531 4537 -497
rect -457 -599 -423 -565
rect 4503 -599 4537 -565
rect -357 -697 -323 -663
rect -289 -697 -255 -663
rect -221 -697 -187 -663
rect -153 -697 -119 -663
rect -85 -697 -51 -663
rect -17 -697 17 -663
rect 51 -697 85 -663
rect 119 -697 153 -663
rect 187 -697 221 -663
rect 255 -697 289 -663
rect 323 -697 357 -663
rect 391 -697 425 -663
rect 459 -697 493 -663
rect 527 -697 561 -663
rect 595 -697 629 -663
rect 663 -697 697 -663
rect 731 -697 765 -663
rect 799 -697 833 -663
rect 867 -697 901 -663
rect 935 -697 969 -663
rect 1003 -697 1037 -663
rect 1071 -697 1105 -663
rect 1139 -697 1173 -663
rect 1207 -697 1241 -663
rect 1275 -697 1309 -663
rect 1343 -697 1377 -663
rect 1411 -697 1445 -663
rect 1479 -697 1513 -663
rect 1547 -697 1581 -663
rect 1615 -697 1649 -663
rect 1683 -697 1717 -663
rect 1751 -697 1785 -663
rect 1819 -697 1853 -663
rect 1887 -697 1921 -663
rect 1955 -697 1989 -663
rect 2023 -697 2057 -663
rect 2091 -697 2125 -663
rect 2159 -697 2193 -663
rect 2227 -697 2261 -663
rect 2295 -697 2329 -663
rect 2363 -697 2397 -663
rect 2431 -697 2465 -663
rect 2499 -697 2533 -663
rect 2567 -697 2601 -663
rect 2635 -697 2669 -663
rect 2703 -697 2737 -663
rect 2771 -697 2805 -663
rect 2839 -697 2873 -663
rect 2907 -697 2941 -663
rect 2975 -697 3009 -663
rect 3043 -697 3077 -663
rect 3111 -697 3145 -663
rect 3179 -697 3213 -663
rect 3247 -697 3281 -663
rect 3315 -697 3349 -663
rect 3383 -697 3417 -663
rect 3451 -697 3485 -663
rect 3519 -697 3553 -663
rect 3587 -697 3621 -663
rect 3655 -697 3689 -663
rect 3723 -697 3757 -663
rect 3791 -697 3825 -663
rect 3859 -697 3893 -663
rect 3927 -697 3961 -663
rect 3995 -697 4029 -663
rect 4063 -697 4097 -663
rect 4131 -697 4165 -663
rect 4199 -697 4233 -663
rect 4267 -697 4301 -663
rect 4335 -697 4369 -663
rect 4403 -697 4437 -663
rect 8123 423 8157 457
rect 8191 423 8225 457
rect 8259 423 8293 457
rect 8327 423 8361 457
rect 8395 423 8429 457
rect 8463 423 8497 457
rect 8531 423 8565 457
rect 8599 423 8633 457
rect 8667 423 8701 457
rect 8735 423 8769 457
rect 8803 423 8837 457
rect 8871 423 8905 457
rect 8939 423 8973 457
rect 9007 423 9041 457
rect 9075 423 9109 457
rect 9143 423 9177 457
rect 9211 423 9245 457
rect 9279 423 9313 457
rect 9347 423 9381 457
rect 9415 423 9449 457
rect 9483 423 9517 457
rect 9551 423 9585 457
rect 9619 423 9653 457
rect 9687 423 9721 457
rect 9755 423 9789 457
rect 9823 423 9857 457
rect 9891 423 9925 457
rect 9959 423 9993 457
rect 10027 423 10061 457
rect 10095 423 10129 457
rect 10163 423 10197 457
rect 10231 423 10265 457
rect 10299 423 10333 457
rect 10367 423 10401 457
rect 10435 423 10469 457
rect 10503 423 10537 457
rect 10571 423 10605 457
rect 10639 423 10673 457
rect 10707 423 10741 457
rect 10775 423 10809 457
rect 10843 423 10877 457
rect 10911 423 10945 457
rect 10979 423 11013 457
rect 11047 423 11081 457
rect 11115 423 11149 457
rect 11183 423 11217 457
rect 11251 423 11285 457
rect 11319 423 11353 457
rect 11387 423 11421 457
rect 11455 423 11489 457
rect 11523 423 11557 457
rect 11591 423 11625 457
rect 11659 423 11693 457
rect 11727 423 11761 457
rect 11795 423 11829 457
rect 11863 423 11897 457
rect 11931 423 11965 457
rect 11999 423 12033 457
rect 12067 423 12101 457
rect 12135 423 12169 457
rect 12203 423 12237 457
rect 12271 423 12305 457
rect 12339 423 12373 457
rect 12407 423 12441 457
rect 12475 423 12509 457
rect 12543 423 12577 457
rect 12611 423 12645 457
rect 12679 423 12713 457
rect 12747 423 12781 457
rect 12815 423 12849 457
rect 12883 423 12917 457
rect 8023 285 8057 319
rect 8023 217 8057 251
rect 8023 149 8057 183
rect 8023 81 8057 115
rect 8023 13 8057 47
rect 8023 -55 8057 -21
rect 8023 -123 8057 -89
rect 8023 -191 8057 -157
rect 8023 -259 8057 -225
rect 8023 -327 8057 -293
rect 8023 -395 8057 -361
rect 8023 -463 8057 -429
rect 8023 -531 8057 -497
rect 12983 285 13017 319
rect 12983 217 13017 251
rect 12983 149 13017 183
rect 12983 81 13017 115
rect 12983 13 13017 47
rect 12983 -55 13017 -21
rect 12983 -123 13017 -89
rect 12983 -191 13017 -157
rect 12983 -259 13017 -225
rect 12983 -327 13017 -293
rect 12983 -395 13017 -361
rect 12983 -463 13017 -429
rect 12983 -531 13017 -497
rect 8023 -599 8057 -565
rect 12983 -599 13017 -565
rect 8123 -697 8157 -663
rect 8191 -697 8225 -663
rect 8259 -697 8293 -663
rect 8327 -697 8361 -663
rect 8395 -697 8429 -663
rect 8463 -697 8497 -663
rect 8531 -697 8565 -663
rect 8599 -697 8633 -663
rect 8667 -697 8701 -663
rect 8735 -697 8769 -663
rect 8803 -697 8837 -663
rect 8871 -697 8905 -663
rect 8939 -697 8973 -663
rect 9007 -697 9041 -663
rect 9075 -697 9109 -663
rect 9143 -697 9177 -663
rect 9211 -697 9245 -663
rect 9279 -697 9313 -663
rect 9347 -697 9381 -663
rect 9415 -697 9449 -663
rect 9483 -697 9517 -663
rect 9551 -697 9585 -663
rect 9619 -697 9653 -663
rect 9687 -697 9721 -663
rect 9755 -697 9789 -663
rect 9823 -697 9857 -663
rect 9891 -697 9925 -663
rect 9959 -697 9993 -663
rect 10027 -697 10061 -663
rect 10095 -697 10129 -663
rect 10163 -697 10197 -663
rect 10231 -697 10265 -663
rect 10299 -697 10333 -663
rect 10367 -697 10401 -663
rect 10435 -697 10469 -663
rect 10503 -697 10537 -663
rect 10571 -697 10605 -663
rect 10639 -697 10673 -663
rect 10707 -697 10741 -663
rect 10775 -697 10809 -663
rect 10843 -697 10877 -663
rect 10911 -697 10945 -663
rect 10979 -697 11013 -663
rect 11047 -697 11081 -663
rect 11115 -697 11149 -663
rect 11183 -697 11217 -663
rect 11251 -697 11285 -663
rect 11319 -697 11353 -663
rect 11387 -697 11421 -663
rect 11455 -697 11489 -663
rect 11523 -697 11557 -663
rect 11591 -697 11625 -663
rect 11659 -697 11693 -663
rect 11727 -697 11761 -663
rect 11795 -697 11829 -663
rect 11863 -697 11897 -663
rect 11931 -697 11965 -663
rect 11999 -697 12033 -663
rect 12067 -697 12101 -663
rect 12135 -697 12169 -663
rect 12203 -697 12237 -663
rect 12271 -697 12305 -663
rect 12339 -697 12373 -663
rect 12407 -697 12441 -663
rect 12475 -697 12509 -663
rect 12543 -697 12577 -663
rect 12611 -697 12645 -663
rect 12679 -697 12713 -663
rect 12747 -697 12781 -663
rect 12815 -697 12849 -663
rect 12883 -697 12917 -663
<< mvnsubdiffcont >>
rect -187 4103 -153 4137
rect -119 4103 -85 4137
rect -51 4103 -17 4137
rect 17 4103 51 4137
rect 85 4103 119 4137
rect 153 4103 187 4137
rect 221 4103 255 4137
rect 289 4103 323 4137
rect 357 4103 391 4137
rect 425 4103 459 4137
rect 493 4103 527 4137
rect 561 4103 595 4137
rect 629 4103 663 4137
rect 697 4103 731 4137
rect 765 4103 799 4137
rect 833 4103 867 4137
rect 901 4103 935 4137
rect 969 4103 1003 4137
rect 1037 4103 1071 4137
rect 1105 4103 1139 4137
rect 1173 4103 1207 4137
rect 1241 4103 1275 4137
rect 1309 4103 1343 4137
rect 1377 4103 1411 4137
rect 1445 4103 1479 4137
rect 1513 4103 1547 4137
rect 1581 4103 1615 4137
rect 1649 4103 1683 4137
rect 1717 4103 1751 4137
rect 1785 4103 1819 4137
rect 1853 4103 1887 4137
rect 1921 4103 1955 4137
rect 1989 4103 2023 4137
rect 2057 4103 2091 4137
rect 2125 4103 2159 4137
rect 2193 4103 2227 4137
rect 2261 4103 2295 4137
rect 2329 4103 2363 4137
rect 2397 4103 2431 4137
rect 2465 4103 2499 4137
rect 2533 4103 2567 4137
rect 2601 4103 2635 4137
rect 2669 4103 2703 4137
rect 2737 4103 2771 4137
rect 2805 4103 2839 4137
rect 2873 4103 2907 4137
rect 2941 4103 2975 4137
rect 3009 4103 3043 4137
rect 3077 4103 3111 4137
rect 3145 4103 3179 4137
rect 3213 4103 3247 4137
rect 3281 4103 3315 4137
rect 3349 4103 3383 4137
rect 3417 4103 3451 4137
rect 3485 4103 3519 4137
rect 3553 4103 3587 4137
rect 3621 4103 3655 4137
rect 3689 4103 3723 4137
rect 3757 4103 3791 4137
rect 3825 4103 3859 4137
rect 3893 4103 3927 4137
rect 3961 4103 3995 4137
rect 4029 4103 4063 4137
rect 4097 4103 4131 4137
rect 4165 4103 4199 4137
rect 4233 4103 4267 4137
rect -297 3989 -263 4023
rect -297 3921 -263 3955
rect 4343 3989 4377 4023
rect 4343 3921 4377 3955
rect -297 3853 -263 3887
rect -297 3785 -263 3819
rect 4343 3853 4377 3887
rect 4343 3785 4377 3819
rect -297 3717 -263 3751
rect 4343 3717 4377 3751
rect -297 3649 -263 3683
rect -297 3581 -263 3615
rect 4343 3649 4377 3683
rect -297 3513 -263 3547
rect -297 3445 -263 3479
rect 4343 3581 4377 3615
rect 4343 3513 4377 3547
rect 4343 3445 4377 3479
rect -297 3377 -263 3411
rect 4343 3377 4377 3411
rect -187 3303 -153 3337
rect -119 3303 -85 3337
rect -51 3303 -17 3337
rect 17 3303 51 3337
rect 85 3303 119 3337
rect 153 3303 187 3337
rect 221 3303 255 3337
rect 289 3303 323 3337
rect 357 3303 391 3337
rect 425 3303 459 3337
rect 493 3303 527 3337
rect 561 3303 595 3337
rect 629 3303 663 3337
rect 697 3303 731 3337
rect 765 3303 799 3337
rect 833 3303 867 3337
rect 901 3303 935 3337
rect 969 3303 1003 3337
rect 1037 3303 1071 3337
rect 1105 3303 1139 3337
rect 1173 3303 1207 3337
rect 1241 3303 1275 3337
rect 1309 3303 1343 3337
rect 1377 3303 1411 3337
rect 1445 3303 1479 3337
rect 1513 3303 1547 3337
rect 1581 3303 1615 3337
rect 1649 3303 1683 3337
rect 1717 3303 1751 3337
rect 1785 3303 1819 3337
rect 1853 3303 1887 3337
rect 1921 3303 1955 3337
rect 1989 3303 2023 3337
rect 2057 3303 2091 3337
rect 2125 3303 2159 3337
rect 2193 3303 2227 3337
rect 2261 3303 2295 3337
rect 2329 3303 2363 3337
rect 2397 3303 2431 3337
rect 2465 3303 2499 3337
rect 2533 3303 2567 3337
rect 2601 3303 2635 3337
rect 2669 3303 2703 3337
rect 2737 3303 2771 3337
rect 2805 3303 2839 3337
rect 2873 3303 2907 3337
rect 2941 3303 2975 3337
rect 3009 3303 3043 3337
rect 3077 3303 3111 3337
rect 3145 3303 3179 3337
rect 3213 3303 3247 3337
rect 3281 3303 3315 3337
rect 3349 3303 3383 3337
rect 3417 3303 3451 3337
rect 3485 3303 3519 3337
rect 3553 3303 3587 3337
rect 3621 3303 3655 3337
rect 3689 3303 3723 3337
rect 3757 3303 3791 3337
rect 3825 3303 3859 3337
rect 3893 3303 3927 3337
rect 3961 3303 3995 3337
rect 4029 3303 4063 3337
rect 4097 3303 4131 3337
rect 4165 3303 4199 3337
rect 4233 3303 4267 3337
rect 8293 4103 8327 4137
rect 8361 4103 8395 4137
rect 8429 4103 8463 4137
rect 8497 4103 8531 4137
rect 8565 4103 8599 4137
rect 8633 4103 8667 4137
rect 8701 4103 8735 4137
rect 8769 4103 8803 4137
rect 8837 4103 8871 4137
rect 8905 4103 8939 4137
rect 8973 4103 9007 4137
rect 9041 4103 9075 4137
rect 9109 4103 9143 4137
rect 9177 4103 9211 4137
rect 9245 4103 9279 4137
rect 9313 4103 9347 4137
rect 9381 4103 9415 4137
rect 9449 4103 9483 4137
rect 9517 4103 9551 4137
rect 9585 4103 9619 4137
rect 9653 4103 9687 4137
rect 9721 4103 9755 4137
rect 9789 4103 9823 4137
rect 9857 4103 9891 4137
rect 9925 4103 9959 4137
rect 9993 4103 10027 4137
rect 10061 4103 10095 4137
rect 10129 4103 10163 4137
rect 10197 4103 10231 4137
rect 10265 4103 10299 4137
rect 10333 4103 10367 4137
rect 10401 4103 10435 4137
rect 10469 4103 10503 4137
rect 10537 4103 10571 4137
rect 10605 4103 10639 4137
rect 10673 4103 10707 4137
rect 10741 4103 10775 4137
rect 10809 4103 10843 4137
rect 10877 4103 10911 4137
rect 10945 4103 10979 4137
rect 11013 4103 11047 4137
rect 11081 4103 11115 4137
rect 11149 4103 11183 4137
rect 11217 4103 11251 4137
rect 11285 4103 11319 4137
rect 11353 4103 11387 4137
rect 11421 4103 11455 4137
rect 11489 4103 11523 4137
rect 11557 4103 11591 4137
rect 11625 4103 11659 4137
rect 11693 4103 11727 4137
rect 11761 4103 11795 4137
rect 11829 4103 11863 4137
rect 11897 4103 11931 4137
rect 11965 4103 11999 4137
rect 12033 4103 12067 4137
rect 12101 4103 12135 4137
rect 12169 4103 12203 4137
rect 12237 4103 12271 4137
rect 12305 4103 12339 4137
rect 12373 4103 12407 4137
rect 12441 4103 12475 4137
rect 12509 4103 12543 4137
rect 12577 4103 12611 4137
rect 12645 4103 12679 4137
rect 12713 4103 12747 4137
rect 8183 3989 8217 4023
rect 8183 3921 8217 3955
rect 12823 3989 12857 4023
rect 12823 3921 12857 3955
rect 8183 3853 8217 3887
rect 8183 3785 8217 3819
rect 12823 3853 12857 3887
rect 12823 3785 12857 3819
rect 8183 3717 8217 3751
rect 12823 3717 12857 3751
rect 8183 3649 8217 3683
rect 8183 3581 8217 3615
rect 12823 3649 12857 3683
rect 8183 3513 8217 3547
rect 8183 3445 8217 3479
rect 12823 3581 12857 3615
rect 12823 3513 12857 3547
rect 12823 3445 12857 3479
rect 8183 3377 8217 3411
rect 12823 3377 12857 3411
rect 8293 3303 8327 3337
rect 8361 3303 8395 3337
rect 8429 3303 8463 3337
rect 8497 3303 8531 3337
rect 8565 3303 8599 3337
rect 8633 3303 8667 3337
rect 8701 3303 8735 3337
rect 8769 3303 8803 3337
rect 8837 3303 8871 3337
rect 8905 3303 8939 3337
rect 8973 3303 9007 3337
rect 9041 3303 9075 3337
rect 9109 3303 9143 3337
rect 9177 3303 9211 3337
rect 9245 3303 9279 3337
rect 9313 3303 9347 3337
rect 9381 3303 9415 3337
rect 9449 3303 9483 3337
rect 9517 3303 9551 3337
rect 9585 3303 9619 3337
rect 9653 3303 9687 3337
rect 9721 3303 9755 3337
rect 9789 3303 9823 3337
rect 9857 3303 9891 3337
rect 9925 3303 9959 3337
rect 9993 3303 10027 3337
rect 10061 3303 10095 3337
rect 10129 3303 10163 3337
rect 10197 3303 10231 3337
rect 10265 3303 10299 3337
rect 10333 3303 10367 3337
rect 10401 3303 10435 3337
rect 10469 3303 10503 3337
rect 10537 3303 10571 3337
rect 10605 3303 10639 3337
rect 10673 3303 10707 3337
rect 10741 3303 10775 3337
rect 10809 3303 10843 3337
rect 10877 3303 10911 3337
rect 10945 3303 10979 3337
rect 11013 3303 11047 3337
rect 11081 3303 11115 3337
rect 11149 3303 11183 3337
rect 11217 3303 11251 3337
rect 11285 3303 11319 3337
rect 11353 3303 11387 3337
rect 11421 3303 11455 3337
rect 11489 3303 11523 3337
rect 11557 3303 11591 3337
rect 11625 3303 11659 3337
rect 11693 3303 11727 3337
rect 11761 3303 11795 3337
rect 11829 3303 11863 3337
rect 11897 3303 11931 3337
rect 11965 3303 11999 3337
rect 12033 3303 12067 3337
rect 12101 3303 12135 3337
rect 12169 3303 12203 3337
rect 12237 3303 12271 3337
rect 12305 3303 12339 3337
rect 12373 3303 12407 3337
rect 12441 3303 12475 3337
rect 12509 3303 12543 3337
rect 12577 3303 12611 3337
rect 12645 3303 12679 3337
rect 12713 3303 12747 3337
rect -187 2823 -153 2857
rect -119 2823 -85 2857
rect -51 2823 -17 2857
rect 17 2823 51 2857
rect 85 2823 119 2857
rect 153 2823 187 2857
rect 221 2823 255 2857
rect 289 2823 323 2857
rect 357 2823 391 2857
rect 425 2823 459 2857
rect 493 2823 527 2857
rect 561 2823 595 2857
rect 629 2823 663 2857
rect 697 2823 731 2857
rect 765 2823 799 2857
rect 833 2823 867 2857
rect 901 2823 935 2857
rect 969 2823 1003 2857
rect 1037 2823 1071 2857
rect 1105 2823 1139 2857
rect 1173 2823 1207 2857
rect 1241 2823 1275 2857
rect 1309 2823 1343 2857
rect 1377 2823 1411 2857
rect 1445 2823 1479 2857
rect 1513 2823 1547 2857
rect 1581 2823 1615 2857
rect 1649 2823 1683 2857
rect 1717 2823 1751 2857
rect 1785 2823 1819 2857
rect 1853 2823 1887 2857
rect 1921 2823 1955 2857
rect 1989 2823 2023 2857
rect 2057 2823 2091 2857
rect 2125 2823 2159 2857
rect 2193 2823 2227 2857
rect 2261 2823 2295 2857
rect 2329 2823 2363 2857
rect 2397 2823 2431 2857
rect 2465 2823 2499 2857
rect 2533 2823 2567 2857
rect 2601 2823 2635 2857
rect 2669 2823 2703 2857
rect 2737 2823 2771 2857
rect 2805 2823 2839 2857
rect 2873 2823 2907 2857
rect 2941 2823 2975 2857
rect 3009 2823 3043 2857
rect 3077 2823 3111 2857
rect 3145 2823 3179 2857
rect 3213 2823 3247 2857
rect 3281 2823 3315 2857
rect 3349 2823 3383 2857
rect 3417 2823 3451 2857
rect 3485 2823 3519 2857
rect 3553 2823 3587 2857
rect 3621 2823 3655 2857
rect 3689 2823 3723 2857
rect 3757 2823 3791 2857
rect 3825 2823 3859 2857
rect 3893 2823 3927 2857
rect 3961 2823 3995 2857
rect 4029 2823 4063 2857
rect 4097 2823 4131 2857
rect 4165 2823 4199 2857
rect 4233 2823 4267 2857
rect -297 2749 -263 2783
rect 4343 2749 4377 2783
rect -297 2681 -263 2715
rect -297 2613 -263 2647
rect -297 2545 -263 2579
rect 4343 2681 4377 2715
rect 4343 2613 4377 2647
rect -297 2477 -263 2511
rect 4343 2545 4377 2579
rect 4343 2477 4377 2511
rect -297 2409 -263 2443
rect 4343 2409 4377 2443
rect -297 2341 -263 2375
rect -297 2273 -263 2307
rect 4343 2341 4377 2375
rect 4343 2273 4377 2307
rect -297 2205 -263 2239
rect -297 2137 -263 2171
rect 4343 2205 4377 2239
rect 4343 2137 4377 2171
rect -187 2023 -153 2057
rect -119 2023 -85 2057
rect -51 2023 -17 2057
rect 17 2023 51 2057
rect 85 2023 119 2057
rect 153 2023 187 2057
rect 221 2023 255 2057
rect 289 2023 323 2057
rect 357 2023 391 2057
rect 425 2023 459 2057
rect 493 2023 527 2057
rect 561 2023 595 2057
rect 629 2023 663 2057
rect 697 2023 731 2057
rect 765 2023 799 2057
rect 833 2023 867 2057
rect 901 2023 935 2057
rect 969 2023 1003 2057
rect 1037 2023 1071 2057
rect 1105 2023 1139 2057
rect 1173 2023 1207 2057
rect 1241 2023 1275 2057
rect 1309 2023 1343 2057
rect 1377 2023 1411 2057
rect 1445 2023 1479 2057
rect 1513 2023 1547 2057
rect 1581 2023 1615 2057
rect 1649 2023 1683 2057
rect 1717 2023 1751 2057
rect 1785 2023 1819 2057
rect 1853 2023 1887 2057
rect 1921 2023 1955 2057
rect 1989 2023 2023 2057
rect 2057 2023 2091 2057
rect 2125 2023 2159 2057
rect 2193 2023 2227 2057
rect 2261 2023 2295 2057
rect 2329 2023 2363 2057
rect 2397 2023 2431 2057
rect 2465 2023 2499 2057
rect 2533 2023 2567 2057
rect 2601 2023 2635 2057
rect 2669 2023 2703 2057
rect 2737 2023 2771 2057
rect 2805 2023 2839 2057
rect 2873 2023 2907 2057
rect 2941 2023 2975 2057
rect 3009 2023 3043 2057
rect 3077 2023 3111 2057
rect 3145 2023 3179 2057
rect 3213 2023 3247 2057
rect 3281 2023 3315 2057
rect 3349 2023 3383 2057
rect 3417 2023 3451 2057
rect 3485 2023 3519 2057
rect 3553 2023 3587 2057
rect 3621 2023 3655 2057
rect 3689 2023 3723 2057
rect 3757 2023 3791 2057
rect 3825 2023 3859 2057
rect 3893 2023 3927 2057
rect 3961 2023 3995 2057
rect 4029 2023 4063 2057
rect 4097 2023 4131 2057
rect 4165 2023 4199 2057
rect 4233 2023 4267 2057
rect 8293 2823 8327 2857
rect 8361 2823 8395 2857
rect 8429 2823 8463 2857
rect 8497 2823 8531 2857
rect 8565 2823 8599 2857
rect 8633 2823 8667 2857
rect 8701 2823 8735 2857
rect 8769 2823 8803 2857
rect 8837 2823 8871 2857
rect 8905 2823 8939 2857
rect 8973 2823 9007 2857
rect 9041 2823 9075 2857
rect 9109 2823 9143 2857
rect 9177 2823 9211 2857
rect 9245 2823 9279 2857
rect 9313 2823 9347 2857
rect 9381 2823 9415 2857
rect 9449 2823 9483 2857
rect 9517 2823 9551 2857
rect 9585 2823 9619 2857
rect 9653 2823 9687 2857
rect 9721 2823 9755 2857
rect 9789 2823 9823 2857
rect 9857 2823 9891 2857
rect 9925 2823 9959 2857
rect 9993 2823 10027 2857
rect 10061 2823 10095 2857
rect 10129 2823 10163 2857
rect 10197 2823 10231 2857
rect 10265 2823 10299 2857
rect 10333 2823 10367 2857
rect 10401 2823 10435 2857
rect 10469 2823 10503 2857
rect 10537 2823 10571 2857
rect 10605 2823 10639 2857
rect 10673 2823 10707 2857
rect 10741 2823 10775 2857
rect 10809 2823 10843 2857
rect 10877 2823 10911 2857
rect 10945 2823 10979 2857
rect 11013 2823 11047 2857
rect 11081 2823 11115 2857
rect 11149 2823 11183 2857
rect 11217 2823 11251 2857
rect 11285 2823 11319 2857
rect 11353 2823 11387 2857
rect 11421 2823 11455 2857
rect 11489 2823 11523 2857
rect 11557 2823 11591 2857
rect 11625 2823 11659 2857
rect 11693 2823 11727 2857
rect 11761 2823 11795 2857
rect 11829 2823 11863 2857
rect 11897 2823 11931 2857
rect 11965 2823 11999 2857
rect 12033 2823 12067 2857
rect 12101 2823 12135 2857
rect 12169 2823 12203 2857
rect 12237 2823 12271 2857
rect 12305 2823 12339 2857
rect 12373 2823 12407 2857
rect 12441 2823 12475 2857
rect 12509 2823 12543 2857
rect 12577 2823 12611 2857
rect 12645 2823 12679 2857
rect 12713 2823 12747 2857
rect 8183 2749 8217 2783
rect 12823 2749 12857 2783
rect 8183 2681 8217 2715
rect 8183 2613 8217 2647
rect 8183 2545 8217 2579
rect 12823 2681 12857 2715
rect 12823 2613 12857 2647
rect 8183 2477 8217 2511
rect 12823 2545 12857 2579
rect 12823 2477 12857 2511
rect 8183 2409 8217 2443
rect 12823 2409 12857 2443
rect 8183 2341 8217 2375
rect 8183 2273 8217 2307
rect 12823 2341 12857 2375
rect 12823 2273 12857 2307
rect 8183 2205 8217 2239
rect 8183 2137 8217 2171
rect 12823 2205 12857 2239
rect 12823 2137 12857 2171
rect 8293 2023 8327 2057
rect 8361 2023 8395 2057
rect 8429 2023 8463 2057
rect 8497 2023 8531 2057
rect 8565 2023 8599 2057
rect 8633 2023 8667 2057
rect 8701 2023 8735 2057
rect 8769 2023 8803 2057
rect 8837 2023 8871 2057
rect 8905 2023 8939 2057
rect 8973 2023 9007 2057
rect 9041 2023 9075 2057
rect 9109 2023 9143 2057
rect 9177 2023 9211 2057
rect 9245 2023 9279 2057
rect 9313 2023 9347 2057
rect 9381 2023 9415 2057
rect 9449 2023 9483 2057
rect 9517 2023 9551 2057
rect 9585 2023 9619 2057
rect 9653 2023 9687 2057
rect 9721 2023 9755 2057
rect 9789 2023 9823 2057
rect 9857 2023 9891 2057
rect 9925 2023 9959 2057
rect 9993 2023 10027 2057
rect 10061 2023 10095 2057
rect 10129 2023 10163 2057
rect 10197 2023 10231 2057
rect 10265 2023 10299 2057
rect 10333 2023 10367 2057
rect 10401 2023 10435 2057
rect 10469 2023 10503 2057
rect 10537 2023 10571 2057
rect 10605 2023 10639 2057
rect 10673 2023 10707 2057
rect 10741 2023 10775 2057
rect 10809 2023 10843 2057
rect 10877 2023 10911 2057
rect 10945 2023 10979 2057
rect 11013 2023 11047 2057
rect 11081 2023 11115 2057
rect 11149 2023 11183 2057
rect 11217 2023 11251 2057
rect 11285 2023 11319 2057
rect 11353 2023 11387 2057
rect 11421 2023 11455 2057
rect 11489 2023 11523 2057
rect 11557 2023 11591 2057
rect 11625 2023 11659 2057
rect 11693 2023 11727 2057
rect 11761 2023 11795 2057
rect 11829 2023 11863 2057
rect 11897 2023 11931 2057
rect 11965 2023 11999 2057
rect 12033 2023 12067 2057
rect 12101 2023 12135 2057
rect 12169 2023 12203 2057
rect 12237 2023 12271 2057
rect 12305 2023 12339 2057
rect 12373 2023 12407 2057
rect 12441 2023 12475 2057
rect 12509 2023 12543 2057
rect 12577 2023 12611 2057
rect 12645 2023 12679 2057
rect 12713 2023 12747 2057
rect -187 1543 -153 1577
rect -119 1543 -85 1577
rect -51 1543 -17 1577
rect 17 1543 51 1577
rect 85 1543 119 1577
rect 153 1543 187 1577
rect 221 1543 255 1577
rect 289 1543 323 1577
rect 357 1543 391 1577
rect 425 1543 459 1577
rect 493 1543 527 1577
rect 561 1543 595 1577
rect 629 1543 663 1577
rect 697 1543 731 1577
rect 765 1543 799 1577
rect 833 1543 867 1577
rect 901 1543 935 1577
rect 969 1543 1003 1577
rect 1037 1543 1071 1577
rect 1105 1543 1139 1577
rect 1173 1543 1207 1577
rect 1241 1543 1275 1577
rect 1309 1543 1343 1577
rect 1377 1543 1411 1577
rect 1445 1543 1479 1577
rect 1513 1543 1547 1577
rect 1581 1543 1615 1577
rect 1649 1543 1683 1577
rect 1717 1543 1751 1577
rect 1785 1543 1819 1577
rect 1853 1543 1887 1577
rect 1921 1543 1955 1577
rect 1989 1543 2023 1577
rect 2057 1543 2091 1577
rect 2125 1543 2159 1577
rect 2193 1543 2227 1577
rect 2261 1543 2295 1577
rect 2329 1543 2363 1577
rect 2397 1543 2431 1577
rect 2465 1543 2499 1577
rect 2533 1543 2567 1577
rect 2601 1543 2635 1577
rect 2669 1543 2703 1577
rect 2737 1543 2771 1577
rect 2805 1543 2839 1577
rect 2873 1543 2907 1577
rect 2941 1543 2975 1577
rect 3009 1543 3043 1577
rect 3077 1543 3111 1577
rect 3145 1543 3179 1577
rect 3213 1543 3247 1577
rect 3281 1543 3315 1577
rect 3349 1543 3383 1577
rect 3417 1543 3451 1577
rect 3485 1543 3519 1577
rect 3553 1543 3587 1577
rect 3621 1543 3655 1577
rect 3689 1543 3723 1577
rect 3757 1543 3791 1577
rect 3825 1543 3859 1577
rect 3893 1543 3927 1577
rect 3961 1543 3995 1577
rect 4029 1543 4063 1577
rect 4097 1543 4131 1577
rect 4165 1543 4199 1577
rect 4233 1543 4267 1577
rect -297 1429 -263 1463
rect -297 1361 -263 1395
rect 4343 1429 4377 1463
rect 4343 1361 4377 1395
rect -297 1293 -263 1327
rect -297 1225 -263 1259
rect 4343 1293 4377 1327
rect 4343 1225 4377 1259
rect -297 1157 -263 1191
rect 4343 1157 4377 1191
rect -297 1089 -263 1123
rect -297 1021 -263 1055
rect 4343 1089 4377 1123
rect -297 953 -263 987
rect -297 885 -263 919
rect 4343 1021 4377 1055
rect 4343 953 4377 987
rect 4343 885 4377 919
rect -297 817 -263 851
rect 4343 817 4377 851
rect -187 743 -153 777
rect -119 743 -85 777
rect -51 743 -17 777
rect 17 743 51 777
rect 85 743 119 777
rect 153 743 187 777
rect 221 743 255 777
rect 289 743 323 777
rect 357 743 391 777
rect 425 743 459 777
rect 493 743 527 777
rect 561 743 595 777
rect 629 743 663 777
rect 697 743 731 777
rect 765 743 799 777
rect 833 743 867 777
rect 901 743 935 777
rect 969 743 1003 777
rect 1037 743 1071 777
rect 1105 743 1139 777
rect 1173 743 1207 777
rect 1241 743 1275 777
rect 1309 743 1343 777
rect 1377 743 1411 777
rect 1445 743 1479 777
rect 1513 743 1547 777
rect 1581 743 1615 777
rect 1649 743 1683 777
rect 1717 743 1751 777
rect 1785 743 1819 777
rect 1853 743 1887 777
rect 1921 743 1955 777
rect 1989 743 2023 777
rect 2057 743 2091 777
rect 2125 743 2159 777
rect 2193 743 2227 777
rect 2261 743 2295 777
rect 2329 743 2363 777
rect 2397 743 2431 777
rect 2465 743 2499 777
rect 2533 743 2567 777
rect 2601 743 2635 777
rect 2669 743 2703 777
rect 2737 743 2771 777
rect 2805 743 2839 777
rect 2873 743 2907 777
rect 2941 743 2975 777
rect 3009 743 3043 777
rect 3077 743 3111 777
rect 3145 743 3179 777
rect 3213 743 3247 777
rect 3281 743 3315 777
rect 3349 743 3383 777
rect 3417 743 3451 777
rect 3485 743 3519 777
rect 3553 743 3587 777
rect 3621 743 3655 777
rect 3689 743 3723 777
rect 3757 743 3791 777
rect 3825 743 3859 777
rect 3893 743 3927 777
rect 3961 743 3995 777
rect 4029 743 4063 777
rect 4097 743 4131 777
rect 4165 743 4199 777
rect 4233 743 4267 777
rect 8293 1543 8327 1577
rect 8361 1543 8395 1577
rect 8429 1543 8463 1577
rect 8497 1543 8531 1577
rect 8565 1543 8599 1577
rect 8633 1543 8667 1577
rect 8701 1543 8735 1577
rect 8769 1543 8803 1577
rect 8837 1543 8871 1577
rect 8905 1543 8939 1577
rect 8973 1543 9007 1577
rect 9041 1543 9075 1577
rect 9109 1543 9143 1577
rect 9177 1543 9211 1577
rect 9245 1543 9279 1577
rect 9313 1543 9347 1577
rect 9381 1543 9415 1577
rect 9449 1543 9483 1577
rect 9517 1543 9551 1577
rect 9585 1543 9619 1577
rect 9653 1543 9687 1577
rect 9721 1543 9755 1577
rect 9789 1543 9823 1577
rect 9857 1543 9891 1577
rect 9925 1543 9959 1577
rect 9993 1543 10027 1577
rect 10061 1543 10095 1577
rect 10129 1543 10163 1577
rect 10197 1543 10231 1577
rect 10265 1543 10299 1577
rect 10333 1543 10367 1577
rect 10401 1543 10435 1577
rect 10469 1543 10503 1577
rect 10537 1543 10571 1577
rect 10605 1543 10639 1577
rect 10673 1543 10707 1577
rect 10741 1543 10775 1577
rect 10809 1543 10843 1577
rect 10877 1543 10911 1577
rect 10945 1543 10979 1577
rect 11013 1543 11047 1577
rect 11081 1543 11115 1577
rect 11149 1543 11183 1577
rect 11217 1543 11251 1577
rect 11285 1543 11319 1577
rect 11353 1543 11387 1577
rect 11421 1543 11455 1577
rect 11489 1543 11523 1577
rect 11557 1543 11591 1577
rect 11625 1543 11659 1577
rect 11693 1543 11727 1577
rect 11761 1543 11795 1577
rect 11829 1543 11863 1577
rect 11897 1543 11931 1577
rect 11965 1543 11999 1577
rect 12033 1543 12067 1577
rect 12101 1543 12135 1577
rect 12169 1543 12203 1577
rect 12237 1543 12271 1577
rect 12305 1543 12339 1577
rect 12373 1543 12407 1577
rect 12441 1543 12475 1577
rect 12509 1543 12543 1577
rect 12577 1543 12611 1577
rect 12645 1543 12679 1577
rect 12713 1543 12747 1577
rect 8183 1429 8217 1463
rect 8183 1361 8217 1395
rect 12823 1429 12857 1463
rect 12823 1361 12857 1395
rect 8183 1293 8217 1327
rect 8183 1225 8217 1259
rect 12823 1293 12857 1327
rect 12823 1225 12857 1259
rect 8183 1157 8217 1191
rect 12823 1157 12857 1191
rect 8183 1089 8217 1123
rect 8183 1021 8217 1055
rect 12823 1089 12857 1123
rect 8183 953 8217 987
rect 8183 885 8217 919
rect 12823 1021 12857 1055
rect 12823 953 12857 987
rect 12823 885 12857 919
rect 8183 817 8217 851
rect 12823 817 12857 851
rect 8293 743 8327 777
rect 8361 743 8395 777
rect 8429 743 8463 777
rect 8497 743 8531 777
rect 8565 743 8599 777
rect 8633 743 8667 777
rect 8701 743 8735 777
rect 8769 743 8803 777
rect 8837 743 8871 777
rect 8905 743 8939 777
rect 8973 743 9007 777
rect 9041 743 9075 777
rect 9109 743 9143 777
rect 9177 743 9211 777
rect 9245 743 9279 777
rect 9313 743 9347 777
rect 9381 743 9415 777
rect 9449 743 9483 777
rect 9517 743 9551 777
rect 9585 743 9619 777
rect 9653 743 9687 777
rect 9721 743 9755 777
rect 9789 743 9823 777
rect 9857 743 9891 777
rect 9925 743 9959 777
rect 9993 743 10027 777
rect 10061 743 10095 777
rect 10129 743 10163 777
rect 10197 743 10231 777
rect 10265 743 10299 777
rect 10333 743 10367 777
rect 10401 743 10435 777
rect 10469 743 10503 777
rect 10537 743 10571 777
rect 10605 743 10639 777
rect 10673 743 10707 777
rect 10741 743 10775 777
rect 10809 743 10843 777
rect 10877 743 10911 777
rect 10945 743 10979 777
rect 11013 743 11047 777
rect 11081 743 11115 777
rect 11149 743 11183 777
rect 11217 743 11251 777
rect 11285 743 11319 777
rect 11353 743 11387 777
rect 11421 743 11455 777
rect 11489 743 11523 777
rect 11557 743 11591 777
rect 11625 743 11659 777
rect 11693 743 11727 777
rect 11761 743 11795 777
rect 11829 743 11863 777
rect 11897 743 11931 777
rect 11965 743 11999 777
rect 12033 743 12067 777
rect 12101 743 12135 777
rect 12169 743 12203 777
rect 12237 743 12271 777
rect 12305 743 12339 777
rect 12373 743 12407 777
rect 12441 743 12475 777
rect 12509 743 12543 777
rect 12577 743 12611 777
rect 12645 743 12679 777
rect 12713 743 12747 777
rect -187 263 -153 297
rect -119 263 -85 297
rect -51 263 -17 297
rect 17 263 51 297
rect 85 263 119 297
rect 153 263 187 297
rect 221 263 255 297
rect 289 263 323 297
rect 357 263 391 297
rect 425 263 459 297
rect 493 263 527 297
rect 561 263 595 297
rect 629 263 663 297
rect 697 263 731 297
rect 765 263 799 297
rect 833 263 867 297
rect 901 263 935 297
rect 969 263 1003 297
rect 1037 263 1071 297
rect 1105 263 1139 297
rect 1173 263 1207 297
rect 1241 263 1275 297
rect 1309 263 1343 297
rect 1377 263 1411 297
rect 1445 263 1479 297
rect 1513 263 1547 297
rect 1581 263 1615 297
rect 1649 263 1683 297
rect 1717 263 1751 297
rect 1785 263 1819 297
rect 1853 263 1887 297
rect 1921 263 1955 297
rect 1989 263 2023 297
rect 2057 263 2091 297
rect 2125 263 2159 297
rect 2193 263 2227 297
rect 2261 263 2295 297
rect 2329 263 2363 297
rect 2397 263 2431 297
rect 2465 263 2499 297
rect 2533 263 2567 297
rect 2601 263 2635 297
rect 2669 263 2703 297
rect 2737 263 2771 297
rect 2805 263 2839 297
rect 2873 263 2907 297
rect 2941 263 2975 297
rect 3009 263 3043 297
rect 3077 263 3111 297
rect 3145 263 3179 297
rect 3213 263 3247 297
rect 3281 263 3315 297
rect 3349 263 3383 297
rect 3417 263 3451 297
rect 3485 263 3519 297
rect 3553 263 3587 297
rect 3621 263 3655 297
rect 3689 263 3723 297
rect 3757 263 3791 297
rect 3825 263 3859 297
rect 3893 263 3927 297
rect 3961 263 3995 297
rect 4029 263 4063 297
rect 4097 263 4131 297
rect 4165 263 4199 297
rect 4233 263 4267 297
rect -297 189 -263 223
rect 4343 189 4377 223
rect -297 121 -263 155
rect -297 53 -263 87
rect -297 -15 -263 19
rect 4343 121 4377 155
rect 4343 53 4377 87
rect -297 -83 -263 -49
rect 4343 -15 4377 19
rect 4343 -83 4377 -49
rect -297 -151 -263 -117
rect 4343 -151 4377 -117
rect -297 -219 -263 -185
rect -297 -287 -263 -253
rect 4343 -219 4377 -185
rect 4343 -287 4377 -253
rect -297 -355 -263 -321
rect -297 -423 -263 -389
rect 4343 -355 4377 -321
rect 4343 -423 4377 -389
rect -187 -537 -153 -503
rect -119 -537 -85 -503
rect -51 -537 -17 -503
rect 17 -537 51 -503
rect 85 -537 119 -503
rect 153 -537 187 -503
rect 221 -537 255 -503
rect 289 -537 323 -503
rect 357 -537 391 -503
rect 425 -537 459 -503
rect 493 -537 527 -503
rect 561 -537 595 -503
rect 629 -537 663 -503
rect 697 -537 731 -503
rect 765 -537 799 -503
rect 833 -537 867 -503
rect 901 -537 935 -503
rect 969 -537 1003 -503
rect 1037 -537 1071 -503
rect 1105 -537 1139 -503
rect 1173 -537 1207 -503
rect 1241 -537 1275 -503
rect 1309 -537 1343 -503
rect 1377 -537 1411 -503
rect 1445 -537 1479 -503
rect 1513 -537 1547 -503
rect 1581 -537 1615 -503
rect 1649 -537 1683 -503
rect 1717 -537 1751 -503
rect 1785 -537 1819 -503
rect 1853 -537 1887 -503
rect 1921 -537 1955 -503
rect 1989 -537 2023 -503
rect 2057 -537 2091 -503
rect 2125 -537 2159 -503
rect 2193 -537 2227 -503
rect 2261 -537 2295 -503
rect 2329 -537 2363 -503
rect 2397 -537 2431 -503
rect 2465 -537 2499 -503
rect 2533 -537 2567 -503
rect 2601 -537 2635 -503
rect 2669 -537 2703 -503
rect 2737 -537 2771 -503
rect 2805 -537 2839 -503
rect 2873 -537 2907 -503
rect 2941 -537 2975 -503
rect 3009 -537 3043 -503
rect 3077 -537 3111 -503
rect 3145 -537 3179 -503
rect 3213 -537 3247 -503
rect 3281 -537 3315 -503
rect 3349 -537 3383 -503
rect 3417 -537 3451 -503
rect 3485 -537 3519 -503
rect 3553 -537 3587 -503
rect 3621 -537 3655 -503
rect 3689 -537 3723 -503
rect 3757 -537 3791 -503
rect 3825 -537 3859 -503
rect 3893 -537 3927 -503
rect 3961 -537 3995 -503
rect 4029 -537 4063 -503
rect 4097 -537 4131 -503
rect 4165 -537 4199 -503
rect 4233 -537 4267 -503
rect 8293 263 8327 297
rect 8361 263 8395 297
rect 8429 263 8463 297
rect 8497 263 8531 297
rect 8565 263 8599 297
rect 8633 263 8667 297
rect 8701 263 8735 297
rect 8769 263 8803 297
rect 8837 263 8871 297
rect 8905 263 8939 297
rect 8973 263 9007 297
rect 9041 263 9075 297
rect 9109 263 9143 297
rect 9177 263 9211 297
rect 9245 263 9279 297
rect 9313 263 9347 297
rect 9381 263 9415 297
rect 9449 263 9483 297
rect 9517 263 9551 297
rect 9585 263 9619 297
rect 9653 263 9687 297
rect 9721 263 9755 297
rect 9789 263 9823 297
rect 9857 263 9891 297
rect 9925 263 9959 297
rect 9993 263 10027 297
rect 10061 263 10095 297
rect 10129 263 10163 297
rect 10197 263 10231 297
rect 10265 263 10299 297
rect 10333 263 10367 297
rect 10401 263 10435 297
rect 10469 263 10503 297
rect 10537 263 10571 297
rect 10605 263 10639 297
rect 10673 263 10707 297
rect 10741 263 10775 297
rect 10809 263 10843 297
rect 10877 263 10911 297
rect 10945 263 10979 297
rect 11013 263 11047 297
rect 11081 263 11115 297
rect 11149 263 11183 297
rect 11217 263 11251 297
rect 11285 263 11319 297
rect 11353 263 11387 297
rect 11421 263 11455 297
rect 11489 263 11523 297
rect 11557 263 11591 297
rect 11625 263 11659 297
rect 11693 263 11727 297
rect 11761 263 11795 297
rect 11829 263 11863 297
rect 11897 263 11931 297
rect 11965 263 11999 297
rect 12033 263 12067 297
rect 12101 263 12135 297
rect 12169 263 12203 297
rect 12237 263 12271 297
rect 12305 263 12339 297
rect 12373 263 12407 297
rect 12441 263 12475 297
rect 12509 263 12543 297
rect 12577 263 12611 297
rect 12645 263 12679 297
rect 12713 263 12747 297
rect 8183 189 8217 223
rect 12823 189 12857 223
rect 8183 121 8217 155
rect 8183 53 8217 87
rect 8183 -15 8217 19
rect 12823 121 12857 155
rect 12823 53 12857 87
rect 8183 -83 8217 -49
rect 12823 -15 12857 19
rect 12823 -83 12857 -49
rect 8183 -151 8217 -117
rect 12823 -151 12857 -117
rect 8183 -219 8217 -185
rect 8183 -287 8217 -253
rect 12823 -219 12857 -185
rect 12823 -287 12857 -253
rect 8183 -355 8217 -321
rect 8183 -423 8217 -389
rect 12823 -355 12857 -321
rect 12823 -423 12857 -389
rect 8293 -537 8327 -503
rect 8361 -537 8395 -503
rect 8429 -537 8463 -503
rect 8497 -537 8531 -503
rect 8565 -537 8599 -503
rect 8633 -537 8667 -503
rect 8701 -537 8735 -503
rect 8769 -537 8803 -503
rect 8837 -537 8871 -503
rect 8905 -537 8939 -503
rect 8973 -537 9007 -503
rect 9041 -537 9075 -503
rect 9109 -537 9143 -503
rect 9177 -537 9211 -503
rect 9245 -537 9279 -503
rect 9313 -537 9347 -503
rect 9381 -537 9415 -503
rect 9449 -537 9483 -503
rect 9517 -537 9551 -503
rect 9585 -537 9619 -503
rect 9653 -537 9687 -503
rect 9721 -537 9755 -503
rect 9789 -537 9823 -503
rect 9857 -537 9891 -503
rect 9925 -537 9959 -503
rect 9993 -537 10027 -503
rect 10061 -537 10095 -503
rect 10129 -537 10163 -503
rect 10197 -537 10231 -503
rect 10265 -537 10299 -503
rect 10333 -537 10367 -503
rect 10401 -537 10435 -503
rect 10469 -537 10503 -503
rect 10537 -537 10571 -503
rect 10605 -537 10639 -503
rect 10673 -537 10707 -503
rect 10741 -537 10775 -503
rect 10809 -537 10843 -503
rect 10877 -537 10911 -503
rect 10945 -537 10979 -503
rect 11013 -537 11047 -503
rect 11081 -537 11115 -503
rect 11149 -537 11183 -503
rect 11217 -537 11251 -503
rect 11285 -537 11319 -503
rect 11353 -537 11387 -503
rect 11421 -537 11455 -503
rect 11489 -537 11523 -503
rect 11557 -537 11591 -503
rect 11625 -537 11659 -503
rect 11693 -537 11727 -503
rect 11761 -537 11795 -503
rect 11829 -537 11863 -503
rect 11897 -537 11931 -503
rect 11965 -537 11999 -503
rect 12033 -537 12067 -503
rect 12101 -537 12135 -503
rect 12169 -537 12203 -503
rect 12237 -537 12271 -503
rect 12305 -537 12339 -503
rect 12373 -537 12407 -503
rect 12441 -537 12475 -503
rect 12509 -537 12543 -503
rect 12577 -537 12611 -503
rect 12645 -537 12679 -503
rect 12713 -537 12747 -503
<< poly >>
rect 40 4000 4040 4040
rect 40 3817 4040 3916
rect 40 3783 85 3817
rect 119 3783 153 3817
rect 187 3783 221 3817
rect 255 3783 289 3817
rect 323 3783 357 3817
rect 391 3783 425 3817
rect 459 3783 493 3817
rect 527 3783 561 3817
rect 595 3783 629 3817
rect 663 3783 697 3817
rect 731 3783 765 3817
rect 799 3783 833 3817
rect 867 3783 901 3817
rect 935 3783 969 3817
rect 1003 3783 1037 3817
rect 1071 3783 1105 3817
rect 1139 3783 1173 3817
rect 1207 3783 1241 3817
rect 1275 3783 1309 3817
rect 1343 3783 1377 3817
rect 1411 3783 1445 3817
rect 1479 3783 1513 3817
rect 1547 3783 1581 3817
rect 1615 3783 1649 3817
rect 1683 3783 1717 3817
rect 1751 3783 1785 3817
rect 1819 3783 1853 3817
rect 1887 3783 1921 3817
rect 1955 3783 1989 3817
rect 2023 3783 2057 3817
rect 2091 3783 2125 3817
rect 2159 3783 2193 3817
rect 2227 3783 2261 3817
rect 2295 3783 2329 3817
rect 2363 3783 2397 3817
rect 2431 3783 2465 3817
rect 2499 3783 2533 3817
rect 2567 3783 2601 3817
rect 2635 3783 2669 3817
rect 2703 3783 2737 3817
rect 2771 3783 2805 3817
rect 2839 3783 2873 3817
rect 2907 3783 2941 3817
rect 2975 3783 3009 3817
rect 3043 3783 3077 3817
rect 3111 3783 3145 3817
rect 3179 3783 3213 3817
rect 3247 3783 3281 3817
rect 3315 3783 3349 3817
rect 3383 3783 3417 3817
rect 3451 3783 3485 3817
rect 3519 3783 3553 3817
rect 3587 3783 3621 3817
rect 3655 3783 3689 3817
rect 3723 3783 3757 3817
rect 3791 3783 3825 3817
rect 3859 3783 3893 3817
rect 3927 3783 3961 3817
rect 3995 3783 4040 3817
rect 40 3760 4040 3783
rect 40 3680 4040 3710
rect 40 3497 4040 3596
rect 40 3463 85 3497
rect 119 3463 153 3497
rect 187 3463 221 3497
rect 255 3463 289 3497
rect 323 3463 357 3497
rect 391 3463 425 3497
rect 459 3463 493 3497
rect 527 3463 561 3497
rect 595 3463 629 3497
rect 663 3463 697 3497
rect 731 3463 765 3497
rect 799 3463 833 3497
rect 867 3463 901 3497
rect 935 3463 969 3497
rect 1003 3463 1037 3497
rect 1071 3463 1105 3497
rect 1139 3463 1173 3497
rect 1207 3463 1241 3497
rect 1275 3463 1309 3497
rect 1343 3463 1377 3497
rect 1411 3463 1445 3497
rect 1479 3463 1513 3497
rect 1547 3463 1581 3497
rect 1615 3463 1649 3497
rect 1683 3463 1717 3497
rect 1751 3463 1785 3497
rect 1819 3463 1853 3497
rect 1887 3463 1921 3497
rect 1955 3463 1989 3497
rect 2023 3463 2057 3497
rect 2091 3463 2125 3497
rect 2159 3463 2193 3497
rect 2227 3463 2261 3497
rect 2295 3463 2329 3497
rect 2363 3463 2397 3497
rect 2431 3463 2465 3497
rect 2499 3463 2533 3497
rect 2567 3463 2601 3497
rect 2635 3463 2669 3497
rect 2703 3463 2737 3497
rect 2771 3463 2805 3497
rect 2839 3463 2873 3497
rect 2907 3463 2941 3497
rect 2975 3463 3009 3497
rect 3043 3463 3077 3497
rect 3111 3463 3145 3497
rect 3179 3463 3213 3497
rect 3247 3463 3281 3497
rect 3315 3463 3349 3497
rect 3383 3463 3417 3497
rect 3451 3463 3485 3497
rect 3519 3463 3553 3497
rect 3587 3463 3621 3497
rect 3655 3463 3689 3497
rect 3723 3463 3757 3497
rect 3791 3463 3825 3497
rect 3859 3463 3893 3497
rect 3927 3463 3961 3497
rect 3995 3463 4040 3497
rect 40 3440 4040 3463
rect 8520 4000 12520 4040
rect 8520 3817 12520 3916
rect 8520 3783 8565 3817
rect 8599 3783 8633 3817
rect 8667 3783 8701 3817
rect 8735 3783 8769 3817
rect 8803 3783 8837 3817
rect 8871 3783 8905 3817
rect 8939 3783 8973 3817
rect 9007 3783 9041 3817
rect 9075 3783 9109 3817
rect 9143 3783 9177 3817
rect 9211 3783 9245 3817
rect 9279 3783 9313 3817
rect 9347 3783 9381 3817
rect 9415 3783 9449 3817
rect 9483 3783 9517 3817
rect 9551 3783 9585 3817
rect 9619 3783 9653 3817
rect 9687 3783 9721 3817
rect 9755 3783 9789 3817
rect 9823 3783 9857 3817
rect 9891 3783 9925 3817
rect 9959 3783 9993 3817
rect 10027 3783 10061 3817
rect 10095 3783 10129 3817
rect 10163 3783 10197 3817
rect 10231 3783 10265 3817
rect 10299 3783 10333 3817
rect 10367 3783 10401 3817
rect 10435 3783 10469 3817
rect 10503 3783 10537 3817
rect 10571 3783 10605 3817
rect 10639 3783 10673 3817
rect 10707 3783 10741 3817
rect 10775 3783 10809 3817
rect 10843 3783 10877 3817
rect 10911 3783 10945 3817
rect 10979 3783 11013 3817
rect 11047 3783 11081 3817
rect 11115 3783 11149 3817
rect 11183 3783 11217 3817
rect 11251 3783 11285 3817
rect 11319 3783 11353 3817
rect 11387 3783 11421 3817
rect 11455 3783 11489 3817
rect 11523 3783 11557 3817
rect 11591 3783 11625 3817
rect 11659 3783 11693 3817
rect 11727 3783 11761 3817
rect 11795 3783 11829 3817
rect 11863 3783 11897 3817
rect 11931 3783 11965 3817
rect 11999 3783 12033 3817
rect 12067 3783 12101 3817
rect 12135 3783 12169 3817
rect 12203 3783 12237 3817
rect 12271 3783 12305 3817
rect 12339 3783 12373 3817
rect 12407 3783 12441 3817
rect 12475 3783 12520 3817
rect 8520 3760 12520 3783
rect 8520 3680 12520 3710
rect 8520 3497 12520 3596
rect 8520 3463 8565 3497
rect 8599 3463 8633 3497
rect 8667 3463 8701 3497
rect 8735 3463 8769 3497
rect 8803 3463 8837 3497
rect 8871 3463 8905 3497
rect 8939 3463 8973 3497
rect 9007 3463 9041 3497
rect 9075 3463 9109 3497
rect 9143 3463 9177 3497
rect 9211 3463 9245 3497
rect 9279 3463 9313 3497
rect 9347 3463 9381 3497
rect 9415 3463 9449 3497
rect 9483 3463 9517 3497
rect 9551 3463 9585 3497
rect 9619 3463 9653 3497
rect 9687 3463 9721 3497
rect 9755 3463 9789 3497
rect 9823 3463 9857 3497
rect 9891 3463 9925 3497
rect 9959 3463 9993 3497
rect 10027 3463 10061 3497
rect 10095 3463 10129 3497
rect 10163 3463 10197 3497
rect 10231 3463 10265 3497
rect 10299 3463 10333 3497
rect 10367 3463 10401 3497
rect 10435 3463 10469 3497
rect 10503 3463 10537 3497
rect 10571 3463 10605 3497
rect 10639 3463 10673 3497
rect 10707 3463 10741 3497
rect 10775 3463 10809 3497
rect 10843 3463 10877 3497
rect 10911 3463 10945 3497
rect 10979 3463 11013 3497
rect 11047 3463 11081 3497
rect 11115 3463 11149 3497
rect 11183 3463 11217 3497
rect 11251 3463 11285 3497
rect 11319 3463 11353 3497
rect 11387 3463 11421 3497
rect 11455 3463 11489 3497
rect 11523 3463 11557 3497
rect 11591 3463 11625 3497
rect 11659 3463 11693 3497
rect 11727 3463 11761 3497
rect 11795 3463 11829 3497
rect 11863 3463 11897 3497
rect 11931 3463 11965 3497
rect 11999 3463 12033 3497
rect 12067 3463 12101 3497
rect 12135 3463 12169 3497
rect 12203 3463 12237 3497
rect 12271 3463 12305 3497
rect 12339 3463 12373 3497
rect 12407 3463 12441 3497
rect 12475 3463 12520 3497
rect 8520 3440 12520 3463
rect 40 2697 4040 2720
rect 40 2663 85 2697
rect 119 2663 153 2697
rect 187 2663 221 2697
rect 255 2663 289 2697
rect 323 2663 357 2697
rect 391 2663 425 2697
rect 459 2663 493 2697
rect 527 2663 561 2697
rect 595 2663 629 2697
rect 663 2663 697 2697
rect 731 2663 765 2697
rect 799 2663 833 2697
rect 867 2663 901 2697
rect 935 2663 969 2697
rect 1003 2663 1037 2697
rect 1071 2663 1105 2697
rect 1139 2663 1173 2697
rect 1207 2663 1241 2697
rect 1275 2663 1309 2697
rect 1343 2663 1377 2697
rect 1411 2663 1445 2697
rect 1479 2663 1513 2697
rect 1547 2663 1581 2697
rect 1615 2663 1649 2697
rect 1683 2663 1717 2697
rect 1751 2663 1785 2697
rect 1819 2663 1853 2697
rect 1887 2663 1921 2697
rect 1955 2663 1989 2697
rect 2023 2663 2057 2697
rect 2091 2663 2125 2697
rect 2159 2663 2193 2697
rect 2227 2663 2261 2697
rect 2295 2663 2329 2697
rect 2363 2663 2397 2697
rect 2431 2663 2465 2697
rect 2499 2663 2533 2697
rect 2567 2663 2601 2697
rect 2635 2663 2669 2697
rect 2703 2663 2737 2697
rect 2771 2663 2805 2697
rect 2839 2663 2873 2697
rect 2907 2663 2941 2697
rect 2975 2663 3009 2697
rect 3043 2663 3077 2697
rect 3111 2663 3145 2697
rect 3179 2663 3213 2697
rect 3247 2663 3281 2697
rect 3315 2663 3349 2697
rect 3383 2663 3417 2697
rect 3451 2663 3485 2697
rect 3519 2663 3553 2697
rect 3587 2663 3621 2697
rect 3655 2663 3689 2697
rect 3723 2663 3757 2697
rect 3791 2663 3825 2697
rect 3859 2663 3893 2697
rect 3927 2663 3961 2697
rect 3995 2663 4040 2697
rect 40 2564 4040 2663
rect 40 2450 4040 2480
rect 40 2377 4040 2400
rect 40 2343 85 2377
rect 119 2343 153 2377
rect 187 2343 221 2377
rect 255 2343 289 2377
rect 323 2343 357 2377
rect 391 2343 425 2377
rect 459 2343 493 2377
rect 527 2343 561 2377
rect 595 2343 629 2377
rect 663 2343 697 2377
rect 731 2343 765 2377
rect 799 2343 833 2377
rect 867 2343 901 2377
rect 935 2343 969 2377
rect 1003 2343 1037 2377
rect 1071 2343 1105 2377
rect 1139 2343 1173 2377
rect 1207 2343 1241 2377
rect 1275 2343 1309 2377
rect 1343 2343 1377 2377
rect 1411 2343 1445 2377
rect 1479 2343 1513 2377
rect 1547 2343 1581 2377
rect 1615 2343 1649 2377
rect 1683 2343 1717 2377
rect 1751 2343 1785 2377
rect 1819 2343 1853 2377
rect 1887 2343 1921 2377
rect 1955 2343 1989 2377
rect 2023 2343 2057 2377
rect 2091 2343 2125 2377
rect 2159 2343 2193 2377
rect 2227 2343 2261 2377
rect 2295 2343 2329 2377
rect 2363 2343 2397 2377
rect 2431 2343 2465 2377
rect 2499 2343 2533 2377
rect 2567 2343 2601 2377
rect 2635 2343 2669 2377
rect 2703 2343 2737 2377
rect 2771 2343 2805 2377
rect 2839 2343 2873 2377
rect 2907 2343 2941 2377
rect 2975 2343 3009 2377
rect 3043 2343 3077 2377
rect 3111 2343 3145 2377
rect 3179 2343 3213 2377
rect 3247 2343 3281 2377
rect 3315 2343 3349 2377
rect 3383 2343 3417 2377
rect 3451 2343 3485 2377
rect 3519 2343 3553 2377
rect 3587 2343 3621 2377
rect 3655 2343 3689 2377
rect 3723 2343 3757 2377
rect 3791 2343 3825 2377
rect 3859 2343 3893 2377
rect 3927 2343 3961 2377
rect 3995 2343 4040 2377
rect 40 2244 4040 2343
rect 40 2120 4040 2160
rect 8520 2697 12520 2720
rect 8520 2663 8565 2697
rect 8599 2663 8633 2697
rect 8667 2663 8701 2697
rect 8735 2663 8769 2697
rect 8803 2663 8837 2697
rect 8871 2663 8905 2697
rect 8939 2663 8973 2697
rect 9007 2663 9041 2697
rect 9075 2663 9109 2697
rect 9143 2663 9177 2697
rect 9211 2663 9245 2697
rect 9279 2663 9313 2697
rect 9347 2663 9381 2697
rect 9415 2663 9449 2697
rect 9483 2663 9517 2697
rect 9551 2663 9585 2697
rect 9619 2663 9653 2697
rect 9687 2663 9721 2697
rect 9755 2663 9789 2697
rect 9823 2663 9857 2697
rect 9891 2663 9925 2697
rect 9959 2663 9993 2697
rect 10027 2663 10061 2697
rect 10095 2663 10129 2697
rect 10163 2663 10197 2697
rect 10231 2663 10265 2697
rect 10299 2663 10333 2697
rect 10367 2663 10401 2697
rect 10435 2663 10469 2697
rect 10503 2663 10537 2697
rect 10571 2663 10605 2697
rect 10639 2663 10673 2697
rect 10707 2663 10741 2697
rect 10775 2663 10809 2697
rect 10843 2663 10877 2697
rect 10911 2663 10945 2697
rect 10979 2663 11013 2697
rect 11047 2663 11081 2697
rect 11115 2663 11149 2697
rect 11183 2663 11217 2697
rect 11251 2663 11285 2697
rect 11319 2663 11353 2697
rect 11387 2663 11421 2697
rect 11455 2663 11489 2697
rect 11523 2663 11557 2697
rect 11591 2663 11625 2697
rect 11659 2663 11693 2697
rect 11727 2663 11761 2697
rect 11795 2663 11829 2697
rect 11863 2663 11897 2697
rect 11931 2663 11965 2697
rect 11999 2663 12033 2697
rect 12067 2663 12101 2697
rect 12135 2663 12169 2697
rect 12203 2663 12237 2697
rect 12271 2663 12305 2697
rect 12339 2663 12373 2697
rect 12407 2663 12441 2697
rect 12475 2663 12520 2697
rect 8520 2564 12520 2663
rect 8520 2450 12520 2480
rect 8520 2377 12520 2400
rect 8520 2343 8565 2377
rect 8599 2343 8633 2377
rect 8667 2343 8701 2377
rect 8735 2343 8769 2377
rect 8803 2343 8837 2377
rect 8871 2343 8905 2377
rect 8939 2343 8973 2377
rect 9007 2343 9041 2377
rect 9075 2343 9109 2377
rect 9143 2343 9177 2377
rect 9211 2343 9245 2377
rect 9279 2343 9313 2377
rect 9347 2343 9381 2377
rect 9415 2343 9449 2377
rect 9483 2343 9517 2377
rect 9551 2343 9585 2377
rect 9619 2343 9653 2377
rect 9687 2343 9721 2377
rect 9755 2343 9789 2377
rect 9823 2343 9857 2377
rect 9891 2343 9925 2377
rect 9959 2343 9993 2377
rect 10027 2343 10061 2377
rect 10095 2343 10129 2377
rect 10163 2343 10197 2377
rect 10231 2343 10265 2377
rect 10299 2343 10333 2377
rect 10367 2343 10401 2377
rect 10435 2343 10469 2377
rect 10503 2343 10537 2377
rect 10571 2343 10605 2377
rect 10639 2343 10673 2377
rect 10707 2343 10741 2377
rect 10775 2343 10809 2377
rect 10843 2343 10877 2377
rect 10911 2343 10945 2377
rect 10979 2343 11013 2377
rect 11047 2343 11081 2377
rect 11115 2343 11149 2377
rect 11183 2343 11217 2377
rect 11251 2343 11285 2377
rect 11319 2343 11353 2377
rect 11387 2343 11421 2377
rect 11455 2343 11489 2377
rect 11523 2343 11557 2377
rect 11591 2343 11625 2377
rect 11659 2343 11693 2377
rect 11727 2343 11761 2377
rect 11795 2343 11829 2377
rect 11863 2343 11897 2377
rect 11931 2343 11965 2377
rect 11999 2343 12033 2377
rect 12067 2343 12101 2377
rect 12135 2343 12169 2377
rect 12203 2343 12237 2377
rect 12271 2343 12305 2377
rect 12339 2343 12373 2377
rect 12407 2343 12441 2377
rect 12475 2343 12520 2377
rect 8520 2244 12520 2343
rect 8520 2120 12520 2160
rect 40 1440 4040 1480
rect 40 1257 4040 1356
rect 40 1223 85 1257
rect 119 1223 153 1257
rect 187 1223 221 1257
rect 255 1223 289 1257
rect 323 1223 357 1257
rect 391 1223 425 1257
rect 459 1223 493 1257
rect 527 1223 561 1257
rect 595 1223 629 1257
rect 663 1223 697 1257
rect 731 1223 765 1257
rect 799 1223 833 1257
rect 867 1223 901 1257
rect 935 1223 969 1257
rect 1003 1223 1037 1257
rect 1071 1223 1105 1257
rect 1139 1223 1173 1257
rect 1207 1223 1241 1257
rect 1275 1223 1309 1257
rect 1343 1223 1377 1257
rect 1411 1223 1445 1257
rect 1479 1223 1513 1257
rect 1547 1223 1581 1257
rect 1615 1223 1649 1257
rect 1683 1223 1717 1257
rect 1751 1223 1785 1257
rect 1819 1223 1853 1257
rect 1887 1223 1921 1257
rect 1955 1223 1989 1257
rect 2023 1223 2057 1257
rect 2091 1223 2125 1257
rect 2159 1223 2193 1257
rect 2227 1223 2261 1257
rect 2295 1223 2329 1257
rect 2363 1223 2397 1257
rect 2431 1223 2465 1257
rect 2499 1223 2533 1257
rect 2567 1223 2601 1257
rect 2635 1223 2669 1257
rect 2703 1223 2737 1257
rect 2771 1223 2805 1257
rect 2839 1223 2873 1257
rect 2907 1223 2941 1257
rect 2975 1223 3009 1257
rect 3043 1223 3077 1257
rect 3111 1223 3145 1257
rect 3179 1223 3213 1257
rect 3247 1223 3281 1257
rect 3315 1223 3349 1257
rect 3383 1223 3417 1257
rect 3451 1223 3485 1257
rect 3519 1223 3553 1257
rect 3587 1223 3621 1257
rect 3655 1223 3689 1257
rect 3723 1223 3757 1257
rect 3791 1223 3825 1257
rect 3859 1223 3893 1257
rect 3927 1223 3961 1257
rect 3995 1223 4040 1257
rect 40 1200 4040 1223
rect 40 1120 4040 1150
rect 40 937 4040 1036
rect 40 903 85 937
rect 119 903 153 937
rect 187 903 221 937
rect 255 903 289 937
rect 323 903 357 937
rect 391 903 425 937
rect 459 903 493 937
rect 527 903 561 937
rect 595 903 629 937
rect 663 903 697 937
rect 731 903 765 937
rect 799 903 833 937
rect 867 903 901 937
rect 935 903 969 937
rect 1003 903 1037 937
rect 1071 903 1105 937
rect 1139 903 1173 937
rect 1207 903 1241 937
rect 1275 903 1309 937
rect 1343 903 1377 937
rect 1411 903 1445 937
rect 1479 903 1513 937
rect 1547 903 1581 937
rect 1615 903 1649 937
rect 1683 903 1717 937
rect 1751 903 1785 937
rect 1819 903 1853 937
rect 1887 903 1921 937
rect 1955 903 1989 937
rect 2023 903 2057 937
rect 2091 903 2125 937
rect 2159 903 2193 937
rect 2227 903 2261 937
rect 2295 903 2329 937
rect 2363 903 2397 937
rect 2431 903 2465 937
rect 2499 903 2533 937
rect 2567 903 2601 937
rect 2635 903 2669 937
rect 2703 903 2737 937
rect 2771 903 2805 937
rect 2839 903 2873 937
rect 2907 903 2941 937
rect 2975 903 3009 937
rect 3043 903 3077 937
rect 3111 903 3145 937
rect 3179 903 3213 937
rect 3247 903 3281 937
rect 3315 903 3349 937
rect 3383 903 3417 937
rect 3451 903 3485 937
rect 3519 903 3553 937
rect 3587 903 3621 937
rect 3655 903 3689 937
rect 3723 903 3757 937
rect 3791 903 3825 937
rect 3859 903 3893 937
rect 3927 903 3961 937
rect 3995 903 4040 937
rect 40 880 4040 903
rect 8520 1440 12520 1480
rect 8520 1257 12520 1356
rect 8520 1223 8565 1257
rect 8599 1223 8633 1257
rect 8667 1223 8701 1257
rect 8735 1223 8769 1257
rect 8803 1223 8837 1257
rect 8871 1223 8905 1257
rect 8939 1223 8973 1257
rect 9007 1223 9041 1257
rect 9075 1223 9109 1257
rect 9143 1223 9177 1257
rect 9211 1223 9245 1257
rect 9279 1223 9313 1257
rect 9347 1223 9381 1257
rect 9415 1223 9449 1257
rect 9483 1223 9517 1257
rect 9551 1223 9585 1257
rect 9619 1223 9653 1257
rect 9687 1223 9721 1257
rect 9755 1223 9789 1257
rect 9823 1223 9857 1257
rect 9891 1223 9925 1257
rect 9959 1223 9993 1257
rect 10027 1223 10061 1257
rect 10095 1223 10129 1257
rect 10163 1223 10197 1257
rect 10231 1223 10265 1257
rect 10299 1223 10333 1257
rect 10367 1223 10401 1257
rect 10435 1223 10469 1257
rect 10503 1223 10537 1257
rect 10571 1223 10605 1257
rect 10639 1223 10673 1257
rect 10707 1223 10741 1257
rect 10775 1223 10809 1257
rect 10843 1223 10877 1257
rect 10911 1223 10945 1257
rect 10979 1223 11013 1257
rect 11047 1223 11081 1257
rect 11115 1223 11149 1257
rect 11183 1223 11217 1257
rect 11251 1223 11285 1257
rect 11319 1223 11353 1257
rect 11387 1223 11421 1257
rect 11455 1223 11489 1257
rect 11523 1223 11557 1257
rect 11591 1223 11625 1257
rect 11659 1223 11693 1257
rect 11727 1223 11761 1257
rect 11795 1223 11829 1257
rect 11863 1223 11897 1257
rect 11931 1223 11965 1257
rect 11999 1223 12033 1257
rect 12067 1223 12101 1257
rect 12135 1223 12169 1257
rect 12203 1223 12237 1257
rect 12271 1223 12305 1257
rect 12339 1223 12373 1257
rect 12407 1223 12441 1257
rect 12475 1223 12520 1257
rect 8520 1200 12520 1223
rect 8520 1120 12520 1150
rect 8520 937 12520 1036
rect 8520 903 8565 937
rect 8599 903 8633 937
rect 8667 903 8701 937
rect 8735 903 8769 937
rect 8803 903 8837 937
rect 8871 903 8905 937
rect 8939 903 8973 937
rect 9007 903 9041 937
rect 9075 903 9109 937
rect 9143 903 9177 937
rect 9211 903 9245 937
rect 9279 903 9313 937
rect 9347 903 9381 937
rect 9415 903 9449 937
rect 9483 903 9517 937
rect 9551 903 9585 937
rect 9619 903 9653 937
rect 9687 903 9721 937
rect 9755 903 9789 937
rect 9823 903 9857 937
rect 9891 903 9925 937
rect 9959 903 9993 937
rect 10027 903 10061 937
rect 10095 903 10129 937
rect 10163 903 10197 937
rect 10231 903 10265 937
rect 10299 903 10333 937
rect 10367 903 10401 937
rect 10435 903 10469 937
rect 10503 903 10537 937
rect 10571 903 10605 937
rect 10639 903 10673 937
rect 10707 903 10741 937
rect 10775 903 10809 937
rect 10843 903 10877 937
rect 10911 903 10945 937
rect 10979 903 11013 937
rect 11047 903 11081 937
rect 11115 903 11149 937
rect 11183 903 11217 937
rect 11251 903 11285 937
rect 11319 903 11353 937
rect 11387 903 11421 937
rect 11455 903 11489 937
rect 11523 903 11557 937
rect 11591 903 11625 937
rect 11659 903 11693 937
rect 11727 903 11761 937
rect 11795 903 11829 937
rect 11863 903 11897 937
rect 11931 903 11965 937
rect 11999 903 12033 937
rect 12067 903 12101 937
rect 12135 903 12169 937
rect 12203 903 12237 937
rect 12271 903 12305 937
rect 12339 903 12373 937
rect 12407 903 12441 937
rect 12475 903 12520 937
rect 8520 880 12520 903
rect 40 137 4040 160
rect 40 103 85 137
rect 119 103 153 137
rect 187 103 221 137
rect 255 103 289 137
rect 323 103 357 137
rect 391 103 425 137
rect 459 103 493 137
rect 527 103 561 137
rect 595 103 629 137
rect 663 103 697 137
rect 731 103 765 137
rect 799 103 833 137
rect 867 103 901 137
rect 935 103 969 137
rect 1003 103 1037 137
rect 1071 103 1105 137
rect 1139 103 1173 137
rect 1207 103 1241 137
rect 1275 103 1309 137
rect 1343 103 1377 137
rect 1411 103 1445 137
rect 1479 103 1513 137
rect 1547 103 1581 137
rect 1615 103 1649 137
rect 1683 103 1717 137
rect 1751 103 1785 137
rect 1819 103 1853 137
rect 1887 103 1921 137
rect 1955 103 1989 137
rect 2023 103 2057 137
rect 2091 103 2125 137
rect 2159 103 2193 137
rect 2227 103 2261 137
rect 2295 103 2329 137
rect 2363 103 2397 137
rect 2431 103 2465 137
rect 2499 103 2533 137
rect 2567 103 2601 137
rect 2635 103 2669 137
rect 2703 103 2737 137
rect 2771 103 2805 137
rect 2839 103 2873 137
rect 2907 103 2941 137
rect 2975 103 3009 137
rect 3043 103 3077 137
rect 3111 103 3145 137
rect 3179 103 3213 137
rect 3247 103 3281 137
rect 3315 103 3349 137
rect 3383 103 3417 137
rect 3451 103 3485 137
rect 3519 103 3553 137
rect 3587 103 3621 137
rect 3655 103 3689 137
rect 3723 103 3757 137
rect 3791 103 3825 137
rect 3859 103 3893 137
rect 3927 103 3961 137
rect 3995 103 4040 137
rect 40 4 4040 103
rect 40 -110 4040 -80
rect 40 -183 4040 -160
rect 40 -217 85 -183
rect 119 -217 153 -183
rect 187 -217 221 -183
rect 255 -217 289 -183
rect 323 -217 357 -183
rect 391 -217 425 -183
rect 459 -217 493 -183
rect 527 -217 561 -183
rect 595 -217 629 -183
rect 663 -217 697 -183
rect 731 -217 765 -183
rect 799 -217 833 -183
rect 867 -217 901 -183
rect 935 -217 969 -183
rect 1003 -217 1037 -183
rect 1071 -217 1105 -183
rect 1139 -217 1173 -183
rect 1207 -217 1241 -183
rect 1275 -217 1309 -183
rect 1343 -217 1377 -183
rect 1411 -217 1445 -183
rect 1479 -217 1513 -183
rect 1547 -217 1581 -183
rect 1615 -217 1649 -183
rect 1683 -217 1717 -183
rect 1751 -217 1785 -183
rect 1819 -217 1853 -183
rect 1887 -217 1921 -183
rect 1955 -217 1989 -183
rect 2023 -217 2057 -183
rect 2091 -217 2125 -183
rect 2159 -217 2193 -183
rect 2227 -217 2261 -183
rect 2295 -217 2329 -183
rect 2363 -217 2397 -183
rect 2431 -217 2465 -183
rect 2499 -217 2533 -183
rect 2567 -217 2601 -183
rect 2635 -217 2669 -183
rect 2703 -217 2737 -183
rect 2771 -217 2805 -183
rect 2839 -217 2873 -183
rect 2907 -217 2941 -183
rect 2975 -217 3009 -183
rect 3043 -217 3077 -183
rect 3111 -217 3145 -183
rect 3179 -217 3213 -183
rect 3247 -217 3281 -183
rect 3315 -217 3349 -183
rect 3383 -217 3417 -183
rect 3451 -217 3485 -183
rect 3519 -217 3553 -183
rect 3587 -217 3621 -183
rect 3655 -217 3689 -183
rect 3723 -217 3757 -183
rect 3791 -217 3825 -183
rect 3859 -217 3893 -183
rect 3927 -217 3961 -183
rect 3995 -217 4040 -183
rect 40 -316 4040 -217
rect 40 -440 4040 -400
rect 8520 137 12520 160
rect 8520 103 8565 137
rect 8599 103 8633 137
rect 8667 103 8701 137
rect 8735 103 8769 137
rect 8803 103 8837 137
rect 8871 103 8905 137
rect 8939 103 8973 137
rect 9007 103 9041 137
rect 9075 103 9109 137
rect 9143 103 9177 137
rect 9211 103 9245 137
rect 9279 103 9313 137
rect 9347 103 9381 137
rect 9415 103 9449 137
rect 9483 103 9517 137
rect 9551 103 9585 137
rect 9619 103 9653 137
rect 9687 103 9721 137
rect 9755 103 9789 137
rect 9823 103 9857 137
rect 9891 103 9925 137
rect 9959 103 9993 137
rect 10027 103 10061 137
rect 10095 103 10129 137
rect 10163 103 10197 137
rect 10231 103 10265 137
rect 10299 103 10333 137
rect 10367 103 10401 137
rect 10435 103 10469 137
rect 10503 103 10537 137
rect 10571 103 10605 137
rect 10639 103 10673 137
rect 10707 103 10741 137
rect 10775 103 10809 137
rect 10843 103 10877 137
rect 10911 103 10945 137
rect 10979 103 11013 137
rect 11047 103 11081 137
rect 11115 103 11149 137
rect 11183 103 11217 137
rect 11251 103 11285 137
rect 11319 103 11353 137
rect 11387 103 11421 137
rect 11455 103 11489 137
rect 11523 103 11557 137
rect 11591 103 11625 137
rect 11659 103 11693 137
rect 11727 103 11761 137
rect 11795 103 11829 137
rect 11863 103 11897 137
rect 11931 103 11965 137
rect 11999 103 12033 137
rect 12067 103 12101 137
rect 12135 103 12169 137
rect 12203 103 12237 137
rect 12271 103 12305 137
rect 12339 103 12373 137
rect 12407 103 12441 137
rect 12475 103 12520 137
rect 8520 4 12520 103
rect 8520 -110 12520 -80
rect 8520 -183 12520 -160
rect 8520 -217 8565 -183
rect 8599 -217 8633 -183
rect 8667 -217 8701 -183
rect 8735 -217 8769 -183
rect 8803 -217 8837 -183
rect 8871 -217 8905 -183
rect 8939 -217 8973 -183
rect 9007 -217 9041 -183
rect 9075 -217 9109 -183
rect 9143 -217 9177 -183
rect 9211 -217 9245 -183
rect 9279 -217 9313 -183
rect 9347 -217 9381 -183
rect 9415 -217 9449 -183
rect 9483 -217 9517 -183
rect 9551 -217 9585 -183
rect 9619 -217 9653 -183
rect 9687 -217 9721 -183
rect 9755 -217 9789 -183
rect 9823 -217 9857 -183
rect 9891 -217 9925 -183
rect 9959 -217 9993 -183
rect 10027 -217 10061 -183
rect 10095 -217 10129 -183
rect 10163 -217 10197 -183
rect 10231 -217 10265 -183
rect 10299 -217 10333 -183
rect 10367 -217 10401 -183
rect 10435 -217 10469 -183
rect 10503 -217 10537 -183
rect 10571 -217 10605 -183
rect 10639 -217 10673 -183
rect 10707 -217 10741 -183
rect 10775 -217 10809 -183
rect 10843 -217 10877 -183
rect 10911 -217 10945 -183
rect 10979 -217 11013 -183
rect 11047 -217 11081 -183
rect 11115 -217 11149 -183
rect 11183 -217 11217 -183
rect 11251 -217 11285 -183
rect 11319 -217 11353 -183
rect 11387 -217 11421 -183
rect 11455 -217 11489 -183
rect 11523 -217 11557 -183
rect 11591 -217 11625 -183
rect 11659 -217 11693 -183
rect 11727 -217 11761 -183
rect 11795 -217 11829 -183
rect 11863 -217 11897 -183
rect 11931 -217 11965 -183
rect 11999 -217 12033 -183
rect 12067 -217 12101 -183
rect 12135 -217 12169 -183
rect 12203 -217 12237 -183
rect 12271 -217 12305 -183
rect 12339 -217 12373 -183
rect 12407 -217 12441 -183
rect 12475 -217 12520 -183
rect 8520 -316 12520 -217
rect 8520 -440 12520 -400
<< polycont >>
rect 85 3783 119 3817
rect 153 3783 187 3817
rect 221 3783 255 3817
rect 289 3783 323 3817
rect 357 3783 391 3817
rect 425 3783 459 3817
rect 493 3783 527 3817
rect 561 3783 595 3817
rect 629 3783 663 3817
rect 697 3783 731 3817
rect 765 3783 799 3817
rect 833 3783 867 3817
rect 901 3783 935 3817
rect 969 3783 1003 3817
rect 1037 3783 1071 3817
rect 1105 3783 1139 3817
rect 1173 3783 1207 3817
rect 1241 3783 1275 3817
rect 1309 3783 1343 3817
rect 1377 3783 1411 3817
rect 1445 3783 1479 3817
rect 1513 3783 1547 3817
rect 1581 3783 1615 3817
rect 1649 3783 1683 3817
rect 1717 3783 1751 3817
rect 1785 3783 1819 3817
rect 1853 3783 1887 3817
rect 1921 3783 1955 3817
rect 1989 3783 2023 3817
rect 2057 3783 2091 3817
rect 2125 3783 2159 3817
rect 2193 3783 2227 3817
rect 2261 3783 2295 3817
rect 2329 3783 2363 3817
rect 2397 3783 2431 3817
rect 2465 3783 2499 3817
rect 2533 3783 2567 3817
rect 2601 3783 2635 3817
rect 2669 3783 2703 3817
rect 2737 3783 2771 3817
rect 2805 3783 2839 3817
rect 2873 3783 2907 3817
rect 2941 3783 2975 3817
rect 3009 3783 3043 3817
rect 3077 3783 3111 3817
rect 3145 3783 3179 3817
rect 3213 3783 3247 3817
rect 3281 3783 3315 3817
rect 3349 3783 3383 3817
rect 3417 3783 3451 3817
rect 3485 3783 3519 3817
rect 3553 3783 3587 3817
rect 3621 3783 3655 3817
rect 3689 3783 3723 3817
rect 3757 3783 3791 3817
rect 3825 3783 3859 3817
rect 3893 3783 3927 3817
rect 3961 3783 3995 3817
rect 85 3463 119 3497
rect 153 3463 187 3497
rect 221 3463 255 3497
rect 289 3463 323 3497
rect 357 3463 391 3497
rect 425 3463 459 3497
rect 493 3463 527 3497
rect 561 3463 595 3497
rect 629 3463 663 3497
rect 697 3463 731 3497
rect 765 3463 799 3497
rect 833 3463 867 3497
rect 901 3463 935 3497
rect 969 3463 1003 3497
rect 1037 3463 1071 3497
rect 1105 3463 1139 3497
rect 1173 3463 1207 3497
rect 1241 3463 1275 3497
rect 1309 3463 1343 3497
rect 1377 3463 1411 3497
rect 1445 3463 1479 3497
rect 1513 3463 1547 3497
rect 1581 3463 1615 3497
rect 1649 3463 1683 3497
rect 1717 3463 1751 3497
rect 1785 3463 1819 3497
rect 1853 3463 1887 3497
rect 1921 3463 1955 3497
rect 1989 3463 2023 3497
rect 2057 3463 2091 3497
rect 2125 3463 2159 3497
rect 2193 3463 2227 3497
rect 2261 3463 2295 3497
rect 2329 3463 2363 3497
rect 2397 3463 2431 3497
rect 2465 3463 2499 3497
rect 2533 3463 2567 3497
rect 2601 3463 2635 3497
rect 2669 3463 2703 3497
rect 2737 3463 2771 3497
rect 2805 3463 2839 3497
rect 2873 3463 2907 3497
rect 2941 3463 2975 3497
rect 3009 3463 3043 3497
rect 3077 3463 3111 3497
rect 3145 3463 3179 3497
rect 3213 3463 3247 3497
rect 3281 3463 3315 3497
rect 3349 3463 3383 3497
rect 3417 3463 3451 3497
rect 3485 3463 3519 3497
rect 3553 3463 3587 3497
rect 3621 3463 3655 3497
rect 3689 3463 3723 3497
rect 3757 3463 3791 3497
rect 3825 3463 3859 3497
rect 3893 3463 3927 3497
rect 3961 3463 3995 3497
rect 8565 3783 8599 3817
rect 8633 3783 8667 3817
rect 8701 3783 8735 3817
rect 8769 3783 8803 3817
rect 8837 3783 8871 3817
rect 8905 3783 8939 3817
rect 8973 3783 9007 3817
rect 9041 3783 9075 3817
rect 9109 3783 9143 3817
rect 9177 3783 9211 3817
rect 9245 3783 9279 3817
rect 9313 3783 9347 3817
rect 9381 3783 9415 3817
rect 9449 3783 9483 3817
rect 9517 3783 9551 3817
rect 9585 3783 9619 3817
rect 9653 3783 9687 3817
rect 9721 3783 9755 3817
rect 9789 3783 9823 3817
rect 9857 3783 9891 3817
rect 9925 3783 9959 3817
rect 9993 3783 10027 3817
rect 10061 3783 10095 3817
rect 10129 3783 10163 3817
rect 10197 3783 10231 3817
rect 10265 3783 10299 3817
rect 10333 3783 10367 3817
rect 10401 3783 10435 3817
rect 10469 3783 10503 3817
rect 10537 3783 10571 3817
rect 10605 3783 10639 3817
rect 10673 3783 10707 3817
rect 10741 3783 10775 3817
rect 10809 3783 10843 3817
rect 10877 3783 10911 3817
rect 10945 3783 10979 3817
rect 11013 3783 11047 3817
rect 11081 3783 11115 3817
rect 11149 3783 11183 3817
rect 11217 3783 11251 3817
rect 11285 3783 11319 3817
rect 11353 3783 11387 3817
rect 11421 3783 11455 3817
rect 11489 3783 11523 3817
rect 11557 3783 11591 3817
rect 11625 3783 11659 3817
rect 11693 3783 11727 3817
rect 11761 3783 11795 3817
rect 11829 3783 11863 3817
rect 11897 3783 11931 3817
rect 11965 3783 11999 3817
rect 12033 3783 12067 3817
rect 12101 3783 12135 3817
rect 12169 3783 12203 3817
rect 12237 3783 12271 3817
rect 12305 3783 12339 3817
rect 12373 3783 12407 3817
rect 12441 3783 12475 3817
rect 8565 3463 8599 3497
rect 8633 3463 8667 3497
rect 8701 3463 8735 3497
rect 8769 3463 8803 3497
rect 8837 3463 8871 3497
rect 8905 3463 8939 3497
rect 8973 3463 9007 3497
rect 9041 3463 9075 3497
rect 9109 3463 9143 3497
rect 9177 3463 9211 3497
rect 9245 3463 9279 3497
rect 9313 3463 9347 3497
rect 9381 3463 9415 3497
rect 9449 3463 9483 3497
rect 9517 3463 9551 3497
rect 9585 3463 9619 3497
rect 9653 3463 9687 3497
rect 9721 3463 9755 3497
rect 9789 3463 9823 3497
rect 9857 3463 9891 3497
rect 9925 3463 9959 3497
rect 9993 3463 10027 3497
rect 10061 3463 10095 3497
rect 10129 3463 10163 3497
rect 10197 3463 10231 3497
rect 10265 3463 10299 3497
rect 10333 3463 10367 3497
rect 10401 3463 10435 3497
rect 10469 3463 10503 3497
rect 10537 3463 10571 3497
rect 10605 3463 10639 3497
rect 10673 3463 10707 3497
rect 10741 3463 10775 3497
rect 10809 3463 10843 3497
rect 10877 3463 10911 3497
rect 10945 3463 10979 3497
rect 11013 3463 11047 3497
rect 11081 3463 11115 3497
rect 11149 3463 11183 3497
rect 11217 3463 11251 3497
rect 11285 3463 11319 3497
rect 11353 3463 11387 3497
rect 11421 3463 11455 3497
rect 11489 3463 11523 3497
rect 11557 3463 11591 3497
rect 11625 3463 11659 3497
rect 11693 3463 11727 3497
rect 11761 3463 11795 3497
rect 11829 3463 11863 3497
rect 11897 3463 11931 3497
rect 11965 3463 11999 3497
rect 12033 3463 12067 3497
rect 12101 3463 12135 3497
rect 12169 3463 12203 3497
rect 12237 3463 12271 3497
rect 12305 3463 12339 3497
rect 12373 3463 12407 3497
rect 12441 3463 12475 3497
rect 85 2663 119 2697
rect 153 2663 187 2697
rect 221 2663 255 2697
rect 289 2663 323 2697
rect 357 2663 391 2697
rect 425 2663 459 2697
rect 493 2663 527 2697
rect 561 2663 595 2697
rect 629 2663 663 2697
rect 697 2663 731 2697
rect 765 2663 799 2697
rect 833 2663 867 2697
rect 901 2663 935 2697
rect 969 2663 1003 2697
rect 1037 2663 1071 2697
rect 1105 2663 1139 2697
rect 1173 2663 1207 2697
rect 1241 2663 1275 2697
rect 1309 2663 1343 2697
rect 1377 2663 1411 2697
rect 1445 2663 1479 2697
rect 1513 2663 1547 2697
rect 1581 2663 1615 2697
rect 1649 2663 1683 2697
rect 1717 2663 1751 2697
rect 1785 2663 1819 2697
rect 1853 2663 1887 2697
rect 1921 2663 1955 2697
rect 1989 2663 2023 2697
rect 2057 2663 2091 2697
rect 2125 2663 2159 2697
rect 2193 2663 2227 2697
rect 2261 2663 2295 2697
rect 2329 2663 2363 2697
rect 2397 2663 2431 2697
rect 2465 2663 2499 2697
rect 2533 2663 2567 2697
rect 2601 2663 2635 2697
rect 2669 2663 2703 2697
rect 2737 2663 2771 2697
rect 2805 2663 2839 2697
rect 2873 2663 2907 2697
rect 2941 2663 2975 2697
rect 3009 2663 3043 2697
rect 3077 2663 3111 2697
rect 3145 2663 3179 2697
rect 3213 2663 3247 2697
rect 3281 2663 3315 2697
rect 3349 2663 3383 2697
rect 3417 2663 3451 2697
rect 3485 2663 3519 2697
rect 3553 2663 3587 2697
rect 3621 2663 3655 2697
rect 3689 2663 3723 2697
rect 3757 2663 3791 2697
rect 3825 2663 3859 2697
rect 3893 2663 3927 2697
rect 3961 2663 3995 2697
rect 85 2343 119 2377
rect 153 2343 187 2377
rect 221 2343 255 2377
rect 289 2343 323 2377
rect 357 2343 391 2377
rect 425 2343 459 2377
rect 493 2343 527 2377
rect 561 2343 595 2377
rect 629 2343 663 2377
rect 697 2343 731 2377
rect 765 2343 799 2377
rect 833 2343 867 2377
rect 901 2343 935 2377
rect 969 2343 1003 2377
rect 1037 2343 1071 2377
rect 1105 2343 1139 2377
rect 1173 2343 1207 2377
rect 1241 2343 1275 2377
rect 1309 2343 1343 2377
rect 1377 2343 1411 2377
rect 1445 2343 1479 2377
rect 1513 2343 1547 2377
rect 1581 2343 1615 2377
rect 1649 2343 1683 2377
rect 1717 2343 1751 2377
rect 1785 2343 1819 2377
rect 1853 2343 1887 2377
rect 1921 2343 1955 2377
rect 1989 2343 2023 2377
rect 2057 2343 2091 2377
rect 2125 2343 2159 2377
rect 2193 2343 2227 2377
rect 2261 2343 2295 2377
rect 2329 2343 2363 2377
rect 2397 2343 2431 2377
rect 2465 2343 2499 2377
rect 2533 2343 2567 2377
rect 2601 2343 2635 2377
rect 2669 2343 2703 2377
rect 2737 2343 2771 2377
rect 2805 2343 2839 2377
rect 2873 2343 2907 2377
rect 2941 2343 2975 2377
rect 3009 2343 3043 2377
rect 3077 2343 3111 2377
rect 3145 2343 3179 2377
rect 3213 2343 3247 2377
rect 3281 2343 3315 2377
rect 3349 2343 3383 2377
rect 3417 2343 3451 2377
rect 3485 2343 3519 2377
rect 3553 2343 3587 2377
rect 3621 2343 3655 2377
rect 3689 2343 3723 2377
rect 3757 2343 3791 2377
rect 3825 2343 3859 2377
rect 3893 2343 3927 2377
rect 3961 2343 3995 2377
rect 8565 2663 8599 2697
rect 8633 2663 8667 2697
rect 8701 2663 8735 2697
rect 8769 2663 8803 2697
rect 8837 2663 8871 2697
rect 8905 2663 8939 2697
rect 8973 2663 9007 2697
rect 9041 2663 9075 2697
rect 9109 2663 9143 2697
rect 9177 2663 9211 2697
rect 9245 2663 9279 2697
rect 9313 2663 9347 2697
rect 9381 2663 9415 2697
rect 9449 2663 9483 2697
rect 9517 2663 9551 2697
rect 9585 2663 9619 2697
rect 9653 2663 9687 2697
rect 9721 2663 9755 2697
rect 9789 2663 9823 2697
rect 9857 2663 9891 2697
rect 9925 2663 9959 2697
rect 9993 2663 10027 2697
rect 10061 2663 10095 2697
rect 10129 2663 10163 2697
rect 10197 2663 10231 2697
rect 10265 2663 10299 2697
rect 10333 2663 10367 2697
rect 10401 2663 10435 2697
rect 10469 2663 10503 2697
rect 10537 2663 10571 2697
rect 10605 2663 10639 2697
rect 10673 2663 10707 2697
rect 10741 2663 10775 2697
rect 10809 2663 10843 2697
rect 10877 2663 10911 2697
rect 10945 2663 10979 2697
rect 11013 2663 11047 2697
rect 11081 2663 11115 2697
rect 11149 2663 11183 2697
rect 11217 2663 11251 2697
rect 11285 2663 11319 2697
rect 11353 2663 11387 2697
rect 11421 2663 11455 2697
rect 11489 2663 11523 2697
rect 11557 2663 11591 2697
rect 11625 2663 11659 2697
rect 11693 2663 11727 2697
rect 11761 2663 11795 2697
rect 11829 2663 11863 2697
rect 11897 2663 11931 2697
rect 11965 2663 11999 2697
rect 12033 2663 12067 2697
rect 12101 2663 12135 2697
rect 12169 2663 12203 2697
rect 12237 2663 12271 2697
rect 12305 2663 12339 2697
rect 12373 2663 12407 2697
rect 12441 2663 12475 2697
rect 8565 2343 8599 2377
rect 8633 2343 8667 2377
rect 8701 2343 8735 2377
rect 8769 2343 8803 2377
rect 8837 2343 8871 2377
rect 8905 2343 8939 2377
rect 8973 2343 9007 2377
rect 9041 2343 9075 2377
rect 9109 2343 9143 2377
rect 9177 2343 9211 2377
rect 9245 2343 9279 2377
rect 9313 2343 9347 2377
rect 9381 2343 9415 2377
rect 9449 2343 9483 2377
rect 9517 2343 9551 2377
rect 9585 2343 9619 2377
rect 9653 2343 9687 2377
rect 9721 2343 9755 2377
rect 9789 2343 9823 2377
rect 9857 2343 9891 2377
rect 9925 2343 9959 2377
rect 9993 2343 10027 2377
rect 10061 2343 10095 2377
rect 10129 2343 10163 2377
rect 10197 2343 10231 2377
rect 10265 2343 10299 2377
rect 10333 2343 10367 2377
rect 10401 2343 10435 2377
rect 10469 2343 10503 2377
rect 10537 2343 10571 2377
rect 10605 2343 10639 2377
rect 10673 2343 10707 2377
rect 10741 2343 10775 2377
rect 10809 2343 10843 2377
rect 10877 2343 10911 2377
rect 10945 2343 10979 2377
rect 11013 2343 11047 2377
rect 11081 2343 11115 2377
rect 11149 2343 11183 2377
rect 11217 2343 11251 2377
rect 11285 2343 11319 2377
rect 11353 2343 11387 2377
rect 11421 2343 11455 2377
rect 11489 2343 11523 2377
rect 11557 2343 11591 2377
rect 11625 2343 11659 2377
rect 11693 2343 11727 2377
rect 11761 2343 11795 2377
rect 11829 2343 11863 2377
rect 11897 2343 11931 2377
rect 11965 2343 11999 2377
rect 12033 2343 12067 2377
rect 12101 2343 12135 2377
rect 12169 2343 12203 2377
rect 12237 2343 12271 2377
rect 12305 2343 12339 2377
rect 12373 2343 12407 2377
rect 12441 2343 12475 2377
rect 85 1223 119 1257
rect 153 1223 187 1257
rect 221 1223 255 1257
rect 289 1223 323 1257
rect 357 1223 391 1257
rect 425 1223 459 1257
rect 493 1223 527 1257
rect 561 1223 595 1257
rect 629 1223 663 1257
rect 697 1223 731 1257
rect 765 1223 799 1257
rect 833 1223 867 1257
rect 901 1223 935 1257
rect 969 1223 1003 1257
rect 1037 1223 1071 1257
rect 1105 1223 1139 1257
rect 1173 1223 1207 1257
rect 1241 1223 1275 1257
rect 1309 1223 1343 1257
rect 1377 1223 1411 1257
rect 1445 1223 1479 1257
rect 1513 1223 1547 1257
rect 1581 1223 1615 1257
rect 1649 1223 1683 1257
rect 1717 1223 1751 1257
rect 1785 1223 1819 1257
rect 1853 1223 1887 1257
rect 1921 1223 1955 1257
rect 1989 1223 2023 1257
rect 2057 1223 2091 1257
rect 2125 1223 2159 1257
rect 2193 1223 2227 1257
rect 2261 1223 2295 1257
rect 2329 1223 2363 1257
rect 2397 1223 2431 1257
rect 2465 1223 2499 1257
rect 2533 1223 2567 1257
rect 2601 1223 2635 1257
rect 2669 1223 2703 1257
rect 2737 1223 2771 1257
rect 2805 1223 2839 1257
rect 2873 1223 2907 1257
rect 2941 1223 2975 1257
rect 3009 1223 3043 1257
rect 3077 1223 3111 1257
rect 3145 1223 3179 1257
rect 3213 1223 3247 1257
rect 3281 1223 3315 1257
rect 3349 1223 3383 1257
rect 3417 1223 3451 1257
rect 3485 1223 3519 1257
rect 3553 1223 3587 1257
rect 3621 1223 3655 1257
rect 3689 1223 3723 1257
rect 3757 1223 3791 1257
rect 3825 1223 3859 1257
rect 3893 1223 3927 1257
rect 3961 1223 3995 1257
rect 85 903 119 937
rect 153 903 187 937
rect 221 903 255 937
rect 289 903 323 937
rect 357 903 391 937
rect 425 903 459 937
rect 493 903 527 937
rect 561 903 595 937
rect 629 903 663 937
rect 697 903 731 937
rect 765 903 799 937
rect 833 903 867 937
rect 901 903 935 937
rect 969 903 1003 937
rect 1037 903 1071 937
rect 1105 903 1139 937
rect 1173 903 1207 937
rect 1241 903 1275 937
rect 1309 903 1343 937
rect 1377 903 1411 937
rect 1445 903 1479 937
rect 1513 903 1547 937
rect 1581 903 1615 937
rect 1649 903 1683 937
rect 1717 903 1751 937
rect 1785 903 1819 937
rect 1853 903 1887 937
rect 1921 903 1955 937
rect 1989 903 2023 937
rect 2057 903 2091 937
rect 2125 903 2159 937
rect 2193 903 2227 937
rect 2261 903 2295 937
rect 2329 903 2363 937
rect 2397 903 2431 937
rect 2465 903 2499 937
rect 2533 903 2567 937
rect 2601 903 2635 937
rect 2669 903 2703 937
rect 2737 903 2771 937
rect 2805 903 2839 937
rect 2873 903 2907 937
rect 2941 903 2975 937
rect 3009 903 3043 937
rect 3077 903 3111 937
rect 3145 903 3179 937
rect 3213 903 3247 937
rect 3281 903 3315 937
rect 3349 903 3383 937
rect 3417 903 3451 937
rect 3485 903 3519 937
rect 3553 903 3587 937
rect 3621 903 3655 937
rect 3689 903 3723 937
rect 3757 903 3791 937
rect 3825 903 3859 937
rect 3893 903 3927 937
rect 3961 903 3995 937
rect 8565 1223 8599 1257
rect 8633 1223 8667 1257
rect 8701 1223 8735 1257
rect 8769 1223 8803 1257
rect 8837 1223 8871 1257
rect 8905 1223 8939 1257
rect 8973 1223 9007 1257
rect 9041 1223 9075 1257
rect 9109 1223 9143 1257
rect 9177 1223 9211 1257
rect 9245 1223 9279 1257
rect 9313 1223 9347 1257
rect 9381 1223 9415 1257
rect 9449 1223 9483 1257
rect 9517 1223 9551 1257
rect 9585 1223 9619 1257
rect 9653 1223 9687 1257
rect 9721 1223 9755 1257
rect 9789 1223 9823 1257
rect 9857 1223 9891 1257
rect 9925 1223 9959 1257
rect 9993 1223 10027 1257
rect 10061 1223 10095 1257
rect 10129 1223 10163 1257
rect 10197 1223 10231 1257
rect 10265 1223 10299 1257
rect 10333 1223 10367 1257
rect 10401 1223 10435 1257
rect 10469 1223 10503 1257
rect 10537 1223 10571 1257
rect 10605 1223 10639 1257
rect 10673 1223 10707 1257
rect 10741 1223 10775 1257
rect 10809 1223 10843 1257
rect 10877 1223 10911 1257
rect 10945 1223 10979 1257
rect 11013 1223 11047 1257
rect 11081 1223 11115 1257
rect 11149 1223 11183 1257
rect 11217 1223 11251 1257
rect 11285 1223 11319 1257
rect 11353 1223 11387 1257
rect 11421 1223 11455 1257
rect 11489 1223 11523 1257
rect 11557 1223 11591 1257
rect 11625 1223 11659 1257
rect 11693 1223 11727 1257
rect 11761 1223 11795 1257
rect 11829 1223 11863 1257
rect 11897 1223 11931 1257
rect 11965 1223 11999 1257
rect 12033 1223 12067 1257
rect 12101 1223 12135 1257
rect 12169 1223 12203 1257
rect 12237 1223 12271 1257
rect 12305 1223 12339 1257
rect 12373 1223 12407 1257
rect 12441 1223 12475 1257
rect 8565 903 8599 937
rect 8633 903 8667 937
rect 8701 903 8735 937
rect 8769 903 8803 937
rect 8837 903 8871 937
rect 8905 903 8939 937
rect 8973 903 9007 937
rect 9041 903 9075 937
rect 9109 903 9143 937
rect 9177 903 9211 937
rect 9245 903 9279 937
rect 9313 903 9347 937
rect 9381 903 9415 937
rect 9449 903 9483 937
rect 9517 903 9551 937
rect 9585 903 9619 937
rect 9653 903 9687 937
rect 9721 903 9755 937
rect 9789 903 9823 937
rect 9857 903 9891 937
rect 9925 903 9959 937
rect 9993 903 10027 937
rect 10061 903 10095 937
rect 10129 903 10163 937
rect 10197 903 10231 937
rect 10265 903 10299 937
rect 10333 903 10367 937
rect 10401 903 10435 937
rect 10469 903 10503 937
rect 10537 903 10571 937
rect 10605 903 10639 937
rect 10673 903 10707 937
rect 10741 903 10775 937
rect 10809 903 10843 937
rect 10877 903 10911 937
rect 10945 903 10979 937
rect 11013 903 11047 937
rect 11081 903 11115 937
rect 11149 903 11183 937
rect 11217 903 11251 937
rect 11285 903 11319 937
rect 11353 903 11387 937
rect 11421 903 11455 937
rect 11489 903 11523 937
rect 11557 903 11591 937
rect 11625 903 11659 937
rect 11693 903 11727 937
rect 11761 903 11795 937
rect 11829 903 11863 937
rect 11897 903 11931 937
rect 11965 903 11999 937
rect 12033 903 12067 937
rect 12101 903 12135 937
rect 12169 903 12203 937
rect 12237 903 12271 937
rect 12305 903 12339 937
rect 12373 903 12407 937
rect 12441 903 12475 937
rect 85 103 119 137
rect 153 103 187 137
rect 221 103 255 137
rect 289 103 323 137
rect 357 103 391 137
rect 425 103 459 137
rect 493 103 527 137
rect 561 103 595 137
rect 629 103 663 137
rect 697 103 731 137
rect 765 103 799 137
rect 833 103 867 137
rect 901 103 935 137
rect 969 103 1003 137
rect 1037 103 1071 137
rect 1105 103 1139 137
rect 1173 103 1207 137
rect 1241 103 1275 137
rect 1309 103 1343 137
rect 1377 103 1411 137
rect 1445 103 1479 137
rect 1513 103 1547 137
rect 1581 103 1615 137
rect 1649 103 1683 137
rect 1717 103 1751 137
rect 1785 103 1819 137
rect 1853 103 1887 137
rect 1921 103 1955 137
rect 1989 103 2023 137
rect 2057 103 2091 137
rect 2125 103 2159 137
rect 2193 103 2227 137
rect 2261 103 2295 137
rect 2329 103 2363 137
rect 2397 103 2431 137
rect 2465 103 2499 137
rect 2533 103 2567 137
rect 2601 103 2635 137
rect 2669 103 2703 137
rect 2737 103 2771 137
rect 2805 103 2839 137
rect 2873 103 2907 137
rect 2941 103 2975 137
rect 3009 103 3043 137
rect 3077 103 3111 137
rect 3145 103 3179 137
rect 3213 103 3247 137
rect 3281 103 3315 137
rect 3349 103 3383 137
rect 3417 103 3451 137
rect 3485 103 3519 137
rect 3553 103 3587 137
rect 3621 103 3655 137
rect 3689 103 3723 137
rect 3757 103 3791 137
rect 3825 103 3859 137
rect 3893 103 3927 137
rect 3961 103 3995 137
rect 85 -217 119 -183
rect 153 -217 187 -183
rect 221 -217 255 -183
rect 289 -217 323 -183
rect 357 -217 391 -183
rect 425 -217 459 -183
rect 493 -217 527 -183
rect 561 -217 595 -183
rect 629 -217 663 -183
rect 697 -217 731 -183
rect 765 -217 799 -183
rect 833 -217 867 -183
rect 901 -217 935 -183
rect 969 -217 1003 -183
rect 1037 -217 1071 -183
rect 1105 -217 1139 -183
rect 1173 -217 1207 -183
rect 1241 -217 1275 -183
rect 1309 -217 1343 -183
rect 1377 -217 1411 -183
rect 1445 -217 1479 -183
rect 1513 -217 1547 -183
rect 1581 -217 1615 -183
rect 1649 -217 1683 -183
rect 1717 -217 1751 -183
rect 1785 -217 1819 -183
rect 1853 -217 1887 -183
rect 1921 -217 1955 -183
rect 1989 -217 2023 -183
rect 2057 -217 2091 -183
rect 2125 -217 2159 -183
rect 2193 -217 2227 -183
rect 2261 -217 2295 -183
rect 2329 -217 2363 -183
rect 2397 -217 2431 -183
rect 2465 -217 2499 -183
rect 2533 -217 2567 -183
rect 2601 -217 2635 -183
rect 2669 -217 2703 -183
rect 2737 -217 2771 -183
rect 2805 -217 2839 -183
rect 2873 -217 2907 -183
rect 2941 -217 2975 -183
rect 3009 -217 3043 -183
rect 3077 -217 3111 -183
rect 3145 -217 3179 -183
rect 3213 -217 3247 -183
rect 3281 -217 3315 -183
rect 3349 -217 3383 -183
rect 3417 -217 3451 -183
rect 3485 -217 3519 -183
rect 3553 -217 3587 -183
rect 3621 -217 3655 -183
rect 3689 -217 3723 -183
rect 3757 -217 3791 -183
rect 3825 -217 3859 -183
rect 3893 -217 3927 -183
rect 3961 -217 3995 -183
rect 8565 103 8599 137
rect 8633 103 8667 137
rect 8701 103 8735 137
rect 8769 103 8803 137
rect 8837 103 8871 137
rect 8905 103 8939 137
rect 8973 103 9007 137
rect 9041 103 9075 137
rect 9109 103 9143 137
rect 9177 103 9211 137
rect 9245 103 9279 137
rect 9313 103 9347 137
rect 9381 103 9415 137
rect 9449 103 9483 137
rect 9517 103 9551 137
rect 9585 103 9619 137
rect 9653 103 9687 137
rect 9721 103 9755 137
rect 9789 103 9823 137
rect 9857 103 9891 137
rect 9925 103 9959 137
rect 9993 103 10027 137
rect 10061 103 10095 137
rect 10129 103 10163 137
rect 10197 103 10231 137
rect 10265 103 10299 137
rect 10333 103 10367 137
rect 10401 103 10435 137
rect 10469 103 10503 137
rect 10537 103 10571 137
rect 10605 103 10639 137
rect 10673 103 10707 137
rect 10741 103 10775 137
rect 10809 103 10843 137
rect 10877 103 10911 137
rect 10945 103 10979 137
rect 11013 103 11047 137
rect 11081 103 11115 137
rect 11149 103 11183 137
rect 11217 103 11251 137
rect 11285 103 11319 137
rect 11353 103 11387 137
rect 11421 103 11455 137
rect 11489 103 11523 137
rect 11557 103 11591 137
rect 11625 103 11659 137
rect 11693 103 11727 137
rect 11761 103 11795 137
rect 11829 103 11863 137
rect 11897 103 11931 137
rect 11965 103 11999 137
rect 12033 103 12067 137
rect 12101 103 12135 137
rect 12169 103 12203 137
rect 12237 103 12271 137
rect 12305 103 12339 137
rect 12373 103 12407 137
rect 12441 103 12475 137
rect 8565 -217 8599 -183
rect 8633 -217 8667 -183
rect 8701 -217 8735 -183
rect 8769 -217 8803 -183
rect 8837 -217 8871 -183
rect 8905 -217 8939 -183
rect 8973 -217 9007 -183
rect 9041 -217 9075 -183
rect 9109 -217 9143 -183
rect 9177 -217 9211 -183
rect 9245 -217 9279 -183
rect 9313 -217 9347 -183
rect 9381 -217 9415 -183
rect 9449 -217 9483 -183
rect 9517 -217 9551 -183
rect 9585 -217 9619 -183
rect 9653 -217 9687 -183
rect 9721 -217 9755 -183
rect 9789 -217 9823 -183
rect 9857 -217 9891 -183
rect 9925 -217 9959 -183
rect 9993 -217 10027 -183
rect 10061 -217 10095 -183
rect 10129 -217 10163 -183
rect 10197 -217 10231 -183
rect 10265 -217 10299 -183
rect 10333 -217 10367 -183
rect 10401 -217 10435 -183
rect 10469 -217 10503 -183
rect 10537 -217 10571 -183
rect 10605 -217 10639 -183
rect 10673 -217 10707 -183
rect 10741 -217 10775 -183
rect 10809 -217 10843 -183
rect 10877 -217 10911 -183
rect 10945 -217 10979 -183
rect 11013 -217 11047 -183
rect 11081 -217 11115 -183
rect 11149 -217 11183 -183
rect 11217 -217 11251 -183
rect 11285 -217 11319 -183
rect 11353 -217 11387 -183
rect 11421 -217 11455 -183
rect 11489 -217 11523 -183
rect 11557 -217 11591 -183
rect 11625 -217 11659 -183
rect 11693 -217 11727 -183
rect 11761 -217 11795 -183
rect 11829 -217 11863 -183
rect 11897 -217 11931 -183
rect 11965 -217 11999 -183
rect 12033 -217 12067 -183
rect 12101 -217 12135 -183
rect 12169 -217 12203 -183
rect 12237 -217 12271 -183
rect 12305 -217 12339 -183
rect 12373 -217 12407 -183
rect 12441 -217 12475 -183
<< locali >>
rect -480 4297 13040 4320
rect -480 4263 -357 4297
rect -323 4263 -289 4297
rect -255 4263 -221 4297
rect -187 4263 -153 4297
rect -119 4263 -85 4297
rect -51 4263 -17 4297
rect 17 4263 51 4297
rect 85 4263 119 4297
rect 153 4263 187 4297
rect 221 4263 255 4297
rect 289 4263 323 4297
rect 357 4263 391 4297
rect 425 4263 459 4297
rect 493 4263 527 4297
rect 561 4263 595 4297
rect 629 4263 663 4297
rect 697 4263 731 4297
rect 765 4263 799 4297
rect 833 4263 867 4297
rect 901 4263 935 4297
rect 969 4263 1003 4297
rect 1037 4263 1071 4297
rect 1105 4263 1139 4297
rect 1173 4263 1207 4297
rect 1241 4263 1275 4297
rect 1309 4263 1343 4297
rect 1377 4263 1411 4297
rect 1445 4263 1479 4297
rect 1513 4263 1547 4297
rect 1581 4263 1615 4297
rect 1649 4263 1683 4297
rect 1717 4263 1751 4297
rect 1785 4263 1819 4297
rect 1853 4263 1887 4297
rect 1921 4263 1955 4297
rect 1989 4263 2023 4297
rect 2057 4263 2091 4297
rect 2125 4263 2159 4297
rect 2193 4263 2227 4297
rect 2261 4263 2295 4297
rect 2329 4263 2363 4297
rect 2397 4263 2431 4297
rect 2465 4263 2499 4297
rect 2533 4263 2567 4297
rect 2601 4263 2635 4297
rect 2669 4263 2703 4297
rect 2737 4263 2771 4297
rect 2805 4263 2839 4297
rect 2873 4263 2907 4297
rect 2941 4263 2975 4297
rect 3009 4263 3043 4297
rect 3077 4263 3111 4297
rect 3145 4263 3179 4297
rect 3213 4263 3247 4297
rect 3281 4263 3315 4297
rect 3349 4263 3383 4297
rect 3417 4263 3451 4297
rect 3485 4263 3519 4297
rect 3553 4263 3587 4297
rect 3621 4263 3655 4297
rect 3689 4263 3723 4297
rect 3757 4263 3791 4297
rect 3825 4263 3859 4297
rect 3893 4263 3927 4297
rect 3961 4263 3995 4297
rect 4029 4263 4063 4297
rect 4097 4263 4131 4297
rect 4165 4263 4199 4297
rect 4233 4263 4267 4297
rect 4301 4263 4335 4297
rect 4369 4263 4403 4297
rect 4437 4263 8123 4297
rect 8157 4263 8191 4297
rect 8225 4263 8259 4297
rect 8293 4263 8327 4297
rect 8361 4263 8395 4297
rect 8429 4263 8463 4297
rect 8497 4263 8531 4297
rect 8565 4263 8599 4297
rect 8633 4263 8667 4297
rect 8701 4263 8735 4297
rect 8769 4263 8803 4297
rect 8837 4263 8871 4297
rect 8905 4263 8939 4297
rect 8973 4263 9007 4297
rect 9041 4263 9075 4297
rect 9109 4263 9143 4297
rect 9177 4263 9211 4297
rect 9245 4263 9279 4297
rect 9313 4263 9347 4297
rect 9381 4263 9415 4297
rect 9449 4263 9483 4297
rect 9517 4263 9551 4297
rect 9585 4263 9619 4297
rect 9653 4263 9687 4297
rect 9721 4263 9755 4297
rect 9789 4263 9823 4297
rect 9857 4263 9891 4297
rect 9925 4263 9959 4297
rect 9993 4263 10027 4297
rect 10061 4263 10095 4297
rect 10129 4263 10163 4297
rect 10197 4263 10231 4297
rect 10265 4263 10299 4297
rect 10333 4263 10367 4297
rect 10401 4263 10435 4297
rect 10469 4263 10503 4297
rect 10537 4263 10571 4297
rect 10605 4263 10639 4297
rect 10673 4263 10707 4297
rect 10741 4263 10775 4297
rect 10809 4263 10843 4297
rect 10877 4263 10911 4297
rect 10945 4263 10979 4297
rect 11013 4263 11047 4297
rect 11081 4263 11115 4297
rect 11149 4263 11183 4297
rect 11217 4263 11251 4297
rect 11285 4263 11319 4297
rect 11353 4263 11387 4297
rect 11421 4263 11455 4297
rect 11489 4263 11523 4297
rect 11557 4263 11591 4297
rect 11625 4263 11659 4297
rect 11693 4263 11727 4297
rect 11761 4263 11795 4297
rect 11829 4263 11863 4297
rect 11897 4263 11931 4297
rect 11965 4263 11999 4297
rect 12033 4263 12067 4297
rect 12101 4263 12135 4297
rect 12169 4263 12203 4297
rect 12237 4263 12271 4297
rect 12305 4263 12339 4297
rect 12373 4263 12407 4297
rect 12441 4263 12475 4297
rect 12509 4263 12543 4297
rect 12577 4263 12611 4297
rect 12645 4263 12679 4297
rect 12713 4263 12747 4297
rect 12781 4263 12815 4297
rect 12849 4263 12883 4297
rect 12917 4263 13040 4297
rect -480 4240 13040 4263
rect -480 4199 -400 4240
rect -480 4165 -457 4199
rect -423 4165 -400 4199
rect -480 4131 -400 4165
rect 4480 4199 4560 4240
rect 4480 4165 4503 4199
rect 4537 4165 4560 4199
rect -480 4097 -457 4131
rect -423 4097 -400 4131
rect -480 4063 -400 4097
rect -480 4029 -457 4063
rect -423 4029 -400 4063
rect -480 3995 -400 4029
rect -480 3961 -457 3995
rect -423 3961 -400 3995
rect -480 3927 -400 3961
rect -480 3893 -457 3927
rect -423 3893 -400 3927
rect -480 3859 -400 3893
rect -480 3825 -457 3859
rect -423 3825 -400 3859
rect -480 3791 -400 3825
rect -480 3757 -457 3791
rect -423 3757 -400 3791
rect -480 3723 -400 3757
rect -480 3689 -457 3723
rect -423 3689 -400 3723
rect -480 3655 -400 3689
rect -480 3621 -457 3655
rect -423 3621 -400 3655
rect -480 3587 -400 3621
rect -480 3553 -457 3587
rect -423 3553 -400 3587
rect -480 3519 -400 3553
rect -480 3485 -457 3519
rect -423 3485 -400 3519
rect -480 3451 -400 3485
rect -480 3417 -457 3451
rect -423 3417 -400 3451
rect -480 3383 -400 3417
rect -480 3349 -457 3383
rect -423 3349 -400 3383
rect -480 3315 -400 3349
rect -480 3281 -457 3315
rect -423 3281 -400 3315
rect -480 3200 -400 3281
rect -320 4137 4400 4160
rect -320 4103 -297 4137
rect -263 4103 -187 4137
rect -153 4103 -119 4137
rect -85 4103 -51 4137
rect -17 4103 17 4137
rect 51 4103 85 4137
rect 119 4103 153 4137
rect 187 4103 221 4137
rect 255 4103 289 4137
rect 323 4103 357 4137
rect 391 4103 425 4137
rect 459 4103 493 4137
rect 527 4103 561 4137
rect 595 4103 629 4137
rect 663 4103 697 4137
rect 731 4103 765 4137
rect 799 4103 833 4137
rect 867 4103 901 4137
rect 935 4103 969 4137
rect 1003 4103 1037 4137
rect 1071 4103 1105 4137
rect 1139 4103 1173 4137
rect 1207 4103 1241 4137
rect 1275 4103 1309 4137
rect 1343 4103 1377 4137
rect 1411 4103 1445 4137
rect 1479 4103 1513 4137
rect 1547 4103 1581 4137
rect 1615 4103 1649 4137
rect 1683 4103 1717 4137
rect 1751 4103 1785 4137
rect 1819 4103 1853 4137
rect 1887 4103 1921 4137
rect 1955 4103 1989 4137
rect 2023 4103 2057 4137
rect 2091 4103 2125 4137
rect 2159 4103 2193 4137
rect 2227 4103 2261 4137
rect 2295 4103 2329 4137
rect 2363 4103 2397 4137
rect 2431 4103 2465 4137
rect 2499 4103 2533 4137
rect 2567 4103 2601 4137
rect 2635 4103 2669 4137
rect 2703 4103 2737 4137
rect 2771 4103 2805 4137
rect 2839 4103 2873 4137
rect 2907 4103 2941 4137
rect 2975 4103 3009 4137
rect 3043 4103 3077 4137
rect 3111 4103 3145 4137
rect 3179 4103 3213 4137
rect 3247 4103 3281 4137
rect 3315 4103 3349 4137
rect 3383 4103 3417 4137
rect 3451 4103 3485 4137
rect 3519 4103 3553 4137
rect 3587 4103 3621 4137
rect 3655 4103 3689 4137
rect 3723 4103 3757 4137
rect 3791 4103 3825 4137
rect 3859 4103 3893 4137
rect 3927 4103 3961 4137
rect 3995 4103 4029 4137
rect 4063 4103 4097 4137
rect 4131 4103 4165 4137
rect 4199 4103 4233 4137
rect 4267 4103 4400 4137
rect -320 4080 4400 4103
rect -320 4023 -240 4080
rect -320 3989 -297 4023
rect -263 3989 -240 4023
rect 4320 4023 4400 4080
rect -320 3955 -240 3989
rect -320 3921 -297 3955
rect -263 3921 -240 3955
rect -320 3887 -240 3921
rect -160 3977 -80 4000
rect -160 3943 -137 3977
rect -103 3943 -80 3977
rect -160 3916 -80 3943
rect 4160 3977 4240 4000
rect 4160 3943 4183 3977
rect 4217 3943 4240 3977
rect 4160 3916 4240 3943
rect 4320 3989 4343 4023
rect 4377 3989 4400 4023
rect 4320 3955 4400 3989
rect 4320 3921 4343 3955
rect 4377 3921 4400 3955
rect -320 3853 -297 3887
rect -263 3853 -240 3887
rect -320 3819 -240 3853
rect 4320 3887 4400 3921
rect 4320 3853 4343 3887
rect 4377 3853 4400 3887
rect -320 3785 -297 3819
rect -263 3785 -240 3819
rect -320 3751 -240 3785
rect 40 3817 4040 3840
rect 40 3783 79 3817
rect 119 3783 151 3817
rect 187 3783 221 3817
rect 257 3783 289 3817
rect 329 3783 357 3817
rect 401 3783 425 3817
rect 473 3783 493 3817
rect 545 3783 561 3817
rect 617 3783 629 3817
rect 689 3783 697 3817
rect 761 3783 765 3817
rect 867 3783 871 3817
rect 935 3783 943 3817
rect 1003 3783 1015 3817
rect 1071 3783 1087 3817
rect 1139 3783 1159 3817
rect 1207 3783 1231 3817
rect 1275 3783 1303 3817
rect 1343 3783 1375 3817
rect 1411 3783 1445 3817
rect 1481 3783 1513 3817
rect 1553 3783 1581 3817
rect 1625 3783 1649 3817
rect 1697 3783 1717 3817
rect 1769 3783 1785 3817
rect 1841 3783 1853 3817
rect 1913 3783 1921 3817
rect 1985 3783 1989 3817
rect 2091 3783 2095 3817
rect 2159 3783 2167 3817
rect 2227 3783 2239 3817
rect 2295 3783 2311 3817
rect 2363 3783 2383 3817
rect 2431 3783 2455 3817
rect 2499 3783 2527 3817
rect 2567 3783 2599 3817
rect 2635 3783 2669 3817
rect 2705 3783 2737 3817
rect 2777 3783 2805 3817
rect 2849 3783 2873 3817
rect 2921 3783 2941 3817
rect 2993 3783 3009 3817
rect 3065 3783 3077 3817
rect 3137 3783 3145 3817
rect 3209 3783 3213 3817
rect 3315 3783 3319 3817
rect 3383 3783 3391 3817
rect 3451 3783 3463 3817
rect 3519 3783 3535 3817
rect 3587 3783 3607 3817
rect 3655 3783 3679 3817
rect 3723 3783 3751 3817
rect 3791 3783 3823 3817
rect 3859 3783 3893 3817
rect 3929 3783 3961 3817
rect 4001 3783 4040 3817
rect 40 3760 4040 3783
rect 4320 3819 4400 3853
rect 4320 3785 4343 3819
rect 4377 3785 4400 3819
rect -320 3717 -297 3751
rect -263 3717 -240 3751
rect -320 3683 -240 3717
rect -320 3649 -297 3683
rect -263 3649 -240 3683
rect 4320 3751 4400 3785
rect 4320 3717 4343 3751
rect 4377 3717 4400 3751
rect 4320 3683 4400 3717
rect -320 3615 -240 3649
rect -320 3581 -297 3615
rect -263 3581 -240 3615
rect -160 3657 -80 3680
rect -160 3623 -137 3657
rect -103 3623 -80 3657
rect -160 3596 -80 3623
rect 4160 3657 4240 3680
rect 4160 3623 4183 3657
rect 4217 3623 4240 3657
rect 4160 3596 4240 3623
rect 4320 3649 4343 3683
rect 4377 3649 4400 3683
rect 4320 3615 4400 3649
rect -320 3547 -240 3581
rect -320 3513 -297 3547
rect -263 3513 -240 3547
rect 4320 3581 4343 3615
rect 4377 3581 4400 3615
rect 4320 3547 4400 3581
rect -320 3479 -240 3513
rect -320 3445 -297 3479
rect -263 3445 -240 3479
rect -320 3411 -240 3445
rect 40 3497 4040 3520
rect 40 3463 79 3497
rect 119 3463 151 3497
rect 187 3463 221 3497
rect 257 3463 289 3497
rect 329 3463 357 3497
rect 401 3463 425 3497
rect 473 3463 493 3497
rect 545 3463 561 3497
rect 617 3463 629 3497
rect 689 3463 697 3497
rect 761 3463 765 3497
rect 867 3463 871 3497
rect 935 3463 943 3497
rect 1003 3463 1015 3497
rect 1071 3463 1087 3497
rect 1139 3463 1159 3497
rect 1207 3463 1231 3497
rect 1275 3463 1303 3497
rect 1343 3463 1375 3497
rect 1411 3463 1445 3497
rect 1481 3463 1513 3497
rect 1553 3463 1581 3497
rect 1625 3463 1649 3497
rect 1697 3463 1717 3497
rect 1769 3463 1785 3497
rect 1841 3463 1853 3497
rect 1913 3463 1921 3497
rect 1985 3463 1989 3497
rect 2091 3463 2095 3497
rect 2159 3463 2167 3497
rect 2227 3463 2239 3497
rect 2295 3463 2311 3497
rect 2363 3463 2383 3497
rect 2431 3463 2455 3497
rect 2499 3463 2527 3497
rect 2567 3463 2599 3497
rect 2635 3463 2669 3497
rect 2705 3463 2737 3497
rect 2777 3463 2805 3497
rect 2849 3463 2873 3497
rect 2921 3463 2941 3497
rect 2993 3463 3009 3497
rect 3065 3463 3077 3497
rect 3137 3463 3145 3497
rect 3209 3463 3213 3497
rect 3315 3463 3319 3497
rect 3383 3463 3391 3497
rect 3451 3463 3463 3497
rect 3519 3463 3535 3497
rect 3587 3463 3607 3497
rect 3655 3463 3679 3497
rect 3723 3463 3751 3497
rect 3791 3463 3823 3497
rect 3859 3463 3893 3497
rect 3929 3463 3961 3497
rect 4001 3463 4040 3497
rect 40 3440 4040 3463
rect 4320 3513 4343 3547
rect 4377 3513 4400 3547
rect 4320 3479 4400 3513
rect 4320 3445 4343 3479
rect 4377 3445 4400 3479
rect -320 3377 -297 3411
rect -263 3377 -240 3411
rect -320 3360 -240 3377
rect 4320 3411 4400 3445
rect 4320 3377 4343 3411
rect 4377 3377 4400 3411
rect 4320 3360 4400 3377
rect -320 3337 4400 3360
rect -320 3303 -187 3337
rect -153 3303 -119 3337
rect -85 3303 -51 3337
rect -17 3303 17 3337
rect 51 3303 85 3337
rect 119 3303 153 3337
rect 187 3303 221 3337
rect 255 3303 289 3337
rect 323 3303 357 3337
rect 391 3303 425 3337
rect 459 3303 493 3337
rect 527 3303 561 3337
rect 595 3303 629 3337
rect 663 3303 697 3337
rect 731 3303 765 3337
rect 799 3303 833 3337
rect 867 3303 901 3337
rect 935 3303 969 3337
rect 1003 3303 1037 3337
rect 1071 3303 1105 3337
rect 1139 3303 1173 3337
rect 1207 3303 1241 3337
rect 1275 3303 1309 3337
rect 1343 3303 1377 3337
rect 1411 3303 1445 3337
rect 1479 3303 1513 3337
rect 1547 3303 1581 3337
rect 1615 3303 1649 3337
rect 1683 3303 1717 3337
rect 1751 3303 1785 3337
rect 1819 3303 1853 3337
rect 1887 3303 1921 3337
rect 1955 3303 1989 3337
rect 2023 3303 2057 3337
rect 2091 3303 2125 3337
rect 2159 3303 2193 3337
rect 2227 3303 2261 3337
rect 2295 3303 2329 3337
rect 2363 3303 2397 3337
rect 2431 3303 2465 3337
rect 2499 3303 2533 3337
rect 2567 3303 2601 3337
rect 2635 3303 2669 3337
rect 2703 3303 2737 3337
rect 2771 3303 2805 3337
rect 2839 3303 2873 3337
rect 2907 3303 2941 3337
rect 2975 3303 3009 3337
rect 3043 3303 3077 3337
rect 3111 3303 3145 3337
rect 3179 3303 3213 3337
rect 3247 3303 3281 3337
rect 3315 3303 3349 3337
rect 3383 3303 3417 3337
rect 3451 3303 3485 3337
rect 3519 3303 3553 3337
rect 3587 3303 3621 3337
rect 3655 3303 3689 3337
rect 3723 3303 3757 3337
rect 3791 3303 3825 3337
rect 3859 3303 3893 3337
rect 3927 3303 3961 3337
rect 3995 3303 4029 3337
rect 4063 3303 4097 3337
rect 4131 3303 4165 3337
rect 4199 3303 4233 3337
rect 4267 3303 4400 3337
rect -320 3280 4400 3303
rect 4480 4131 4560 4165
rect 4480 4097 4503 4131
rect 4537 4097 4560 4131
rect 4480 4063 4560 4097
rect 4480 4029 4503 4063
rect 4537 4029 4560 4063
rect 4480 3995 4560 4029
rect 4480 3961 4503 3995
rect 4537 3961 4560 3995
rect 4480 3927 4560 3961
rect 4480 3893 4503 3927
rect 4537 3893 4560 3927
rect 4480 3859 4560 3893
rect 4480 3825 4503 3859
rect 4537 3825 4560 3859
rect 4480 3791 4560 3825
rect 4480 3757 4503 3791
rect 4537 3757 4560 3791
rect 4480 3723 4560 3757
rect 4480 3689 4503 3723
rect 4537 3689 4560 3723
rect 4480 3655 4560 3689
rect 4480 3621 4503 3655
rect 4537 3621 4560 3655
rect 4480 3587 4560 3621
rect 4480 3553 4503 3587
rect 4537 3553 4560 3587
rect 4480 3519 4560 3553
rect 4480 3485 4503 3519
rect 4537 3485 4560 3519
rect 4480 3451 4560 3485
rect 4480 3417 4503 3451
rect 4537 3417 4560 3451
rect 4480 3383 4560 3417
rect 4480 3349 4503 3383
rect 4537 3349 4560 3383
rect 4480 3315 4560 3349
rect 4480 3281 4503 3315
rect 4537 3281 4560 3315
rect 4480 3200 4560 3281
rect -480 3177 4560 3200
rect -480 3143 -357 3177
rect -323 3143 -289 3177
rect -255 3143 -221 3177
rect -187 3143 -153 3177
rect -119 3143 -85 3177
rect -51 3143 -17 3177
rect 17 3143 51 3177
rect 85 3143 119 3177
rect 153 3143 187 3177
rect 221 3143 255 3177
rect 289 3143 323 3177
rect 357 3143 391 3177
rect 425 3143 459 3177
rect 493 3143 527 3177
rect 561 3143 595 3177
rect 629 3143 663 3177
rect 697 3143 731 3177
rect 765 3143 799 3177
rect 833 3143 867 3177
rect 901 3143 935 3177
rect 969 3143 1003 3177
rect 1037 3143 1071 3177
rect 1105 3143 1139 3177
rect 1173 3143 1207 3177
rect 1241 3143 1275 3177
rect 1309 3143 1343 3177
rect 1377 3143 1411 3177
rect 1445 3143 1479 3177
rect 1513 3143 1547 3177
rect 1581 3143 1615 3177
rect 1649 3143 1683 3177
rect 1717 3143 1751 3177
rect 1785 3143 1819 3177
rect 1853 3143 1887 3177
rect 1921 3143 1955 3177
rect 1989 3143 2023 3177
rect 2057 3143 2091 3177
rect 2125 3143 2159 3177
rect 2193 3143 2227 3177
rect 2261 3143 2295 3177
rect 2329 3143 2363 3177
rect 2397 3143 2431 3177
rect 2465 3143 2499 3177
rect 2533 3143 2567 3177
rect 2601 3143 2635 3177
rect 2669 3143 2703 3177
rect 2737 3143 2771 3177
rect 2805 3143 2839 3177
rect 2873 3143 2907 3177
rect 2941 3143 2975 3177
rect 3009 3143 3043 3177
rect 3077 3143 3111 3177
rect 3145 3143 3179 3177
rect 3213 3143 3247 3177
rect 3281 3143 3315 3177
rect 3349 3143 3383 3177
rect 3417 3143 3451 3177
rect 3485 3143 3519 3177
rect 3553 3143 3587 3177
rect 3621 3143 3655 3177
rect 3689 3143 3723 3177
rect 3757 3143 3791 3177
rect 3825 3143 3859 3177
rect 3893 3143 3927 3177
rect 3961 3143 3995 3177
rect 4029 3143 4063 3177
rect 4097 3143 4131 3177
rect 4165 3143 4199 3177
rect 4233 3143 4267 3177
rect 4301 3143 4335 3177
rect 4369 3143 4403 3177
rect 4437 3143 4560 3177
rect -480 3120 4560 3143
rect -480 3040 -400 3120
rect 4480 3040 4560 3120
rect -480 3017 4560 3040
rect -480 2983 -357 3017
rect -323 2983 -289 3017
rect -255 2983 -221 3017
rect -187 2983 -153 3017
rect -119 2983 -85 3017
rect -51 2983 -17 3017
rect 17 2983 51 3017
rect 85 2983 119 3017
rect 153 2983 187 3017
rect 221 2983 255 3017
rect 289 2983 323 3017
rect 357 2983 391 3017
rect 425 2983 459 3017
rect 493 2983 527 3017
rect 561 2983 595 3017
rect 629 2983 663 3017
rect 697 2983 731 3017
rect 765 2983 799 3017
rect 833 2983 867 3017
rect 901 2983 935 3017
rect 969 2983 1003 3017
rect 1037 2983 1071 3017
rect 1105 2983 1139 3017
rect 1173 2983 1207 3017
rect 1241 2983 1275 3017
rect 1309 2983 1343 3017
rect 1377 2983 1411 3017
rect 1445 2983 1479 3017
rect 1513 2983 1547 3017
rect 1581 2983 1615 3017
rect 1649 2983 1683 3017
rect 1717 2983 1751 3017
rect 1785 2983 1819 3017
rect 1853 2983 1887 3017
rect 1921 2983 1955 3017
rect 1989 2983 2023 3017
rect 2057 2983 2091 3017
rect 2125 2983 2159 3017
rect 2193 2983 2227 3017
rect 2261 2983 2295 3017
rect 2329 2983 2363 3017
rect 2397 2983 2431 3017
rect 2465 2983 2499 3017
rect 2533 2983 2567 3017
rect 2601 2983 2635 3017
rect 2669 2983 2703 3017
rect 2737 2983 2771 3017
rect 2805 2983 2839 3017
rect 2873 2983 2907 3017
rect 2941 2983 2975 3017
rect 3009 2983 3043 3017
rect 3077 2983 3111 3017
rect 3145 2983 3179 3017
rect 3213 2983 3247 3017
rect 3281 2983 3315 3017
rect 3349 2983 3383 3017
rect 3417 2983 3451 3017
rect 3485 2983 3519 3017
rect 3553 2983 3587 3017
rect 3621 2983 3655 3017
rect 3689 2983 3723 3017
rect 3757 2983 3791 3017
rect 3825 2983 3859 3017
rect 3893 2983 3927 3017
rect 3961 2983 3995 3017
rect 4029 2983 4063 3017
rect 4097 2983 4131 3017
rect 4165 2983 4199 3017
rect 4233 2983 4267 3017
rect 4301 2983 4335 3017
rect 4369 2983 4403 3017
rect 4437 2983 4560 3017
rect -480 2960 4560 2983
rect -480 2879 -400 2960
rect -480 2845 -457 2879
rect -423 2845 -400 2879
rect -480 2811 -400 2845
rect -480 2777 -457 2811
rect -423 2777 -400 2811
rect -480 2743 -400 2777
rect -480 2709 -457 2743
rect -423 2709 -400 2743
rect -480 2675 -400 2709
rect -480 2641 -457 2675
rect -423 2641 -400 2675
rect -480 2607 -400 2641
rect -480 2573 -457 2607
rect -423 2573 -400 2607
rect -480 2539 -400 2573
rect -480 2505 -457 2539
rect -423 2505 -400 2539
rect -480 2471 -400 2505
rect -480 2437 -457 2471
rect -423 2437 -400 2471
rect -480 2403 -400 2437
rect -480 2369 -457 2403
rect -423 2369 -400 2403
rect -480 2335 -400 2369
rect -480 2301 -457 2335
rect -423 2301 -400 2335
rect -480 2267 -400 2301
rect -480 2233 -457 2267
rect -423 2233 -400 2267
rect -480 2199 -400 2233
rect -480 2165 -457 2199
rect -423 2165 -400 2199
rect -480 2131 -400 2165
rect -480 2097 -457 2131
rect -423 2097 -400 2131
rect -480 2063 -400 2097
rect -480 2029 -457 2063
rect -423 2029 -400 2063
rect -480 1995 -400 2029
rect -320 2857 4400 2880
rect -320 2823 -187 2857
rect -153 2823 -119 2857
rect -85 2823 -51 2857
rect -17 2823 17 2857
rect 51 2823 85 2857
rect 119 2823 153 2857
rect 187 2823 221 2857
rect 255 2823 289 2857
rect 323 2823 357 2857
rect 391 2823 425 2857
rect 459 2823 493 2857
rect 527 2823 561 2857
rect 595 2823 629 2857
rect 663 2823 697 2857
rect 731 2823 765 2857
rect 799 2823 833 2857
rect 867 2823 901 2857
rect 935 2823 969 2857
rect 1003 2823 1037 2857
rect 1071 2823 1105 2857
rect 1139 2823 1173 2857
rect 1207 2823 1241 2857
rect 1275 2823 1309 2857
rect 1343 2823 1377 2857
rect 1411 2823 1445 2857
rect 1479 2823 1513 2857
rect 1547 2823 1581 2857
rect 1615 2823 1649 2857
rect 1683 2823 1717 2857
rect 1751 2823 1785 2857
rect 1819 2823 1853 2857
rect 1887 2823 1921 2857
rect 1955 2823 1989 2857
rect 2023 2823 2057 2857
rect 2091 2823 2125 2857
rect 2159 2823 2193 2857
rect 2227 2823 2261 2857
rect 2295 2823 2329 2857
rect 2363 2823 2397 2857
rect 2431 2823 2465 2857
rect 2499 2823 2533 2857
rect 2567 2823 2601 2857
rect 2635 2823 2669 2857
rect 2703 2823 2737 2857
rect 2771 2823 2805 2857
rect 2839 2823 2873 2857
rect 2907 2823 2941 2857
rect 2975 2823 3009 2857
rect 3043 2823 3077 2857
rect 3111 2823 3145 2857
rect 3179 2823 3213 2857
rect 3247 2823 3281 2857
rect 3315 2823 3349 2857
rect 3383 2823 3417 2857
rect 3451 2823 3485 2857
rect 3519 2823 3553 2857
rect 3587 2823 3621 2857
rect 3655 2823 3689 2857
rect 3723 2823 3757 2857
rect 3791 2823 3825 2857
rect 3859 2823 3893 2857
rect 3927 2823 3961 2857
rect 3995 2823 4029 2857
rect 4063 2823 4097 2857
rect 4131 2823 4165 2857
rect 4217 2823 4233 2857
rect 4267 2823 4400 2857
rect -320 2800 4400 2823
rect -320 2783 -240 2800
rect -320 2749 -297 2783
rect -263 2749 -240 2783
rect -320 2715 -240 2749
rect 4320 2783 4400 2800
rect 4320 2749 4343 2783
rect 4377 2749 4400 2783
rect -320 2681 -297 2715
rect -263 2681 -240 2715
rect -320 2647 -240 2681
rect -320 2613 -297 2647
rect -263 2613 -240 2647
rect 40 2697 4040 2720
rect 40 2663 79 2697
rect 119 2663 151 2697
rect 187 2663 221 2697
rect 257 2663 289 2697
rect 329 2663 357 2697
rect 401 2663 425 2697
rect 473 2663 493 2697
rect 545 2663 561 2697
rect 617 2663 629 2697
rect 689 2663 697 2697
rect 761 2663 765 2697
rect 867 2663 871 2697
rect 935 2663 943 2697
rect 1003 2663 1015 2697
rect 1071 2663 1087 2697
rect 1139 2663 1159 2697
rect 1207 2663 1231 2697
rect 1275 2663 1303 2697
rect 1343 2663 1375 2697
rect 1411 2663 1445 2697
rect 1481 2663 1513 2697
rect 1553 2663 1581 2697
rect 1625 2663 1649 2697
rect 1697 2663 1717 2697
rect 1769 2663 1785 2697
rect 1841 2663 1853 2697
rect 1913 2663 1921 2697
rect 1985 2663 1989 2697
rect 2091 2663 2095 2697
rect 2159 2663 2167 2697
rect 2227 2663 2239 2697
rect 2295 2663 2311 2697
rect 2363 2663 2383 2697
rect 2431 2663 2455 2697
rect 2499 2663 2527 2697
rect 2567 2663 2599 2697
rect 2635 2663 2669 2697
rect 2705 2663 2737 2697
rect 2777 2663 2805 2697
rect 2849 2663 2873 2697
rect 2921 2663 2941 2697
rect 2993 2663 3009 2697
rect 3065 2663 3077 2697
rect 3137 2663 3145 2697
rect 3209 2663 3213 2697
rect 3315 2663 3319 2697
rect 3383 2663 3391 2697
rect 3451 2663 3463 2697
rect 3519 2663 3535 2697
rect 3587 2663 3607 2697
rect 3655 2663 3679 2697
rect 3723 2663 3751 2697
rect 3791 2663 3823 2697
rect 3859 2663 3893 2697
rect 3929 2663 3961 2697
rect 4001 2663 4040 2697
rect 40 2640 4040 2663
rect 4320 2715 4400 2749
rect 4320 2681 4343 2715
rect 4377 2681 4400 2715
rect 4320 2647 4400 2681
rect -320 2579 -240 2613
rect -320 2545 -297 2579
rect -263 2545 -240 2579
rect 4320 2613 4343 2647
rect 4377 2613 4400 2647
rect 4320 2579 4400 2613
rect -320 2511 -240 2545
rect -320 2477 -297 2511
rect -263 2477 -240 2511
rect -160 2537 -80 2564
rect -160 2503 -137 2537
rect -103 2503 -80 2537
rect -160 2480 -80 2503
rect 4160 2537 4240 2564
rect 4160 2503 4183 2537
rect 4217 2503 4240 2537
rect 4160 2480 4240 2503
rect 4320 2545 4343 2579
rect 4377 2545 4400 2579
rect 4320 2511 4400 2545
rect -320 2443 -240 2477
rect -320 2409 -297 2443
rect -263 2409 -240 2443
rect -320 2375 -240 2409
rect 4320 2477 4343 2511
rect 4377 2477 4400 2511
rect 4320 2443 4400 2477
rect 4320 2409 4343 2443
rect 4377 2409 4400 2443
rect -320 2341 -297 2375
rect -263 2341 -240 2375
rect -320 2307 -240 2341
rect 40 2377 4040 2400
rect 40 2343 79 2377
rect 119 2343 151 2377
rect 187 2343 221 2377
rect 257 2343 289 2377
rect 329 2343 357 2377
rect 401 2343 425 2377
rect 473 2343 493 2377
rect 545 2343 561 2377
rect 617 2343 629 2377
rect 689 2343 697 2377
rect 761 2343 765 2377
rect 867 2343 871 2377
rect 935 2343 943 2377
rect 1003 2343 1015 2377
rect 1071 2343 1087 2377
rect 1139 2343 1159 2377
rect 1207 2343 1231 2377
rect 1275 2343 1303 2377
rect 1343 2343 1375 2377
rect 1411 2343 1445 2377
rect 1481 2343 1513 2377
rect 1553 2343 1581 2377
rect 1625 2343 1649 2377
rect 1697 2343 1717 2377
rect 1769 2343 1785 2377
rect 1841 2343 1853 2377
rect 1913 2343 1921 2377
rect 1985 2343 1989 2377
rect 2091 2343 2095 2377
rect 2159 2343 2167 2377
rect 2227 2343 2239 2377
rect 2295 2343 2311 2377
rect 2363 2343 2383 2377
rect 2431 2343 2455 2377
rect 2499 2343 2527 2377
rect 2567 2343 2599 2377
rect 2635 2343 2669 2377
rect 2705 2343 2737 2377
rect 2777 2343 2805 2377
rect 2849 2343 2873 2377
rect 2921 2343 2941 2377
rect 2993 2343 3009 2377
rect 3065 2343 3077 2377
rect 3137 2343 3145 2377
rect 3209 2343 3213 2377
rect 3315 2343 3319 2377
rect 3383 2343 3391 2377
rect 3451 2343 3463 2377
rect 3519 2343 3535 2377
rect 3587 2343 3607 2377
rect 3655 2343 3679 2377
rect 3723 2343 3751 2377
rect 3791 2343 3823 2377
rect 3859 2343 3893 2377
rect 3929 2343 3961 2377
rect 4001 2343 4040 2377
rect 40 2320 4040 2343
rect 4320 2375 4400 2409
rect 4320 2341 4343 2375
rect 4377 2341 4400 2375
rect -320 2273 -297 2307
rect -263 2273 -240 2307
rect -320 2239 -240 2273
rect 4320 2307 4400 2341
rect 4320 2273 4343 2307
rect 4377 2273 4400 2307
rect -320 2205 -297 2239
rect -263 2205 -240 2239
rect -320 2171 -240 2205
rect -320 2137 -297 2171
rect -263 2137 -240 2171
rect -160 2217 -80 2244
rect -160 2183 -137 2217
rect -103 2183 -80 2217
rect -160 2160 -80 2183
rect 4160 2217 4240 2244
rect 4160 2183 4183 2217
rect 4217 2183 4240 2217
rect 4160 2160 4240 2183
rect 4320 2239 4400 2273
rect 4320 2205 4343 2239
rect 4377 2205 4400 2239
rect 4320 2171 4400 2205
rect -320 2080 -240 2137
rect 4320 2137 4343 2171
rect 4377 2137 4400 2171
rect 4320 2080 4400 2137
rect -320 2057 4400 2080
rect -320 2023 -187 2057
rect -153 2023 -119 2057
rect -85 2023 -51 2057
rect -17 2023 17 2057
rect 51 2023 85 2057
rect 119 2023 153 2057
rect 187 2023 221 2057
rect 255 2023 289 2057
rect 323 2023 357 2057
rect 391 2023 425 2057
rect 459 2023 493 2057
rect 527 2023 561 2057
rect 595 2023 629 2057
rect 663 2023 697 2057
rect 731 2023 765 2057
rect 799 2023 833 2057
rect 867 2023 901 2057
rect 935 2023 969 2057
rect 1003 2023 1037 2057
rect 1071 2023 1105 2057
rect 1139 2023 1173 2057
rect 1207 2023 1241 2057
rect 1275 2023 1309 2057
rect 1343 2023 1377 2057
rect 1411 2023 1445 2057
rect 1479 2023 1513 2057
rect 1547 2023 1581 2057
rect 1615 2023 1649 2057
rect 1683 2023 1717 2057
rect 1751 2023 1785 2057
rect 1819 2023 1853 2057
rect 1887 2023 1921 2057
rect 1955 2023 1989 2057
rect 2023 2023 2057 2057
rect 2091 2023 2125 2057
rect 2159 2023 2193 2057
rect 2227 2023 2261 2057
rect 2295 2023 2329 2057
rect 2363 2023 2397 2057
rect 2431 2023 2465 2057
rect 2499 2023 2533 2057
rect 2567 2023 2601 2057
rect 2635 2023 2669 2057
rect 2703 2023 2737 2057
rect 2771 2023 2805 2057
rect 2839 2023 2873 2057
rect 2907 2023 2941 2057
rect 2975 2023 3009 2057
rect 3043 2023 3077 2057
rect 3111 2023 3145 2057
rect 3179 2023 3213 2057
rect 3247 2023 3281 2057
rect 3315 2023 3349 2057
rect 3383 2023 3417 2057
rect 3451 2023 3485 2057
rect 3519 2023 3553 2057
rect 3587 2023 3621 2057
rect 3655 2023 3689 2057
rect 3723 2023 3757 2057
rect 3791 2023 3825 2057
rect 3859 2023 3893 2057
rect 3927 2023 3961 2057
rect 3995 2023 4029 2057
rect 4063 2023 4097 2057
rect 4131 2023 4165 2057
rect 4199 2023 4233 2057
rect 4267 2023 4400 2057
rect -320 2000 4400 2023
rect 4480 2879 4560 2960
rect 4480 2845 4503 2879
rect 4537 2845 4560 2879
rect 4480 2811 4560 2845
rect 4480 2777 4503 2811
rect 4537 2777 4560 2811
rect 4480 2743 4560 2777
rect 4480 2709 4503 2743
rect 4537 2709 4560 2743
rect 4480 2675 4560 2709
rect 4480 2641 4503 2675
rect 4537 2641 4560 2675
rect 4480 2607 4560 2641
rect 4480 2573 4503 2607
rect 4537 2573 4560 2607
rect 4480 2539 4560 2573
rect 4480 2505 4503 2539
rect 4537 2505 4560 2539
rect 4480 2471 4560 2505
rect 4480 2437 4503 2471
rect 4537 2437 4560 2471
rect 4480 2403 4560 2437
rect 4480 2369 4503 2403
rect 4537 2369 4560 2403
rect 4480 2335 4560 2369
rect 4480 2301 4503 2335
rect 4537 2301 4560 2335
rect 4480 2267 4560 2301
rect 4480 2233 4503 2267
rect 4537 2233 4560 2267
rect 4480 2199 4560 2233
rect 4480 2165 4503 2199
rect 4537 2165 4560 2199
rect 4480 2131 4560 2165
rect 4480 2097 4503 2131
rect 4537 2097 4560 2131
rect 4480 2063 4560 2097
rect 4480 2029 4503 2063
rect 4537 2029 4560 2063
rect -480 1961 -457 1995
rect -423 1961 -400 1995
rect -480 1920 -400 1961
rect 4480 1995 4560 2029
rect 4480 1961 4503 1995
rect 4537 1961 4560 1995
rect 4480 1920 4560 1961
rect -480 1897 4560 1920
rect -480 1863 -357 1897
rect -323 1863 -289 1897
rect -255 1863 -221 1897
rect -187 1863 -153 1897
rect -119 1863 -85 1897
rect -51 1863 -17 1897
rect 17 1863 51 1897
rect 85 1863 119 1897
rect 153 1863 187 1897
rect 221 1863 255 1897
rect 289 1863 323 1897
rect 357 1863 391 1897
rect 425 1863 459 1897
rect 493 1863 527 1897
rect 561 1863 595 1897
rect 629 1863 663 1897
rect 697 1863 731 1897
rect 765 1863 799 1897
rect 833 1863 867 1897
rect 901 1863 935 1897
rect 969 1863 1003 1897
rect 1037 1863 1071 1897
rect 1105 1863 1139 1897
rect 1173 1863 1207 1897
rect 1241 1863 1275 1897
rect 1309 1863 1343 1897
rect 1377 1863 1411 1897
rect 1445 1863 1479 1897
rect 1513 1863 1547 1897
rect 1581 1863 1615 1897
rect 1649 1863 1683 1897
rect 1717 1863 1751 1897
rect 1785 1863 1819 1897
rect 1853 1863 1887 1897
rect 1921 1863 1955 1897
rect 1989 1863 2023 1897
rect 2057 1863 2091 1897
rect 2125 1863 2159 1897
rect 2193 1863 2227 1897
rect 2261 1863 2295 1897
rect 2329 1863 2363 1897
rect 2397 1863 2431 1897
rect 2465 1863 2499 1897
rect 2533 1863 2567 1897
rect 2601 1863 2635 1897
rect 2669 1863 2703 1897
rect 2737 1863 2771 1897
rect 2805 1863 2839 1897
rect 2873 1863 2907 1897
rect 2941 1863 2975 1897
rect 3009 1863 3043 1897
rect 3077 1863 3111 1897
rect 3145 1863 3179 1897
rect 3213 1863 3247 1897
rect 3281 1863 3315 1897
rect 3349 1863 3383 1897
rect 3417 1863 3451 1897
rect 3485 1863 3519 1897
rect 3553 1863 3587 1897
rect 3621 1863 3655 1897
rect 3689 1863 3723 1897
rect 3757 1863 3791 1897
rect 3825 1863 3859 1897
rect 3893 1863 3927 1897
rect 3961 1863 3995 1897
rect 4029 1863 4063 1897
rect 4097 1863 4131 1897
rect 4165 1863 4199 1897
rect 4233 1863 4267 1897
rect 4301 1863 4335 1897
rect 4369 1863 4403 1897
rect 4437 1863 4560 1897
rect -480 1840 4560 1863
rect -480 1817 -160 1840
rect -480 1783 -297 1817
rect -263 1783 -160 1817
rect -480 1760 -160 1783
rect 4480 1760 4560 1840
rect -480 1737 4560 1760
rect -480 1703 -357 1737
rect -323 1703 -289 1737
rect -255 1703 -221 1737
rect -187 1703 -153 1737
rect -119 1703 -85 1737
rect -51 1703 -17 1737
rect 17 1703 51 1737
rect 85 1703 119 1737
rect 153 1703 187 1737
rect 221 1703 255 1737
rect 289 1703 323 1737
rect 357 1703 391 1737
rect 425 1703 459 1737
rect 493 1703 527 1737
rect 561 1703 595 1737
rect 629 1703 663 1737
rect 697 1703 731 1737
rect 765 1703 799 1737
rect 833 1703 867 1737
rect 901 1703 935 1737
rect 969 1703 1003 1737
rect 1037 1703 1071 1737
rect 1105 1703 1139 1737
rect 1173 1703 1207 1737
rect 1241 1703 1275 1737
rect 1309 1703 1343 1737
rect 1377 1703 1411 1737
rect 1445 1703 1479 1737
rect 1513 1703 1547 1737
rect 1581 1703 1615 1737
rect 1649 1703 1683 1737
rect 1717 1703 1751 1737
rect 1785 1703 1819 1737
rect 1853 1703 1887 1737
rect 1921 1703 1955 1737
rect 1989 1703 2023 1737
rect 2057 1703 2091 1737
rect 2125 1703 2159 1737
rect 2193 1703 2227 1737
rect 2261 1703 2295 1737
rect 2329 1703 2363 1737
rect 2397 1703 2431 1737
rect 2465 1703 2499 1737
rect 2533 1703 2567 1737
rect 2601 1703 2635 1737
rect 2669 1703 2703 1737
rect 2737 1703 2771 1737
rect 2805 1703 2839 1737
rect 2873 1703 2907 1737
rect 2941 1703 2975 1737
rect 3009 1703 3043 1737
rect 3077 1703 3111 1737
rect 3145 1703 3179 1737
rect 3213 1703 3247 1737
rect 3281 1703 3315 1737
rect 3349 1703 3383 1737
rect 3417 1703 3451 1737
rect 3485 1703 3519 1737
rect 3553 1703 3587 1737
rect 3621 1703 3655 1737
rect 3689 1703 3723 1737
rect 3757 1703 3791 1737
rect 3825 1703 3859 1737
rect 3893 1703 3927 1737
rect 3961 1703 3995 1737
rect 4029 1703 4063 1737
rect 4097 1703 4131 1737
rect 4165 1703 4199 1737
rect 4233 1703 4267 1737
rect 4301 1703 4335 1737
rect 4369 1703 4403 1737
rect 4437 1703 4560 1737
rect -480 1680 4560 1703
rect -480 1639 -400 1680
rect -480 1605 -457 1639
rect -423 1605 -400 1639
rect -480 1571 -400 1605
rect 4480 1639 4560 1680
rect 4480 1605 4503 1639
rect 4537 1605 4560 1639
rect -480 1537 -457 1571
rect -423 1537 -400 1571
rect -480 1503 -400 1537
rect -480 1469 -457 1503
rect -423 1469 -400 1503
rect -480 1435 -400 1469
rect -480 1401 -457 1435
rect -423 1401 -400 1435
rect -480 1367 -400 1401
rect -480 1333 -457 1367
rect -423 1333 -400 1367
rect -480 1299 -400 1333
rect -480 1265 -457 1299
rect -423 1265 -400 1299
rect -480 1231 -400 1265
rect -480 1197 -457 1231
rect -423 1197 -400 1231
rect -480 1163 -400 1197
rect -480 1129 -457 1163
rect -423 1129 -400 1163
rect -480 1095 -400 1129
rect -480 1061 -457 1095
rect -423 1061 -400 1095
rect -480 1027 -400 1061
rect -480 993 -457 1027
rect -423 993 -400 1027
rect -480 959 -400 993
rect -480 925 -457 959
rect -423 925 -400 959
rect -480 891 -400 925
rect -480 857 -457 891
rect -423 857 -400 891
rect -480 823 -400 857
rect -480 789 -457 823
rect -423 789 -400 823
rect -480 755 -400 789
rect -480 721 -457 755
rect -423 721 -400 755
rect -480 640 -400 721
rect -320 1577 4400 1600
rect -320 1543 -187 1577
rect -153 1543 -119 1577
rect -85 1543 -51 1577
rect -17 1543 17 1577
rect 51 1543 85 1577
rect 119 1543 153 1577
rect 187 1543 221 1577
rect 255 1543 289 1577
rect 323 1543 357 1577
rect 391 1543 425 1577
rect 459 1543 493 1577
rect 527 1543 561 1577
rect 595 1543 629 1577
rect 663 1543 697 1577
rect 731 1543 765 1577
rect 799 1543 833 1577
rect 867 1543 901 1577
rect 935 1543 969 1577
rect 1003 1543 1037 1577
rect 1071 1543 1105 1577
rect 1139 1543 1173 1577
rect 1207 1543 1241 1577
rect 1275 1543 1309 1577
rect 1343 1543 1377 1577
rect 1411 1543 1445 1577
rect 1479 1543 1513 1577
rect 1547 1543 1581 1577
rect 1615 1543 1649 1577
rect 1683 1543 1717 1577
rect 1751 1543 1785 1577
rect 1819 1543 1853 1577
rect 1887 1543 1921 1577
rect 1955 1543 1989 1577
rect 2023 1543 2057 1577
rect 2091 1543 2125 1577
rect 2159 1543 2193 1577
rect 2227 1543 2261 1577
rect 2295 1543 2329 1577
rect 2363 1543 2397 1577
rect 2431 1543 2465 1577
rect 2499 1543 2533 1577
rect 2567 1543 2601 1577
rect 2635 1543 2669 1577
rect 2703 1543 2737 1577
rect 2771 1543 2805 1577
rect 2839 1543 2873 1577
rect 2907 1543 2941 1577
rect 2975 1543 3009 1577
rect 3043 1543 3077 1577
rect 3111 1543 3145 1577
rect 3179 1543 3213 1577
rect 3247 1543 3281 1577
rect 3315 1543 3349 1577
rect 3383 1543 3417 1577
rect 3451 1543 3485 1577
rect 3519 1543 3553 1577
rect 3587 1543 3621 1577
rect 3655 1543 3689 1577
rect 3723 1543 3757 1577
rect 3791 1543 3825 1577
rect 3859 1543 3893 1577
rect 3927 1543 3961 1577
rect 3995 1543 4029 1577
rect 4063 1543 4097 1577
rect 4131 1543 4165 1577
rect 4199 1543 4233 1577
rect 4267 1543 4400 1577
rect -320 1520 4400 1543
rect -320 1463 -240 1520
rect -320 1429 -297 1463
rect -263 1429 -240 1463
rect 4320 1463 4400 1520
rect -320 1395 -240 1429
rect -320 1361 -297 1395
rect -263 1361 -240 1395
rect -320 1327 -240 1361
rect -160 1417 -80 1440
rect -160 1383 -137 1417
rect -103 1383 -80 1417
rect -160 1356 -80 1383
rect 4160 1417 4240 1440
rect 4160 1383 4183 1417
rect 4217 1383 4240 1417
rect 4160 1356 4240 1383
rect 4320 1429 4343 1463
rect 4377 1429 4400 1463
rect 4320 1395 4400 1429
rect 4320 1361 4343 1395
rect 4377 1361 4400 1395
rect -320 1293 -297 1327
rect -263 1293 -240 1327
rect -320 1259 -240 1293
rect 4320 1327 4400 1361
rect 4320 1293 4343 1327
rect 4377 1293 4400 1327
rect -320 1225 -297 1259
rect -263 1225 -240 1259
rect -320 1191 -240 1225
rect 40 1257 4040 1280
rect 40 1223 79 1257
rect 119 1223 151 1257
rect 187 1223 221 1257
rect 257 1223 289 1257
rect 329 1223 357 1257
rect 401 1223 425 1257
rect 473 1223 493 1257
rect 545 1223 561 1257
rect 617 1223 629 1257
rect 689 1223 697 1257
rect 761 1223 765 1257
rect 867 1223 871 1257
rect 935 1223 943 1257
rect 1003 1223 1015 1257
rect 1071 1223 1087 1257
rect 1139 1223 1159 1257
rect 1207 1223 1231 1257
rect 1275 1223 1303 1257
rect 1343 1223 1375 1257
rect 1411 1223 1445 1257
rect 1481 1223 1513 1257
rect 1553 1223 1581 1257
rect 1625 1223 1649 1257
rect 1697 1223 1717 1257
rect 1769 1223 1785 1257
rect 1841 1223 1853 1257
rect 1913 1223 1921 1257
rect 1985 1223 1989 1257
rect 2091 1223 2095 1257
rect 2159 1223 2167 1257
rect 2227 1223 2239 1257
rect 2295 1223 2311 1257
rect 2363 1223 2383 1257
rect 2431 1223 2455 1257
rect 2499 1223 2527 1257
rect 2567 1223 2599 1257
rect 2635 1223 2669 1257
rect 2705 1223 2737 1257
rect 2777 1223 2805 1257
rect 2849 1223 2873 1257
rect 2921 1223 2941 1257
rect 2993 1223 3009 1257
rect 3065 1223 3077 1257
rect 3137 1223 3145 1257
rect 3209 1223 3213 1257
rect 3315 1223 3319 1257
rect 3383 1223 3391 1257
rect 3451 1223 3463 1257
rect 3519 1223 3535 1257
rect 3587 1223 3607 1257
rect 3655 1223 3679 1257
rect 3723 1223 3751 1257
rect 3791 1223 3823 1257
rect 3859 1223 3893 1257
rect 3929 1223 3961 1257
rect 4001 1223 4040 1257
rect 40 1200 4040 1223
rect 4320 1259 4400 1293
rect 4320 1225 4343 1259
rect 4377 1225 4400 1259
rect -320 1157 -297 1191
rect -263 1157 -240 1191
rect -320 1123 -240 1157
rect -320 1089 -297 1123
rect -263 1089 -240 1123
rect 4320 1191 4400 1225
rect 4320 1157 4343 1191
rect 4377 1157 4400 1191
rect 4320 1123 4400 1157
rect -320 1055 -240 1089
rect -320 1021 -297 1055
rect -263 1021 -240 1055
rect -160 1097 -80 1120
rect -160 1063 -137 1097
rect -103 1063 -80 1097
rect -160 1036 -80 1063
rect 4160 1097 4240 1120
rect 4160 1063 4183 1097
rect 4217 1063 4240 1097
rect 4160 1036 4240 1063
rect 4320 1089 4343 1123
rect 4377 1089 4400 1123
rect 4320 1055 4400 1089
rect -320 987 -240 1021
rect -320 953 -297 987
rect -263 953 -240 987
rect 4320 1021 4343 1055
rect 4377 1021 4400 1055
rect 4320 987 4400 1021
rect -320 919 -240 953
rect -320 885 -297 919
rect -263 885 -240 919
rect -320 851 -240 885
rect 40 937 4040 960
rect 40 903 79 937
rect 119 903 151 937
rect 187 903 221 937
rect 257 903 289 937
rect 329 903 357 937
rect 401 903 425 937
rect 473 903 493 937
rect 545 903 561 937
rect 617 903 629 937
rect 689 903 697 937
rect 761 903 765 937
rect 867 903 871 937
rect 935 903 943 937
rect 1003 903 1015 937
rect 1071 903 1087 937
rect 1139 903 1159 937
rect 1207 903 1231 937
rect 1275 903 1303 937
rect 1343 903 1375 937
rect 1411 903 1445 937
rect 1481 903 1513 937
rect 1553 903 1581 937
rect 1625 903 1649 937
rect 1697 903 1717 937
rect 1769 903 1785 937
rect 1841 903 1853 937
rect 1913 903 1921 937
rect 1985 903 1989 937
rect 2091 903 2095 937
rect 2159 903 2167 937
rect 2227 903 2239 937
rect 2295 903 2311 937
rect 2363 903 2383 937
rect 2431 903 2455 937
rect 2499 903 2527 937
rect 2567 903 2599 937
rect 2635 903 2669 937
rect 2705 903 2737 937
rect 2777 903 2805 937
rect 2849 903 2873 937
rect 2921 903 2941 937
rect 2993 903 3009 937
rect 3065 903 3077 937
rect 3137 903 3145 937
rect 3209 903 3213 937
rect 3315 903 3319 937
rect 3383 903 3391 937
rect 3451 903 3463 937
rect 3519 903 3535 937
rect 3587 903 3607 937
rect 3655 903 3679 937
rect 3723 903 3751 937
rect 3791 903 3823 937
rect 3859 903 3893 937
rect 3929 903 3961 937
rect 4001 903 4040 937
rect 40 880 4040 903
rect 4320 953 4343 987
rect 4377 953 4400 987
rect 4320 919 4400 953
rect 4320 885 4343 919
rect 4377 885 4400 919
rect -320 817 -297 851
rect -263 817 -240 851
rect -320 800 -240 817
rect 4320 851 4400 885
rect 4320 817 4343 851
rect 4377 817 4400 851
rect 4320 800 4400 817
rect -320 777 4400 800
rect -320 743 -187 777
rect -153 743 -119 777
rect -85 743 -51 777
rect -17 743 17 777
rect 51 743 85 777
rect 119 743 153 777
rect 187 743 221 777
rect 255 743 289 777
rect 323 743 357 777
rect 391 743 425 777
rect 459 743 493 777
rect 527 743 561 777
rect 595 743 629 777
rect 663 743 697 777
rect 731 743 765 777
rect 799 743 833 777
rect 867 743 901 777
rect 935 743 969 777
rect 1003 743 1037 777
rect 1071 743 1105 777
rect 1139 743 1173 777
rect 1207 743 1241 777
rect 1275 743 1309 777
rect 1343 743 1377 777
rect 1411 743 1445 777
rect 1479 743 1513 777
rect 1547 743 1581 777
rect 1615 743 1649 777
rect 1683 743 1717 777
rect 1751 743 1785 777
rect 1819 743 1853 777
rect 1887 743 1921 777
rect 1955 743 1989 777
rect 2023 743 2057 777
rect 2091 743 2125 777
rect 2159 743 2193 777
rect 2227 743 2261 777
rect 2295 743 2329 777
rect 2363 743 2397 777
rect 2431 743 2465 777
rect 2499 743 2533 777
rect 2567 743 2601 777
rect 2635 743 2669 777
rect 2703 743 2737 777
rect 2771 743 2805 777
rect 2839 743 2873 777
rect 2907 743 2941 777
rect 2975 743 3009 777
rect 3043 743 3077 777
rect 3111 743 3145 777
rect 3179 743 3213 777
rect 3247 743 3281 777
rect 3315 743 3349 777
rect 3383 743 3417 777
rect 3451 743 3485 777
rect 3519 743 3553 777
rect 3587 743 3621 777
rect 3655 743 3689 777
rect 3723 743 3757 777
rect 3791 743 3825 777
rect 3859 743 3893 777
rect 3927 743 3961 777
rect 3995 743 4029 777
rect 4063 743 4097 777
rect 4131 743 4165 777
rect 4217 743 4233 777
rect 4267 743 4400 777
rect -320 720 4400 743
rect 4480 1571 4560 1605
rect 4480 1537 4503 1571
rect 4537 1537 4560 1571
rect 4480 1503 4560 1537
rect 4480 1469 4503 1503
rect 4537 1469 4560 1503
rect 4480 1435 4560 1469
rect 4480 1401 4503 1435
rect 4537 1401 4560 1435
rect 4480 1367 4560 1401
rect 4480 1333 4503 1367
rect 4537 1333 4560 1367
rect 4480 1299 4560 1333
rect 4480 1265 4503 1299
rect 4537 1265 4560 1299
rect 4480 1231 4560 1265
rect 4480 1197 4503 1231
rect 4537 1197 4560 1231
rect 4480 1163 4560 1197
rect 4480 1129 4503 1163
rect 4537 1129 4560 1163
rect 4480 1095 4560 1129
rect 4480 1061 4503 1095
rect 4537 1061 4560 1095
rect 4480 1027 4560 1061
rect 4480 993 4503 1027
rect 4537 993 4560 1027
rect 4480 959 4560 993
rect 4480 925 4503 959
rect 4537 925 4560 959
rect 4480 891 4560 925
rect 4480 857 4503 891
rect 4537 857 4560 891
rect 4480 823 4560 857
rect 4480 789 4503 823
rect 4537 789 4560 823
rect 4480 755 4560 789
rect 4480 721 4503 755
rect 4537 721 4560 755
rect 4480 640 4560 721
rect -480 617 4560 640
rect -480 583 -357 617
rect -323 583 -289 617
rect -255 583 -221 617
rect -187 583 -153 617
rect -119 583 -85 617
rect -51 583 -17 617
rect 17 583 51 617
rect 85 583 119 617
rect 153 583 187 617
rect 221 583 255 617
rect 289 583 323 617
rect 357 583 391 617
rect 425 583 459 617
rect 493 583 527 617
rect 561 583 595 617
rect 629 583 663 617
rect 697 583 731 617
rect 765 583 799 617
rect 833 583 867 617
rect 901 583 935 617
rect 969 583 1003 617
rect 1037 583 1071 617
rect 1105 583 1139 617
rect 1173 583 1207 617
rect 1241 583 1275 617
rect 1309 583 1343 617
rect 1377 583 1411 617
rect 1445 583 1479 617
rect 1513 583 1547 617
rect 1581 583 1615 617
rect 1649 583 1683 617
rect 1717 583 1751 617
rect 1785 583 1819 617
rect 1853 583 1887 617
rect 1921 583 1955 617
rect 1989 583 2023 617
rect 2057 583 2091 617
rect 2125 583 2159 617
rect 2193 583 2227 617
rect 2261 583 2295 617
rect 2329 583 2363 617
rect 2397 583 2431 617
rect 2465 583 2499 617
rect 2533 583 2567 617
rect 2601 583 2635 617
rect 2669 583 2703 617
rect 2737 583 2771 617
rect 2805 583 2839 617
rect 2873 583 2907 617
rect 2941 583 2975 617
rect 3009 583 3043 617
rect 3077 583 3111 617
rect 3145 583 3179 617
rect 3213 583 3247 617
rect 3281 583 3315 617
rect 3349 583 3383 617
rect 3417 583 3451 617
rect 3485 583 3519 617
rect 3553 583 3587 617
rect 3621 583 3655 617
rect 3689 583 3723 617
rect 3757 583 3791 617
rect 3825 583 3859 617
rect 3893 583 3927 617
rect 3961 583 3995 617
rect 4029 583 4063 617
rect 4097 583 4131 617
rect 4165 583 4199 617
rect 4233 583 4267 617
rect 4301 583 4335 617
rect 4369 583 4403 617
rect 4437 583 4560 617
rect -480 560 4560 583
rect -480 480 -400 560
rect 4480 480 4560 560
rect -480 457 4560 480
rect -480 423 -357 457
rect -323 423 -289 457
rect -255 423 -221 457
rect -187 423 -153 457
rect -119 423 -85 457
rect -51 423 -17 457
rect 17 423 51 457
rect 85 423 119 457
rect 153 423 187 457
rect 221 423 255 457
rect 289 423 323 457
rect 357 423 391 457
rect 425 423 459 457
rect 493 423 527 457
rect 561 423 595 457
rect 629 423 663 457
rect 697 423 731 457
rect 765 423 799 457
rect 833 423 867 457
rect 901 423 935 457
rect 969 423 1003 457
rect 1037 423 1071 457
rect 1105 423 1139 457
rect 1173 423 1207 457
rect 1241 423 1275 457
rect 1309 423 1343 457
rect 1377 423 1411 457
rect 1445 423 1479 457
rect 1513 423 1547 457
rect 1581 423 1615 457
rect 1649 423 1683 457
rect 1717 423 1751 457
rect 1785 423 1819 457
rect 1853 423 1887 457
rect 1921 423 1955 457
rect 1989 423 2023 457
rect 2057 423 2091 457
rect 2125 423 2159 457
rect 2193 423 2227 457
rect 2261 423 2295 457
rect 2329 423 2363 457
rect 2397 423 2431 457
rect 2465 423 2499 457
rect 2533 423 2567 457
rect 2601 423 2635 457
rect 2669 423 2703 457
rect 2737 423 2771 457
rect 2805 423 2839 457
rect 2873 423 2907 457
rect 2941 423 2975 457
rect 3009 423 3043 457
rect 3077 423 3111 457
rect 3145 423 3179 457
rect 3213 423 3247 457
rect 3281 423 3315 457
rect 3349 423 3383 457
rect 3417 423 3451 457
rect 3485 423 3519 457
rect 3553 423 3587 457
rect 3621 423 3655 457
rect 3689 423 3723 457
rect 3757 423 3791 457
rect 3825 423 3859 457
rect 3893 423 3927 457
rect 3961 423 3995 457
rect 4029 423 4063 457
rect 4097 423 4131 457
rect 4165 423 4199 457
rect 4233 423 4267 457
rect 4301 423 4335 457
rect 4369 423 4403 457
rect 4437 423 4560 457
rect -480 400 4560 423
rect -480 319 -400 400
rect -480 285 -457 319
rect -423 285 -400 319
rect -480 251 -400 285
rect -480 217 -457 251
rect -423 217 -400 251
rect -480 183 -400 217
rect -480 149 -457 183
rect -423 149 -400 183
rect -480 115 -400 149
rect -480 81 -457 115
rect -423 81 -400 115
rect -480 47 -400 81
rect -480 13 -457 47
rect -423 13 -400 47
rect -480 -21 -400 13
rect -480 -55 -457 -21
rect -423 -55 -400 -21
rect -480 -89 -400 -55
rect -480 -123 -457 -89
rect -423 -123 -400 -89
rect -480 -157 -400 -123
rect -480 -191 -457 -157
rect -423 -191 -400 -157
rect -480 -225 -400 -191
rect -480 -259 -457 -225
rect -423 -259 -400 -225
rect -480 -293 -400 -259
rect -480 -327 -457 -293
rect -423 -327 -400 -293
rect -480 -361 -400 -327
rect -480 -395 -457 -361
rect -423 -395 -400 -361
rect -480 -429 -400 -395
rect -480 -463 -457 -429
rect -423 -463 -400 -429
rect -480 -497 -400 -463
rect -480 -531 -457 -497
rect -423 -531 -400 -497
rect -480 -565 -400 -531
rect -320 297 4400 320
rect -320 263 -187 297
rect -153 263 -119 297
rect -85 263 -51 297
rect -17 263 17 297
rect 51 263 85 297
rect 119 263 153 297
rect 187 263 221 297
rect 255 263 289 297
rect 323 263 357 297
rect 391 263 425 297
rect 459 263 493 297
rect 527 263 561 297
rect 595 263 629 297
rect 663 263 697 297
rect 731 263 765 297
rect 799 263 833 297
rect 867 263 901 297
rect 935 263 969 297
rect 1003 263 1037 297
rect 1071 263 1105 297
rect 1139 263 1173 297
rect 1207 263 1241 297
rect 1275 263 1309 297
rect 1343 263 1377 297
rect 1411 263 1445 297
rect 1479 263 1513 297
rect 1547 263 1581 297
rect 1615 263 1649 297
rect 1683 263 1717 297
rect 1751 263 1785 297
rect 1819 263 1853 297
rect 1887 263 1921 297
rect 1955 263 1989 297
rect 2023 263 2057 297
rect 2091 263 2125 297
rect 2159 263 2193 297
rect 2227 263 2261 297
rect 2295 263 2329 297
rect 2363 263 2397 297
rect 2431 263 2465 297
rect 2499 263 2533 297
rect 2567 263 2601 297
rect 2635 263 2669 297
rect 2703 263 2737 297
rect 2771 263 2805 297
rect 2839 263 2873 297
rect 2907 263 2941 297
rect 2975 263 3009 297
rect 3043 263 3077 297
rect 3111 263 3145 297
rect 3179 263 3213 297
rect 3247 263 3281 297
rect 3315 263 3349 297
rect 3383 263 3417 297
rect 3451 263 3485 297
rect 3519 263 3553 297
rect 3587 263 3621 297
rect 3655 263 3689 297
rect 3723 263 3757 297
rect 3791 263 3825 297
rect 3859 263 3893 297
rect 3927 263 3961 297
rect 3995 263 4029 297
rect 4063 263 4097 297
rect 4131 263 4165 297
rect 4199 263 4233 297
rect 4267 263 4400 297
rect -320 240 4400 263
rect -320 223 -240 240
rect -320 189 -297 223
rect -263 189 -240 223
rect -320 155 -240 189
rect 4320 223 4400 240
rect 4320 189 4343 223
rect 4377 189 4400 223
rect -320 121 -297 155
rect -263 121 -240 155
rect -320 87 -240 121
rect -320 53 -297 87
rect -263 53 -240 87
rect 40 137 4040 160
rect 40 103 79 137
rect 119 103 151 137
rect 187 103 221 137
rect 257 103 289 137
rect 329 103 357 137
rect 401 103 425 137
rect 473 103 493 137
rect 545 103 561 137
rect 617 103 629 137
rect 689 103 697 137
rect 761 103 765 137
rect 867 103 871 137
rect 935 103 943 137
rect 1003 103 1015 137
rect 1071 103 1087 137
rect 1139 103 1159 137
rect 1207 103 1231 137
rect 1275 103 1303 137
rect 1343 103 1375 137
rect 1411 103 1445 137
rect 1481 103 1513 137
rect 1553 103 1581 137
rect 1625 103 1649 137
rect 1697 103 1717 137
rect 1769 103 1785 137
rect 1841 103 1853 137
rect 1913 103 1921 137
rect 1985 103 1989 137
rect 2091 103 2095 137
rect 2159 103 2167 137
rect 2227 103 2239 137
rect 2295 103 2311 137
rect 2363 103 2383 137
rect 2431 103 2455 137
rect 2499 103 2527 137
rect 2567 103 2599 137
rect 2635 103 2669 137
rect 2705 103 2737 137
rect 2777 103 2805 137
rect 2849 103 2873 137
rect 2921 103 2941 137
rect 2993 103 3009 137
rect 3065 103 3077 137
rect 3137 103 3145 137
rect 3209 103 3213 137
rect 3315 103 3319 137
rect 3383 103 3391 137
rect 3451 103 3463 137
rect 3519 103 3535 137
rect 3587 103 3607 137
rect 3655 103 3679 137
rect 3723 103 3751 137
rect 3791 103 3823 137
rect 3859 103 3893 137
rect 3929 103 3961 137
rect 4001 103 4040 137
rect 40 80 4040 103
rect 4320 155 4400 189
rect 4320 121 4343 155
rect 4377 121 4400 155
rect 4320 87 4400 121
rect -320 19 -240 53
rect -320 -15 -297 19
rect -263 -15 -240 19
rect 4320 53 4343 87
rect 4377 53 4400 87
rect 4320 19 4400 53
rect -320 -49 -240 -15
rect -320 -83 -297 -49
rect -263 -83 -240 -49
rect -160 -23 -80 4
rect -160 -57 -137 -23
rect -103 -57 -80 -23
rect -160 -80 -80 -57
rect 4160 -23 4240 4
rect 4160 -57 4183 -23
rect 4217 -57 4240 -23
rect 4160 -80 4240 -57
rect 4320 -15 4343 19
rect 4377 -15 4400 19
rect 4320 -49 4400 -15
rect -320 -117 -240 -83
rect -320 -151 -297 -117
rect -263 -151 -240 -117
rect -320 -185 -240 -151
rect 4320 -83 4343 -49
rect 4377 -83 4400 -49
rect 4320 -117 4400 -83
rect 4320 -151 4343 -117
rect 4377 -151 4400 -117
rect -320 -219 -297 -185
rect -263 -219 -240 -185
rect -320 -253 -240 -219
rect 40 -183 4040 -160
rect 40 -217 79 -183
rect 119 -217 151 -183
rect 187 -217 221 -183
rect 257 -217 289 -183
rect 329 -217 357 -183
rect 401 -217 425 -183
rect 473 -217 493 -183
rect 545 -217 561 -183
rect 617 -217 629 -183
rect 689 -217 697 -183
rect 761 -217 765 -183
rect 867 -217 871 -183
rect 935 -217 943 -183
rect 1003 -217 1015 -183
rect 1071 -217 1087 -183
rect 1139 -217 1159 -183
rect 1207 -217 1231 -183
rect 1275 -217 1303 -183
rect 1343 -217 1375 -183
rect 1411 -217 1445 -183
rect 1481 -217 1513 -183
rect 1553 -217 1581 -183
rect 1625 -217 1649 -183
rect 1697 -217 1717 -183
rect 1769 -217 1785 -183
rect 1841 -217 1853 -183
rect 1913 -217 1921 -183
rect 1985 -217 1989 -183
rect 2091 -217 2095 -183
rect 2159 -217 2167 -183
rect 2227 -217 2239 -183
rect 2295 -217 2311 -183
rect 2363 -217 2383 -183
rect 2431 -217 2455 -183
rect 2499 -217 2527 -183
rect 2567 -217 2599 -183
rect 2635 -217 2669 -183
rect 2705 -217 2737 -183
rect 2777 -217 2805 -183
rect 2849 -217 2873 -183
rect 2921 -217 2941 -183
rect 2993 -217 3009 -183
rect 3065 -217 3077 -183
rect 3137 -217 3145 -183
rect 3209 -217 3213 -183
rect 3315 -217 3319 -183
rect 3383 -217 3391 -183
rect 3451 -217 3463 -183
rect 3519 -217 3535 -183
rect 3587 -217 3607 -183
rect 3655 -217 3679 -183
rect 3723 -217 3751 -183
rect 3791 -217 3823 -183
rect 3859 -217 3893 -183
rect 3929 -217 3961 -183
rect 4001 -217 4040 -183
rect 40 -240 4040 -217
rect 4320 -185 4400 -151
rect 4320 -219 4343 -185
rect 4377 -219 4400 -185
rect -320 -287 -297 -253
rect -263 -287 -240 -253
rect -320 -321 -240 -287
rect 4320 -253 4400 -219
rect 4320 -287 4343 -253
rect 4377 -287 4400 -253
rect -320 -355 -297 -321
rect -263 -355 -240 -321
rect -320 -389 -240 -355
rect -320 -423 -297 -389
rect -263 -423 -240 -389
rect -160 -343 -80 -316
rect -160 -377 -137 -343
rect -103 -377 -80 -343
rect -160 -400 -80 -377
rect 4160 -343 4240 -316
rect 4160 -377 4183 -343
rect 4217 -377 4240 -343
rect 4160 -400 4240 -377
rect 4320 -321 4400 -287
rect 4320 -355 4343 -321
rect 4377 -355 4400 -321
rect 4320 -389 4400 -355
rect -320 -480 -240 -423
rect 4320 -423 4343 -389
rect 4377 -423 4400 -389
rect 4320 -480 4400 -423
rect -320 -503 4400 -480
rect -320 -537 -297 -503
rect -263 -537 -187 -503
rect -153 -537 -119 -503
rect -85 -537 -51 -503
rect -17 -537 17 -503
rect 51 -537 85 -503
rect 119 -537 153 -503
rect 187 -537 221 -503
rect 255 -537 289 -503
rect 323 -537 357 -503
rect 391 -537 425 -503
rect 459 -537 493 -503
rect 527 -537 561 -503
rect 595 -537 629 -503
rect 663 -537 697 -503
rect 731 -537 765 -503
rect 799 -537 833 -503
rect 867 -537 901 -503
rect 935 -537 969 -503
rect 1003 -537 1037 -503
rect 1071 -537 1105 -503
rect 1139 -537 1173 -503
rect 1207 -537 1241 -503
rect 1275 -537 1309 -503
rect 1343 -537 1377 -503
rect 1411 -537 1445 -503
rect 1479 -537 1513 -503
rect 1547 -537 1581 -503
rect 1615 -537 1649 -503
rect 1683 -537 1717 -503
rect 1751 -537 1785 -503
rect 1819 -537 1853 -503
rect 1887 -537 1921 -503
rect 1955 -537 1989 -503
rect 2023 -537 2057 -503
rect 2091 -537 2125 -503
rect 2159 -537 2193 -503
rect 2227 -537 2261 -503
rect 2295 -537 2329 -503
rect 2363 -537 2397 -503
rect 2431 -537 2465 -503
rect 2499 -537 2533 -503
rect 2567 -537 2601 -503
rect 2635 -537 2669 -503
rect 2703 -537 2737 -503
rect 2771 -537 2805 -503
rect 2839 -537 2873 -503
rect 2907 -537 2941 -503
rect 2975 -537 3009 -503
rect 3043 -537 3077 -503
rect 3111 -537 3145 -503
rect 3179 -537 3213 -503
rect 3247 -537 3281 -503
rect 3315 -537 3349 -503
rect 3383 -537 3417 -503
rect 3451 -537 3485 -503
rect 3519 -537 3553 -503
rect 3587 -537 3621 -503
rect 3655 -537 3689 -503
rect 3723 -537 3757 -503
rect 3791 -537 3825 -503
rect 3859 -537 3893 -503
rect 3927 -537 3961 -503
rect 3995 -537 4029 -503
rect 4063 -537 4097 -503
rect 4131 -537 4165 -503
rect 4199 -537 4233 -503
rect 4267 -537 4400 -503
rect -320 -560 4400 -537
rect 4480 319 4560 400
rect 4480 285 4503 319
rect 4537 285 4560 319
rect 4480 251 4560 285
rect 4480 217 4503 251
rect 4537 217 4560 251
rect 4480 183 4560 217
rect 4480 149 4503 183
rect 4537 149 4560 183
rect 4480 115 4560 149
rect 4480 81 4503 115
rect 4537 81 4560 115
rect 4480 47 4560 81
rect 4480 13 4503 47
rect 4537 13 4560 47
rect 4480 -21 4560 13
rect 4480 -55 4503 -21
rect 4537 -55 4560 -21
rect 4480 -89 4560 -55
rect 4480 -123 4503 -89
rect 4537 -123 4560 -89
rect 4480 -157 4560 -123
rect 4480 -191 4503 -157
rect 4537 -191 4560 -157
rect 4480 -225 4560 -191
rect 4480 -259 4503 -225
rect 4537 -259 4560 -225
rect 4480 -293 4560 -259
rect 4480 -327 4503 -293
rect 4537 -327 4560 -293
rect 4480 -361 4560 -327
rect 4480 -395 4503 -361
rect 4537 -395 4560 -361
rect 4480 -429 4560 -395
rect 4480 -463 4503 -429
rect 4537 -463 4560 -429
rect 4480 -497 4560 -463
rect 4480 -531 4503 -497
rect 4537 -531 4560 -497
rect -480 -599 -457 -565
rect -423 -599 -400 -565
rect -480 -640 -400 -599
rect 4480 -565 4560 -531
rect 4480 -599 4503 -565
rect 4537 -599 4560 -565
rect 4480 -640 4560 -599
rect 8000 4199 8080 4240
rect 8000 4165 8023 4199
rect 8057 4165 8080 4199
rect 8000 4131 8080 4165
rect 12960 4199 13040 4240
rect 12960 4165 12983 4199
rect 13017 4165 13040 4199
rect 8000 4097 8023 4131
rect 8057 4097 8080 4131
rect 8000 4063 8080 4097
rect 8000 4029 8023 4063
rect 8057 4029 8080 4063
rect 8000 3995 8080 4029
rect 8000 3961 8023 3995
rect 8057 3961 8080 3995
rect 8000 3927 8080 3961
rect 8000 3893 8023 3927
rect 8057 3893 8080 3927
rect 8000 3859 8080 3893
rect 8000 3825 8023 3859
rect 8057 3825 8080 3859
rect 8000 3791 8080 3825
rect 8000 3757 8023 3791
rect 8057 3757 8080 3791
rect 8000 3723 8080 3757
rect 8000 3689 8023 3723
rect 8057 3689 8080 3723
rect 8000 3655 8080 3689
rect 8000 3621 8023 3655
rect 8057 3621 8080 3655
rect 8000 3587 8080 3621
rect 8000 3553 8023 3587
rect 8057 3553 8080 3587
rect 8000 3519 8080 3553
rect 8000 3485 8023 3519
rect 8057 3485 8080 3519
rect 8000 3451 8080 3485
rect 8000 3417 8023 3451
rect 8057 3417 8080 3451
rect 8000 3383 8080 3417
rect 8000 3349 8023 3383
rect 8057 3349 8080 3383
rect 8000 3315 8080 3349
rect 8000 3281 8023 3315
rect 8057 3281 8080 3315
rect 8000 3200 8080 3281
rect 8160 4137 12880 4160
rect 8160 4103 8293 4137
rect 8327 4103 8361 4137
rect 8395 4103 8429 4137
rect 8463 4103 8497 4137
rect 8531 4103 8565 4137
rect 8599 4103 8633 4137
rect 8667 4103 8701 4137
rect 8735 4103 8769 4137
rect 8803 4103 8837 4137
rect 8871 4103 8905 4137
rect 8939 4103 8973 4137
rect 9007 4103 9041 4137
rect 9075 4103 9109 4137
rect 9143 4103 9177 4137
rect 9211 4103 9245 4137
rect 9279 4103 9313 4137
rect 9347 4103 9381 4137
rect 9415 4103 9449 4137
rect 9483 4103 9517 4137
rect 9551 4103 9585 4137
rect 9619 4103 9653 4137
rect 9687 4103 9721 4137
rect 9755 4103 9789 4137
rect 9823 4103 9857 4137
rect 9891 4103 9925 4137
rect 9959 4103 9993 4137
rect 10027 4103 10061 4137
rect 10095 4103 10129 4137
rect 10163 4103 10197 4137
rect 10231 4103 10265 4137
rect 10299 4103 10333 4137
rect 10367 4103 10401 4137
rect 10435 4103 10469 4137
rect 10503 4103 10537 4137
rect 10571 4103 10605 4137
rect 10639 4103 10673 4137
rect 10707 4103 10741 4137
rect 10775 4103 10809 4137
rect 10843 4103 10877 4137
rect 10911 4103 10945 4137
rect 10979 4103 11013 4137
rect 11047 4103 11081 4137
rect 11115 4103 11149 4137
rect 11183 4103 11217 4137
rect 11251 4103 11285 4137
rect 11319 4103 11353 4137
rect 11387 4103 11421 4137
rect 11455 4103 11489 4137
rect 11523 4103 11557 4137
rect 11591 4103 11625 4137
rect 11659 4103 11693 4137
rect 11727 4103 11761 4137
rect 11795 4103 11829 4137
rect 11863 4103 11897 4137
rect 11931 4103 11965 4137
rect 11999 4103 12033 4137
rect 12067 4103 12101 4137
rect 12135 4103 12169 4137
rect 12203 4103 12237 4137
rect 12271 4103 12305 4137
rect 12339 4103 12373 4137
rect 12407 4103 12441 4137
rect 12475 4103 12509 4137
rect 12543 4103 12577 4137
rect 12611 4103 12645 4137
rect 12679 4103 12713 4137
rect 12747 4103 12823 4137
rect 12857 4103 12880 4137
rect 8160 4080 12880 4103
rect 8160 4023 8240 4080
rect 8160 3989 8183 4023
rect 8217 3989 8240 4023
rect 12800 4023 12880 4080
rect 8160 3955 8240 3989
rect 8160 3921 8183 3955
rect 8217 3921 8240 3955
rect 8160 3887 8240 3921
rect 8320 3977 8400 4000
rect 8320 3943 8343 3977
rect 8377 3943 8400 3977
rect 8320 3916 8400 3943
rect 12640 3977 12720 4000
rect 12640 3943 12663 3977
rect 12697 3943 12720 3977
rect 12640 3916 12720 3943
rect 12800 3989 12823 4023
rect 12857 3989 12880 4023
rect 12800 3955 12880 3989
rect 12800 3921 12823 3955
rect 12857 3921 12880 3955
rect 8160 3853 8183 3887
rect 8217 3853 8240 3887
rect 8160 3819 8240 3853
rect 12800 3887 12880 3921
rect 12800 3853 12823 3887
rect 12857 3853 12880 3887
rect 8160 3785 8183 3819
rect 8217 3785 8240 3819
rect 8160 3751 8240 3785
rect 8520 3817 12520 3840
rect 8520 3783 8559 3817
rect 8599 3783 8631 3817
rect 8667 3783 8701 3817
rect 8737 3783 8769 3817
rect 8809 3783 8837 3817
rect 8881 3783 8905 3817
rect 8953 3783 8973 3817
rect 9025 3783 9041 3817
rect 9097 3783 9109 3817
rect 9169 3783 9177 3817
rect 9241 3783 9245 3817
rect 9347 3783 9351 3817
rect 9415 3783 9423 3817
rect 9483 3783 9495 3817
rect 9551 3783 9567 3817
rect 9619 3783 9639 3817
rect 9687 3783 9711 3817
rect 9755 3783 9783 3817
rect 9823 3783 9855 3817
rect 9891 3783 9925 3817
rect 9961 3783 9993 3817
rect 10033 3783 10061 3817
rect 10105 3783 10129 3817
rect 10177 3783 10197 3817
rect 10249 3783 10265 3817
rect 10321 3783 10333 3817
rect 10393 3783 10401 3817
rect 10465 3783 10469 3817
rect 10571 3783 10575 3817
rect 10639 3783 10647 3817
rect 10707 3783 10719 3817
rect 10775 3783 10791 3817
rect 10843 3783 10863 3817
rect 10911 3783 10935 3817
rect 10979 3783 11007 3817
rect 11047 3783 11079 3817
rect 11115 3783 11149 3817
rect 11185 3783 11217 3817
rect 11257 3783 11285 3817
rect 11329 3783 11353 3817
rect 11401 3783 11421 3817
rect 11473 3783 11489 3817
rect 11545 3783 11557 3817
rect 11617 3783 11625 3817
rect 11689 3783 11693 3817
rect 11795 3783 11799 3817
rect 11863 3783 11871 3817
rect 11931 3783 11943 3817
rect 11999 3783 12015 3817
rect 12067 3783 12087 3817
rect 12135 3783 12159 3817
rect 12203 3783 12231 3817
rect 12271 3783 12303 3817
rect 12339 3783 12373 3817
rect 12409 3783 12441 3817
rect 12481 3783 12520 3817
rect 8520 3760 12520 3783
rect 12800 3819 12880 3853
rect 12800 3785 12823 3819
rect 12857 3785 12880 3819
rect 8160 3717 8183 3751
rect 8217 3717 8240 3751
rect 8160 3683 8240 3717
rect 8160 3649 8183 3683
rect 8217 3649 8240 3683
rect 12800 3751 12880 3785
rect 12800 3717 12823 3751
rect 12857 3717 12880 3751
rect 12800 3683 12880 3717
rect 8160 3615 8240 3649
rect 8160 3581 8183 3615
rect 8217 3581 8240 3615
rect 8320 3657 8400 3680
rect 8320 3623 8343 3657
rect 8377 3623 8400 3657
rect 8320 3596 8400 3623
rect 12640 3657 12720 3680
rect 12640 3623 12663 3657
rect 12697 3623 12720 3657
rect 12640 3596 12720 3623
rect 12800 3649 12823 3683
rect 12857 3649 12880 3683
rect 12800 3615 12880 3649
rect 8160 3547 8240 3581
rect 8160 3513 8183 3547
rect 8217 3513 8240 3547
rect 12800 3581 12823 3615
rect 12857 3581 12880 3615
rect 12800 3547 12880 3581
rect 8160 3479 8240 3513
rect 8160 3445 8183 3479
rect 8217 3445 8240 3479
rect 8160 3411 8240 3445
rect 8520 3497 12520 3520
rect 8520 3463 8559 3497
rect 8599 3463 8631 3497
rect 8667 3463 8701 3497
rect 8737 3463 8769 3497
rect 8809 3463 8837 3497
rect 8881 3463 8905 3497
rect 8953 3463 8973 3497
rect 9025 3463 9041 3497
rect 9097 3463 9109 3497
rect 9169 3463 9177 3497
rect 9241 3463 9245 3497
rect 9347 3463 9351 3497
rect 9415 3463 9423 3497
rect 9483 3463 9495 3497
rect 9551 3463 9567 3497
rect 9619 3463 9639 3497
rect 9687 3463 9711 3497
rect 9755 3463 9783 3497
rect 9823 3463 9855 3497
rect 9891 3463 9925 3497
rect 9961 3463 9993 3497
rect 10033 3463 10061 3497
rect 10105 3463 10129 3497
rect 10177 3463 10197 3497
rect 10249 3463 10265 3497
rect 10321 3463 10333 3497
rect 10393 3463 10401 3497
rect 10465 3463 10469 3497
rect 10571 3463 10575 3497
rect 10639 3463 10647 3497
rect 10707 3463 10719 3497
rect 10775 3463 10791 3497
rect 10843 3463 10863 3497
rect 10911 3463 10935 3497
rect 10979 3463 11007 3497
rect 11047 3463 11079 3497
rect 11115 3463 11149 3497
rect 11185 3463 11217 3497
rect 11257 3463 11285 3497
rect 11329 3463 11353 3497
rect 11401 3463 11421 3497
rect 11473 3463 11489 3497
rect 11545 3463 11557 3497
rect 11617 3463 11625 3497
rect 11689 3463 11693 3497
rect 11795 3463 11799 3497
rect 11863 3463 11871 3497
rect 11931 3463 11943 3497
rect 11999 3463 12015 3497
rect 12067 3463 12087 3497
rect 12135 3463 12159 3497
rect 12203 3463 12231 3497
rect 12271 3463 12303 3497
rect 12339 3463 12373 3497
rect 12409 3463 12441 3497
rect 12481 3463 12520 3497
rect 8520 3440 12520 3463
rect 12800 3513 12823 3547
rect 12857 3513 12880 3547
rect 12800 3479 12880 3513
rect 12800 3445 12823 3479
rect 12857 3445 12880 3479
rect 8160 3377 8183 3411
rect 8217 3377 8240 3411
rect 8160 3360 8240 3377
rect 12800 3411 12880 3445
rect 12800 3377 12823 3411
rect 12857 3377 12880 3411
rect 12800 3360 12880 3377
rect 8160 3337 12880 3360
rect 8160 3303 8293 3337
rect 8327 3303 8361 3337
rect 8395 3303 8429 3337
rect 8463 3303 8497 3337
rect 8531 3303 8565 3337
rect 8599 3303 8633 3337
rect 8667 3303 8701 3337
rect 8735 3303 8769 3337
rect 8803 3303 8837 3337
rect 8871 3303 8905 3337
rect 8939 3303 8973 3337
rect 9007 3303 9041 3337
rect 9075 3303 9109 3337
rect 9143 3303 9177 3337
rect 9211 3303 9245 3337
rect 9279 3303 9313 3337
rect 9347 3303 9381 3337
rect 9415 3303 9449 3337
rect 9483 3303 9517 3337
rect 9551 3303 9585 3337
rect 9619 3303 9653 3337
rect 9687 3303 9721 3337
rect 9755 3303 9789 3337
rect 9823 3303 9857 3337
rect 9891 3303 9925 3337
rect 9959 3303 9993 3337
rect 10027 3303 10061 3337
rect 10095 3303 10129 3337
rect 10163 3303 10197 3337
rect 10231 3303 10265 3337
rect 10299 3303 10333 3337
rect 10367 3303 10401 3337
rect 10435 3303 10469 3337
rect 10503 3303 10537 3337
rect 10571 3303 10605 3337
rect 10639 3303 10673 3337
rect 10707 3303 10741 3337
rect 10775 3303 10809 3337
rect 10843 3303 10877 3337
rect 10911 3303 10945 3337
rect 10979 3303 11013 3337
rect 11047 3303 11081 3337
rect 11115 3303 11149 3337
rect 11183 3303 11217 3337
rect 11251 3303 11285 3337
rect 11319 3303 11353 3337
rect 11387 3303 11421 3337
rect 11455 3303 11489 3337
rect 11523 3303 11557 3337
rect 11591 3303 11625 3337
rect 11659 3303 11693 3337
rect 11727 3303 11761 3337
rect 11795 3303 11829 3337
rect 11863 3303 11897 3337
rect 11931 3303 11965 3337
rect 11999 3303 12033 3337
rect 12067 3303 12101 3337
rect 12135 3303 12169 3337
rect 12203 3303 12237 3337
rect 12271 3303 12305 3337
rect 12339 3303 12373 3337
rect 12407 3303 12441 3337
rect 12475 3303 12509 3337
rect 12543 3303 12577 3337
rect 12611 3303 12645 3337
rect 12679 3303 12713 3337
rect 12747 3303 12880 3337
rect 8160 3280 12880 3303
rect 12960 4131 13040 4165
rect 12960 4097 12983 4131
rect 13017 4097 13040 4131
rect 12960 4063 13040 4097
rect 12960 4029 12983 4063
rect 13017 4029 13040 4063
rect 12960 3995 13040 4029
rect 12960 3961 12983 3995
rect 13017 3961 13040 3995
rect 12960 3927 13040 3961
rect 12960 3893 12983 3927
rect 13017 3893 13040 3927
rect 12960 3859 13040 3893
rect 12960 3825 12983 3859
rect 13017 3825 13040 3859
rect 12960 3791 13040 3825
rect 12960 3757 12983 3791
rect 13017 3757 13040 3791
rect 12960 3723 13040 3757
rect 12960 3689 12983 3723
rect 13017 3689 13040 3723
rect 12960 3655 13040 3689
rect 12960 3621 12983 3655
rect 13017 3621 13040 3655
rect 12960 3587 13040 3621
rect 12960 3553 12983 3587
rect 13017 3553 13040 3587
rect 12960 3519 13040 3553
rect 12960 3485 12983 3519
rect 13017 3485 13040 3519
rect 12960 3451 13040 3485
rect 12960 3417 12983 3451
rect 13017 3417 13040 3451
rect 12960 3383 13040 3417
rect 12960 3349 12983 3383
rect 13017 3349 13040 3383
rect 12960 3315 13040 3349
rect 12960 3281 12983 3315
rect 13017 3281 13040 3315
rect 12960 3200 13040 3281
rect 8000 3177 13040 3200
rect 8000 3143 8123 3177
rect 8157 3143 8191 3177
rect 8225 3143 8259 3177
rect 8293 3143 8327 3177
rect 8361 3143 8395 3177
rect 8429 3143 8463 3177
rect 8497 3143 8531 3177
rect 8565 3143 8599 3177
rect 8633 3143 8667 3177
rect 8701 3143 8735 3177
rect 8769 3143 8803 3177
rect 8837 3143 8871 3177
rect 8905 3143 8939 3177
rect 8973 3143 9007 3177
rect 9041 3143 9075 3177
rect 9109 3143 9143 3177
rect 9177 3143 9211 3177
rect 9245 3143 9279 3177
rect 9313 3143 9347 3177
rect 9381 3143 9415 3177
rect 9449 3143 9483 3177
rect 9517 3143 9551 3177
rect 9585 3143 9619 3177
rect 9653 3143 9687 3177
rect 9721 3143 9755 3177
rect 9789 3143 9823 3177
rect 9857 3143 9891 3177
rect 9925 3143 9959 3177
rect 9993 3143 10027 3177
rect 10061 3143 10095 3177
rect 10129 3143 10163 3177
rect 10197 3143 10231 3177
rect 10265 3143 10299 3177
rect 10333 3143 10367 3177
rect 10401 3143 10435 3177
rect 10469 3143 10503 3177
rect 10537 3143 10571 3177
rect 10605 3143 10639 3177
rect 10673 3143 10707 3177
rect 10741 3143 10775 3177
rect 10809 3143 10843 3177
rect 10877 3143 10911 3177
rect 10945 3143 10979 3177
rect 11013 3143 11047 3177
rect 11081 3143 11115 3177
rect 11149 3143 11183 3177
rect 11217 3143 11251 3177
rect 11285 3143 11319 3177
rect 11353 3143 11387 3177
rect 11421 3143 11455 3177
rect 11489 3143 11523 3177
rect 11557 3143 11591 3177
rect 11625 3143 11659 3177
rect 11693 3143 11727 3177
rect 11761 3143 11795 3177
rect 11829 3143 11863 3177
rect 11897 3143 11931 3177
rect 11965 3143 11999 3177
rect 12033 3143 12067 3177
rect 12101 3143 12135 3177
rect 12169 3143 12203 3177
rect 12237 3143 12271 3177
rect 12305 3143 12339 3177
rect 12373 3143 12407 3177
rect 12441 3143 12475 3177
rect 12509 3143 12543 3177
rect 12577 3143 12611 3177
rect 12645 3143 12679 3177
rect 12713 3143 12747 3177
rect 12781 3143 12815 3177
rect 12849 3143 12883 3177
rect 12917 3143 13040 3177
rect 8000 3120 13040 3143
rect 8000 3040 8080 3120
rect 12960 3040 13040 3120
rect 8000 3017 13040 3040
rect 8000 2983 8123 3017
rect 8157 2983 8191 3017
rect 8225 2983 8259 3017
rect 8293 2983 8327 3017
rect 8361 2983 8395 3017
rect 8429 2983 8463 3017
rect 8497 2983 8531 3017
rect 8565 2983 8599 3017
rect 8633 2983 8667 3017
rect 8701 2983 8735 3017
rect 8769 2983 8803 3017
rect 8837 2983 8871 3017
rect 8905 2983 8939 3017
rect 8973 2983 9007 3017
rect 9041 2983 9075 3017
rect 9109 2983 9143 3017
rect 9177 2983 9211 3017
rect 9245 2983 9279 3017
rect 9313 2983 9347 3017
rect 9381 2983 9415 3017
rect 9449 2983 9483 3017
rect 9517 2983 9551 3017
rect 9585 2983 9619 3017
rect 9653 2983 9687 3017
rect 9721 2983 9755 3017
rect 9789 2983 9823 3017
rect 9857 2983 9891 3017
rect 9925 2983 9959 3017
rect 9993 2983 10027 3017
rect 10061 2983 10095 3017
rect 10129 2983 10163 3017
rect 10197 2983 10231 3017
rect 10265 2983 10299 3017
rect 10333 2983 10367 3017
rect 10401 2983 10435 3017
rect 10469 2983 10503 3017
rect 10537 2983 10571 3017
rect 10605 2983 10639 3017
rect 10673 2983 10707 3017
rect 10741 2983 10775 3017
rect 10809 2983 10843 3017
rect 10877 2983 10911 3017
rect 10945 2983 10979 3017
rect 11013 2983 11047 3017
rect 11081 2983 11115 3017
rect 11149 2983 11183 3017
rect 11217 2983 11251 3017
rect 11285 2983 11319 3017
rect 11353 2983 11387 3017
rect 11421 2983 11455 3017
rect 11489 2983 11523 3017
rect 11557 2983 11591 3017
rect 11625 2983 11659 3017
rect 11693 2983 11727 3017
rect 11761 2983 11795 3017
rect 11829 2983 11863 3017
rect 11897 2983 11931 3017
rect 11965 2983 11999 3017
rect 12033 2983 12067 3017
rect 12101 2983 12135 3017
rect 12169 2983 12203 3017
rect 12237 2983 12271 3017
rect 12305 2983 12339 3017
rect 12373 2983 12407 3017
rect 12441 2983 12475 3017
rect 12509 2983 12543 3017
rect 12577 2983 12611 3017
rect 12645 2983 12679 3017
rect 12713 2983 12747 3017
rect 12781 2983 12815 3017
rect 12849 2983 12883 3017
rect 12917 2983 13040 3017
rect 8000 2960 13040 2983
rect 8000 2879 8080 2960
rect 8000 2845 8023 2879
rect 8057 2845 8080 2879
rect 8000 2811 8080 2845
rect 8000 2777 8023 2811
rect 8057 2777 8080 2811
rect 8000 2743 8080 2777
rect 8000 2709 8023 2743
rect 8057 2709 8080 2743
rect 8000 2675 8080 2709
rect 8000 2641 8023 2675
rect 8057 2641 8080 2675
rect 8000 2607 8080 2641
rect 8000 2573 8023 2607
rect 8057 2573 8080 2607
rect 8000 2539 8080 2573
rect 8000 2505 8023 2539
rect 8057 2505 8080 2539
rect 8000 2471 8080 2505
rect 8000 2437 8023 2471
rect 8057 2437 8080 2471
rect 8000 2403 8080 2437
rect 8000 2369 8023 2403
rect 8057 2369 8080 2403
rect 8000 2335 8080 2369
rect 8000 2301 8023 2335
rect 8057 2301 8080 2335
rect 8000 2267 8080 2301
rect 8000 2233 8023 2267
rect 8057 2233 8080 2267
rect 8000 2199 8080 2233
rect 8000 2165 8023 2199
rect 8057 2165 8080 2199
rect 8000 2131 8080 2165
rect 8000 2097 8023 2131
rect 8057 2097 8080 2131
rect 8000 2063 8080 2097
rect 8000 2029 8023 2063
rect 8057 2029 8080 2063
rect 8000 1995 8080 2029
rect 8160 2857 12880 2880
rect 8160 2823 8293 2857
rect 8327 2823 8343 2857
rect 8395 2823 8429 2857
rect 8463 2823 8497 2857
rect 8531 2823 8565 2857
rect 8599 2823 8633 2857
rect 8667 2823 8701 2857
rect 8735 2823 8769 2857
rect 8803 2823 8837 2857
rect 8871 2823 8905 2857
rect 8939 2823 8973 2857
rect 9007 2823 9041 2857
rect 9075 2823 9109 2857
rect 9143 2823 9177 2857
rect 9211 2823 9245 2857
rect 9279 2823 9313 2857
rect 9347 2823 9381 2857
rect 9415 2823 9449 2857
rect 9483 2823 9517 2857
rect 9551 2823 9585 2857
rect 9619 2823 9653 2857
rect 9687 2823 9721 2857
rect 9755 2823 9789 2857
rect 9823 2823 9857 2857
rect 9891 2823 9925 2857
rect 9959 2823 9993 2857
rect 10027 2823 10061 2857
rect 10095 2823 10129 2857
rect 10163 2823 10197 2857
rect 10231 2823 10265 2857
rect 10299 2823 10333 2857
rect 10367 2823 10401 2857
rect 10435 2823 10469 2857
rect 10503 2823 10537 2857
rect 10571 2823 10605 2857
rect 10639 2823 10673 2857
rect 10707 2823 10741 2857
rect 10775 2823 10809 2857
rect 10843 2823 10877 2857
rect 10911 2823 10945 2857
rect 10979 2823 11013 2857
rect 11047 2823 11081 2857
rect 11115 2823 11149 2857
rect 11183 2823 11217 2857
rect 11251 2823 11285 2857
rect 11319 2823 11353 2857
rect 11387 2823 11421 2857
rect 11455 2823 11489 2857
rect 11523 2823 11557 2857
rect 11591 2823 11625 2857
rect 11659 2823 11693 2857
rect 11727 2823 11761 2857
rect 11795 2823 11829 2857
rect 11863 2823 11897 2857
rect 11931 2823 11965 2857
rect 11999 2823 12033 2857
rect 12067 2823 12101 2857
rect 12135 2823 12169 2857
rect 12203 2823 12237 2857
rect 12271 2823 12305 2857
rect 12339 2823 12373 2857
rect 12407 2823 12441 2857
rect 12475 2823 12509 2857
rect 12543 2823 12577 2857
rect 12611 2823 12645 2857
rect 12679 2823 12713 2857
rect 12747 2823 12880 2857
rect 8160 2800 12880 2823
rect 8160 2783 8240 2800
rect 8160 2749 8183 2783
rect 8217 2749 8240 2783
rect 8160 2715 8240 2749
rect 12800 2783 12880 2800
rect 12800 2749 12823 2783
rect 12857 2749 12880 2783
rect 8160 2681 8183 2715
rect 8217 2681 8240 2715
rect 8160 2647 8240 2681
rect 8160 2613 8183 2647
rect 8217 2613 8240 2647
rect 8520 2697 12520 2720
rect 8520 2663 8559 2697
rect 8599 2663 8631 2697
rect 8667 2663 8701 2697
rect 8737 2663 8769 2697
rect 8809 2663 8837 2697
rect 8881 2663 8905 2697
rect 8953 2663 8973 2697
rect 9025 2663 9041 2697
rect 9097 2663 9109 2697
rect 9169 2663 9177 2697
rect 9241 2663 9245 2697
rect 9347 2663 9351 2697
rect 9415 2663 9423 2697
rect 9483 2663 9495 2697
rect 9551 2663 9567 2697
rect 9619 2663 9639 2697
rect 9687 2663 9711 2697
rect 9755 2663 9783 2697
rect 9823 2663 9855 2697
rect 9891 2663 9925 2697
rect 9961 2663 9993 2697
rect 10033 2663 10061 2697
rect 10105 2663 10129 2697
rect 10177 2663 10197 2697
rect 10249 2663 10265 2697
rect 10321 2663 10333 2697
rect 10393 2663 10401 2697
rect 10465 2663 10469 2697
rect 10571 2663 10575 2697
rect 10639 2663 10647 2697
rect 10707 2663 10719 2697
rect 10775 2663 10791 2697
rect 10843 2663 10863 2697
rect 10911 2663 10935 2697
rect 10979 2663 11007 2697
rect 11047 2663 11079 2697
rect 11115 2663 11149 2697
rect 11185 2663 11217 2697
rect 11257 2663 11285 2697
rect 11329 2663 11353 2697
rect 11401 2663 11421 2697
rect 11473 2663 11489 2697
rect 11545 2663 11557 2697
rect 11617 2663 11625 2697
rect 11689 2663 11693 2697
rect 11795 2663 11799 2697
rect 11863 2663 11871 2697
rect 11931 2663 11943 2697
rect 11999 2663 12015 2697
rect 12067 2663 12087 2697
rect 12135 2663 12159 2697
rect 12203 2663 12231 2697
rect 12271 2663 12303 2697
rect 12339 2663 12373 2697
rect 12409 2663 12441 2697
rect 12481 2663 12520 2697
rect 8520 2640 12520 2663
rect 12800 2715 12880 2749
rect 12800 2681 12823 2715
rect 12857 2681 12880 2715
rect 12800 2647 12880 2681
rect 8160 2579 8240 2613
rect 8160 2545 8183 2579
rect 8217 2545 8240 2579
rect 12800 2613 12823 2647
rect 12857 2613 12880 2647
rect 12800 2579 12880 2613
rect 8160 2511 8240 2545
rect 8160 2477 8183 2511
rect 8217 2477 8240 2511
rect 8320 2537 8400 2564
rect 8320 2503 8343 2537
rect 8377 2503 8400 2537
rect 8320 2480 8400 2503
rect 12640 2537 12720 2564
rect 12640 2503 12663 2537
rect 12697 2503 12720 2537
rect 12640 2480 12720 2503
rect 12800 2545 12823 2579
rect 12857 2545 12880 2579
rect 12800 2511 12880 2545
rect 8160 2443 8240 2477
rect 8160 2409 8183 2443
rect 8217 2409 8240 2443
rect 8160 2375 8240 2409
rect 12800 2477 12823 2511
rect 12857 2477 12880 2511
rect 12800 2443 12880 2477
rect 12800 2409 12823 2443
rect 12857 2409 12880 2443
rect 8160 2341 8183 2375
rect 8217 2341 8240 2375
rect 8160 2307 8240 2341
rect 8520 2377 12520 2400
rect 8520 2343 8559 2377
rect 8599 2343 8631 2377
rect 8667 2343 8701 2377
rect 8737 2343 8769 2377
rect 8809 2343 8837 2377
rect 8881 2343 8905 2377
rect 8953 2343 8973 2377
rect 9025 2343 9041 2377
rect 9097 2343 9109 2377
rect 9169 2343 9177 2377
rect 9241 2343 9245 2377
rect 9347 2343 9351 2377
rect 9415 2343 9423 2377
rect 9483 2343 9495 2377
rect 9551 2343 9567 2377
rect 9619 2343 9639 2377
rect 9687 2343 9711 2377
rect 9755 2343 9783 2377
rect 9823 2343 9855 2377
rect 9891 2343 9925 2377
rect 9961 2343 9993 2377
rect 10033 2343 10061 2377
rect 10105 2343 10129 2377
rect 10177 2343 10197 2377
rect 10249 2343 10265 2377
rect 10321 2343 10333 2377
rect 10393 2343 10401 2377
rect 10465 2343 10469 2377
rect 10571 2343 10575 2377
rect 10639 2343 10647 2377
rect 10707 2343 10719 2377
rect 10775 2343 10791 2377
rect 10843 2343 10863 2377
rect 10911 2343 10935 2377
rect 10979 2343 11007 2377
rect 11047 2343 11079 2377
rect 11115 2343 11149 2377
rect 11185 2343 11217 2377
rect 11257 2343 11285 2377
rect 11329 2343 11353 2377
rect 11401 2343 11421 2377
rect 11473 2343 11489 2377
rect 11545 2343 11557 2377
rect 11617 2343 11625 2377
rect 11689 2343 11693 2377
rect 11795 2343 11799 2377
rect 11863 2343 11871 2377
rect 11931 2343 11943 2377
rect 11999 2343 12015 2377
rect 12067 2343 12087 2377
rect 12135 2343 12159 2377
rect 12203 2343 12231 2377
rect 12271 2343 12303 2377
rect 12339 2343 12373 2377
rect 12409 2343 12441 2377
rect 12481 2343 12520 2377
rect 8520 2320 12520 2343
rect 12800 2375 12880 2409
rect 12800 2341 12823 2375
rect 12857 2341 12880 2375
rect 8160 2273 8183 2307
rect 8217 2273 8240 2307
rect 8160 2239 8240 2273
rect 12800 2307 12880 2341
rect 12800 2273 12823 2307
rect 12857 2273 12880 2307
rect 8160 2205 8183 2239
rect 8217 2205 8240 2239
rect 8160 2171 8240 2205
rect 8160 2137 8183 2171
rect 8217 2137 8240 2171
rect 8320 2217 8400 2244
rect 8320 2183 8343 2217
rect 8377 2183 8400 2217
rect 8320 2160 8400 2183
rect 12640 2217 12720 2244
rect 12640 2183 12663 2217
rect 12697 2183 12720 2217
rect 12640 2160 12720 2183
rect 12800 2239 12880 2273
rect 12800 2205 12823 2239
rect 12857 2205 12880 2239
rect 12800 2171 12880 2205
rect 8160 2080 8240 2137
rect 12800 2137 12823 2171
rect 12857 2137 12880 2171
rect 12800 2080 12880 2137
rect 8160 2057 12880 2080
rect 8160 2023 8293 2057
rect 8327 2023 8361 2057
rect 8395 2023 8429 2057
rect 8463 2023 8497 2057
rect 8531 2023 8565 2057
rect 8599 2023 8633 2057
rect 8667 2023 8701 2057
rect 8735 2023 8769 2057
rect 8803 2023 8837 2057
rect 8871 2023 8905 2057
rect 8939 2023 8973 2057
rect 9007 2023 9041 2057
rect 9075 2023 9109 2057
rect 9143 2023 9177 2057
rect 9211 2023 9245 2057
rect 9279 2023 9313 2057
rect 9347 2023 9381 2057
rect 9415 2023 9449 2057
rect 9483 2023 9517 2057
rect 9551 2023 9585 2057
rect 9619 2023 9653 2057
rect 9687 2023 9721 2057
rect 9755 2023 9789 2057
rect 9823 2023 9857 2057
rect 9891 2023 9925 2057
rect 9959 2023 9993 2057
rect 10027 2023 10061 2057
rect 10095 2023 10129 2057
rect 10163 2023 10197 2057
rect 10231 2023 10265 2057
rect 10299 2023 10333 2057
rect 10367 2023 10401 2057
rect 10435 2023 10469 2057
rect 10503 2023 10537 2057
rect 10571 2023 10605 2057
rect 10639 2023 10673 2057
rect 10707 2023 10741 2057
rect 10775 2023 10809 2057
rect 10843 2023 10877 2057
rect 10911 2023 10945 2057
rect 10979 2023 11013 2057
rect 11047 2023 11081 2057
rect 11115 2023 11149 2057
rect 11183 2023 11217 2057
rect 11251 2023 11285 2057
rect 11319 2023 11353 2057
rect 11387 2023 11421 2057
rect 11455 2023 11489 2057
rect 11523 2023 11557 2057
rect 11591 2023 11625 2057
rect 11659 2023 11693 2057
rect 11727 2023 11761 2057
rect 11795 2023 11829 2057
rect 11863 2023 11897 2057
rect 11931 2023 11965 2057
rect 11999 2023 12033 2057
rect 12067 2023 12101 2057
rect 12135 2023 12169 2057
rect 12203 2023 12237 2057
rect 12271 2023 12305 2057
rect 12339 2023 12373 2057
rect 12407 2023 12441 2057
rect 12475 2023 12509 2057
rect 12543 2023 12577 2057
rect 12611 2023 12645 2057
rect 12679 2023 12713 2057
rect 12747 2023 12880 2057
rect 8160 2000 12880 2023
rect 12960 2879 13040 2960
rect 12960 2845 12983 2879
rect 13017 2845 13040 2879
rect 12960 2811 13040 2845
rect 12960 2777 12983 2811
rect 13017 2777 13040 2811
rect 12960 2743 13040 2777
rect 12960 2709 12983 2743
rect 13017 2709 13040 2743
rect 12960 2675 13040 2709
rect 12960 2641 12983 2675
rect 13017 2641 13040 2675
rect 12960 2607 13040 2641
rect 12960 2573 12983 2607
rect 13017 2573 13040 2607
rect 12960 2539 13040 2573
rect 12960 2505 12983 2539
rect 13017 2505 13040 2539
rect 12960 2471 13040 2505
rect 12960 2437 12983 2471
rect 13017 2437 13040 2471
rect 12960 2403 13040 2437
rect 12960 2369 12983 2403
rect 13017 2369 13040 2403
rect 12960 2335 13040 2369
rect 12960 2301 12983 2335
rect 13017 2301 13040 2335
rect 12960 2267 13040 2301
rect 12960 2233 12983 2267
rect 13017 2233 13040 2267
rect 12960 2199 13040 2233
rect 12960 2165 12983 2199
rect 13017 2165 13040 2199
rect 12960 2131 13040 2165
rect 12960 2097 12983 2131
rect 13017 2097 13040 2131
rect 12960 2063 13040 2097
rect 12960 2029 12983 2063
rect 13017 2029 13040 2063
rect 8000 1961 8023 1995
rect 8057 1961 8080 1995
rect 8000 1920 8080 1961
rect 12960 1995 13040 2029
rect 12960 1961 12983 1995
rect 13017 1961 13040 1995
rect 12960 1920 13040 1961
rect 8000 1897 13040 1920
rect 8000 1863 8123 1897
rect 8157 1863 8191 1897
rect 8225 1863 8259 1897
rect 8293 1863 8327 1897
rect 8361 1863 8395 1897
rect 8429 1863 8463 1897
rect 8497 1863 8531 1897
rect 8565 1863 8599 1897
rect 8633 1863 8667 1897
rect 8701 1863 8735 1897
rect 8769 1863 8803 1897
rect 8837 1863 8871 1897
rect 8905 1863 8939 1897
rect 8973 1863 9007 1897
rect 9041 1863 9075 1897
rect 9109 1863 9143 1897
rect 9177 1863 9211 1897
rect 9245 1863 9279 1897
rect 9313 1863 9347 1897
rect 9381 1863 9415 1897
rect 9449 1863 9483 1897
rect 9517 1863 9551 1897
rect 9585 1863 9619 1897
rect 9653 1863 9687 1897
rect 9721 1863 9755 1897
rect 9789 1863 9823 1897
rect 9857 1863 9891 1897
rect 9925 1863 9959 1897
rect 9993 1863 10027 1897
rect 10061 1863 10095 1897
rect 10129 1863 10163 1897
rect 10197 1863 10231 1897
rect 10265 1863 10299 1897
rect 10333 1863 10367 1897
rect 10401 1863 10435 1897
rect 10469 1863 10503 1897
rect 10537 1863 10571 1897
rect 10605 1863 10639 1897
rect 10673 1863 10707 1897
rect 10741 1863 10775 1897
rect 10809 1863 10843 1897
rect 10877 1863 10911 1897
rect 10945 1863 10979 1897
rect 11013 1863 11047 1897
rect 11081 1863 11115 1897
rect 11149 1863 11183 1897
rect 11217 1863 11251 1897
rect 11285 1863 11319 1897
rect 11353 1863 11387 1897
rect 11421 1863 11455 1897
rect 11489 1863 11523 1897
rect 11557 1863 11591 1897
rect 11625 1863 11659 1897
rect 11693 1863 11727 1897
rect 11761 1863 11795 1897
rect 11829 1863 11863 1897
rect 11897 1863 11931 1897
rect 11965 1863 11999 1897
rect 12033 1863 12067 1897
rect 12101 1863 12135 1897
rect 12169 1863 12203 1897
rect 12237 1863 12271 1897
rect 12305 1863 12339 1897
rect 12373 1863 12407 1897
rect 12441 1863 12475 1897
rect 12509 1863 12543 1897
rect 12577 1863 12611 1897
rect 12645 1863 12679 1897
rect 12713 1863 12747 1897
rect 12781 1863 12815 1897
rect 12849 1863 12883 1897
rect 12917 1863 13040 1897
rect 8000 1840 13040 1863
rect 8000 1760 8080 1840
rect 12720 1817 13040 1840
rect 12720 1783 12823 1817
rect 12857 1783 13040 1817
rect 12720 1760 13040 1783
rect 8000 1737 13040 1760
rect 8000 1703 8123 1737
rect 8157 1703 8191 1737
rect 8225 1703 8259 1737
rect 8293 1703 8327 1737
rect 8361 1703 8395 1737
rect 8429 1703 8463 1737
rect 8497 1703 8531 1737
rect 8565 1703 8599 1737
rect 8633 1703 8667 1737
rect 8701 1703 8735 1737
rect 8769 1703 8803 1737
rect 8837 1703 8871 1737
rect 8905 1703 8939 1737
rect 8973 1703 9007 1737
rect 9041 1703 9075 1737
rect 9109 1703 9143 1737
rect 9177 1703 9211 1737
rect 9245 1703 9279 1737
rect 9313 1703 9347 1737
rect 9381 1703 9415 1737
rect 9449 1703 9483 1737
rect 9517 1703 9551 1737
rect 9585 1703 9619 1737
rect 9653 1703 9687 1737
rect 9721 1703 9755 1737
rect 9789 1703 9823 1737
rect 9857 1703 9891 1737
rect 9925 1703 9959 1737
rect 9993 1703 10027 1737
rect 10061 1703 10095 1737
rect 10129 1703 10163 1737
rect 10197 1703 10231 1737
rect 10265 1703 10299 1737
rect 10333 1703 10367 1737
rect 10401 1703 10435 1737
rect 10469 1703 10503 1737
rect 10537 1703 10571 1737
rect 10605 1703 10639 1737
rect 10673 1703 10707 1737
rect 10741 1703 10775 1737
rect 10809 1703 10843 1737
rect 10877 1703 10911 1737
rect 10945 1703 10979 1737
rect 11013 1703 11047 1737
rect 11081 1703 11115 1737
rect 11149 1703 11183 1737
rect 11217 1703 11251 1737
rect 11285 1703 11319 1737
rect 11353 1703 11387 1737
rect 11421 1703 11455 1737
rect 11489 1703 11523 1737
rect 11557 1703 11591 1737
rect 11625 1703 11659 1737
rect 11693 1703 11727 1737
rect 11761 1703 11795 1737
rect 11829 1703 11863 1737
rect 11897 1703 11931 1737
rect 11965 1703 11999 1737
rect 12033 1703 12067 1737
rect 12101 1703 12135 1737
rect 12169 1703 12203 1737
rect 12237 1703 12271 1737
rect 12305 1703 12339 1737
rect 12373 1703 12407 1737
rect 12441 1703 12475 1737
rect 12509 1703 12543 1737
rect 12577 1703 12611 1737
rect 12645 1703 12679 1737
rect 12713 1703 12747 1737
rect 12781 1703 12815 1737
rect 12849 1703 12883 1737
rect 12917 1703 13040 1737
rect 8000 1680 13040 1703
rect 8000 1639 8080 1680
rect 8000 1605 8023 1639
rect 8057 1605 8080 1639
rect 8000 1571 8080 1605
rect 12960 1639 13040 1680
rect 12960 1605 12983 1639
rect 13017 1605 13040 1639
rect 8000 1537 8023 1571
rect 8057 1537 8080 1571
rect 8000 1503 8080 1537
rect 8000 1469 8023 1503
rect 8057 1469 8080 1503
rect 8000 1435 8080 1469
rect 8000 1401 8023 1435
rect 8057 1401 8080 1435
rect 8000 1367 8080 1401
rect 8000 1333 8023 1367
rect 8057 1333 8080 1367
rect 8000 1299 8080 1333
rect 8000 1265 8023 1299
rect 8057 1265 8080 1299
rect 8000 1231 8080 1265
rect 8000 1197 8023 1231
rect 8057 1197 8080 1231
rect 8000 1163 8080 1197
rect 8000 1129 8023 1163
rect 8057 1129 8080 1163
rect 8000 1095 8080 1129
rect 8000 1061 8023 1095
rect 8057 1061 8080 1095
rect 8000 1027 8080 1061
rect 8000 993 8023 1027
rect 8057 993 8080 1027
rect 8000 959 8080 993
rect 8000 925 8023 959
rect 8057 925 8080 959
rect 8000 891 8080 925
rect 8000 857 8023 891
rect 8057 857 8080 891
rect 8000 823 8080 857
rect 8000 789 8023 823
rect 8057 789 8080 823
rect 8000 755 8080 789
rect 8000 721 8023 755
rect 8057 721 8080 755
rect 8000 640 8080 721
rect 8160 1577 12880 1600
rect 8160 1543 8293 1577
rect 8327 1543 8361 1577
rect 8395 1543 8429 1577
rect 8463 1543 8497 1577
rect 8531 1543 8565 1577
rect 8599 1543 8633 1577
rect 8667 1543 8701 1577
rect 8735 1543 8769 1577
rect 8803 1543 8837 1577
rect 8871 1543 8905 1577
rect 8939 1543 8973 1577
rect 9007 1543 9041 1577
rect 9075 1543 9109 1577
rect 9143 1543 9177 1577
rect 9211 1543 9245 1577
rect 9279 1543 9313 1577
rect 9347 1543 9381 1577
rect 9415 1543 9449 1577
rect 9483 1543 9517 1577
rect 9551 1543 9585 1577
rect 9619 1543 9653 1577
rect 9687 1543 9721 1577
rect 9755 1543 9789 1577
rect 9823 1543 9857 1577
rect 9891 1543 9925 1577
rect 9959 1543 9993 1577
rect 10027 1543 10061 1577
rect 10095 1543 10129 1577
rect 10163 1543 10197 1577
rect 10231 1543 10265 1577
rect 10299 1543 10333 1577
rect 10367 1543 10401 1577
rect 10435 1543 10469 1577
rect 10503 1543 10537 1577
rect 10571 1543 10605 1577
rect 10639 1543 10673 1577
rect 10707 1543 10741 1577
rect 10775 1543 10809 1577
rect 10843 1543 10877 1577
rect 10911 1543 10945 1577
rect 10979 1543 11013 1577
rect 11047 1543 11081 1577
rect 11115 1543 11149 1577
rect 11183 1543 11217 1577
rect 11251 1543 11285 1577
rect 11319 1543 11353 1577
rect 11387 1543 11421 1577
rect 11455 1543 11489 1577
rect 11523 1543 11557 1577
rect 11591 1543 11625 1577
rect 11659 1543 11693 1577
rect 11727 1543 11761 1577
rect 11795 1543 11829 1577
rect 11863 1543 11897 1577
rect 11931 1543 11965 1577
rect 11999 1543 12033 1577
rect 12067 1543 12101 1577
rect 12135 1543 12169 1577
rect 12203 1543 12237 1577
rect 12271 1543 12305 1577
rect 12339 1543 12373 1577
rect 12407 1543 12441 1577
rect 12475 1543 12509 1577
rect 12543 1543 12577 1577
rect 12611 1543 12645 1577
rect 12679 1543 12713 1577
rect 12747 1543 12880 1577
rect 8160 1520 12880 1543
rect 8160 1463 8240 1520
rect 8160 1429 8183 1463
rect 8217 1429 8240 1463
rect 12800 1463 12880 1520
rect 8160 1395 8240 1429
rect 8160 1361 8183 1395
rect 8217 1361 8240 1395
rect 8160 1327 8240 1361
rect 8320 1417 8400 1440
rect 8320 1383 8343 1417
rect 8377 1383 8400 1417
rect 8320 1356 8400 1383
rect 12640 1417 12720 1440
rect 12640 1383 12663 1417
rect 12697 1383 12720 1417
rect 12640 1356 12720 1383
rect 12800 1429 12823 1463
rect 12857 1429 12880 1463
rect 12800 1395 12880 1429
rect 12800 1361 12823 1395
rect 12857 1361 12880 1395
rect 8160 1293 8183 1327
rect 8217 1293 8240 1327
rect 8160 1259 8240 1293
rect 12800 1327 12880 1361
rect 12800 1293 12823 1327
rect 12857 1293 12880 1327
rect 8160 1225 8183 1259
rect 8217 1225 8240 1259
rect 8160 1191 8240 1225
rect 8520 1257 12520 1280
rect 8520 1223 8559 1257
rect 8599 1223 8631 1257
rect 8667 1223 8701 1257
rect 8737 1223 8769 1257
rect 8809 1223 8837 1257
rect 8881 1223 8905 1257
rect 8953 1223 8973 1257
rect 9025 1223 9041 1257
rect 9097 1223 9109 1257
rect 9169 1223 9177 1257
rect 9241 1223 9245 1257
rect 9347 1223 9351 1257
rect 9415 1223 9423 1257
rect 9483 1223 9495 1257
rect 9551 1223 9567 1257
rect 9619 1223 9639 1257
rect 9687 1223 9711 1257
rect 9755 1223 9783 1257
rect 9823 1223 9855 1257
rect 9891 1223 9925 1257
rect 9961 1223 9993 1257
rect 10033 1223 10061 1257
rect 10105 1223 10129 1257
rect 10177 1223 10197 1257
rect 10249 1223 10265 1257
rect 10321 1223 10333 1257
rect 10393 1223 10401 1257
rect 10465 1223 10469 1257
rect 10571 1223 10575 1257
rect 10639 1223 10647 1257
rect 10707 1223 10719 1257
rect 10775 1223 10791 1257
rect 10843 1223 10863 1257
rect 10911 1223 10935 1257
rect 10979 1223 11007 1257
rect 11047 1223 11079 1257
rect 11115 1223 11149 1257
rect 11185 1223 11217 1257
rect 11257 1223 11285 1257
rect 11329 1223 11353 1257
rect 11401 1223 11421 1257
rect 11473 1223 11489 1257
rect 11545 1223 11557 1257
rect 11617 1223 11625 1257
rect 11689 1223 11693 1257
rect 11795 1223 11799 1257
rect 11863 1223 11871 1257
rect 11931 1223 11943 1257
rect 11999 1223 12015 1257
rect 12067 1223 12087 1257
rect 12135 1223 12159 1257
rect 12203 1223 12231 1257
rect 12271 1223 12303 1257
rect 12339 1223 12373 1257
rect 12409 1223 12441 1257
rect 12481 1223 12520 1257
rect 8520 1200 12520 1223
rect 12800 1259 12880 1293
rect 12800 1225 12823 1259
rect 12857 1225 12880 1259
rect 8160 1157 8183 1191
rect 8217 1157 8240 1191
rect 8160 1123 8240 1157
rect 8160 1089 8183 1123
rect 8217 1089 8240 1123
rect 12800 1191 12880 1225
rect 12800 1157 12823 1191
rect 12857 1157 12880 1191
rect 12800 1123 12880 1157
rect 8160 1055 8240 1089
rect 8160 1021 8183 1055
rect 8217 1021 8240 1055
rect 8320 1097 8400 1120
rect 8320 1063 8343 1097
rect 8377 1063 8400 1097
rect 8320 1036 8400 1063
rect 12640 1097 12720 1120
rect 12640 1063 12663 1097
rect 12697 1063 12720 1097
rect 12640 1036 12720 1063
rect 12800 1089 12823 1123
rect 12857 1089 12880 1123
rect 12800 1055 12880 1089
rect 8160 987 8240 1021
rect 8160 953 8183 987
rect 8217 953 8240 987
rect 12800 1021 12823 1055
rect 12857 1021 12880 1055
rect 12800 987 12880 1021
rect 8160 919 8240 953
rect 8160 885 8183 919
rect 8217 885 8240 919
rect 8160 851 8240 885
rect 8520 937 12520 960
rect 8520 903 8559 937
rect 8599 903 8631 937
rect 8667 903 8701 937
rect 8737 903 8769 937
rect 8809 903 8837 937
rect 8881 903 8905 937
rect 8953 903 8973 937
rect 9025 903 9041 937
rect 9097 903 9109 937
rect 9169 903 9177 937
rect 9241 903 9245 937
rect 9347 903 9351 937
rect 9415 903 9423 937
rect 9483 903 9495 937
rect 9551 903 9567 937
rect 9619 903 9639 937
rect 9687 903 9711 937
rect 9755 903 9783 937
rect 9823 903 9855 937
rect 9891 903 9925 937
rect 9961 903 9993 937
rect 10033 903 10061 937
rect 10105 903 10129 937
rect 10177 903 10197 937
rect 10249 903 10265 937
rect 10321 903 10333 937
rect 10393 903 10401 937
rect 10465 903 10469 937
rect 10571 903 10575 937
rect 10639 903 10647 937
rect 10707 903 10719 937
rect 10775 903 10791 937
rect 10843 903 10863 937
rect 10911 903 10935 937
rect 10979 903 11007 937
rect 11047 903 11079 937
rect 11115 903 11149 937
rect 11185 903 11217 937
rect 11257 903 11285 937
rect 11329 903 11353 937
rect 11401 903 11421 937
rect 11473 903 11489 937
rect 11545 903 11557 937
rect 11617 903 11625 937
rect 11689 903 11693 937
rect 11795 903 11799 937
rect 11863 903 11871 937
rect 11931 903 11943 937
rect 11999 903 12015 937
rect 12067 903 12087 937
rect 12135 903 12159 937
rect 12203 903 12231 937
rect 12271 903 12303 937
rect 12339 903 12373 937
rect 12409 903 12441 937
rect 12481 903 12520 937
rect 8520 880 12520 903
rect 12800 953 12823 987
rect 12857 953 12880 987
rect 12800 919 12880 953
rect 12800 885 12823 919
rect 12857 885 12880 919
rect 8160 817 8183 851
rect 8217 817 8240 851
rect 8160 800 8240 817
rect 12800 851 12880 885
rect 12800 817 12823 851
rect 12857 817 12880 851
rect 12800 800 12880 817
rect 8160 777 12880 800
rect 8160 743 8293 777
rect 8327 743 8343 777
rect 8395 743 8429 777
rect 8463 743 8497 777
rect 8531 743 8565 777
rect 8599 743 8633 777
rect 8667 743 8701 777
rect 8735 743 8769 777
rect 8803 743 8837 777
rect 8871 743 8905 777
rect 8939 743 8973 777
rect 9007 743 9041 777
rect 9075 743 9109 777
rect 9143 743 9177 777
rect 9211 743 9245 777
rect 9279 743 9313 777
rect 9347 743 9381 777
rect 9415 743 9449 777
rect 9483 743 9517 777
rect 9551 743 9585 777
rect 9619 743 9653 777
rect 9687 743 9721 777
rect 9755 743 9789 777
rect 9823 743 9857 777
rect 9891 743 9925 777
rect 9959 743 9993 777
rect 10027 743 10061 777
rect 10095 743 10129 777
rect 10163 743 10197 777
rect 10231 743 10265 777
rect 10299 743 10333 777
rect 10367 743 10401 777
rect 10435 743 10469 777
rect 10503 743 10537 777
rect 10571 743 10605 777
rect 10639 743 10673 777
rect 10707 743 10741 777
rect 10775 743 10809 777
rect 10843 743 10877 777
rect 10911 743 10945 777
rect 10979 743 11013 777
rect 11047 743 11081 777
rect 11115 743 11149 777
rect 11183 743 11217 777
rect 11251 743 11285 777
rect 11319 743 11353 777
rect 11387 743 11421 777
rect 11455 743 11489 777
rect 11523 743 11557 777
rect 11591 743 11625 777
rect 11659 743 11693 777
rect 11727 743 11761 777
rect 11795 743 11829 777
rect 11863 743 11897 777
rect 11931 743 11965 777
rect 11999 743 12033 777
rect 12067 743 12101 777
rect 12135 743 12169 777
rect 12203 743 12237 777
rect 12271 743 12305 777
rect 12339 743 12373 777
rect 12407 743 12441 777
rect 12475 743 12509 777
rect 12543 743 12577 777
rect 12611 743 12645 777
rect 12679 743 12713 777
rect 12747 743 12880 777
rect 8160 720 12880 743
rect 12960 1571 13040 1605
rect 12960 1537 12983 1571
rect 13017 1537 13040 1571
rect 12960 1503 13040 1537
rect 12960 1469 12983 1503
rect 13017 1469 13040 1503
rect 12960 1435 13040 1469
rect 12960 1401 12983 1435
rect 13017 1401 13040 1435
rect 12960 1367 13040 1401
rect 12960 1333 12983 1367
rect 13017 1333 13040 1367
rect 12960 1299 13040 1333
rect 12960 1265 12983 1299
rect 13017 1265 13040 1299
rect 12960 1231 13040 1265
rect 12960 1197 12983 1231
rect 13017 1197 13040 1231
rect 12960 1163 13040 1197
rect 12960 1129 12983 1163
rect 13017 1129 13040 1163
rect 12960 1095 13040 1129
rect 12960 1061 12983 1095
rect 13017 1061 13040 1095
rect 12960 1027 13040 1061
rect 12960 993 12983 1027
rect 13017 993 13040 1027
rect 12960 959 13040 993
rect 12960 925 12983 959
rect 13017 925 13040 959
rect 12960 891 13040 925
rect 12960 857 12983 891
rect 13017 857 13040 891
rect 12960 823 13040 857
rect 12960 789 12983 823
rect 13017 789 13040 823
rect 12960 755 13040 789
rect 12960 721 12983 755
rect 13017 721 13040 755
rect 12960 640 13040 721
rect 8000 617 13040 640
rect 8000 583 8123 617
rect 8157 583 8191 617
rect 8225 583 8259 617
rect 8293 583 8327 617
rect 8361 583 8395 617
rect 8429 583 8463 617
rect 8497 583 8531 617
rect 8565 583 8599 617
rect 8633 583 8667 617
rect 8701 583 8735 617
rect 8769 583 8803 617
rect 8837 583 8871 617
rect 8905 583 8939 617
rect 8973 583 9007 617
rect 9041 583 9075 617
rect 9109 583 9143 617
rect 9177 583 9211 617
rect 9245 583 9279 617
rect 9313 583 9347 617
rect 9381 583 9415 617
rect 9449 583 9483 617
rect 9517 583 9551 617
rect 9585 583 9619 617
rect 9653 583 9687 617
rect 9721 583 9755 617
rect 9789 583 9823 617
rect 9857 583 9891 617
rect 9925 583 9959 617
rect 9993 583 10027 617
rect 10061 583 10095 617
rect 10129 583 10163 617
rect 10197 583 10231 617
rect 10265 583 10299 617
rect 10333 583 10367 617
rect 10401 583 10435 617
rect 10469 583 10503 617
rect 10537 583 10571 617
rect 10605 583 10639 617
rect 10673 583 10707 617
rect 10741 583 10775 617
rect 10809 583 10843 617
rect 10877 583 10911 617
rect 10945 583 10979 617
rect 11013 583 11047 617
rect 11081 583 11115 617
rect 11149 583 11183 617
rect 11217 583 11251 617
rect 11285 583 11319 617
rect 11353 583 11387 617
rect 11421 583 11455 617
rect 11489 583 11523 617
rect 11557 583 11591 617
rect 11625 583 11659 617
rect 11693 583 11727 617
rect 11761 583 11795 617
rect 11829 583 11863 617
rect 11897 583 11931 617
rect 11965 583 11999 617
rect 12033 583 12067 617
rect 12101 583 12135 617
rect 12169 583 12203 617
rect 12237 583 12271 617
rect 12305 583 12339 617
rect 12373 583 12407 617
rect 12441 583 12475 617
rect 12509 583 12543 617
rect 12577 583 12611 617
rect 12645 583 12679 617
rect 12713 583 12747 617
rect 12781 583 12815 617
rect 12849 583 12883 617
rect 12917 583 13040 617
rect 8000 560 13040 583
rect 8000 480 8080 560
rect 12960 480 13040 560
rect 8000 457 13040 480
rect 8000 423 8123 457
rect 8157 423 8191 457
rect 8225 423 8259 457
rect 8293 423 8327 457
rect 8361 423 8395 457
rect 8429 423 8463 457
rect 8497 423 8531 457
rect 8565 423 8599 457
rect 8633 423 8667 457
rect 8701 423 8735 457
rect 8769 423 8803 457
rect 8837 423 8871 457
rect 8905 423 8939 457
rect 8973 423 9007 457
rect 9041 423 9075 457
rect 9109 423 9143 457
rect 9177 423 9211 457
rect 9245 423 9279 457
rect 9313 423 9347 457
rect 9381 423 9415 457
rect 9449 423 9483 457
rect 9517 423 9551 457
rect 9585 423 9619 457
rect 9653 423 9687 457
rect 9721 423 9755 457
rect 9789 423 9823 457
rect 9857 423 9891 457
rect 9925 423 9959 457
rect 9993 423 10027 457
rect 10061 423 10095 457
rect 10129 423 10163 457
rect 10197 423 10231 457
rect 10265 423 10299 457
rect 10333 423 10367 457
rect 10401 423 10435 457
rect 10469 423 10503 457
rect 10537 423 10571 457
rect 10605 423 10639 457
rect 10673 423 10707 457
rect 10741 423 10775 457
rect 10809 423 10843 457
rect 10877 423 10911 457
rect 10945 423 10979 457
rect 11013 423 11047 457
rect 11081 423 11115 457
rect 11149 423 11183 457
rect 11217 423 11251 457
rect 11285 423 11319 457
rect 11353 423 11387 457
rect 11421 423 11455 457
rect 11489 423 11523 457
rect 11557 423 11591 457
rect 11625 423 11659 457
rect 11693 423 11727 457
rect 11761 423 11795 457
rect 11829 423 11863 457
rect 11897 423 11931 457
rect 11965 423 11999 457
rect 12033 423 12067 457
rect 12101 423 12135 457
rect 12169 423 12203 457
rect 12237 423 12271 457
rect 12305 423 12339 457
rect 12373 423 12407 457
rect 12441 423 12475 457
rect 12509 423 12543 457
rect 12577 423 12611 457
rect 12645 423 12679 457
rect 12713 423 12747 457
rect 12781 423 12815 457
rect 12849 423 12883 457
rect 12917 423 13040 457
rect 8000 400 13040 423
rect 8000 319 8080 400
rect 8000 285 8023 319
rect 8057 285 8080 319
rect 8000 251 8080 285
rect 8000 217 8023 251
rect 8057 217 8080 251
rect 8000 183 8080 217
rect 8000 149 8023 183
rect 8057 149 8080 183
rect 8000 115 8080 149
rect 8000 81 8023 115
rect 8057 81 8080 115
rect 8000 47 8080 81
rect 8000 13 8023 47
rect 8057 13 8080 47
rect 8000 -21 8080 13
rect 8000 -55 8023 -21
rect 8057 -55 8080 -21
rect 8000 -89 8080 -55
rect 8000 -123 8023 -89
rect 8057 -123 8080 -89
rect 8000 -157 8080 -123
rect 8000 -191 8023 -157
rect 8057 -191 8080 -157
rect 8000 -225 8080 -191
rect 8000 -259 8023 -225
rect 8057 -259 8080 -225
rect 8000 -293 8080 -259
rect 8000 -327 8023 -293
rect 8057 -327 8080 -293
rect 8000 -361 8080 -327
rect 8000 -395 8023 -361
rect 8057 -395 8080 -361
rect 8000 -429 8080 -395
rect 8000 -463 8023 -429
rect 8057 -463 8080 -429
rect 8000 -497 8080 -463
rect 8000 -531 8023 -497
rect 8057 -531 8080 -497
rect 8000 -565 8080 -531
rect 8160 297 12880 320
rect 8160 263 8293 297
rect 8327 263 8361 297
rect 8395 263 8429 297
rect 8463 263 8497 297
rect 8531 263 8565 297
rect 8599 263 8633 297
rect 8667 263 8701 297
rect 8735 263 8769 297
rect 8803 263 8837 297
rect 8871 263 8905 297
rect 8939 263 8973 297
rect 9007 263 9041 297
rect 9075 263 9109 297
rect 9143 263 9177 297
rect 9211 263 9245 297
rect 9279 263 9313 297
rect 9347 263 9381 297
rect 9415 263 9449 297
rect 9483 263 9517 297
rect 9551 263 9585 297
rect 9619 263 9653 297
rect 9687 263 9721 297
rect 9755 263 9789 297
rect 9823 263 9857 297
rect 9891 263 9925 297
rect 9959 263 9993 297
rect 10027 263 10061 297
rect 10095 263 10129 297
rect 10163 263 10197 297
rect 10231 263 10265 297
rect 10299 263 10333 297
rect 10367 263 10401 297
rect 10435 263 10469 297
rect 10503 263 10537 297
rect 10571 263 10605 297
rect 10639 263 10673 297
rect 10707 263 10741 297
rect 10775 263 10809 297
rect 10843 263 10877 297
rect 10911 263 10945 297
rect 10979 263 11013 297
rect 11047 263 11081 297
rect 11115 263 11149 297
rect 11183 263 11217 297
rect 11251 263 11285 297
rect 11319 263 11353 297
rect 11387 263 11421 297
rect 11455 263 11489 297
rect 11523 263 11557 297
rect 11591 263 11625 297
rect 11659 263 11693 297
rect 11727 263 11761 297
rect 11795 263 11829 297
rect 11863 263 11897 297
rect 11931 263 11965 297
rect 11999 263 12033 297
rect 12067 263 12101 297
rect 12135 263 12169 297
rect 12203 263 12237 297
rect 12271 263 12305 297
rect 12339 263 12373 297
rect 12407 263 12441 297
rect 12475 263 12509 297
rect 12543 263 12577 297
rect 12611 263 12645 297
rect 12679 263 12713 297
rect 12747 263 12880 297
rect 8160 240 12880 263
rect 8160 223 8240 240
rect 8160 189 8183 223
rect 8217 189 8240 223
rect 8160 155 8240 189
rect 12800 223 12880 240
rect 12800 189 12823 223
rect 12857 189 12880 223
rect 8160 121 8183 155
rect 8217 121 8240 155
rect 8160 87 8240 121
rect 8160 53 8183 87
rect 8217 53 8240 87
rect 8520 137 12520 160
rect 8520 103 8559 137
rect 8599 103 8631 137
rect 8667 103 8701 137
rect 8737 103 8769 137
rect 8809 103 8837 137
rect 8881 103 8905 137
rect 8953 103 8973 137
rect 9025 103 9041 137
rect 9097 103 9109 137
rect 9169 103 9177 137
rect 9241 103 9245 137
rect 9347 103 9351 137
rect 9415 103 9423 137
rect 9483 103 9495 137
rect 9551 103 9567 137
rect 9619 103 9639 137
rect 9687 103 9711 137
rect 9755 103 9783 137
rect 9823 103 9855 137
rect 9891 103 9925 137
rect 9961 103 9993 137
rect 10033 103 10061 137
rect 10105 103 10129 137
rect 10177 103 10197 137
rect 10249 103 10265 137
rect 10321 103 10333 137
rect 10393 103 10401 137
rect 10465 103 10469 137
rect 10571 103 10575 137
rect 10639 103 10647 137
rect 10707 103 10719 137
rect 10775 103 10791 137
rect 10843 103 10863 137
rect 10911 103 10935 137
rect 10979 103 11007 137
rect 11047 103 11079 137
rect 11115 103 11149 137
rect 11185 103 11217 137
rect 11257 103 11285 137
rect 11329 103 11353 137
rect 11401 103 11421 137
rect 11473 103 11489 137
rect 11545 103 11557 137
rect 11617 103 11625 137
rect 11689 103 11693 137
rect 11795 103 11799 137
rect 11863 103 11871 137
rect 11931 103 11943 137
rect 11999 103 12015 137
rect 12067 103 12087 137
rect 12135 103 12159 137
rect 12203 103 12231 137
rect 12271 103 12303 137
rect 12339 103 12373 137
rect 12409 103 12441 137
rect 12481 103 12520 137
rect 8520 80 12520 103
rect 12800 155 12880 189
rect 12800 121 12823 155
rect 12857 121 12880 155
rect 12800 87 12880 121
rect 8160 19 8240 53
rect 8160 -15 8183 19
rect 8217 -15 8240 19
rect 12800 53 12823 87
rect 12857 53 12880 87
rect 12800 19 12880 53
rect 8160 -49 8240 -15
rect 8160 -83 8183 -49
rect 8217 -83 8240 -49
rect 8320 -23 8400 4
rect 8320 -57 8343 -23
rect 8377 -57 8400 -23
rect 8320 -80 8400 -57
rect 12640 -23 12720 4
rect 12640 -57 12663 -23
rect 12697 -57 12720 -23
rect 12640 -80 12720 -57
rect 12800 -15 12823 19
rect 12857 -15 12880 19
rect 12800 -49 12880 -15
rect 8160 -117 8240 -83
rect 8160 -151 8183 -117
rect 8217 -151 8240 -117
rect 8160 -185 8240 -151
rect 12800 -83 12823 -49
rect 12857 -83 12880 -49
rect 12800 -117 12880 -83
rect 12800 -151 12823 -117
rect 12857 -151 12880 -117
rect 8160 -219 8183 -185
rect 8217 -219 8240 -185
rect 8160 -253 8240 -219
rect 8520 -183 12520 -160
rect 8520 -217 8559 -183
rect 8599 -217 8631 -183
rect 8667 -217 8701 -183
rect 8737 -217 8769 -183
rect 8809 -217 8837 -183
rect 8881 -217 8905 -183
rect 8953 -217 8973 -183
rect 9025 -217 9041 -183
rect 9097 -217 9109 -183
rect 9169 -217 9177 -183
rect 9241 -217 9245 -183
rect 9347 -217 9351 -183
rect 9415 -217 9423 -183
rect 9483 -217 9495 -183
rect 9551 -217 9567 -183
rect 9619 -217 9639 -183
rect 9687 -217 9711 -183
rect 9755 -217 9783 -183
rect 9823 -217 9855 -183
rect 9891 -217 9925 -183
rect 9961 -217 9993 -183
rect 10033 -217 10061 -183
rect 10105 -217 10129 -183
rect 10177 -217 10197 -183
rect 10249 -217 10265 -183
rect 10321 -217 10333 -183
rect 10393 -217 10401 -183
rect 10465 -217 10469 -183
rect 10571 -217 10575 -183
rect 10639 -217 10647 -183
rect 10707 -217 10719 -183
rect 10775 -217 10791 -183
rect 10843 -217 10863 -183
rect 10911 -217 10935 -183
rect 10979 -217 11007 -183
rect 11047 -217 11079 -183
rect 11115 -217 11149 -183
rect 11185 -217 11217 -183
rect 11257 -217 11285 -183
rect 11329 -217 11353 -183
rect 11401 -217 11421 -183
rect 11473 -217 11489 -183
rect 11545 -217 11557 -183
rect 11617 -217 11625 -183
rect 11689 -217 11693 -183
rect 11795 -217 11799 -183
rect 11863 -217 11871 -183
rect 11931 -217 11943 -183
rect 11999 -217 12015 -183
rect 12067 -217 12087 -183
rect 12135 -217 12159 -183
rect 12203 -217 12231 -183
rect 12271 -217 12303 -183
rect 12339 -217 12373 -183
rect 12409 -217 12441 -183
rect 12481 -217 12520 -183
rect 8520 -240 12520 -217
rect 12800 -185 12880 -151
rect 12800 -219 12823 -185
rect 12857 -219 12880 -185
rect 8160 -287 8183 -253
rect 8217 -287 8240 -253
rect 8160 -321 8240 -287
rect 12800 -253 12880 -219
rect 12800 -287 12823 -253
rect 12857 -287 12880 -253
rect 8160 -355 8183 -321
rect 8217 -355 8240 -321
rect 8160 -389 8240 -355
rect 8160 -423 8183 -389
rect 8217 -423 8240 -389
rect 8320 -343 8400 -316
rect 8320 -377 8343 -343
rect 8377 -377 8400 -343
rect 8320 -400 8400 -377
rect 12640 -343 12720 -316
rect 12640 -377 12663 -343
rect 12697 -377 12720 -343
rect 12640 -400 12720 -377
rect 12800 -321 12880 -287
rect 12800 -355 12823 -321
rect 12857 -355 12880 -321
rect 12800 -389 12880 -355
rect 8160 -480 8240 -423
rect 12800 -423 12823 -389
rect 12857 -423 12880 -389
rect 12800 -480 12880 -423
rect 8160 -503 12880 -480
rect 8160 -537 8293 -503
rect 8327 -537 8361 -503
rect 8395 -537 8429 -503
rect 8463 -537 8497 -503
rect 8531 -537 8565 -503
rect 8599 -537 8633 -503
rect 8667 -537 8701 -503
rect 8735 -537 8769 -503
rect 8803 -537 8837 -503
rect 8871 -537 8905 -503
rect 8939 -537 8973 -503
rect 9007 -537 9041 -503
rect 9075 -537 9109 -503
rect 9143 -537 9177 -503
rect 9211 -537 9245 -503
rect 9279 -537 9313 -503
rect 9347 -537 9381 -503
rect 9415 -537 9449 -503
rect 9483 -537 9517 -503
rect 9551 -537 9585 -503
rect 9619 -537 9653 -503
rect 9687 -537 9721 -503
rect 9755 -537 9789 -503
rect 9823 -537 9857 -503
rect 9891 -537 9925 -503
rect 9959 -537 9993 -503
rect 10027 -537 10061 -503
rect 10095 -537 10129 -503
rect 10163 -537 10197 -503
rect 10231 -537 10265 -503
rect 10299 -537 10333 -503
rect 10367 -537 10401 -503
rect 10435 -537 10469 -503
rect 10503 -537 10537 -503
rect 10571 -537 10605 -503
rect 10639 -537 10673 -503
rect 10707 -537 10741 -503
rect 10775 -537 10809 -503
rect 10843 -537 10877 -503
rect 10911 -537 10945 -503
rect 10979 -537 11013 -503
rect 11047 -537 11081 -503
rect 11115 -537 11149 -503
rect 11183 -537 11217 -503
rect 11251 -537 11285 -503
rect 11319 -537 11353 -503
rect 11387 -537 11421 -503
rect 11455 -537 11489 -503
rect 11523 -537 11557 -503
rect 11591 -537 11625 -503
rect 11659 -537 11693 -503
rect 11727 -537 11761 -503
rect 11795 -537 11829 -503
rect 11863 -537 11897 -503
rect 11931 -537 11965 -503
rect 11999 -537 12033 -503
rect 12067 -537 12101 -503
rect 12135 -537 12169 -503
rect 12203 -537 12237 -503
rect 12271 -537 12305 -503
rect 12339 -537 12373 -503
rect 12407 -537 12441 -503
rect 12475 -537 12509 -503
rect 12543 -537 12577 -503
rect 12611 -537 12645 -503
rect 12679 -537 12713 -503
rect 12747 -537 12823 -503
rect 12857 -537 12880 -503
rect 8160 -560 12880 -537
rect 12960 319 13040 400
rect 12960 285 12983 319
rect 13017 285 13040 319
rect 12960 251 13040 285
rect 12960 217 12983 251
rect 13017 217 13040 251
rect 12960 183 13040 217
rect 12960 149 12983 183
rect 13017 149 13040 183
rect 12960 115 13040 149
rect 12960 81 12983 115
rect 13017 81 13040 115
rect 12960 47 13040 81
rect 12960 13 12983 47
rect 13017 13 13040 47
rect 12960 -21 13040 13
rect 12960 -55 12983 -21
rect 13017 -55 13040 -21
rect 12960 -89 13040 -55
rect 12960 -123 12983 -89
rect 13017 -123 13040 -89
rect 12960 -157 13040 -123
rect 12960 -191 12983 -157
rect 13017 -191 13040 -157
rect 12960 -225 13040 -191
rect 12960 -259 12983 -225
rect 13017 -259 13040 -225
rect 12960 -293 13040 -259
rect 12960 -327 12983 -293
rect 13017 -327 13040 -293
rect 12960 -361 13040 -327
rect 12960 -395 12983 -361
rect 13017 -395 13040 -361
rect 12960 -429 13040 -395
rect 12960 -463 12983 -429
rect 13017 -463 13040 -429
rect 12960 -497 13040 -463
rect 12960 -531 12983 -497
rect 13017 -531 13040 -497
rect 8000 -599 8023 -565
rect 8057 -599 8080 -565
rect 8000 -640 8080 -599
rect 12960 -565 13040 -531
rect 12960 -599 12983 -565
rect 13017 -599 13040 -565
rect 12960 -640 13040 -599
rect -480 -663 13040 -640
rect -480 -697 -357 -663
rect -323 -697 -289 -663
rect -255 -697 -221 -663
rect -187 -697 -153 -663
rect -119 -697 -85 -663
rect -51 -697 -17 -663
rect 17 -697 51 -663
rect 85 -697 119 -663
rect 153 -697 187 -663
rect 221 -697 255 -663
rect 289 -697 323 -663
rect 357 -697 391 -663
rect 425 -697 459 -663
rect 493 -697 527 -663
rect 561 -697 595 -663
rect 629 -697 663 -663
rect 697 -697 731 -663
rect 765 -697 799 -663
rect 833 -697 867 -663
rect 901 -697 935 -663
rect 969 -697 1003 -663
rect 1037 -697 1071 -663
rect 1105 -697 1139 -663
rect 1173 -697 1207 -663
rect 1241 -697 1275 -663
rect 1309 -697 1343 -663
rect 1377 -697 1411 -663
rect 1445 -697 1479 -663
rect 1513 -697 1547 -663
rect 1581 -697 1615 -663
rect 1649 -697 1683 -663
rect 1717 -697 1751 -663
rect 1785 -697 1819 -663
rect 1853 -697 1887 -663
rect 1921 -697 1955 -663
rect 1989 -697 2023 -663
rect 2057 -697 2091 -663
rect 2125 -697 2159 -663
rect 2193 -697 2227 -663
rect 2261 -697 2295 -663
rect 2329 -697 2363 -663
rect 2397 -697 2431 -663
rect 2465 -697 2499 -663
rect 2533 -697 2567 -663
rect 2601 -697 2635 -663
rect 2669 -697 2703 -663
rect 2737 -697 2771 -663
rect 2805 -697 2839 -663
rect 2873 -697 2907 -663
rect 2941 -697 2975 -663
rect 3009 -697 3043 -663
rect 3077 -697 3111 -663
rect 3145 -697 3179 -663
rect 3213 -697 3247 -663
rect 3281 -697 3315 -663
rect 3349 -697 3383 -663
rect 3417 -697 3451 -663
rect 3485 -697 3519 -663
rect 3553 -697 3587 -663
rect 3621 -697 3655 -663
rect 3689 -697 3723 -663
rect 3757 -697 3791 -663
rect 3825 -697 3859 -663
rect 3893 -697 3927 -663
rect 3961 -697 3995 -663
rect 4029 -697 4063 -663
rect 4097 -697 4131 -663
rect 4165 -697 4199 -663
rect 4233 -697 4267 -663
rect 4301 -697 4335 -663
rect 4369 -697 4403 -663
rect 4437 -697 8123 -663
rect 8157 -697 8191 -663
rect 8225 -697 8259 -663
rect 8293 -697 8327 -663
rect 8361 -697 8395 -663
rect 8429 -697 8463 -663
rect 8497 -697 8531 -663
rect 8565 -697 8599 -663
rect 8633 -697 8667 -663
rect 8701 -697 8735 -663
rect 8769 -697 8803 -663
rect 8837 -697 8871 -663
rect 8905 -697 8939 -663
rect 8973 -697 9007 -663
rect 9041 -697 9075 -663
rect 9109 -697 9143 -663
rect 9177 -697 9211 -663
rect 9245 -697 9279 -663
rect 9313 -697 9347 -663
rect 9381 -697 9415 -663
rect 9449 -697 9483 -663
rect 9517 -697 9551 -663
rect 9585 -697 9619 -663
rect 9653 -697 9687 -663
rect 9721 -697 9755 -663
rect 9789 -697 9823 -663
rect 9857 -697 9891 -663
rect 9925 -697 9959 -663
rect 9993 -697 10027 -663
rect 10061 -697 10095 -663
rect 10129 -697 10163 -663
rect 10197 -697 10231 -663
rect 10265 -697 10299 -663
rect 10333 -697 10367 -663
rect 10401 -697 10435 -663
rect 10469 -697 10503 -663
rect 10537 -697 10571 -663
rect 10605 -697 10639 -663
rect 10673 -697 10707 -663
rect 10741 -697 10775 -663
rect 10809 -697 10843 -663
rect 10877 -697 10911 -663
rect 10945 -697 10979 -663
rect 11013 -697 11047 -663
rect 11081 -697 11115 -663
rect 11149 -697 11183 -663
rect 11217 -697 11251 -663
rect 11285 -697 11319 -663
rect 11353 -697 11387 -663
rect 11421 -697 11455 -663
rect 11489 -697 11523 -663
rect 11557 -697 11591 -663
rect 11625 -697 11659 -663
rect 11693 -697 11727 -663
rect 11761 -697 11795 -663
rect 11829 -697 11863 -663
rect 11897 -697 11931 -663
rect 11965 -697 11999 -663
rect 12033 -697 12067 -663
rect 12101 -697 12135 -663
rect 12169 -697 12203 -663
rect 12237 -697 12271 -663
rect 12305 -697 12339 -663
rect 12373 -697 12407 -663
rect 12441 -697 12475 -663
rect 12509 -697 12543 -663
rect 12577 -697 12611 -663
rect 12645 -697 12679 -663
rect 12713 -697 12747 -663
rect 12781 -697 12815 -663
rect 12849 -697 12883 -663
rect 12917 -697 13040 -663
rect -480 -720 13040 -697
<< viali >>
rect -297 4103 -263 4137
rect -137 3943 -103 3977
rect 4183 3943 4217 3977
rect 79 3783 85 3817
rect 85 3783 113 3817
rect 151 3783 153 3817
rect 153 3783 185 3817
rect 223 3783 255 3817
rect 255 3783 257 3817
rect 295 3783 323 3817
rect 323 3783 329 3817
rect 367 3783 391 3817
rect 391 3783 401 3817
rect 439 3783 459 3817
rect 459 3783 473 3817
rect 511 3783 527 3817
rect 527 3783 545 3817
rect 583 3783 595 3817
rect 595 3783 617 3817
rect 655 3783 663 3817
rect 663 3783 689 3817
rect 727 3783 731 3817
rect 731 3783 761 3817
rect 799 3783 833 3817
rect 871 3783 901 3817
rect 901 3783 905 3817
rect 943 3783 969 3817
rect 969 3783 977 3817
rect 1015 3783 1037 3817
rect 1037 3783 1049 3817
rect 1087 3783 1105 3817
rect 1105 3783 1121 3817
rect 1159 3783 1173 3817
rect 1173 3783 1193 3817
rect 1231 3783 1241 3817
rect 1241 3783 1265 3817
rect 1303 3783 1309 3817
rect 1309 3783 1337 3817
rect 1375 3783 1377 3817
rect 1377 3783 1409 3817
rect 1447 3783 1479 3817
rect 1479 3783 1481 3817
rect 1519 3783 1547 3817
rect 1547 3783 1553 3817
rect 1591 3783 1615 3817
rect 1615 3783 1625 3817
rect 1663 3783 1683 3817
rect 1683 3783 1697 3817
rect 1735 3783 1751 3817
rect 1751 3783 1769 3817
rect 1807 3783 1819 3817
rect 1819 3783 1841 3817
rect 1879 3783 1887 3817
rect 1887 3783 1913 3817
rect 1951 3783 1955 3817
rect 1955 3783 1985 3817
rect 2023 3783 2057 3817
rect 2095 3783 2125 3817
rect 2125 3783 2129 3817
rect 2167 3783 2193 3817
rect 2193 3783 2201 3817
rect 2239 3783 2261 3817
rect 2261 3783 2273 3817
rect 2311 3783 2329 3817
rect 2329 3783 2345 3817
rect 2383 3783 2397 3817
rect 2397 3783 2417 3817
rect 2455 3783 2465 3817
rect 2465 3783 2489 3817
rect 2527 3783 2533 3817
rect 2533 3783 2561 3817
rect 2599 3783 2601 3817
rect 2601 3783 2633 3817
rect 2671 3783 2703 3817
rect 2703 3783 2705 3817
rect 2743 3783 2771 3817
rect 2771 3783 2777 3817
rect 2815 3783 2839 3817
rect 2839 3783 2849 3817
rect 2887 3783 2907 3817
rect 2907 3783 2921 3817
rect 2959 3783 2975 3817
rect 2975 3783 2993 3817
rect 3031 3783 3043 3817
rect 3043 3783 3065 3817
rect 3103 3783 3111 3817
rect 3111 3783 3137 3817
rect 3175 3783 3179 3817
rect 3179 3783 3209 3817
rect 3247 3783 3281 3817
rect 3319 3783 3349 3817
rect 3349 3783 3353 3817
rect 3391 3783 3417 3817
rect 3417 3783 3425 3817
rect 3463 3783 3485 3817
rect 3485 3783 3497 3817
rect 3535 3783 3553 3817
rect 3553 3783 3569 3817
rect 3607 3783 3621 3817
rect 3621 3783 3641 3817
rect 3679 3783 3689 3817
rect 3689 3783 3713 3817
rect 3751 3783 3757 3817
rect 3757 3783 3785 3817
rect 3823 3783 3825 3817
rect 3825 3783 3857 3817
rect 3895 3783 3927 3817
rect 3927 3783 3929 3817
rect 3967 3783 3995 3817
rect 3995 3783 4001 3817
rect -137 3623 -103 3657
rect 4183 3623 4217 3657
rect 79 3463 85 3497
rect 85 3463 113 3497
rect 151 3463 153 3497
rect 153 3463 185 3497
rect 223 3463 255 3497
rect 255 3463 257 3497
rect 295 3463 323 3497
rect 323 3463 329 3497
rect 367 3463 391 3497
rect 391 3463 401 3497
rect 439 3463 459 3497
rect 459 3463 473 3497
rect 511 3463 527 3497
rect 527 3463 545 3497
rect 583 3463 595 3497
rect 595 3463 617 3497
rect 655 3463 663 3497
rect 663 3463 689 3497
rect 727 3463 731 3497
rect 731 3463 761 3497
rect 799 3463 833 3497
rect 871 3463 901 3497
rect 901 3463 905 3497
rect 943 3463 969 3497
rect 969 3463 977 3497
rect 1015 3463 1037 3497
rect 1037 3463 1049 3497
rect 1087 3463 1105 3497
rect 1105 3463 1121 3497
rect 1159 3463 1173 3497
rect 1173 3463 1193 3497
rect 1231 3463 1241 3497
rect 1241 3463 1265 3497
rect 1303 3463 1309 3497
rect 1309 3463 1337 3497
rect 1375 3463 1377 3497
rect 1377 3463 1409 3497
rect 1447 3463 1479 3497
rect 1479 3463 1481 3497
rect 1519 3463 1547 3497
rect 1547 3463 1553 3497
rect 1591 3463 1615 3497
rect 1615 3463 1625 3497
rect 1663 3463 1683 3497
rect 1683 3463 1697 3497
rect 1735 3463 1751 3497
rect 1751 3463 1769 3497
rect 1807 3463 1819 3497
rect 1819 3463 1841 3497
rect 1879 3463 1887 3497
rect 1887 3463 1913 3497
rect 1951 3463 1955 3497
rect 1955 3463 1985 3497
rect 2023 3463 2057 3497
rect 2095 3463 2125 3497
rect 2125 3463 2129 3497
rect 2167 3463 2193 3497
rect 2193 3463 2201 3497
rect 2239 3463 2261 3497
rect 2261 3463 2273 3497
rect 2311 3463 2329 3497
rect 2329 3463 2345 3497
rect 2383 3463 2397 3497
rect 2397 3463 2417 3497
rect 2455 3463 2465 3497
rect 2465 3463 2489 3497
rect 2527 3463 2533 3497
rect 2533 3463 2561 3497
rect 2599 3463 2601 3497
rect 2601 3463 2633 3497
rect 2671 3463 2703 3497
rect 2703 3463 2705 3497
rect 2743 3463 2771 3497
rect 2771 3463 2777 3497
rect 2815 3463 2839 3497
rect 2839 3463 2849 3497
rect 2887 3463 2907 3497
rect 2907 3463 2921 3497
rect 2959 3463 2975 3497
rect 2975 3463 2993 3497
rect 3031 3463 3043 3497
rect 3043 3463 3065 3497
rect 3103 3463 3111 3497
rect 3111 3463 3137 3497
rect 3175 3463 3179 3497
rect 3179 3463 3209 3497
rect 3247 3463 3281 3497
rect 3319 3463 3349 3497
rect 3349 3463 3353 3497
rect 3391 3463 3417 3497
rect 3417 3463 3425 3497
rect 3463 3463 3485 3497
rect 3485 3463 3497 3497
rect 3535 3463 3553 3497
rect 3553 3463 3569 3497
rect 3607 3463 3621 3497
rect 3621 3463 3641 3497
rect 3679 3463 3689 3497
rect 3689 3463 3713 3497
rect 3751 3463 3757 3497
rect 3757 3463 3785 3497
rect 3823 3463 3825 3497
rect 3825 3463 3857 3497
rect 3895 3463 3927 3497
rect 3927 3463 3929 3497
rect 3967 3463 3995 3497
rect 3995 3463 4001 3497
rect 4183 2823 4199 2857
rect 4199 2823 4217 2857
rect 79 2663 85 2697
rect 85 2663 113 2697
rect 151 2663 153 2697
rect 153 2663 185 2697
rect 223 2663 255 2697
rect 255 2663 257 2697
rect 295 2663 323 2697
rect 323 2663 329 2697
rect 367 2663 391 2697
rect 391 2663 401 2697
rect 439 2663 459 2697
rect 459 2663 473 2697
rect 511 2663 527 2697
rect 527 2663 545 2697
rect 583 2663 595 2697
rect 595 2663 617 2697
rect 655 2663 663 2697
rect 663 2663 689 2697
rect 727 2663 731 2697
rect 731 2663 761 2697
rect 799 2663 833 2697
rect 871 2663 901 2697
rect 901 2663 905 2697
rect 943 2663 969 2697
rect 969 2663 977 2697
rect 1015 2663 1037 2697
rect 1037 2663 1049 2697
rect 1087 2663 1105 2697
rect 1105 2663 1121 2697
rect 1159 2663 1173 2697
rect 1173 2663 1193 2697
rect 1231 2663 1241 2697
rect 1241 2663 1265 2697
rect 1303 2663 1309 2697
rect 1309 2663 1337 2697
rect 1375 2663 1377 2697
rect 1377 2663 1409 2697
rect 1447 2663 1479 2697
rect 1479 2663 1481 2697
rect 1519 2663 1547 2697
rect 1547 2663 1553 2697
rect 1591 2663 1615 2697
rect 1615 2663 1625 2697
rect 1663 2663 1683 2697
rect 1683 2663 1697 2697
rect 1735 2663 1751 2697
rect 1751 2663 1769 2697
rect 1807 2663 1819 2697
rect 1819 2663 1841 2697
rect 1879 2663 1887 2697
rect 1887 2663 1913 2697
rect 1951 2663 1955 2697
rect 1955 2663 1985 2697
rect 2023 2663 2057 2697
rect 2095 2663 2125 2697
rect 2125 2663 2129 2697
rect 2167 2663 2193 2697
rect 2193 2663 2201 2697
rect 2239 2663 2261 2697
rect 2261 2663 2273 2697
rect 2311 2663 2329 2697
rect 2329 2663 2345 2697
rect 2383 2663 2397 2697
rect 2397 2663 2417 2697
rect 2455 2663 2465 2697
rect 2465 2663 2489 2697
rect 2527 2663 2533 2697
rect 2533 2663 2561 2697
rect 2599 2663 2601 2697
rect 2601 2663 2633 2697
rect 2671 2663 2703 2697
rect 2703 2663 2705 2697
rect 2743 2663 2771 2697
rect 2771 2663 2777 2697
rect 2815 2663 2839 2697
rect 2839 2663 2849 2697
rect 2887 2663 2907 2697
rect 2907 2663 2921 2697
rect 2959 2663 2975 2697
rect 2975 2663 2993 2697
rect 3031 2663 3043 2697
rect 3043 2663 3065 2697
rect 3103 2663 3111 2697
rect 3111 2663 3137 2697
rect 3175 2663 3179 2697
rect 3179 2663 3209 2697
rect 3247 2663 3281 2697
rect 3319 2663 3349 2697
rect 3349 2663 3353 2697
rect 3391 2663 3417 2697
rect 3417 2663 3425 2697
rect 3463 2663 3485 2697
rect 3485 2663 3497 2697
rect 3535 2663 3553 2697
rect 3553 2663 3569 2697
rect 3607 2663 3621 2697
rect 3621 2663 3641 2697
rect 3679 2663 3689 2697
rect 3689 2663 3713 2697
rect 3751 2663 3757 2697
rect 3757 2663 3785 2697
rect 3823 2663 3825 2697
rect 3825 2663 3857 2697
rect 3895 2663 3927 2697
rect 3927 2663 3929 2697
rect 3967 2663 3995 2697
rect 3995 2663 4001 2697
rect -137 2503 -103 2537
rect 4183 2503 4217 2537
rect 79 2343 85 2377
rect 85 2343 113 2377
rect 151 2343 153 2377
rect 153 2343 185 2377
rect 223 2343 255 2377
rect 255 2343 257 2377
rect 295 2343 323 2377
rect 323 2343 329 2377
rect 367 2343 391 2377
rect 391 2343 401 2377
rect 439 2343 459 2377
rect 459 2343 473 2377
rect 511 2343 527 2377
rect 527 2343 545 2377
rect 583 2343 595 2377
rect 595 2343 617 2377
rect 655 2343 663 2377
rect 663 2343 689 2377
rect 727 2343 731 2377
rect 731 2343 761 2377
rect 799 2343 833 2377
rect 871 2343 901 2377
rect 901 2343 905 2377
rect 943 2343 969 2377
rect 969 2343 977 2377
rect 1015 2343 1037 2377
rect 1037 2343 1049 2377
rect 1087 2343 1105 2377
rect 1105 2343 1121 2377
rect 1159 2343 1173 2377
rect 1173 2343 1193 2377
rect 1231 2343 1241 2377
rect 1241 2343 1265 2377
rect 1303 2343 1309 2377
rect 1309 2343 1337 2377
rect 1375 2343 1377 2377
rect 1377 2343 1409 2377
rect 1447 2343 1479 2377
rect 1479 2343 1481 2377
rect 1519 2343 1547 2377
rect 1547 2343 1553 2377
rect 1591 2343 1615 2377
rect 1615 2343 1625 2377
rect 1663 2343 1683 2377
rect 1683 2343 1697 2377
rect 1735 2343 1751 2377
rect 1751 2343 1769 2377
rect 1807 2343 1819 2377
rect 1819 2343 1841 2377
rect 1879 2343 1887 2377
rect 1887 2343 1913 2377
rect 1951 2343 1955 2377
rect 1955 2343 1985 2377
rect 2023 2343 2057 2377
rect 2095 2343 2125 2377
rect 2125 2343 2129 2377
rect 2167 2343 2193 2377
rect 2193 2343 2201 2377
rect 2239 2343 2261 2377
rect 2261 2343 2273 2377
rect 2311 2343 2329 2377
rect 2329 2343 2345 2377
rect 2383 2343 2397 2377
rect 2397 2343 2417 2377
rect 2455 2343 2465 2377
rect 2465 2343 2489 2377
rect 2527 2343 2533 2377
rect 2533 2343 2561 2377
rect 2599 2343 2601 2377
rect 2601 2343 2633 2377
rect 2671 2343 2703 2377
rect 2703 2343 2705 2377
rect 2743 2343 2771 2377
rect 2771 2343 2777 2377
rect 2815 2343 2839 2377
rect 2839 2343 2849 2377
rect 2887 2343 2907 2377
rect 2907 2343 2921 2377
rect 2959 2343 2975 2377
rect 2975 2343 2993 2377
rect 3031 2343 3043 2377
rect 3043 2343 3065 2377
rect 3103 2343 3111 2377
rect 3111 2343 3137 2377
rect 3175 2343 3179 2377
rect 3179 2343 3209 2377
rect 3247 2343 3281 2377
rect 3319 2343 3349 2377
rect 3349 2343 3353 2377
rect 3391 2343 3417 2377
rect 3417 2343 3425 2377
rect 3463 2343 3485 2377
rect 3485 2343 3497 2377
rect 3535 2343 3553 2377
rect 3553 2343 3569 2377
rect 3607 2343 3621 2377
rect 3621 2343 3641 2377
rect 3679 2343 3689 2377
rect 3689 2343 3713 2377
rect 3751 2343 3757 2377
rect 3757 2343 3785 2377
rect 3823 2343 3825 2377
rect 3825 2343 3857 2377
rect 3895 2343 3927 2377
rect 3927 2343 3929 2377
rect 3967 2343 3995 2377
rect 3995 2343 4001 2377
rect -137 2183 -103 2217
rect 4183 2183 4217 2217
rect -297 1783 -263 1817
rect -137 1383 -103 1417
rect 4183 1383 4217 1417
rect 79 1223 85 1257
rect 85 1223 113 1257
rect 151 1223 153 1257
rect 153 1223 185 1257
rect 223 1223 255 1257
rect 255 1223 257 1257
rect 295 1223 323 1257
rect 323 1223 329 1257
rect 367 1223 391 1257
rect 391 1223 401 1257
rect 439 1223 459 1257
rect 459 1223 473 1257
rect 511 1223 527 1257
rect 527 1223 545 1257
rect 583 1223 595 1257
rect 595 1223 617 1257
rect 655 1223 663 1257
rect 663 1223 689 1257
rect 727 1223 731 1257
rect 731 1223 761 1257
rect 799 1223 833 1257
rect 871 1223 901 1257
rect 901 1223 905 1257
rect 943 1223 969 1257
rect 969 1223 977 1257
rect 1015 1223 1037 1257
rect 1037 1223 1049 1257
rect 1087 1223 1105 1257
rect 1105 1223 1121 1257
rect 1159 1223 1173 1257
rect 1173 1223 1193 1257
rect 1231 1223 1241 1257
rect 1241 1223 1265 1257
rect 1303 1223 1309 1257
rect 1309 1223 1337 1257
rect 1375 1223 1377 1257
rect 1377 1223 1409 1257
rect 1447 1223 1479 1257
rect 1479 1223 1481 1257
rect 1519 1223 1547 1257
rect 1547 1223 1553 1257
rect 1591 1223 1615 1257
rect 1615 1223 1625 1257
rect 1663 1223 1683 1257
rect 1683 1223 1697 1257
rect 1735 1223 1751 1257
rect 1751 1223 1769 1257
rect 1807 1223 1819 1257
rect 1819 1223 1841 1257
rect 1879 1223 1887 1257
rect 1887 1223 1913 1257
rect 1951 1223 1955 1257
rect 1955 1223 1985 1257
rect 2023 1223 2057 1257
rect 2095 1223 2125 1257
rect 2125 1223 2129 1257
rect 2167 1223 2193 1257
rect 2193 1223 2201 1257
rect 2239 1223 2261 1257
rect 2261 1223 2273 1257
rect 2311 1223 2329 1257
rect 2329 1223 2345 1257
rect 2383 1223 2397 1257
rect 2397 1223 2417 1257
rect 2455 1223 2465 1257
rect 2465 1223 2489 1257
rect 2527 1223 2533 1257
rect 2533 1223 2561 1257
rect 2599 1223 2601 1257
rect 2601 1223 2633 1257
rect 2671 1223 2703 1257
rect 2703 1223 2705 1257
rect 2743 1223 2771 1257
rect 2771 1223 2777 1257
rect 2815 1223 2839 1257
rect 2839 1223 2849 1257
rect 2887 1223 2907 1257
rect 2907 1223 2921 1257
rect 2959 1223 2975 1257
rect 2975 1223 2993 1257
rect 3031 1223 3043 1257
rect 3043 1223 3065 1257
rect 3103 1223 3111 1257
rect 3111 1223 3137 1257
rect 3175 1223 3179 1257
rect 3179 1223 3209 1257
rect 3247 1223 3281 1257
rect 3319 1223 3349 1257
rect 3349 1223 3353 1257
rect 3391 1223 3417 1257
rect 3417 1223 3425 1257
rect 3463 1223 3485 1257
rect 3485 1223 3497 1257
rect 3535 1223 3553 1257
rect 3553 1223 3569 1257
rect 3607 1223 3621 1257
rect 3621 1223 3641 1257
rect 3679 1223 3689 1257
rect 3689 1223 3713 1257
rect 3751 1223 3757 1257
rect 3757 1223 3785 1257
rect 3823 1223 3825 1257
rect 3825 1223 3857 1257
rect 3895 1223 3927 1257
rect 3927 1223 3929 1257
rect 3967 1223 3995 1257
rect 3995 1223 4001 1257
rect -137 1063 -103 1097
rect 4183 1063 4217 1097
rect 79 903 85 937
rect 85 903 113 937
rect 151 903 153 937
rect 153 903 185 937
rect 223 903 255 937
rect 255 903 257 937
rect 295 903 323 937
rect 323 903 329 937
rect 367 903 391 937
rect 391 903 401 937
rect 439 903 459 937
rect 459 903 473 937
rect 511 903 527 937
rect 527 903 545 937
rect 583 903 595 937
rect 595 903 617 937
rect 655 903 663 937
rect 663 903 689 937
rect 727 903 731 937
rect 731 903 761 937
rect 799 903 833 937
rect 871 903 901 937
rect 901 903 905 937
rect 943 903 969 937
rect 969 903 977 937
rect 1015 903 1037 937
rect 1037 903 1049 937
rect 1087 903 1105 937
rect 1105 903 1121 937
rect 1159 903 1173 937
rect 1173 903 1193 937
rect 1231 903 1241 937
rect 1241 903 1265 937
rect 1303 903 1309 937
rect 1309 903 1337 937
rect 1375 903 1377 937
rect 1377 903 1409 937
rect 1447 903 1479 937
rect 1479 903 1481 937
rect 1519 903 1547 937
rect 1547 903 1553 937
rect 1591 903 1615 937
rect 1615 903 1625 937
rect 1663 903 1683 937
rect 1683 903 1697 937
rect 1735 903 1751 937
rect 1751 903 1769 937
rect 1807 903 1819 937
rect 1819 903 1841 937
rect 1879 903 1887 937
rect 1887 903 1913 937
rect 1951 903 1955 937
rect 1955 903 1985 937
rect 2023 903 2057 937
rect 2095 903 2125 937
rect 2125 903 2129 937
rect 2167 903 2193 937
rect 2193 903 2201 937
rect 2239 903 2261 937
rect 2261 903 2273 937
rect 2311 903 2329 937
rect 2329 903 2345 937
rect 2383 903 2397 937
rect 2397 903 2417 937
rect 2455 903 2465 937
rect 2465 903 2489 937
rect 2527 903 2533 937
rect 2533 903 2561 937
rect 2599 903 2601 937
rect 2601 903 2633 937
rect 2671 903 2703 937
rect 2703 903 2705 937
rect 2743 903 2771 937
rect 2771 903 2777 937
rect 2815 903 2839 937
rect 2839 903 2849 937
rect 2887 903 2907 937
rect 2907 903 2921 937
rect 2959 903 2975 937
rect 2975 903 2993 937
rect 3031 903 3043 937
rect 3043 903 3065 937
rect 3103 903 3111 937
rect 3111 903 3137 937
rect 3175 903 3179 937
rect 3179 903 3209 937
rect 3247 903 3281 937
rect 3319 903 3349 937
rect 3349 903 3353 937
rect 3391 903 3417 937
rect 3417 903 3425 937
rect 3463 903 3485 937
rect 3485 903 3497 937
rect 3535 903 3553 937
rect 3553 903 3569 937
rect 3607 903 3621 937
rect 3621 903 3641 937
rect 3679 903 3689 937
rect 3689 903 3713 937
rect 3751 903 3757 937
rect 3757 903 3785 937
rect 3823 903 3825 937
rect 3825 903 3857 937
rect 3895 903 3927 937
rect 3927 903 3929 937
rect 3967 903 3995 937
rect 3995 903 4001 937
rect 4183 743 4199 777
rect 4199 743 4217 777
rect 79 103 85 137
rect 85 103 113 137
rect 151 103 153 137
rect 153 103 185 137
rect 223 103 255 137
rect 255 103 257 137
rect 295 103 323 137
rect 323 103 329 137
rect 367 103 391 137
rect 391 103 401 137
rect 439 103 459 137
rect 459 103 473 137
rect 511 103 527 137
rect 527 103 545 137
rect 583 103 595 137
rect 595 103 617 137
rect 655 103 663 137
rect 663 103 689 137
rect 727 103 731 137
rect 731 103 761 137
rect 799 103 833 137
rect 871 103 901 137
rect 901 103 905 137
rect 943 103 969 137
rect 969 103 977 137
rect 1015 103 1037 137
rect 1037 103 1049 137
rect 1087 103 1105 137
rect 1105 103 1121 137
rect 1159 103 1173 137
rect 1173 103 1193 137
rect 1231 103 1241 137
rect 1241 103 1265 137
rect 1303 103 1309 137
rect 1309 103 1337 137
rect 1375 103 1377 137
rect 1377 103 1409 137
rect 1447 103 1479 137
rect 1479 103 1481 137
rect 1519 103 1547 137
rect 1547 103 1553 137
rect 1591 103 1615 137
rect 1615 103 1625 137
rect 1663 103 1683 137
rect 1683 103 1697 137
rect 1735 103 1751 137
rect 1751 103 1769 137
rect 1807 103 1819 137
rect 1819 103 1841 137
rect 1879 103 1887 137
rect 1887 103 1913 137
rect 1951 103 1955 137
rect 1955 103 1985 137
rect 2023 103 2057 137
rect 2095 103 2125 137
rect 2125 103 2129 137
rect 2167 103 2193 137
rect 2193 103 2201 137
rect 2239 103 2261 137
rect 2261 103 2273 137
rect 2311 103 2329 137
rect 2329 103 2345 137
rect 2383 103 2397 137
rect 2397 103 2417 137
rect 2455 103 2465 137
rect 2465 103 2489 137
rect 2527 103 2533 137
rect 2533 103 2561 137
rect 2599 103 2601 137
rect 2601 103 2633 137
rect 2671 103 2703 137
rect 2703 103 2705 137
rect 2743 103 2771 137
rect 2771 103 2777 137
rect 2815 103 2839 137
rect 2839 103 2849 137
rect 2887 103 2907 137
rect 2907 103 2921 137
rect 2959 103 2975 137
rect 2975 103 2993 137
rect 3031 103 3043 137
rect 3043 103 3065 137
rect 3103 103 3111 137
rect 3111 103 3137 137
rect 3175 103 3179 137
rect 3179 103 3209 137
rect 3247 103 3281 137
rect 3319 103 3349 137
rect 3349 103 3353 137
rect 3391 103 3417 137
rect 3417 103 3425 137
rect 3463 103 3485 137
rect 3485 103 3497 137
rect 3535 103 3553 137
rect 3553 103 3569 137
rect 3607 103 3621 137
rect 3621 103 3641 137
rect 3679 103 3689 137
rect 3689 103 3713 137
rect 3751 103 3757 137
rect 3757 103 3785 137
rect 3823 103 3825 137
rect 3825 103 3857 137
rect 3895 103 3927 137
rect 3927 103 3929 137
rect 3967 103 3995 137
rect 3995 103 4001 137
rect -137 -57 -103 -23
rect 4183 -57 4217 -23
rect 79 -217 85 -183
rect 85 -217 113 -183
rect 151 -217 153 -183
rect 153 -217 185 -183
rect 223 -217 255 -183
rect 255 -217 257 -183
rect 295 -217 323 -183
rect 323 -217 329 -183
rect 367 -217 391 -183
rect 391 -217 401 -183
rect 439 -217 459 -183
rect 459 -217 473 -183
rect 511 -217 527 -183
rect 527 -217 545 -183
rect 583 -217 595 -183
rect 595 -217 617 -183
rect 655 -217 663 -183
rect 663 -217 689 -183
rect 727 -217 731 -183
rect 731 -217 761 -183
rect 799 -217 833 -183
rect 871 -217 901 -183
rect 901 -217 905 -183
rect 943 -217 969 -183
rect 969 -217 977 -183
rect 1015 -217 1037 -183
rect 1037 -217 1049 -183
rect 1087 -217 1105 -183
rect 1105 -217 1121 -183
rect 1159 -217 1173 -183
rect 1173 -217 1193 -183
rect 1231 -217 1241 -183
rect 1241 -217 1265 -183
rect 1303 -217 1309 -183
rect 1309 -217 1337 -183
rect 1375 -217 1377 -183
rect 1377 -217 1409 -183
rect 1447 -217 1479 -183
rect 1479 -217 1481 -183
rect 1519 -217 1547 -183
rect 1547 -217 1553 -183
rect 1591 -217 1615 -183
rect 1615 -217 1625 -183
rect 1663 -217 1683 -183
rect 1683 -217 1697 -183
rect 1735 -217 1751 -183
rect 1751 -217 1769 -183
rect 1807 -217 1819 -183
rect 1819 -217 1841 -183
rect 1879 -217 1887 -183
rect 1887 -217 1913 -183
rect 1951 -217 1955 -183
rect 1955 -217 1985 -183
rect 2023 -217 2057 -183
rect 2095 -217 2125 -183
rect 2125 -217 2129 -183
rect 2167 -217 2193 -183
rect 2193 -217 2201 -183
rect 2239 -217 2261 -183
rect 2261 -217 2273 -183
rect 2311 -217 2329 -183
rect 2329 -217 2345 -183
rect 2383 -217 2397 -183
rect 2397 -217 2417 -183
rect 2455 -217 2465 -183
rect 2465 -217 2489 -183
rect 2527 -217 2533 -183
rect 2533 -217 2561 -183
rect 2599 -217 2601 -183
rect 2601 -217 2633 -183
rect 2671 -217 2703 -183
rect 2703 -217 2705 -183
rect 2743 -217 2771 -183
rect 2771 -217 2777 -183
rect 2815 -217 2839 -183
rect 2839 -217 2849 -183
rect 2887 -217 2907 -183
rect 2907 -217 2921 -183
rect 2959 -217 2975 -183
rect 2975 -217 2993 -183
rect 3031 -217 3043 -183
rect 3043 -217 3065 -183
rect 3103 -217 3111 -183
rect 3111 -217 3137 -183
rect 3175 -217 3179 -183
rect 3179 -217 3209 -183
rect 3247 -217 3281 -183
rect 3319 -217 3349 -183
rect 3349 -217 3353 -183
rect 3391 -217 3417 -183
rect 3417 -217 3425 -183
rect 3463 -217 3485 -183
rect 3485 -217 3497 -183
rect 3535 -217 3553 -183
rect 3553 -217 3569 -183
rect 3607 -217 3621 -183
rect 3621 -217 3641 -183
rect 3679 -217 3689 -183
rect 3689 -217 3713 -183
rect 3751 -217 3757 -183
rect 3757 -217 3785 -183
rect 3823 -217 3825 -183
rect 3825 -217 3857 -183
rect 3895 -217 3927 -183
rect 3927 -217 3929 -183
rect 3967 -217 3995 -183
rect 3995 -217 4001 -183
rect -137 -377 -103 -343
rect 4183 -377 4217 -343
rect -297 -537 -263 -503
rect 12823 4103 12857 4137
rect 8343 3943 8377 3977
rect 12663 3943 12697 3977
rect 8559 3783 8565 3817
rect 8565 3783 8593 3817
rect 8631 3783 8633 3817
rect 8633 3783 8665 3817
rect 8703 3783 8735 3817
rect 8735 3783 8737 3817
rect 8775 3783 8803 3817
rect 8803 3783 8809 3817
rect 8847 3783 8871 3817
rect 8871 3783 8881 3817
rect 8919 3783 8939 3817
rect 8939 3783 8953 3817
rect 8991 3783 9007 3817
rect 9007 3783 9025 3817
rect 9063 3783 9075 3817
rect 9075 3783 9097 3817
rect 9135 3783 9143 3817
rect 9143 3783 9169 3817
rect 9207 3783 9211 3817
rect 9211 3783 9241 3817
rect 9279 3783 9313 3817
rect 9351 3783 9381 3817
rect 9381 3783 9385 3817
rect 9423 3783 9449 3817
rect 9449 3783 9457 3817
rect 9495 3783 9517 3817
rect 9517 3783 9529 3817
rect 9567 3783 9585 3817
rect 9585 3783 9601 3817
rect 9639 3783 9653 3817
rect 9653 3783 9673 3817
rect 9711 3783 9721 3817
rect 9721 3783 9745 3817
rect 9783 3783 9789 3817
rect 9789 3783 9817 3817
rect 9855 3783 9857 3817
rect 9857 3783 9889 3817
rect 9927 3783 9959 3817
rect 9959 3783 9961 3817
rect 9999 3783 10027 3817
rect 10027 3783 10033 3817
rect 10071 3783 10095 3817
rect 10095 3783 10105 3817
rect 10143 3783 10163 3817
rect 10163 3783 10177 3817
rect 10215 3783 10231 3817
rect 10231 3783 10249 3817
rect 10287 3783 10299 3817
rect 10299 3783 10321 3817
rect 10359 3783 10367 3817
rect 10367 3783 10393 3817
rect 10431 3783 10435 3817
rect 10435 3783 10465 3817
rect 10503 3783 10537 3817
rect 10575 3783 10605 3817
rect 10605 3783 10609 3817
rect 10647 3783 10673 3817
rect 10673 3783 10681 3817
rect 10719 3783 10741 3817
rect 10741 3783 10753 3817
rect 10791 3783 10809 3817
rect 10809 3783 10825 3817
rect 10863 3783 10877 3817
rect 10877 3783 10897 3817
rect 10935 3783 10945 3817
rect 10945 3783 10969 3817
rect 11007 3783 11013 3817
rect 11013 3783 11041 3817
rect 11079 3783 11081 3817
rect 11081 3783 11113 3817
rect 11151 3783 11183 3817
rect 11183 3783 11185 3817
rect 11223 3783 11251 3817
rect 11251 3783 11257 3817
rect 11295 3783 11319 3817
rect 11319 3783 11329 3817
rect 11367 3783 11387 3817
rect 11387 3783 11401 3817
rect 11439 3783 11455 3817
rect 11455 3783 11473 3817
rect 11511 3783 11523 3817
rect 11523 3783 11545 3817
rect 11583 3783 11591 3817
rect 11591 3783 11617 3817
rect 11655 3783 11659 3817
rect 11659 3783 11689 3817
rect 11727 3783 11761 3817
rect 11799 3783 11829 3817
rect 11829 3783 11833 3817
rect 11871 3783 11897 3817
rect 11897 3783 11905 3817
rect 11943 3783 11965 3817
rect 11965 3783 11977 3817
rect 12015 3783 12033 3817
rect 12033 3783 12049 3817
rect 12087 3783 12101 3817
rect 12101 3783 12121 3817
rect 12159 3783 12169 3817
rect 12169 3783 12193 3817
rect 12231 3783 12237 3817
rect 12237 3783 12265 3817
rect 12303 3783 12305 3817
rect 12305 3783 12337 3817
rect 12375 3783 12407 3817
rect 12407 3783 12409 3817
rect 12447 3783 12475 3817
rect 12475 3783 12481 3817
rect 8343 3623 8377 3657
rect 12663 3623 12697 3657
rect 8559 3463 8565 3497
rect 8565 3463 8593 3497
rect 8631 3463 8633 3497
rect 8633 3463 8665 3497
rect 8703 3463 8735 3497
rect 8735 3463 8737 3497
rect 8775 3463 8803 3497
rect 8803 3463 8809 3497
rect 8847 3463 8871 3497
rect 8871 3463 8881 3497
rect 8919 3463 8939 3497
rect 8939 3463 8953 3497
rect 8991 3463 9007 3497
rect 9007 3463 9025 3497
rect 9063 3463 9075 3497
rect 9075 3463 9097 3497
rect 9135 3463 9143 3497
rect 9143 3463 9169 3497
rect 9207 3463 9211 3497
rect 9211 3463 9241 3497
rect 9279 3463 9313 3497
rect 9351 3463 9381 3497
rect 9381 3463 9385 3497
rect 9423 3463 9449 3497
rect 9449 3463 9457 3497
rect 9495 3463 9517 3497
rect 9517 3463 9529 3497
rect 9567 3463 9585 3497
rect 9585 3463 9601 3497
rect 9639 3463 9653 3497
rect 9653 3463 9673 3497
rect 9711 3463 9721 3497
rect 9721 3463 9745 3497
rect 9783 3463 9789 3497
rect 9789 3463 9817 3497
rect 9855 3463 9857 3497
rect 9857 3463 9889 3497
rect 9927 3463 9959 3497
rect 9959 3463 9961 3497
rect 9999 3463 10027 3497
rect 10027 3463 10033 3497
rect 10071 3463 10095 3497
rect 10095 3463 10105 3497
rect 10143 3463 10163 3497
rect 10163 3463 10177 3497
rect 10215 3463 10231 3497
rect 10231 3463 10249 3497
rect 10287 3463 10299 3497
rect 10299 3463 10321 3497
rect 10359 3463 10367 3497
rect 10367 3463 10393 3497
rect 10431 3463 10435 3497
rect 10435 3463 10465 3497
rect 10503 3463 10537 3497
rect 10575 3463 10605 3497
rect 10605 3463 10609 3497
rect 10647 3463 10673 3497
rect 10673 3463 10681 3497
rect 10719 3463 10741 3497
rect 10741 3463 10753 3497
rect 10791 3463 10809 3497
rect 10809 3463 10825 3497
rect 10863 3463 10877 3497
rect 10877 3463 10897 3497
rect 10935 3463 10945 3497
rect 10945 3463 10969 3497
rect 11007 3463 11013 3497
rect 11013 3463 11041 3497
rect 11079 3463 11081 3497
rect 11081 3463 11113 3497
rect 11151 3463 11183 3497
rect 11183 3463 11185 3497
rect 11223 3463 11251 3497
rect 11251 3463 11257 3497
rect 11295 3463 11319 3497
rect 11319 3463 11329 3497
rect 11367 3463 11387 3497
rect 11387 3463 11401 3497
rect 11439 3463 11455 3497
rect 11455 3463 11473 3497
rect 11511 3463 11523 3497
rect 11523 3463 11545 3497
rect 11583 3463 11591 3497
rect 11591 3463 11617 3497
rect 11655 3463 11659 3497
rect 11659 3463 11689 3497
rect 11727 3463 11761 3497
rect 11799 3463 11829 3497
rect 11829 3463 11833 3497
rect 11871 3463 11897 3497
rect 11897 3463 11905 3497
rect 11943 3463 11965 3497
rect 11965 3463 11977 3497
rect 12015 3463 12033 3497
rect 12033 3463 12049 3497
rect 12087 3463 12101 3497
rect 12101 3463 12121 3497
rect 12159 3463 12169 3497
rect 12169 3463 12193 3497
rect 12231 3463 12237 3497
rect 12237 3463 12265 3497
rect 12303 3463 12305 3497
rect 12305 3463 12337 3497
rect 12375 3463 12407 3497
rect 12407 3463 12409 3497
rect 12447 3463 12475 3497
rect 12475 3463 12481 3497
rect 8343 2823 8361 2857
rect 8361 2823 8377 2857
rect 8559 2663 8565 2697
rect 8565 2663 8593 2697
rect 8631 2663 8633 2697
rect 8633 2663 8665 2697
rect 8703 2663 8735 2697
rect 8735 2663 8737 2697
rect 8775 2663 8803 2697
rect 8803 2663 8809 2697
rect 8847 2663 8871 2697
rect 8871 2663 8881 2697
rect 8919 2663 8939 2697
rect 8939 2663 8953 2697
rect 8991 2663 9007 2697
rect 9007 2663 9025 2697
rect 9063 2663 9075 2697
rect 9075 2663 9097 2697
rect 9135 2663 9143 2697
rect 9143 2663 9169 2697
rect 9207 2663 9211 2697
rect 9211 2663 9241 2697
rect 9279 2663 9313 2697
rect 9351 2663 9381 2697
rect 9381 2663 9385 2697
rect 9423 2663 9449 2697
rect 9449 2663 9457 2697
rect 9495 2663 9517 2697
rect 9517 2663 9529 2697
rect 9567 2663 9585 2697
rect 9585 2663 9601 2697
rect 9639 2663 9653 2697
rect 9653 2663 9673 2697
rect 9711 2663 9721 2697
rect 9721 2663 9745 2697
rect 9783 2663 9789 2697
rect 9789 2663 9817 2697
rect 9855 2663 9857 2697
rect 9857 2663 9889 2697
rect 9927 2663 9959 2697
rect 9959 2663 9961 2697
rect 9999 2663 10027 2697
rect 10027 2663 10033 2697
rect 10071 2663 10095 2697
rect 10095 2663 10105 2697
rect 10143 2663 10163 2697
rect 10163 2663 10177 2697
rect 10215 2663 10231 2697
rect 10231 2663 10249 2697
rect 10287 2663 10299 2697
rect 10299 2663 10321 2697
rect 10359 2663 10367 2697
rect 10367 2663 10393 2697
rect 10431 2663 10435 2697
rect 10435 2663 10465 2697
rect 10503 2663 10537 2697
rect 10575 2663 10605 2697
rect 10605 2663 10609 2697
rect 10647 2663 10673 2697
rect 10673 2663 10681 2697
rect 10719 2663 10741 2697
rect 10741 2663 10753 2697
rect 10791 2663 10809 2697
rect 10809 2663 10825 2697
rect 10863 2663 10877 2697
rect 10877 2663 10897 2697
rect 10935 2663 10945 2697
rect 10945 2663 10969 2697
rect 11007 2663 11013 2697
rect 11013 2663 11041 2697
rect 11079 2663 11081 2697
rect 11081 2663 11113 2697
rect 11151 2663 11183 2697
rect 11183 2663 11185 2697
rect 11223 2663 11251 2697
rect 11251 2663 11257 2697
rect 11295 2663 11319 2697
rect 11319 2663 11329 2697
rect 11367 2663 11387 2697
rect 11387 2663 11401 2697
rect 11439 2663 11455 2697
rect 11455 2663 11473 2697
rect 11511 2663 11523 2697
rect 11523 2663 11545 2697
rect 11583 2663 11591 2697
rect 11591 2663 11617 2697
rect 11655 2663 11659 2697
rect 11659 2663 11689 2697
rect 11727 2663 11761 2697
rect 11799 2663 11829 2697
rect 11829 2663 11833 2697
rect 11871 2663 11897 2697
rect 11897 2663 11905 2697
rect 11943 2663 11965 2697
rect 11965 2663 11977 2697
rect 12015 2663 12033 2697
rect 12033 2663 12049 2697
rect 12087 2663 12101 2697
rect 12101 2663 12121 2697
rect 12159 2663 12169 2697
rect 12169 2663 12193 2697
rect 12231 2663 12237 2697
rect 12237 2663 12265 2697
rect 12303 2663 12305 2697
rect 12305 2663 12337 2697
rect 12375 2663 12407 2697
rect 12407 2663 12409 2697
rect 12447 2663 12475 2697
rect 12475 2663 12481 2697
rect 8343 2503 8377 2537
rect 12663 2503 12697 2537
rect 8559 2343 8565 2377
rect 8565 2343 8593 2377
rect 8631 2343 8633 2377
rect 8633 2343 8665 2377
rect 8703 2343 8735 2377
rect 8735 2343 8737 2377
rect 8775 2343 8803 2377
rect 8803 2343 8809 2377
rect 8847 2343 8871 2377
rect 8871 2343 8881 2377
rect 8919 2343 8939 2377
rect 8939 2343 8953 2377
rect 8991 2343 9007 2377
rect 9007 2343 9025 2377
rect 9063 2343 9075 2377
rect 9075 2343 9097 2377
rect 9135 2343 9143 2377
rect 9143 2343 9169 2377
rect 9207 2343 9211 2377
rect 9211 2343 9241 2377
rect 9279 2343 9313 2377
rect 9351 2343 9381 2377
rect 9381 2343 9385 2377
rect 9423 2343 9449 2377
rect 9449 2343 9457 2377
rect 9495 2343 9517 2377
rect 9517 2343 9529 2377
rect 9567 2343 9585 2377
rect 9585 2343 9601 2377
rect 9639 2343 9653 2377
rect 9653 2343 9673 2377
rect 9711 2343 9721 2377
rect 9721 2343 9745 2377
rect 9783 2343 9789 2377
rect 9789 2343 9817 2377
rect 9855 2343 9857 2377
rect 9857 2343 9889 2377
rect 9927 2343 9959 2377
rect 9959 2343 9961 2377
rect 9999 2343 10027 2377
rect 10027 2343 10033 2377
rect 10071 2343 10095 2377
rect 10095 2343 10105 2377
rect 10143 2343 10163 2377
rect 10163 2343 10177 2377
rect 10215 2343 10231 2377
rect 10231 2343 10249 2377
rect 10287 2343 10299 2377
rect 10299 2343 10321 2377
rect 10359 2343 10367 2377
rect 10367 2343 10393 2377
rect 10431 2343 10435 2377
rect 10435 2343 10465 2377
rect 10503 2343 10537 2377
rect 10575 2343 10605 2377
rect 10605 2343 10609 2377
rect 10647 2343 10673 2377
rect 10673 2343 10681 2377
rect 10719 2343 10741 2377
rect 10741 2343 10753 2377
rect 10791 2343 10809 2377
rect 10809 2343 10825 2377
rect 10863 2343 10877 2377
rect 10877 2343 10897 2377
rect 10935 2343 10945 2377
rect 10945 2343 10969 2377
rect 11007 2343 11013 2377
rect 11013 2343 11041 2377
rect 11079 2343 11081 2377
rect 11081 2343 11113 2377
rect 11151 2343 11183 2377
rect 11183 2343 11185 2377
rect 11223 2343 11251 2377
rect 11251 2343 11257 2377
rect 11295 2343 11319 2377
rect 11319 2343 11329 2377
rect 11367 2343 11387 2377
rect 11387 2343 11401 2377
rect 11439 2343 11455 2377
rect 11455 2343 11473 2377
rect 11511 2343 11523 2377
rect 11523 2343 11545 2377
rect 11583 2343 11591 2377
rect 11591 2343 11617 2377
rect 11655 2343 11659 2377
rect 11659 2343 11689 2377
rect 11727 2343 11761 2377
rect 11799 2343 11829 2377
rect 11829 2343 11833 2377
rect 11871 2343 11897 2377
rect 11897 2343 11905 2377
rect 11943 2343 11965 2377
rect 11965 2343 11977 2377
rect 12015 2343 12033 2377
rect 12033 2343 12049 2377
rect 12087 2343 12101 2377
rect 12101 2343 12121 2377
rect 12159 2343 12169 2377
rect 12169 2343 12193 2377
rect 12231 2343 12237 2377
rect 12237 2343 12265 2377
rect 12303 2343 12305 2377
rect 12305 2343 12337 2377
rect 12375 2343 12407 2377
rect 12407 2343 12409 2377
rect 12447 2343 12475 2377
rect 12475 2343 12481 2377
rect 8343 2183 8377 2217
rect 12663 2183 12697 2217
rect 12823 1783 12857 1817
rect 8343 1383 8377 1417
rect 12663 1383 12697 1417
rect 8559 1223 8565 1257
rect 8565 1223 8593 1257
rect 8631 1223 8633 1257
rect 8633 1223 8665 1257
rect 8703 1223 8735 1257
rect 8735 1223 8737 1257
rect 8775 1223 8803 1257
rect 8803 1223 8809 1257
rect 8847 1223 8871 1257
rect 8871 1223 8881 1257
rect 8919 1223 8939 1257
rect 8939 1223 8953 1257
rect 8991 1223 9007 1257
rect 9007 1223 9025 1257
rect 9063 1223 9075 1257
rect 9075 1223 9097 1257
rect 9135 1223 9143 1257
rect 9143 1223 9169 1257
rect 9207 1223 9211 1257
rect 9211 1223 9241 1257
rect 9279 1223 9313 1257
rect 9351 1223 9381 1257
rect 9381 1223 9385 1257
rect 9423 1223 9449 1257
rect 9449 1223 9457 1257
rect 9495 1223 9517 1257
rect 9517 1223 9529 1257
rect 9567 1223 9585 1257
rect 9585 1223 9601 1257
rect 9639 1223 9653 1257
rect 9653 1223 9673 1257
rect 9711 1223 9721 1257
rect 9721 1223 9745 1257
rect 9783 1223 9789 1257
rect 9789 1223 9817 1257
rect 9855 1223 9857 1257
rect 9857 1223 9889 1257
rect 9927 1223 9959 1257
rect 9959 1223 9961 1257
rect 9999 1223 10027 1257
rect 10027 1223 10033 1257
rect 10071 1223 10095 1257
rect 10095 1223 10105 1257
rect 10143 1223 10163 1257
rect 10163 1223 10177 1257
rect 10215 1223 10231 1257
rect 10231 1223 10249 1257
rect 10287 1223 10299 1257
rect 10299 1223 10321 1257
rect 10359 1223 10367 1257
rect 10367 1223 10393 1257
rect 10431 1223 10435 1257
rect 10435 1223 10465 1257
rect 10503 1223 10537 1257
rect 10575 1223 10605 1257
rect 10605 1223 10609 1257
rect 10647 1223 10673 1257
rect 10673 1223 10681 1257
rect 10719 1223 10741 1257
rect 10741 1223 10753 1257
rect 10791 1223 10809 1257
rect 10809 1223 10825 1257
rect 10863 1223 10877 1257
rect 10877 1223 10897 1257
rect 10935 1223 10945 1257
rect 10945 1223 10969 1257
rect 11007 1223 11013 1257
rect 11013 1223 11041 1257
rect 11079 1223 11081 1257
rect 11081 1223 11113 1257
rect 11151 1223 11183 1257
rect 11183 1223 11185 1257
rect 11223 1223 11251 1257
rect 11251 1223 11257 1257
rect 11295 1223 11319 1257
rect 11319 1223 11329 1257
rect 11367 1223 11387 1257
rect 11387 1223 11401 1257
rect 11439 1223 11455 1257
rect 11455 1223 11473 1257
rect 11511 1223 11523 1257
rect 11523 1223 11545 1257
rect 11583 1223 11591 1257
rect 11591 1223 11617 1257
rect 11655 1223 11659 1257
rect 11659 1223 11689 1257
rect 11727 1223 11761 1257
rect 11799 1223 11829 1257
rect 11829 1223 11833 1257
rect 11871 1223 11897 1257
rect 11897 1223 11905 1257
rect 11943 1223 11965 1257
rect 11965 1223 11977 1257
rect 12015 1223 12033 1257
rect 12033 1223 12049 1257
rect 12087 1223 12101 1257
rect 12101 1223 12121 1257
rect 12159 1223 12169 1257
rect 12169 1223 12193 1257
rect 12231 1223 12237 1257
rect 12237 1223 12265 1257
rect 12303 1223 12305 1257
rect 12305 1223 12337 1257
rect 12375 1223 12407 1257
rect 12407 1223 12409 1257
rect 12447 1223 12475 1257
rect 12475 1223 12481 1257
rect 8343 1063 8377 1097
rect 12663 1063 12697 1097
rect 8559 903 8565 937
rect 8565 903 8593 937
rect 8631 903 8633 937
rect 8633 903 8665 937
rect 8703 903 8735 937
rect 8735 903 8737 937
rect 8775 903 8803 937
rect 8803 903 8809 937
rect 8847 903 8871 937
rect 8871 903 8881 937
rect 8919 903 8939 937
rect 8939 903 8953 937
rect 8991 903 9007 937
rect 9007 903 9025 937
rect 9063 903 9075 937
rect 9075 903 9097 937
rect 9135 903 9143 937
rect 9143 903 9169 937
rect 9207 903 9211 937
rect 9211 903 9241 937
rect 9279 903 9313 937
rect 9351 903 9381 937
rect 9381 903 9385 937
rect 9423 903 9449 937
rect 9449 903 9457 937
rect 9495 903 9517 937
rect 9517 903 9529 937
rect 9567 903 9585 937
rect 9585 903 9601 937
rect 9639 903 9653 937
rect 9653 903 9673 937
rect 9711 903 9721 937
rect 9721 903 9745 937
rect 9783 903 9789 937
rect 9789 903 9817 937
rect 9855 903 9857 937
rect 9857 903 9889 937
rect 9927 903 9959 937
rect 9959 903 9961 937
rect 9999 903 10027 937
rect 10027 903 10033 937
rect 10071 903 10095 937
rect 10095 903 10105 937
rect 10143 903 10163 937
rect 10163 903 10177 937
rect 10215 903 10231 937
rect 10231 903 10249 937
rect 10287 903 10299 937
rect 10299 903 10321 937
rect 10359 903 10367 937
rect 10367 903 10393 937
rect 10431 903 10435 937
rect 10435 903 10465 937
rect 10503 903 10537 937
rect 10575 903 10605 937
rect 10605 903 10609 937
rect 10647 903 10673 937
rect 10673 903 10681 937
rect 10719 903 10741 937
rect 10741 903 10753 937
rect 10791 903 10809 937
rect 10809 903 10825 937
rect 10863 903 10877 937
rect 10877 903 10897 937
rect 10935 903 10945 937
rect 10945 903 10969 937
rect 11007 903 11013 937
rect 11013 903 11041 937
rect 11079 903 11081 937
rect 11081 903 11113 937
rect 11151 903 11183 937
rect 11183 903 11185 937
rect 11223 903 11251 937
rect 11251 903 11257 937
rect 11295 903 11319 937
rect 11319 903 11329 937
rect 11367 903 11387 937
rect 11387 903 11401 937
rect 11439 903 11455 937
rect 11455 903 11473 937
rect 11511 903 11523 937
rect 11523 903 11545 937
rect 11583 903 11591 937
rect 11591 903 11617 937
rect 11655 903 11659 937
rect 11659 903 11689 937
rect 11727 903 11761 937
rect 11799 903 11829 937
rect 11829 903 11833 937
rect 11871 903 11897 937
rect 11897 903 11905 937
rect 11943 903 11965 937
rect 11965 903 11977 937
rect 12015 903 12033 937
rect 12033 903 12049 937
rect 12087 903 12101 937
rect 12101 903 12121 937
rect 12159 903 12169 937
rect 12169 903 12193 937
rect 12231 903 12237 937
rect 12237 903 12265 937
rect 12303 903 12305 937
rect 12305 903 12337 937
rect 12375 903 12407 937
rect 12407 903 12409 937
rect 12447 903 12475 937
rect 12475 903 12481 937
rect 8343 743 8361 777
rect 8361 743 8377 777
rect 8559 103 8565 137
rect 8565 103 8593 137
rect 8631 103 8633 137
rect 8633 103 8665 137
rect 8703 103 8735 137
rect 8735 103 8737 137
rect 8775 103 8803 137
rect 8803 103 8809 137
rect 8847 103 8871 137
rect 8871 103 8881 137
rect 8919 103 8939 137
rect 8939 103 8953 137
rect 8991 103 9007 137
rect 9007 103 9025 137
rect 9063 103 9075 137
rect 9075 103 9097 137
rect 9135 103 9143 137
rect 9143 103 9169 137
rect 9207 103 9211 137
rect 9211 103 9241 137
rect 9279 103 9313 137
rect 9351 103 9381 137
rect 9381 103 9385 137
rect 9423 103 9449 137
rect 9449 103 9457 137
rect 9495 103 9517 137
rect 9517 103 9529 137
rect 9567 103 9585 137
rect 9585 103 9601 137
rect 9639 103 9653 137
rect 9653 103 9673 137
rect 9711 103 9721 137
rect 9721 103 9745 137
rect 9783 103 9789 137
rect 9789 103 9817 137
rect 9855 103 9857 137
rect 9857 103 9889 137
rect 9927 103 9959 137
rect 9959 103 9961 137
rect 9999 103 10027 137
rect 10027 103 10033 137
rect 10071 103 10095 137
rect 10095 103 10105 137
rect 10143 103 10163 137
rect 10163 103 10177 137
rect 10215 103 10231 137
rect 10231 103 10249 137
rect 10287 103 10299 137
rect 10299 103 10321 137
rect 10359 103 10367 137
rect 10367 103 10393 137
rect 10431 103 10435 137
rect 10435 103 10465 137
rect 10503 103 10537 137
rect 10575 103 10605 137
rect 10605 103 10609 137
rect 10647 103 10673 137
rect 10673 103 10681 137
rect 10719 103 10741 137
rect 10741 103 10753 137
rect 10791 103 10809 137
rect 10809 103 10825 137
rect 10863 103 10877 137
rect 10877 103 10897 137
rect 10935 103 10945 137
rect 10945 103 10969 137
rect 11007 103 11013 137
rect 11013 103 11041 137
rect 11079 103 11081 137
rect 11081 103 11113 137
rect 11151 103 11183 137
rect 11183 103 11185 137
rect 11223 103 11251 137
rect 11251 103 11257 137
rect 11295 103 11319 137
rect 11319 103 11329 137
rect 11367 103 11387 137
rect 11387 103 11401 137
rect 11439 103 11455 137
rect 11455 103 11473 137
rect 11511 103 11523 137
rect 11523 103 11545 137
rect 11583 103 11591 137
rect 11591 103 11617 137
rect 11655 103 11659 137
rect 11659 103 11689 137
rect 11727 103 11761 137
rect 11799 103 11829 137
rect 11829 103 11833 137
rect 11871 103 11897 137
rect 11897 103 11905 137
rect 11943 103 11965 137
rect 11965 103 11977 137
rect 12015 103 12033 137
rect 12033 103 12049 137
rect 12087 103 12101 137
rect 12101 103 12121 137
rect 12159 103 12169 137
rect 12169 103 12193 137
rect 12231 103 12237 137
rect 12237 103 12265 137
rect 12303 103 12305 137
rect 12305 103 12337 137
rect 12375 103 12407 137
rect 12407 103 12409 137
rect 12447 103 12475 137
rect 12475 103 12481 137
rect 8343 -57 8377 -23
rect 12663 -57 12697 -23
rect 8559 -217 8565 -183
rect 8565 -217 8593 -183
rect 8631 -217 8633 -183
rect 8633 -217 8665 -183
rect 8703 -217 8735 -183
rect 8735 -217 8737 -183
rect 8775 -217 8803 -183
rect 8803 -217 8809 -183
rect 8847 -217 8871 -183
rect 8871 -217 8881 -183
rect 8919 -217 8939 -183
rect 8939 -217 8953 -183
rect 8991 -217 9007 -183
rect 9007 -217 9025 -183
rect 9063 -217 9075 -183
rect 9075 -217 9097 -183
rect 9135 -217 9143 -183
rect 9143 -217 9169 -183
rect 9207 -217 9211 -183
rect 9211 -217 9241 -183
rect 9279 -217 9313 -183
rect 9351 -217 9381 -183
rect 9381 -217 9385 -183
rect 9423 -217 9449 -183
rect 9449 -217 9457 -183
rect 9495 -217 9517 -183
rect 9517 -217 9529 -183
rect 9567 -217 9585 -183
rect 9585 -217 9601 -183
rect 9639 -217 9653 -183
rect 9653 -217 9673 -183
rect 9711 -217 9721 -183
rect 9721 -217 9745 -183
rect 9783 -217 9789 -183
rect 9789 -217 9817 -183
rect 9855 -217 9857 -183
rect 9857 -217 9889 -183
rect 9927 -217 9959 -183
rect 9959 -217 9961 -183
rect 9999 -217 10027 -183
rect 10027 -217 10033 -183
rect 10071 -217 10095 -183
rect 10095 -217 10105 -183
rect 10143 -217 10163 -183
rect 10163 -217 10177 -183
rect 10215 -217 10231 -183
rect 10231 -217 10249 -183
rect 10287 -217 10299 -183
rect 10299 -217 10321 -183
rect 10359 -217 10367 -183
rect 10367 -217 10393 -183
rect 10431 -217 10435 -183
rect 10435 -217 10465 -183
rect 10503 -217 10537 -183
rect 10575 -217 10605 -183
rect 10605 -217 10609 -183
rect 10647 -217 10673 -183
rect 10673 -217 10681 -183
rect 10719 -217 10741 -183
rect 10741 -217 10753 -183
rect 10791 -217 10809 -183
rect 10809 -217 10825 -183
rect 10863 -217 10877 -183
rect 10877 -217 10897 -183
rect 10935 -217 10945 -183
rect 10945 -217 10969 -183
rect 11007 -217 11013 -183
rect 11013 -217 11041 -183
rect 11079 -217 11081 -183
rect 11081 -217 11113 -183
rect 11151 -217 11183 -183
rect 11183 -217 11185 -183
rect 11223 -217 11251 -183
rect 11251 -217 11257 -183
rect 11295 -217 11319 -183
rect 11319 -217 11329 -183
rect 11367 -217 11387 -183
rect 11387 -217 11401 -183
rect 11439 -217 11455 -183
rect 11455 -217 11473 -183
rect 11511 -217 11523 -183
rect 11523 -217 11545 -183
rect 11583 -217 11591 -183
rect 11591 -217 11617 -183
rect 11655 -217 11659 -183
rect 11659 -217 11689 -183
rect 11727 -217 11761 -183
rect 11799 -217 11829 -183
rect 11829 -217 11833 -183
rect 11871 -217 11897 -183
rect 11897 -217 11905 -183
rect 11943 -217 11965 -183
rect 11965 -217 11977 -183
rect 12015 -217 12033 -183
rect 12033 -217 12049 -183
rect 12087 -217 12101 -183
rect 12101 -217 12121 -183
rect 12159 -217 12169 -183
rect 12169 -217 12193 -183
rect 12231 -217 12237 -183
rect 12237 -217 12265 -183
rect 12303 -217 12305 -183
rect 12305 -217 12337 -183
rect 12375 -217 12407 -183
rect 12407 -217 12409 -183
rect 12447 -217 12475 -183
rect 12475 -217 12481 -183
rect 8343 -377 8377 -343
rect 12663 -377 12697 -343
rect 12823 -537 12857 -503
<< metal1 >>
rect -320 4146 -240 4160
rect -320 4094 -306 4146
rect -254 4094 -240 4146
rect -320 4080 -240 4094
rect 12800 4146 12880 4160
rect 12800 4094 12814 4146
rect 12866 4094 12880 4146
rect 12800 4080 12880 4094
rect -160 3977 -80 4000
rect -160 3943 -137 3977
rect -103 3943 -80 3977
rect -160 3657 -80 3943
rect 4160 3977 4240 4000
rect 4160 3943 4183 3977
rect 4217 3943 4240 3977
rect 40 3826 4040 3840
rect 40 3774 62 3826
rect 114 3774 126 3826
rect 178 3817 190 3826
rect 242 3817 254 3826
rect 306 3817 318 3826
rect 370 3817 382 3826
rect 434 3817 446 3826
rect 185 3783 190 3817
rect 434 3783 439 3817
rect 178 3774 190 3783
rect 242 3774 254 3783
rect 306 3774 318 3783
rect 370 3774 382 3783
rect 434 3774 446 3783
rect 498 3774 510 3826
rect 562 3774 574 3826
rect 626 3774 638 3826
rect 690 3774 702 3826
rect 754 3817 766 3826
rect 818 3817 830 3826
rect 882 3817 894 3826
rect 946 3817 958 3826
rect 1010 3817 1022 3826
rect 761 3783 766 3817
rect 1010 3783 1015 3817
rect 754 3774 766 3783
rect 818 3774 830 3783
rect 882 3774 894 3783
rect 946 3774 958 3783
rect 1010 3774 1022 3783
rect 1074 3774 1086 3826
rect 1138 3774 1150 3826
rect 1202 3774 1214 3826
rect 1266 3774 1278 3826
rect 1330 3817 1342 3826
rect 1394 3817 1406 3826
rect 1458 3817 1470 3826
rect 1522 3817 1534 3826
rect 1586 3817 1598 3826
rect 1337 3783 1342 3817
rect 1586 3783 1591 3817
rect 1330 3774 1342 3783
rect 1394 3774 1406 3783
rect 1458 3774 1470 3783
rect 1522 3774 1534 3783
rect 1586 3774 1598 3783
rect 1650 3774 1662 3826
rect 1714 3774 1726 3826
rect 1778 3774 1790 3826
rect 1842 3774 1854 3826
rect 1906 3817 1918 3826
rect 1970 3817 1982 3826
rect 2034 3817 2046 3826
rect 2098 3817 2110 3826
rect 2162 3817 2174 3826
rect 1913 3783 1918 3817
rect 2162 3783 2167 3817
rect 1906 3774 1918 3783
rect 1970 3774 1982 3783
rect 2034 3774 2046 3783
rect 2098 3774 2110 3783
rect 2162 3774 2174 3783
rect 2226 3774 2238 3826
rect 2290 3774 2302 3826
rect 2354 3774 2366 3826
rect 2418 3774 2430 3826
rect 2482 3817 2494 3826
rect 2546 3817 2558 3826
rect 2610 3817 2622 3826
rect 2674 3817 2686 3826
rect 2738 3817 2750 3826
rect 2489 3783 2494 3817
rect 2738 3783 2743 3817
rect 2482 3774 2494 3783
rect 2546 3774 2558 3783
rect 2610 3774 2622 3783
rect 2674 3774 2686 3783
rect 2738 3774 2750 3783
rect 2802 3774 2814 3826
rect 2866 3774 2878 3826
rect 2930 3774 2942 3826
rect 2994 3774 3006 3826
rect 3058 3817 3070 3826
rect 3122 3817 3134 3826
rect 3186 3817 3198 3826
rect 3250 3817 3262 3826
rect 3314 3817 3326 3826
rect 3065 3783 3070 3817
rect 3314 3783 3319 3817
rect 3058 3774 3070 3783
rect 3122 3774 3134 3783
rect 3186 3774 3198 3783
rect 3250 3774 3262 3783
rect 3314 3774 3326 3783
rect 3378 3774 3390 3826
rect 3442 3774 3454 3826
rect 3506 3774 3518 3826
rect 3570 3774 3582 3826
rect 3634 3817 3646 3826
rect 3698 3817 3710 3826
rect 3762 3817 3774 3826
rect 3826 3817 3838 3826
rect 3890 3817 3902 3826
rect 3641 3783 3646 3817
rect 3890 3783 3895 3817
rect 3634 3774 3646 3783
rect 3698 3774 3710 3783
rect 3762 3774 3774 3783
rect 3826 3774 3838 3783
rect 3890 3774 3902 3783
rect 3954 3774 3966 3826
rect 4018 3774 4040 3826
rect 40 3760 4040 3774
rect -160 3623 -137 3657
rect -103 3623 -80 3657
rect -160 3506 -80 3623
rect 4160 3657 4240 3943
rect 4160 3623 4183 3657
rect 4217 3623 4240 3657
rect -160 3454 -146 3506
rect -94 3454 -80 3506
rect -160 2537 -80 3454
rect 40 3506 4040 3520
rect 40 3454 62 3506
rect 114 3454 126 3506
rect 178 3497 190 3506
rect 242 3497 254 3506
rect 306 3497 318 3506
rect 370 3497 382 3506
rect 434 3497 446 3506
rect 185 3463 190 3497
rect 434 3463 439 3497
rect 178 3454 190 3463
rect 242 3454 254 3463
rect 306 3454 318 3463
rect 370 3454 382 3463
rect 434 3454 446 3463
rect 498 3454 510 3506
rect 562 3454 574 3506
rect 626 3454 638 3506
rect 690 3454 702 3506
rect 754 3497 766 3506
rect 818 3497 830 3506
rect 882 3497 894 3506
rect 946 3497 958 3506
rect 1010 3497 1022 3506
rect 761 3463 766 3497
rect 1010 3463 1015 3497
rect 754 3454 766 3463
rect 818 3454 830 3463
rect 882 3454 894 3463
rect 946 3454 958 3463
rect 1010 3454 1022 3463
rect 1074 3454 1086 3506
rect 1138 3454 1150 3506
rect 1202 3454 1214 3506
rect 1266 3454 1278 3506
rect 1330 3497 1342 3506
rect 1394 3497 1406 3506
rect 1458 3497 1470 3506
rect 1522 3497 1534 3506
rect 1586 3497 1598 3506
rect 1337 3463 1342 3497
rect 1586 3463 1591 3497
rect 1330 3454 1342 3463
rect 1394 3454 1406 3463
rect 1458 3454 1470 3463
rect 1522 3454 1534 3463
rect 1586 3454 1598 3463
rect 1650 3454 1662 3506
rect 1714 3454 1726 3506
rect 1778 3454 1790 3506
rect 1842 3454 1854 3506
rect 1906 3497 1918 3506
rect 1970 3497 1982 3506
rect 2034 3497 2046 3506
rect 2098 3497 2110 3506
rect 2162 3497 2174 3506
rect 1913 3463 1918 3497
rect 2162 3463 2167 3497
rect 1906 3454 1918 3463
rect 1970 3454 1982 3463
rect 2034 3454 2046 3463
rect 2098 3454 2110 3463
rect 2162 3454 2174 3463
rect 2226 3454 2238 3506
rect 2290 3454 2302 3506
rect 2354 3454 2366 3506
rect 2418 3454 2430 3506
rect 2482 3497 2494 3506
rect 2546 3497 2558 3506
rect 2610 3497 2622 3506
rect 2674 3497 2686 3506
rect 2738 3497 2750 3506
rect 2489 3463 2494 3497
rect 2738 3463 2743 3497
rect 2482 3454 2494 3463
rect 2546 3454 2558 3463
rect 2610 3454 2622 3463
rect 2674 3454 2686 3463
rect 2738 3454 2750 3463
rect 2802 3454 2814 3506
rect 2866 3454 2878 3506
rect 2930 3454 2942 3506
rect 2994 3454 3006 3506
rect 3058 3497 3070 3506
rect 3122 3497 3134 3506
rect 3186 3497 3198 3506
rect 3250 3497 3262 3506
rect 3314 3497 3326 3506
rect 3065 3463 3070 3497
rect 3314 3463 3319 3497
rect 3058 3454 3070 3463
rect 3122 3454 3134 3463
rect 3186 3454 3198 3463
rect 3250 3454 3262 3463
rect 3314 3454 3326 3463
rect 3378 3454 3390 3506
rect 3442 3454 3454 3506
rect 3506 3454 3518 3506
rect 3570 3454 3582 3506
rect 3634 3497 3646 3506
rect 3698 3497 3710 3506
rect 3762 3497 3774 3506
rect 3826 3497 3838 3506
rect 3890 3497 3902 3506
rect 3641 3463 3646 3497
rect 3890 3463 3895 3497
rect 3634 3454 3646 3463
rect 3698 3454 3710 3463
rect 3762 3454 3774 3463
rect 3826 3454 3838 3463
rect 3890 3454 3902 3463
rect 3954 3454 3966 3506
rect 4018 3454 4040 3506
rect 40 3440 4040 3454
rect 4160 2857 4240 3623
rect 4160 2823 4183 2857
rect 4217 2823 4240 2857
rect 40 2706 4040 2720
rect 40 2654 62 2706
rect 114 2654 126 2706
rect 178 2697 190 2706
rect 242 2697 254 2706
rect 306 2697 318 2706
rect 370 2697 382 2706
rect 434 2697 446 2706
rect 185 2663 190 2697
rect 434 2663 439 2697
rect 178 2654 190 2663
rect 242 2654 254 2663
rect 306 2654 318 2663
rect 370 2654 382 2663
rect 434 2654 446 2663
rect 498 2654 510 2706
rect 562 2654 574 2706
rect 626 2654 638 2706
rect 690 2654 702 2706
rect 754 2697 766 2706
rect 818 2697 830 2706
rect 882 2697 894 2706
rect 946 2697 958 2706
rect 1010 2697 1022 2706
rect 761 2663 766 2697
rect 1010 2663 1015 2697
rect 754 2654 766 2663
rect 818 2654 830 2663
rect 882 2654 894 2663
rect 946 2654 958 2663
rect 1010 2654 1022 2663
rect 1074 2654 1086 2706
rect 1138 2654 1150 2706
rect 1202 2654 1214 2706
rect 1266 2654 1278 2706
rect 1330 2697 1342 2706
rect 1394 2697 1406 2706
rect 1458 2697 1470 2706
rect 1522 2697 1534 2706
rect 1586 2697 1598 2706
rect 1337 2663 1342 2697
rect 1586 2663 1591 2697
rect 1330 2654 1342 2663
rect 1394 2654 1406 2663
rect 1458 2654 1470 2663
rect 1522 2654 1534 2663
rect 1586 2654 1598 2663
rect 1650 2654 1662 2706
rect 1714 2654 1726 2706
rect 1778 2654 1790 2706
rect 1842 2654 1854 2706
rect 1906 2697 1918 2706
rect 1970 2697 1982 2706
rect 2034 2697 2046 2706
rect 2098 2697 2110 2706
rect 2162 2697 2174 2706
rect 1913 2663 1918 2697
rect 2162 2663 2167 2697
rect 1906 2654 1918 2663
rect 1970 2654 1982 2663
rect 2034 2654 2046 2663
rect 2098 2654 2110 2663
rect 2162 2654 2174 2663
rect 2226 2654 2238 2706
rect 2290 2654 2302 2706
rect 2354 2654 2366 2706
rect 2418 2654 2430 2706
rect 2482 2697 2494 2706
rect 2546 2697 2558 2706
rect 2610 2697 2622 2706
rect 2674 2697 2686 2706
rect 2738 2697 2750 2706
rect 2489 2663 2494 2697
rect 2738 2663 2743 2697
rect 2482 2654 2494 2663
rect 2546 2654 2558 2663
rect 2610 2654 2622 2663
rect 2674 2654 2686 2663
rect 2738 2654 2750 2663
rect 2802 2654 2814 2706
rect 2866 2654 2878 2706
rect 2930 2654 2942 2706
rect 2994 2654 3006 2706
rect 3058 2697 3070 2706
rect 3122 2697 3134 2706
rect 3186 2697 3198 2706
rect 3250 2697 3262 2706
rect 3314 2697 3326 2706
rect 3065 2663 3070 2697
rect 3314 2663 3319 2697
rect 3058 2654 3070 2663
rect 3122 2654 3134 2663
rect 3186 2654 3198 2663
rect 3250 2654 3262 2663
rect 3314 2654 3326 2663
rect 3378 2654 3390 2706
rect 3442 2654 3454 2706
rect 3506 2654 3518 2706
rect 3570 2654 3582 2706
rect 3634 2697 3646 2706
rect 3698 2697 3710 2706
rect 3762 2697 3774 2706
rect 3826 2697 3838 2706
rect 3890 2697 3902 2706
rect 3641 2663 3646 2697
rect 3890 2663 3895 2697
rect 3634 2654 3646 2663
rect 3698 2654 3710 2663
rect 3762 2654 3774 2663
rect 3826 2654 3838 2663
rect 3890 2654 3902 2663
rect 3954 2654 3966 2706
rect 4018 2654 4040 2706
rect 40 2640 4040 2654
rect 4160 2706 4240 2823
rect 4160 2654 4174 2706
rect 4226 2654 4240 2706
rect -160 2503 -137 2537
rect -103 2503 -80 2537
rect -160 2217 -80 2503
rect 4160 2537 4240 2654
rect 4160 2503 4183 2537
rect 4217 2503 4240 2537
rect 40 2386 4040 2400
rect 40 2334 62 2386
rect 114 2334 126 2386
rect 178 2377 190 2386
rect 242 2377 254 2386
rect 306 2377 318 2386
rect 370 2377 382 2386
rect 434 2377 446 2386
rect 185 2343 190 2377
rect 434 2343 439 2377
rect 178 2334 190 2343
rect 242 2334 254 2343
rect 306 2334 318 2343
rect 370 2334 382 2343
rect 434 2334 446 2343
rect 498 2334 510 2386
rect 562 2334 574 2386
rect 626 2334 638 2386
rect 690 2334 702 2386
rect 754 2377 766 2386
rect 818 2377 830 2386
rect 882 2377 894 2386
rect 946 2377 958 2386
rect 1010 2377 1022 2386
rect 761 2343 766 2377
rect 1010 2343 1015 2377
rect 754 2334 766 2343
rect 818 2334 830 2343
rect 882 2334 894 2343
rect 946 2334 958 2343
rect 1010 2334 1022 2343
rect 1074 2334 1086 2386
rect 1138 2334 1150 2386
rect 1202 2334 1214 2386
rect 1266 2334 1278 2386
rect 1330 2377 1342 2386
rect 1394 2377 1406 2386
rect 1458 2377 1470 2386
rect 1522 2377 1534 2386
rect 1586 2377 1598 2386
rect 1337 2343 1342 2377
rect 1586 2343 1591 2377
rect 1330 2334 1342 2343
rect 1394 2334 1406 2343
rect 1458 2334 1470 2343
rect 1522 2334 1534 2343
rect 1586 2334 1598 2343
rect 1650 2334 1662 2386
rect 1714 2334 1726 2386
rect 1778 2334 1790 2386
rect 1842 2334 1854 2386
rect 1906 2377 1918 2386
rect 1970 2377 1982 2386
rect 2034 2377 2046 2386
rect 2098 2377 2110 2386
rect 2162 2377 2174 2386
rect 1913 2343 1918 2377
rect 2162 2343 2167 2377
rect 1906 2334 1918 2343
rect 1970 2334 1982 2343
rect 2034 2334 2046 2343
rect 2098 2334 2110 2343
rect 2162 2334 2174 2343
rect 2226 2334 2238 2386
rect 2290 2334 2302 2386
rect 2354 2334 2366 2386
rect 2418 2334 2430 2386
rect 2482 2377 2494 2386
rect 2546 2377 2558 2386
rect 2610 2377 2622 2386
rect 2674 2377 2686 2386
rect 2738 2377 2750 2386
rect 2489 2343 2494 2377
rect 2738 2343 2743 2377
rect 2482 2334 2494 2343
rect 2546 2334 2558 2343
rect 2610 2334 2622 2343
rect 2674 2334 2686 2343
rect 2738 2334 2750 2343
rect 2802 2334 2814 2386
rect 2866 2334 2878 2386
rect 2930 2334 2942 2386
rect 2994 2334 3006 2386
rect 3058 2377 3070 2386
rect 3122 2377 3134 2386
rect 3186 2377 3198 2386
rect 3250 2377 3262 2386
rect 3314 2377 3326 2386
rect 3065 2343 3070 2377
rect 3314 2343 3319 2377
rect 3058 2334 3070 2343
rect 3122 2334 3134 2343
rect 3186 2334 3198 2343
rect 3250 2334 3262 2343
rect 3314 2334 3326 2343
rect 3378 2334 3390 2386
rect 3442 2334 3454 2386
rect 3506 2334 3518 2386
rect 3570 2334 3582 2386
rect 3634 2377 3646 2386
rect 3698 2377 3710 2386
rect 3762 2377 3774 2386
rect 3826 2377 3838 2386
rect 3890 2377 3902 2386
rect 3641 2343 3646 2377
rect 3890 2343 3895 2377
rect 3634 2334 3646 2343
rect 3698 2334 3710 2343
rect 3762 2334 3774 2343
rect 3826 2334 3838 2343
rect 3890 2334 3902 2343
rect 3954 2334 3966 2386
rect 4018 2334 4040 2386
rect 40 2320 4040 2334
rect -160 2183 -137 2217
rect -103 2183 -80 2217
rect -160 2160 -80 2183
rect 4160 2217 4240 2503
rect 4160 2183 4183 2217
rect 4217 2183 4240 2217
rect 4160 2160 4240 2183
rect 8320 3977 8400 4000
rect 8320 3943 8343 3977
rect 8377 3943 8400 3977
rect 8320 3657 8400 3943
rect 12640 3977 12720 4000
rect 12640 3943 12663 3977
rect 12697 3943 12720 3977
rect 8520 3826 12520 3840
rect 8520 3774 8542 3826
rect 8594 3774 8606 3826
rect 8658 3817 8670 3826
rect 8722 3817 8734 3826
rect 8786 3817 8798 3826
rect 8850 3817 8862 3826
rect 8914 3817 8926 3826
rect 8665 3783 8670 3817
rect 8914 3783 8919 3817
rect 8658 3774 8670 3783
rect 8722 3774 8734 3783
rect 8786 3774 8798 3783
rect 8850 3774 8862 3783
rect 8914 3774 8926 3783
rect 8978 3774 8990 3826
rect 9042 3774 9054 3826
rect 9106 3774 9118 3826
rect 9170 3774 9182 3826
rect 9234 3817 9246 3826
rect 9298 3817 9310 3826
rect 9362 3817 9374 3826
rect 9426 3817 9438 3826
rect 9490 3817 9502 3826
rect 9241 3783 9246 3817
rect 9490 3783 9495 3817
rect 9234 3774 9246 3783
rect 9298 3774 9310 3783
rect 9362 3774 9374 3783
rect 9426 3774 9438 3783
rect 9490 3774 9502 3783
rect 9554 3774 9566 3826
rect 9618 3774 9630 3826
rect 9682 3774 9694 3826
rect 9746 3774 9758 3826
rect 9810 3817 9822 3826
rect 9874 3817 9886 3826
rect 9938 3817 9950 3826
rect 10002 3817 10014 3826
rect 10066 3817 10078 3826
rect 9817 3783 9822 3817
rect 10066 3783 10071 3817
rect 9810 3774 9822 3783
rect 9874 3774 9886 3783
rect 9938 3774 9950 3783
rect 10002 3774 10014 3783
rect 10066 3774 10078 3783
rect 10130 3774 10142 3826
rect 10194 3774 10206 3826
rect 10258 3774 10270 3826
rect 10322 3774 10334 3826
rect 10386 3817 10398 3826
rect 10450 3817 10462 3826
rect 10514 3817 10526 3826
rect 10578 3817 10590 3826
rect 10642 3817 10654 3826
rect 10393 3783 10398 3817
rect 10642 3783 10647 3817
rect 10386 3774 10398 3783
rect 10450 3774 10462 3783
rect 10514 3774 10526 3783
rect 10578 3774 10590 3783
rect 10642 3774 10654 3783
rect 10706 3774 10718 3826
rect 10770 3774 10782 3826
rect 10834 3774 10846 3826
rect 10898 3774 10910 3826
rect 10962 3817 10974 3826
rect 11026 3817 11038 3826
rect 11090 3817 11102 3826
rect 11154 3817 11166 3826
rect 11218 3817 11230 3826
rect 10969 3783 10974 3817
rect 11218 3783 11223 3817
rect 10962 3774 10974 3783
rect 11026 3774 11038 3783
rect 11090 3774 11102 3783
rect 11154 3774 11166 3783
rect 11218 3774 11230 3783
rect 11282 3774 11294 3826
rect 11346 3774 11358 3826
rect 11410 3774 11422 3826
rect 11474 3774 11486 3826
rect 11538 3817 11550 3826
rect 11602 3817 11614 3826
rect 11666 3817 11678 3826
rect 11730 3817 11742 3826
rect 11794 3817 11806 3826
rect 11545 3783 11550 3817
rect 11794 3783 11799 3817
rect 11538 3774 11550 3783
rect 11602 3774 11614 3783
rect 11666 3774 11678 3783
rect 11730 3774 11742 3783
rect 11794 3774 11806 3783
rect 11858 3774 11870 3826
rect 11922 3774 11934 3826
rect 11986 3774 11998 3826
rect 12050 3774 12062 3826
rect 12114 3817 12126 3826
rect 12178 3817 12190 3826
rect 12242 3817 12254 3826
rect 12306 3817 12318 3826
rect 12370 3817 12382 3826
rect 12121 3783 12126 3817
rect 12370 3783 12375 3817
rect 12114 3774 12126 3783
rect 12178 3774 12190 3783
rect 12242 3774 12254 3783
rect 12306 3774 12318 3783
rect 12370 3774 12382 3783
rect 12434 3774 12446 3826
rect 12498 3774 12520 3826
rect 8520 3760 12520 3774
rect 8320 3623 8343 3657
rect 8377 3623 8400 3657
rect 8320 2857 8400 3623
rect 12640 3657 12720 3943
rect 12640 3623 12663 3657
rect 12697 3623 12720 3657
rect 8520 3506 12520 3520
rect 8520 3454 8542 3506
rect 8594 3454 8606 3506
rect 8658 3497 8670 3506
rect 8722 3497 8734 3506
rect 8786 3497 8798 3506
rect 8850 3497 8862 3506
rect 8914 3497 8926 3506
rect 8665 3463 8670 3497
rect 8914 3463 8919 3497
rect 8658 3454 8670 3463
rect 8722 3454 8734 3463
rect 8786 3454 8798 3463
rect 8850 3454 8862 3463
rect 8914 3454 8926 3463
rect 8978 3454 8990 3506
rect 9042 3454 9054 3506
rect 9106 3454 9118 3506
rect 9170 3454 9182 3506
rect 9234 3497 9246 3506
rect 9298 3497 9310 3506
rect 9362 3497 9374 3506
rect 9426 3497 9438 3506
rect 9490 3497 9502 3506
rect 9241 3463 9246 3497
rect 9490 3463 9495 3497
rect 9234 3454 9246 3463
rect 9298 3454 9310 3463
rect 9362 3454 9374 3463
rect 9426 3454 9438 3463
rect 9490 3454 9502 3463
rect 9554 3454 9566 3506
rect 9618 3454 9630 3506
rect 9682 3454 9694 3506
rect 9746 3454 9758 3506
rect 9810 3497 9822 3506
rect 9874 3497 9886 3506
rect 9938 3497 9950 3506
rect 10002 3497 10014 3506
rect 10066 3497 10078 3506
rect 9817 3463 9822 3497
rect 10066 3463 10071 3497
rect 9810 3454 9822 3463
rect 9874 3454 9886 3463
rect 9938 3454 9950 3463
rect 10002 3454 10014 3463
rect 10066 3454 10078 3463
rect 10130 3454 10142 3506
rect 10194 3454 10206 3506
rect 10258 3454 10270 3506
rect 10322 3454 10334 3506
rect 10386 3497 10398 3506
rect 10450 3497 10462 3506
rect 10514 3497 10526 3506
rect 10578 3497 10590 3506
rect 10642 3497 10654 3506
rect 10393 3463 10398 3497
rect 10642 3463 10647 3497
rect 10386 3454 10398 3463
rect 10450 3454 10462 3463
rect 10514 3454 10526 3463
rect 10578 3454 10590 3463
rect 10642 3454 10654 3463
rect 10706 3454 10718 3506
rect 10770 3454 10782 3506
rect 10834 3454 10846 3506
rect 10898 3454 10910 3506
rect 10962 3497 10974 3506
rect 11026 3497 11038 3506
rect 11090 3497 11102 3506
rect 11154 3497 11166 3506
rect 11218 3497 11230 3506
rect 10969 3463 10974 3497
rect 11218 3463 11223 3497
rect 10962 3454 10974 3463
rect 11026 3454 11038 3463
rect 11090 3454 11102 3463
rect 11154 3454 11166 3463
rect 11218 3454 11230 3463
rect 11282 3454 11294 3506
rect 11346 3454 11358 3506
rect 11410 3454 11422 3506
rect 11474 3454 11486 3506
rect 11538 3497 11550 3506
rect 11602 3497 11614 3506
rect 11666 3497 11678 3506
rect 11730 3497 11742 3506
rect 11794 3497 11806 3506
rect 11545 3463 11550 3497
rect 11794 3463 11799 3497
rect 11538 3454 11550 3463
rect 11602 3454 11614 3463
rect 11666 3454 11678 3463
rect 11730 3454 11742 3463
rect 11794 3454 11806 3463
rect 11858 3454 11870 3506
rect 11922 3454 11934 3506
rect 11986 3454 11998 3506
rect 12050 3454 12062 3506
rect 12114 3497 12126 3506
rect 12178 3497 12190 3506
rect 12242 3497 12254 3506
rect 12306 3497 12318 3506
rect 12370 3497 12382 3506
rect 12121 3463 12126 3497
rect 12370 3463 12375 3497
rect 12114 3454 12126 3463
rect 12178 3454 12190 3463
rect 12242 3454 12254 3463
rect 12306 3454 12318 3463
rect 12370 3454 12382 3463
rect 12434 3454 12446 3506
rect 12498 3454 12520 3506
rect 8520 3440 12520 3454
rect 12640 3506 12720 3623
rect 12640 3454 12654 3506
rect 12706 3454 12720 3506
rect 8320 2823 8343 2857
rect 8377 2823 8400 2857
rect 8320 2706 8400 2823
rect 8320 2654 8334 2706
rect 8386 2654 8400 2706
rect 8320 2537 8400 2654
rect 8520 2706 12520 2720
rect 8520 2654 8542 2706
rect 8594 2654 8606 2706
rect 8658 2697 8670 2706
rect 8722 2697 8734 2706
rect 8786 2697 8798 2706
rect 8850 2697 8862 2706
rect 8914 2697 8926 2706
rect 8665 2663 8670 2697
rect 8914 2663 8919 2697
rect 8658 2654 8670 2663
rect 8722 2654 8734 2663
rect 8786 2654 8798 2663
rect 8850 2654 8862 2663
rect 8914 2654 8926 2663
rect 8978 2654 8990 2706
rect 9042 2654 9054 2706
rect 9106 2654 9118 2706
rect 9170 2654 9182 2706
rect 9234 2697 9246 2706
rect 9298 2697 9310 2706
rect 9362 2697 9374 2706
rect 9426 2697 9438 2706
rect 9490 2697 9502 2706
rect 9241 2663 9246 2697
rect 9490 2663 9495 2697
rect 9234 2654 9246 2663
rect 9298 2654 9310 2663
rect 9362 2654 9374 2663
rect 9426 2654 9438 2663
rect 9490 2654 9502 2663
rect 9554 2654 9566 2706
rect 9618 2654 9630 2706
rect 9682 2654 9694 2706
rect 9746 2654 9758 2706
rect 9810 2697 9822 2706
rect 9874 2697 9886 2706
rect 9938 2697 9950 2706
rect 10002 2697 10014 2706
rect 10066 2697 10078 2706
rect 9817 2663 9822 2697
rect 10066 2663 10071 2697
rect 9810 2654 9822 2663
rect 9874 2654 9886 2663
rect 9938 2654 9950 2663
rect 10002 2654 10014 2663
rect 10066 2654 10078 2663
rect 10130 2654 10142 2706
rect 10194 2654 10206 2706
rect 10258 2654 10270 2706
rect 10322 2654 10334 2706
rect 10386 2697 10398 2706
rect 10450 2697 10462 2706
rect 10514 2697 10526 2706
rect 10578 2697 10590 2706
rect 10642 2697 10654 2706
rect 10393 2663 10398 2697
rect 10642 2663 10647 2697
rect 10386 2654 10398 2663
rect 10450 2654 10462 2663
rect 10514 2654 10526 2663
rect 10578 2654 10590 2663
rect 10642 2654 10654 2663
rect 10706 2654 10718 2706
rect 10770 2654 10782 2706
rect 10834 2654 10846 2706
rect 10898 2654 10910 2706
rect 10962 2697 10974 2706
rect 11026 2697 11038 2706
rect 11090 2697 11102 2706
rect 11154 2697 11166 2706
rect 11218 2697 11230 2706
rect 10969 2663 10974 2697
rect 11218 2663 11223 2697
rect 10962 2654 10974 2663
rect 11026 2654 11038 2663
rect 11090 2654 11102 2663
rect 11154 2654 11166 2663
rect 11218 2654 11230 2663
rect 11282 2654 11294 2706
rect 11346 2654 11358 2706
rect 11410 2654 11422 2706
rect 11474 2654 11486 2706
rect 11538 2697 11550 2706
rect 11602 2697 11614 2706
rect 11666 2697 11678 2706
rect 11730 2697 11742 2706
rect 11794 2697 11806 2706
rect 11545 2663 11550 2697
rect 11794 2663 11799 2697
rect 11538 2654 11550 2663
rect 11602 2654 11614 2663
rect 11666 2654 11678 2663
rect 11730 2654 11742 2663
rect 11794 2654 11806 2663
rect 11858 2654 11870 2706
rect 11922 2654 11934 2706
rect 11986 2654 11998 2706
rect 12050 2654 12062 2706
rect 12114 2697 12126 2706
rect 12178 2697 12190 2706
rect 12242 2697 12254 2706
rect 12306 2697 12318 2706
rect 12370 2697 12382 2706
rect 12121 2663 12126 2697
rect 12370 2663 12375 2697
rect 12114 2654 12126 2663
rect 12178 2654 12190 2663
rect 12242 2654 12254 2663
rect 12306 2654 12318 2663
rect 12370 2654 12382 2663
rect 12434 2654 12446 2706
rect 12498 2654 12520 2706
rect 8520 2640 12520 2654
rect 8320 2503 8343 2537
rect 8377 2503 8400 2537
rect 8320 2217 8400 2503
rect 12640 2537 12720 3454
rect 12640 2503 12663 2537
rect 12697 2503 12720 2537
rect 8520 2386 12520 2400
rect 8520 2334 8542 2386
rect 8594 2334 8606 2386
rect 8658 2377 8670 2386
rect 8722 2377 8734 2386
rect 8786 2377 8798 2386
rect 8850 2377 8862 2386
rect 8914 2377 8926 2386
rect 8665 2343 8670 2377
rect 8914 2343 8919 2377
rect 8658 2334 8670 2343
rect 8722 2334 8734 2343
rect 8786 2334 8798 2343
rect 8850 2334 8862 2343
rect 8914 2334 8926 2343
rect 8978 2334 8990 2386
rect 9042 2334 9054 2386
rect 9106 2334 9118 2386
rect 9170 2334 9182 2386
rect 9234 2377 9246 2386
rect 9298 2377 9310 2386
rect 9362 2377 9374 2386
rect 9426 2377 9438 2386
rect 9490 2377 9502 2386
rect 9241 2343 9246 2377
rect 9490 2343 9495 2377
rect 9234 2334 9246 2343
rect 9298 2334 9310 2343
rect 9362 2334 9374 2343
rect 9426 2334 9438 2343
rect 9490 2334 9502 2343
rect 9554 2334 9566 2386
rect 9618 2334 9630 2386
rect 9682 2334 9694 2386
rect 9746 2334 9758 2386
rect 9810 2377 9822 2386
rect 9874 2377 9886 2386
rect 9938 2377 9950 2386
rect 10002 2377 10014 2386
rect 10066 2377 10078 2386
rect 9817 2343 9822 2377
rect 10066 2343 10071 2377
rect 9810 2334 9822 2343
rect 9874 2334 9886 2343
rect 9938 2334 9950 2343
rect 10002 2334 10014 2343
rect 10066 2334 10078 2343
rect 10130 2334 10142 2386
rect 10194 2334 10206 2386
rect 10258 2334 10270 2386
rect 10322 2334 10334 2386
rect 10386 2377 10398 2386
rect 10450 2377 10462 2386
rect 10514 2377 10526 2386
rect 10578 2377 10590 2386
rect 10642 2377 10654 2386
rect 10393 2343 10398 2377
rect 10642 2343 10647 2377
rect 10386 2334 10398 2343
rect 10450 2334 10462 2343
rect 10514 2334 10526 2343
rect 10578 2334 10590 2343
rect 10642 2334 10654 2343
rect 10706 2334 10718 2386
rect 10770 2334 10782 2386
rect 10834 2334 10846 2386
rect 10898 2334 10910 2386
rect 10962 2377 10974 2386
rect 11026 2377 11038 2386
rect 11090 2377 11102 2386
rect 11154 2377 11166 2386
rect 11218 2377 11230 2386
rect 10969 2343 10974 2377
rect 11218 2343 11223 2377
rect 10962 2334 10974 2343
rect 11026 2334 11038 2343
rect 11090 2334 11102 2343
rect 11154 2334 11166 2343
rect 11218 2334 11230 2343
rect 11282 2334 11294 2386
rect 11346 2334 11358 2386
rect 11410 2334 11422 2386
rect 11474 2334 11486 2386
rect 11538 2377 11550 2386
rect 11602 2377 11614 2386
rect 11666 2377 11678 2386
rect 11730 2377 11742 2386
rect 11794 2377 11806 2386
rect 11545 2343 11550 2377
rect 11794 2343 11799 2377
rect 11538 2334 11550 2343
rect 11602 2334 11614 2343
rect 11666 2334 11678 2343
rect 11730 2334 11742 2343
rect 11794 2334 11806 2343
rect 11858 2334 11870 2386
rect 11922 2334 11934 2386
rect 11986 2334 11998 2386
rect 12050 2334 12062 2386
rect 12114 2377 12126 2386
rect 12178 2377 12190 2386
rect 12242 2377 12254 2386
rect 12306 2377 12318 2386
rect 12370 2377 12382 2386
rect 12121 2343 12126 2377
rect 12370 2343 12375 2377
rect 12114 2334 12126 2343
rect 12178 2334 12190 2343
rect 12242 2334 12254 2343
rect 12306 2334 12318 2343
rect 12370 2334 12382 2343
rect 12434 2334 12446 2386
rect 12498 2334 12520 2386
rect 8520 2320 12520 2334
rect 8320 2183 8343 2217
rect 8377 2183 8400 2217
rect 8320 2160 8400 2183
rect 12640 2217 12720 2503
rect 12640 2183 12663 2217
rect 12697 2183 12720 2217
rect 12640 2160 12720 2183
rect -400 1826 -160 1920
rect -400 1774 -306 1826
rect -254 1774 -160 1826
rect -400 1680 -160 1774
rect 12720 1826 12960 1920
rect 12720 1774 12814 1826
rect 12866 1774 12960 1826
rect 12720 1680 12960 1774
rect -160 1417 -80 1440
rect -160 1383 -137 1417
rect -103 1383 -80 1417
rect -160 1097 -80 1383
rect 4160 1417 4240 1440
rect 4160 1383 4183 1417
rect 4217 1383 4240 1417
rect 40 1266 4040 1280
rect 40 1214 62 1266
rect 114 1214 126 1266
rect 178 1257 190 1266
rect 242 1257 254 1266
rect 306 1257 318 1266
rect 370 1257 382 1266
rect 434 1257 446 1266
rect 185 1223 190 1257
rect 434 1223 439 1257
rect 178 1214 190 1223
rect 242 1214 254 1223
rect 306 1214 318 1223
rect 370 1214 382 1223
rect 434 1214 446 1223
rect 498 1214 510 1266
rect 562 1214 574 1266
rect 626 1214 638 1266
rect 690 1214 702 1266
rect 754 1257 766 1266
rect 818 1257 830 1266
rect 882 1257 894 1266
rect 946 1257 958 1266
rect 1010 1257 1022 1266
rect 761 1223 766 1257
rect 1010 1223 1015 1257
rect 754 1214 766 1223
rect 818 1214 830 1223
rect 882 1214 894 1223
rect 946 1214 958 1223
rect 1010 1214 1022 1223
rect 1074 1214 1086 1266
rect 1138 1214 1150 1266
rect 1202 1214 1214 1266
rect 1266 1214 1278 1266
rect 1330 1257 1342 1266
rect 1394 1257 1406 1266
rect 1458 1257 1470 1266
rect 1522 1257 1534 1266
rect 1586 1257 1598 1266
rect 1337 1223 1342 1257
rect 1586 1223 1591 1257
rect 1330 1214 1342 1223
rect 1394 1214 1406 1223
rect 1458 1214 1470 1223
rect 1522 1214 1534 1223
rect 1586 1214 1598 1223
rect 1650 1214 1662 1266
rect 1714 1214 1726 1266
rect 1778 1214 1790 1266
rect 1842 1214 1854 1266
rect 1906 1257 1918 1266
rect 1970 1257 1982 1266
rect 2034 1257 2046 1266
rect 2098 1257 2110 1266
rect 2162 1257 2174 1266
rect 1913 1223 1918 1257
rect 2162 1223 2167 1257
rect 1906 1214 1918 1223
rect 1970 1214 1982 1223
rect 2034 1214 2046 1223
rect 2098 1214 2110 1223
rect 2162 1214 2174 1223
rect 2226 1214 2238 1266
rect 2290 1214 2302 1266
rect 2354 1214 2366 1266
rect 2418 1214 2430 1266
rect 2482 1257 2494 1266
rect 2546 1257 2558 1266
rect 2610 1257 2622 1266
rect 2674 1257 2686 1266
rect 2738 1257 2750 1266
rect 2489 1223 2494 1257
rect 2738 1223 2743 1257
rect 2482 1214 2494 1223
rect 2546 1214 2558 1223
rect 2610 1214 2622 1223
rect 2674 1214 2686 1223
rect 2738 1214 2750 1223
rect 2802 1214 2814 1266
rect 2866 1214 2878 1266
rect 2930 1214 2942 1266
rect 2994 1214 3006 1266
rect 3058 1257 3070 1266
rect 3122 1257 3134 1266
rect 3186 1257 3198 1266
rect 3250 1257 3262 1266
rect 3314 1257 3326 1266
rect 3065 1223 3070 1257
rect 3314 1223 3319 1257
rect 3058 1214 3070 1223
rect 3122 1214 3134 1223
rect 3186 1214 3198 1223
rect 3250 1214 3262 1223
rect 3314 1214 3326 1223
rect 3378 1214 3390 1266
rect 3442 1214 3454 1266
rect 3506 1214 3518 1266
rect 3570 1214 3582 1266
rect 3634 1257 3646 1266
rect 3698 1257 3710 1266
rect 3762 1257 3774 1266
rect 3826 1257 3838 1266
rect 3890 1257 3902 1266
rect 3641 1223 3646 1257
rect 3890 1223 3895 1257
rect 3634 1214 3646 1223
rect 3698 1214 3710 1223
rect 3762 1214 3774 1223
rect 3826 1214 3838 1223
rect 3890 1214 3902 1223
rect 3954 1214 3966 1266
rect 4018 1214 4040 1266
rect 40 1200 4040 1214
rect -160 1063 -137 1097
rect -103 1063 -80 1097
rect -160 146 -80 1063
rect 4160 1097 4240 1383
rect 4160 1063 4183 1097
rect 4217 1063 4240 1097
rect 40 946 4040 960
rect 40 894 62 946
rect 114 894 126 946
rect 178 937 190 946
rect 242 937 254 946
rect 306 937 318 946
rect 370 937 382 946
rect 434 937 446 946
rect 185 903 190 937
rect 434 903 439 937
rect 178 894 190 903
rect 242 894 254 903
rect 306 894 318 903
rect 370 894 382 903
rect 434 894 446 903
rect 498 894 510 946
rect 562 894 574 946
rect 626 894 638 946
rect 690 894 702 946
rect 754 937 766 946
rect 818 937 830 946
rect 882 937 894 946
rect 946 937 958 946
rect 1010 937 1022 946
rect 761 903 766 937
rect 1010 903 1015 937
rect 754 894 766 903
rect 818 894 830 903
rect 882 894 894 903
rect 946 894 958 903
rect 1010 894 1022 903
rect 1074 894 1086 946
rect 1138 894 1150 946
rect 1202 894 1214 946
rect 1266 894 1278 946
rect 1330 937 1342 946
rect 1394 937 1406 946
rect 1458 937 1470 946
rect 1522 937 1534 946
rect 1586 937 1598 946
rect 1337 903 1342 937
rect 1586 903 1591 937
rect 1330 894 1342 903
rect 1394 894 1406 903
rect 1458 894 1470 903
rect 1522 894 1534 903
rect 1586 894 1598 903
rect 1650 894 1662 946
rect 1714 894 1726 946
rect 1778 894 1790 946
rect 1842 894 1854 946
rect 1906 937 1918 946
rect 1970 937 1982 946
rect 2034 937 2046 946
rect 2098 937 2110 946
rect 2162 937 2174 946
rect 1913 903 1918 937
rect 2162 903 2167 937
rect 1906 894 1918 903
rect 1970 894 1982 903
rect 2034 894 2046 903
rect 2098 894 2110 903
rect 2162 894 2174 903
rect 2226 894 2238 946
rect 2290 894 2302 946
rect 2354 894 2366 946
rect 2418 894 2430 946
rect 2482 937 2494 946
rect 2546 937 2558 946
rect 2610 937 2622 946
rect 2674 937 2686 946
rect 2738 937 2750 946
rect 2489 903 2494 937
rect 2738 903 2743 937
rect 2482 894 2494 903
rect 2546 894 2558 903
rect 2610 894 2622 903
rect 2674 894 2686 903
rect 2738 894 2750 903
rect 2802 894 2814 946
rect 2866 894 2878 946
rect 2930 894 2942 946
rect 2994 894 3006 946
rect 3058 937 3070 946
rect 3122 937 3134 946
rect 3186 937 3198 946
rect 3250 937 3262 946
rect 3314 937 3326 946
rect 3065 903 3070 937
rect 3314 903 3319 937
rect 3058 894 3070 903
rect 3122 894 3134 903
rect 3186 894 3198 903
rect 3250 894 3262 903
rect 3314 894 3326 903
rect 3378 894 3390 946
rect 3442 894 3454 946
rect 3506 894 3518 946
rect 3570 894 3582 946
rect 3634 937 3646 946
rect 3698 937 3710 946
rect 3762 937 3774 946
rect 3826 937 3838 946
rect 3890 937 3902 946
rect 3641 903 3646 937
rect 3890 903 3895 937
rect 3634 894 3646 903
rect 3698 894 3710 903
rect 3762 894 3774 903
rect 3826 894 3838 903
rect 3890 894 3902 903
rect 3954 894 3966 946
rect 4018 894 4040 946
rect 40 880 4040 894
rect 4160 946 4240 1063
rect 4160 894 4174 946
rect 4226 894 4240 946
rect 4160 777 4240 894
rect 4160 743 4183 777
rect 4217 743 4240 777
rect -160 94 -146 146
rect -94 94 -80 146
rect -160 -23 -80 94
rect 40 146 4040 160
rect 40 94 62 146
rect 114 94 126 146
rect 178 137 190 146
rect 242 137 254 146
rect 306 137 318 146
rect 370 137 382 146
rect 434 137 446 146
rect 185 103 190 137
rect 434 103 439 137
rect 178 94 190 103
rect 242 94 254 103
rect 306 94 318 103
rect 370 94 382 103
rect 434 94 446 103
rect 498 94 510 146
rect 562 94 574 146
rect 626 94 638 146
rect 690 94 702 146
rect 754 137 766 146
rect 818 137 830 146
rect 882 137 894 146
rect 946 137 958 146
rect 1010 137 1022 146
rect 761 103 766 137
rect 1010 103 1015 137
rect 754 94 766 103
rect 818 94 830 103
rect 882 94 894 103
rect 946 94 958 103
rect 1010 94 1022 103
rect 1074 94 1086 146
rect 1138 94 1150 146
rect 1202 94 1214 146
rect 1266 94 1278 146
rect 1330 137 1342 146
rect 1394 137 1406 146
rect 1458 137 1470 146
rect 1522 137 1534 146
rect 1586 137 1598 146
rect 1337 103 1342 137
rect 1586 103 1591 137
rect 1330 94 1342 103
rect 1394 94 1406 103
rect 1458 94 1470 103
rect 1522 94 1534 103
rect 1586 94 1598 103
rect 1650 94 1662 146
rect 1714 94 1726 146
rect 1778 94 1790 146
rect 1842 94 1854 146
rect 1906 137 1918 146
rect 1970 137 1982 146
rect 2034 137 2046 146
rect 2098 137 2110 146
rect 2162 137 2174 146
rect 1913 103 1918 137
rect 2162 103 2167 137
rect 1906 94 1918 103
rect 1970 94 1982 103
rect 2034 94 2046 103
rect 2098 94 2110 103
rect 2162 94 2174 103
rect 2226 94 2238 146
rect 2290 94 2302 146
rect 2354 94 2366 146
rect 2418 94 2430 146
rect 2482 137 2494 146
rect 2546 137 2558 146
rect 2610 137 2622 146
rect 2674 137 2686 146
rect 2738 137 2750 146
rect 2489 103 2494 137
rect 2738 103 2743 137
rect 2482 94 2494 103
rect 2546 94 2558 103
rect 2610 94 2622 103
rect 2674 94 2686 103
rect 2738 94 2750 103
rect 2802 94 2814 146
rect 2866 94 2878 146
rect 2930 94 2942 146
rect 2994 94 3006 146
rect 3058 137 3070 146
rect 3122 137 3134 146
rect 3186 137 3198 146
rect 3250 137 3262 146
rect 3314 137 3326 146
rect 3065 103 3070 137
rect 3314 103 3319 137
rect 3058 94 3070 103
rect 3122 94 3134 103
rect 3186 94 3198 103
rect 3250 94 3262 103
rect 3314 94 3326 103
rect 3378 94 3390 146
rect 3442 94 3454 146
rect 3506 94 3518 146
rect 3570 94 3582 146
rect 3634 137 3646 146
rect 3698 137 3710 146
rect 3762 137 3774 146
rect 3826 137 3838 146
rect 3890 137 3902 146
rect 3641 103 3646 137
rect 3890 103 3895 137
rect 3634 94 3646 103
rect 3698 94 3710 103
rect 3762 94 3774 103
rect 3826 94 3838 103
rect 3890 94 3902 103
rect 3954 94 3966 146
rect 4018 94 4040 146
rect 40 80 4040 94
rect -160 -57 -137 -23
rect -103 -57 -80 -23
rect -160 -343 -80 -57
rect 4160 -23 4240 743
rect 4160 -57 4183 -23
rect 4217 -57 4240 -23
rect 40 -174 4040 -160
rect 40 -226 62 -174
rect 114 -226 126 -174
rect 178 -183 190 -174
rect 242 -183 254 -174
rect 306 -183 318 -174
rect 370 -183 382 -174
rect 434 -183 446 -174
rect 185 -217 190 -183
rect 434 -217 439 -183
rect 178 -226 190 -217
rect 242 -226 254 -217
rect 306 -226 318 -217
rect 370 -226 382 -217
rect 434 -226 446 -217
rect 498 -226 510 -174
rect 562 -226 574 -174
rect 626 -226 638 -174
rect 690 -226 702 -174
rect 754 -183 766 -174
rect 818 -183 830 -174
rect 882 -183 894 -174
rect 946 -183 958 -174
rect 1010 -183 1022 -174
rect 761 -217 766 -183
rect 1010 -217 1015 -183
rect 754 -226 766 -217
rect 818 -226 830 -217
rect 882 -226 894 -217
rect 946 -226 958 -217
rect 1010 -226 1022 -217
rect 1074 -226 1086 -174
rect 1138 -226 1150 -174
rect 1202 -226 1214 -174
rect 1266 -226 1278 -174
rect 1330 -183 1342 -174
rect 1394 -183 1406 -174
rect 1458 -183 1470 -174
rect 1522 -183 1534 -174
rect 1586 -183 1598 -174
rect 1337 -217 1342 -183
rect 1586 -217 1591 -183
rect 1330 -226 1342 -217
rect 1394 -226 1406 -217
rect 1458 -226 1470 -217
rect 1522 -226 1534 -217
rect 1586 -226 1598 -217
rect 1650 -226 1662 -174
rect 1714 -226 1726 -174
rect 1778 -226 1790 -174
rect 1842 -226 1854 -174
rect 1906 -183 1918 -174
rect 1970 -183 1982 -174
rect 2034 -183 2046 -174
rect 2098 -183 2110 -174
rect 2162 -183 2174 -174
rect 1913 -217 1918 -183
rect 2162 -217 2167 -183
rect 1906 -226 1918 -217
rect 1970 -226 1982 -217
rect 2034 -226 2046 -217
rect 2098 -226 2110 -217
rect 2162 -226 2174 -217
rect 2226 -226 2238 -174
rect 2290 -226 2302 -174
rect 2354 -226 2366 -174
rect 2418 -226 2430 -174
rect 2482 -183 2494 -174
rect 2546 -183 2558 -174
rect 2610 -183 2622 -174
rect 2674 -183 2686 -174
rect 2738 -183 2750 -174
rect 2489 -217 2494 -183
rect 2738 -217 2743 -183
rect 2482 -226 2494 -217
rect 2546 -226 2558 -217
rect 2610 -226 2622 -217
rect 2674 -226 2686 -217
rect 2738 -226 2750 -217
rect 2802 -226 2814 -174
rect 2866 -226 2878 -174
rect 2930 -226 2942 -174
rect 2994 -226 3006 -174
rect 3058 -183 3070 -174
rect 3122 -183 3134 -174
rect 3186 -183 3198 -174
rect 3250 -183 3262 -174
rect 3314 -183 3326 -174
rect 3065 -217 3070 -183
rect 3314 -217 3319 -183
rect 3058 -226 3070 -217
rect 3122 -226 3134 -217
rect 3186 -226 3198 -217
rect 3250 -226 3262 -217
rect 3314 -226 3326 -217
rect 3378 -226 3390 -174
rect 3442 -226 3454 -174
rect 3506 -226 3518 -174
rect 3570 -226 3582 -174
rect 3634 -183 3646 -174
rect 3698 -183 3710 -174
rect 3762 -183 3774 -174
rect 3826 -183 3838 -174
rect 3890 -183 3902 -174
rect 3641 -217 3646 -183
rect 3890 -217 3895 -183
rect 3634 -226 3646 -217
rect 3698 -226 3710 -217
rect 3762 -226 3774 -217
rect 3826 -226 3838 -217
rect 3890 -226 3902 -217
rect 3954 -226 3966 -174
rect 4018 -226 4040 -174
rect 40 -240 4040 -226
rect -160 -377 -137 -343
rect -103 -377 -80 -343
rect -160 -400 -80 -377
rect 4160 -343 4240 -57
rect 4160 -377 4183 -343
rect 4217 -377 4240 -343
rect 4160 -400 4240 -377
rect 8320 1417 8400 1440
rect 8320 1383 8343 1417
rect 8377 1383 8400 1417
rect 8320 1097 8400 1383
rect 12640 1417 12720 1440
rect 12640 1383 12663 1417
rect 12697 1383 12720 1417
rect 8520 1266 12520 1280
rect 8520 1214 8542 1266
rect 8594 1214 8606 1266
rect 8658 1257 8670 1266
rect 8722 1257 8734 1266
rect 8786 1257 8798 1266
rect 8850 1257 8862 1266
rect 8914 1257 8926 1266
rect 8665 1223 8670 1257
rect 8914 1223 8919 1257
rect 8658 1214 8670 1223
rect 8722 1214 8734 1223
rect 8786 1214 8798 1223
rect 8850 1214 8862 1223
rect 8914 1214 8926 1223
rect 8978 1214 8990 1266
rect 9042 1214 9054 1266
rect 9106 1214 9118 1266
rect 9170 1214 9182 1266
rect 9234 1257 9246 1266
rect 9298 1257 9310 1266
rect 9362 1257 9374 1266
rect 9426 1257 9438 1266
rect 9490 1257 9502 1266
rect 9241 1223 9246 1257
rect 9490 1223 9495 1257
rect 9234 1214 9246 1223
rect 9298 1214 9310 1223
rect 9362 1214 9374 1223
rect 9426 1214 9438 1223
rect 9490 1214 9502 1223
rect 9554 1214 9566 1266
rect 9618 1214 9630 1266
rect 9682 1214 9694 1266
rect 9746 1214 9758 1266
rect 9810 1257 9822 1266
rect 9874 1257 9886 1266
rect 9938 1257 9950 1266
rect 10002 1257 10014 1266
rect 10066 1257 10078 1266
rect 9817 1223 9822 1257
rect 10066 1223 10071 1257
rect 9810 1214 9822 1223
rect 9874 1214 9886 1223
rect 9938 1214 9950 1223
rect 10002 1214 10014 1223
rect 10066 1214 10078 1223
rect 10130 1214 10142 1266
rect 10194 1214 10206 1266
rect 10258 1214 10270 1266
rect 10322 1214 10334 1266
rect 10386 1257 10398 1266
rect 10450 1257 10462 1266
rect 10514 1257 10526 1266
rect 10578 1257 10590 1266
rect 10642 1257 10654 1266
rect 10393 1223 10398 1257
rect 10642 1223 10647 1257
rect 10386 1214 10398 1223
rect 10450 1214 10462 1223
rect 10514 1214 10526 1223
rect 10578 1214 10590 1223
rect 10642 1214 10654 1223
rect 10706 1214 10718 1266
rect 10770 1214 10782 1266
rect 10834 1214 10846 1266
rect 10898 1214 10910 1266
rect 10962 1257 10974 1266
rect 11026 1257 11038 1266
rect 11090 1257 11102 1266
rect 11154 1257 11166 1266
rect 11218 1257 11230 1266
rect 10969 1223 10974 1257
rect 11218 1223 11223 1257
rect 10962 1214 10974 1223
rect 11026 1214 11038 1223
rect 11090 1214 11102 1223
rect 11154 1214 11166 1223
rect 11218 1214 11230 1223
rect 11282 1214 11294 1266
rect 11346 1214 11358 1266
rect 11410 1214 11422 1266
rect 11474 1214 11486 1266
rect 11538 1257 11550 1266
rect 11602 1257 11614 1266
rect 11666 1257 11678 1266
rect 11730 1257 11742 1266
rect 11794 1257 11806 1266
rect 11545 1223 11550 1257
rect 11794 1223 11799 1257
rect 11538 1214 11550 1223
rect 11602 1214 11614 1223
rect 11666 1214 11678 1223
rect 11730 1214 11742 1223
rect 11794 1214 11806 1223
rect 11858 1214 11870 1266
rect 11922 1214 11934 1266
rect 11986 1214 11998 1266
rect 12050 1214 12062 1266
rect 12114 1257 12126 1266
rect 12178 1257 12190 1266
rect 12242 1257 12254 1266
rect 12306 1257 12318 1266
rect 12370 1257 12382 1266
rect 12121 1223 12126 1257
rect 12370 1223 12375 1257
rect 12114 1214 12126 1223
rect 12178 1214 12190 1223
rect 12242 1214 12254 1223
rect 12306 1214 12318 1223
rect 12370 1214 12382 1223
rect 12434 1214 12446 1266
rect 12498 1214 12520 1266
rect 8520 1200 12520 1214
rect 8320 1063 8343 1097
rect 8377 1063 8400 1097
rect 8320 946 8400 1063
rect 12640 1097 12720 1383
rect 12640 1063 12663 1097
rect 12697 1063 12720 1097
rect 8320 894 8334 946
rect 8386 894 8400 946
rect 8320 777 8400 894
rect 8520 946 12520 960
rect 8520 894 8542 946
rect 8594 894 8606 946
rect 8658 937 8670 946
rect 8722 937 8734 946
rect 8786 937 8798 946
rect 8850 937 8862 946
rect 8914 937 8926 946
rect 8665 903 8670 937
rect 8914 903 8919 937
rect 8658 894 8670 903
rect 8722 894 8734 903
rect 8786 894 8798 903
rect 8850 894 8862 903
rect 8914 894 8926 903
rect 8978 894 8990 946
rect 9042 894 9054 946
rect 9106 894 9118 946
rect 9170 894 9182 946
rect 9234 937 9246 946
rect 9298 937 9310 946
rect 9362 937 9374 946
rect 9426 937 9438 946
rect 9490 937 9502 946
rect 9241 903 9246 937
rect 9490 903 9495 937
rect 9234 894 9246 903
rect 9298 894 9310 903
rect 9362 894 9374 903
rect 9426 894 9438 903
rect 9490 894 9502 903
rect 9554 894 9566 946
rect 9618 894 9630 946
rect 9682 894 9694 946
rect 9746 894 9758 946
rect 9810 937 9822 946
rect 9874 937 9886 946
rect 9938 937 9950 946
rect 10002 937 10014 946
rect 10066 937 10078 946
rect 9817 903 9822 937
rect 10066 903 10071 937
rect 9810 894 9822 903
rect 9874 894 9886 903
rect 9938 894 9950 903
rect 10002 894 10014 903
rect 10066 894 10078 903
rect 10130 894 10142 946
rect 10194 894 10206 946
rect 10258 894 10270 946
rect 10322 894 10334 946
rect 10386 937 10398 946
rect 10450 937 10462 946
rect 10514 937 10526 946
rect 10578 937 10590 946
rect 10642 937 10654 946
rect 10393 903 10398 937
rect 10642 903 10647 937
rect 10386 894 10398 903
rect 10450 894 10462 903
rect 10514 894 10526 903
rect 10578 894 10590 903
rect 10642 894 10654 903
rect 10706 894 10718 946
rect 10770 894 10782 946
rect 10834 894 10846 946
rect 10898 894 10910 946
rect 10962 937 10974 946
rect 11026 937 11038 946
rect 11090 937 11102 946
rect 11154 937 11166 946
rect 11218 937 11230 946
rect 10969 903 10974 937
rect 11218 903 11223 937
rect 10962 894 10974 903
rect 11026 894 11038 903
rect 11090 894 11102 903
rect 11154 894 11166 903
rect 11218 894 11230 903
rect 11282 894 11294 946
rect 11346 894 11358 946
rect 11410 894 11422 946
rect 11474 894 11486 946
rect 11538 937 11550 946
rect 11602 937 11614 946
rect 11666 937 11678 946
rect 11730 937 11742 946
rect 11794 937 11806 946
rect 11545 903 11550 937
rect 11794 903 11799 937
rect 11538 894 11550 903
rect 11602 894 11614 903
rect 11666 894 11678 903
rect 11730 894 11742 903
rect 11794 894 11806 903
rect 11858 894 11870 946
rect 11922 894 11934 946
rect 11986 894 11998 946
rect 12050 894 12062 946
rect 12114 937 12126 946
rect 12178 937 12190 946
rect 12242 937 12254 946
rect 12306 937 12318 946
rect 12370 937 12382 946
rect 12121 903 12126 937
rect 12370 903 12375 937
rect 12114 894 12126 903
rect 12178 894 12190 903
rect 12242 894 12254 903
rect 12306 894 12318 903
rect 12370 894 12382 903
rect 12434 894 12446 946
rect 12498 894 12520 946
rect 8520 880 12520 894
rect 8320 743 8343 777
rect 8377 743 8400 777
rect 8320 -23 8400 743
rect 8520 146 12520 160
rect 8520 94 8542 146
rect 8594 94 8606 146
rect 8658 137 8670 146
rect 8722 137 8734 146
rect 8786 137 8798 146
rect 8850 137 8862 146
rect 8914 137 8926 146
rect 8665 103 8670 137
rect 8914 103 8919 137
rect 8658 94 8670 103
rect 8722 94 8734 103
rect 8786 94 8798 103
rect 8850 94 8862 103
rect 8914 94 8926 103
rect 8978 94 8990 146
rect 9042 94 9054 146
rect 9106 94 9118 146
rect 9170 94 9182 146
rect 9234 137 9246 146
rect 9298 137 9310 146
rect 9362 137 9374 146
rect 9426 137 9438 146
rect 9490 137 9502 146
rect 9241 103 9246 137
rect 9490 103 9495 137
rect 9234 94 9246 103
rect 9298 94 9310 103
rect 9362 94 9374 103
rect 9426 94 9438 103
rect 9490 94 9502 103
rect 9554 94 9566 146
rect 9618 94 9630 146
rect 9682 94 9694 146
rect 9746 94 9758 146
rect 9810 137 9822 146
rect 9874 137 9886 146
rect 9938 137 9950 146
rect 10002 137 10014 146
rect 10066 137 10078 146
rect 9817 103 9822 137
rect 10066 103 10071 137
rect 9810 94 9822 103
rect 9874 94 9886 103
rect 9938 94 9950 103
rect 10002 94 10014 103
rect 10066 94 10078 103
rect 10130 94 10142 146
rect 10194 94 10206 146
rect 10258 94 10270 146
rect 10322 94 10334 146
rect 10386 137 10398 146
rect 10450 137 10462 146
rect 10514 137 10526 146
rect 10578 137 10590 146
rect 10642 137 10654 146
rect 10393 103 10398 137
rect 10642 103 10647 137
rect 10386 94 10398 103
rect 10450 94 10462 103
rect 10514 94 10526 103
rect 10578 94 10590 103
rect 10642 94 10654 103
rect 10706 94 10718 146
rect 10770 94 10782 146
rect 10834 94 10846 146
rect 10898 94 10910 146
rect 10962 137 10974 146
rect 11026 137 11038 146
rect 11090 137 11102 146
rect 11154 137 11166 146
rect 11218 137 11230 146
rect 10969 103 10974 137
rect 11218 103 11223 137
rect 10962 94 10974 103
rect 11026 94 11038 103
rect 11090 94 11102 103
rect 11154 94 11166 103
rect 11218 94 11230 103
rect 11282 94 11294 146
rect 11346 94 11358 146
rect 11410 94 11422 146
rect 11474 94 11486 146
rect 11538 137 11550 146
rect 11602 137 11614 146
rect 11666 137 11678 146
rect 11730 137 11742 146
rect 11794 137 11806 146
rect 11545 103 11550 137
rect 11794 103 11799 137
rect 11538 94 11550 103
rect 11602 94 11614 103
rect 11666 94 11678 103
rect 11730 94 11742 103
rect 11794 94 11806 103
rect 11858 94 11870 146
rect 11922 94 11934 146
rect 11986 94 11998 146
rect 12050 94 12062 146
rect 12114 137 12126 146
rect 12178 137 12190 146
rect 12242 137 12254 146
rect 12306 137 12318 146
rect 12370 137 12382 146
rect 12121 103 12126 137
rect 12370 103 12375 137
rect 12114 94 12126 103
rect 12178 94 12190 103
rect 12242 94 12254 103
rect 12306 94 12318 103
rect 12370 94 12382 103
rect 12434 94 12446 146
rect 12498 94 12520 146
rect 8520 80 12520 94
rect 12640 146 12720 1063
rect 12640 94 12654 146
rect 12706 94 12720 146
rect 8320 -57 8343 -23
rect 8377 -57 8400 -23
rect 8320 -343 8400 -57
rect 12640 -23 12720 94
rect 12640 -57 12663 -23
rect 12697 -57 12720 -23
rect 8520 -174 12520 -160
rect 8520 -226 8542 -174
rect 8594 -226 8606 -174
rect 8658 -183 8670 -174
rect 8722 -183 8734 -174
rect 8786 -183 8798 -174
rect 8850 -183 8862 -174
rect 8914 -183 8926 -174
rect 8665 -217 8670 -183
rect 8914 -217 8919 -183
rect 8658 -226 8670 -217
rect 8722 -226 8734 -217
rect 8786 -226 8798 -217
rect 8850 -226 8862 -217
rect 8914 -226 8926 -217
rect 8978 -226 8990 -174
rect 9042 -226 9054 -174
rect 9106 -226 9118 -174
rect 9170 -226 9182 -174
rect 9234 -183 9246 -174
rect 9298 -183 9310 -174
rect 9362 -183 9374 -174
rect 9426 -183 9438 -174
rect 9490 -183 9502 -174
rect 9241 -217 9246 -183
rect 9490 -217 9495 -183
rect 9234 -226 9246 -217
rect 9298 -226 9310 -217
rect 9362 -226 9374 -217
rect 9426 -226 9438 -217
rect 9490 -226 9502 -217
rect 9554 -226 9566 -174
rect 9618 -226 9630 -174
rect 9682 -226 9694 -174
rect 9746 -226 9758 -174
rect 9810 -183 9822 -174
rect 9874 -183 9886 -174
rect 9938 -183 9950 -174
rect 10002 -183 10014 -174
rect 10066 -183 10078 -174
rect 9817 -217 9822 -183
rect 10066 -217 10071 -183
rect 9810 -226 9822 -217
rect 9874 -226 9886 -217
rect 9938 -226 9950 -217
rect 10002 -226 10014 -217
rect 10066 -226 10078 -217
rect 10130 -226 10142 -174
rect 10194 -226 10206 -174
rect 10258 -226 10270 -174
rect 10322 -226 10334 -174
rect 10386 -183 10398 -174
rect 10450 -183 10462 -174
rect 10514 -183 10526 -174
rect 10578 -183 10590 -174
rect 10642 -183 10654 -174
rect 10393 -217 10398 -183
rect 10642 -217 10647 -183
rect 10386 -226 10398 -217
rect 10450 -226 10462 -217
rect 10514 -226 10526 -217
rect 10578 -226 10590 -217
rect 10642 -226 10654 -217
rect 10706 -226 10718 -174
rect 10770 -226 10782 -174
rect 10834 -226 10846 -174
rect 10898 -226 10910 -174
rect 10962 -183 10974 -174
rect 11026 -183 11038 -174
rect 11090 -183 11102 -174
rect 11154 -183 11166 -174
rect 11218 -183 11230 -174
rect 10969 -217 10974 -183
rect 11218 -217 11223 -183
rect 10962 -226 10974 -217
rect 11026 -226 11038 -217
rect 11090 -226 11102 -217
rect 11154 -226 11166 -217
rect 11218 -226 11230 -217
rect 11282 -226 11294 -174
rect 11346 -226 11358 -174
rect 11410 -226 11422 -174
rect 11474 -226 11486 -174
rect 11538 -183 11550 -174
rect 11602 -183 11614 -174
rect 11666 -183 11678 -174
rect 11730 -183 11742 -174
rect 11794 -183 11806 -174
rect 11545 -217 11550 -183
rect 11794 -217 11799 -183
rect 11538 -226 11550 -217
rect 11602 -226 11614 -217
rect 11666 -226 11678 -217
rect 11730 -226 11742 -217
rect 11794 -226 11806 -217
rect 11858 -226 11870 -174
rect 11922 -226 11934 -174
rect 11986 -226 11998 -174
rect 12050 -226 12062 -174
rect 12114 -183 12126 -174
rect 12178 -183 12190 -174
rect 12242 -183 12254 -174
rect 12306 -183 12318 -174
rect 12370 -183 12382 -174
rect 12121 -217 12126 -183
rect 12370 -217 12375 -183
rect 12114 -226 12126 -217
rect 12178 -226 12190 -217
rect 12242 -226 12254 -217
rect 12306 -226 12318 -217
rect 12370 -226 12382 -217
rect 12434 -226 12446 -174
rect 12498 -226 12520 -174
rect 8520 -240 12520 -226
rect 8320 -377 8343 -343
rect 8377 -377 8400 -343
rect 8320 -400 8400 -377
rect 12640 -343 12720 -57
rect 12640 -377 12663 -343
rect 12697 -377 12720 -343
rect 12640 -400 12720 -377
rect -320 -494 -240 -480
rect -320 -546 -306 -494
rect -254 -546 -240 -494
rect -320 -560 -240 -546
rect 12800 -494 12880 -480
rect 12800 -546 12814 -494
rect 12866 -546 12880 -494
rect 12800 -560 12880 -546
<< via1 >>
rect -306 4137 -254 4146
rect -306 4103 -297 4137
rect -297 4103 -263 4137
rect -263 4103 -254 4137
rect -306 4094 -254 4103
rect 12814 4137 12866 4146
rect 12814 4103 12823 4137
rect 12823 4103 12857 4137
rect 12857 4103 12866 4137
rect 12814 4094 12866 4103
rect 62 3817 114 3826
rect 62 3783 79 3817
rect 79 3783 113 3817
rect 113 3783 114 3817
rect 62 3774 114 3783
rect 126 3817 178 3826
rect 190 3817 242 3826
rect 254 3817 306 3826
rect 318 3817 370 3826
rect 382 3817 434 3826
rect 446 3817 498 3826
rect 126 3783 151 3817
rect 151 3783 178 3817
rect 190 3783 223 3817
rect 223 3783 242 3817
rect 254 3783 257 3817
rect 257 3783 295 3817
rect 295 3783 306 3817
rect 318 3783 329 3817
rect 329 3783 367 3817
rect 367 3783 370 3817
rect 382 3783 401 3817
rect 401 3783 434 3817
rect 446 3783 473 3817
rect 473 3783 498 3817
rect 126 3774 178 3783
rect 190 3774 242 3783
rect 254 3774 306 3783
rect 318 3774 370 3783
rect 382 3774 434 3783
rect 446 3774 498 3783
rect 510 3817 562 3826
rect 510 3783 511 3817
rect 511 3783 545 3817
rect 545 3783 562 3817
rect 510 3774 562 3783
rect 574 3817 626 3826
rect 574 3783 583 3817
rect 583 3783 617 3817
rect 617 3783 626 3817
rect 574 3774 626 3783
rect 638 3817 690 3826
rect 638 3783 655 3817
rect 655 3783 689 3817
rect 689 3783 690 3817
rect 638 3774 690 3783
rect 702 3817 754 3826
rect 766 3817 818 3826
rect 830 3817 882 3826
rect 894 3817 946 3826
rect 958 3817 1010 3826
rect 1022 3817 1074 3826
rect 702 3783 727 3817
rect 727 3783 754 3817
rect 766 3783 799 3817
rect 799 3783 818 3817
rect 830 3783 833 3817
rect 833 3783 871 3817
rect 871 3783 882 3817
rect 894 3783 905 3817
rect 905 3783 943 3817
rect 943 3783 946 3817
rect 958 3783 977 3817
rect 977 3783 1010 3817
rect 1022 3783 1049 3817
rect 1049 3783 1074 3817
rect 702 3774 754 3783
rect 766 3774 818 3783
rect 830 3774 882 3783
rect 894 3774 946 3783
rect 958 3774 1010 3783
rect 1022 3774 1074 3783
rect 1086 3817 1138 3826
rect 1086 3783 1087 3817
rect 1087 3783 1121 3817
rect 1121 3783 1138 3817
rect 1086 3774 1138 3783
rect 1150 3817 1202 3826
rect 1150 3783 1159 3817
rect 1159 3783 1193 3817
rect 1193 3783 1202 3817
rect 1150 3774 1202 3783
rect 1214 3817 1266 3826
rect 1214 3783 1231 3817
rect 1231 3783 1265 3817
rect 1265 3783 1266 3817
rect 1214 3774 1266 3783
rect 1278 3817 1330 3826
rect 1342 3817 1394 3826
rect 1406 3817 1458 3826
rect 1470 3817 1522 3826
rect 1534 3817 1586 3826
rect 1598 3817 1650 3826
rect 1278 3783 1303 3817
rect 1303 3783 1330 3817
rect 1342 3783 1375 3817
rect 1375 3783 1394 3817
rect 1406 3783 1409 3817
rect 1409 3783 1447 3817
rect 1447 3783 1458 3817
rect 1470 3783 1481 3817
rect 1481 3783 1519 3817
rect 1519 3783 1522 3817
rect 1534 3783 1553 3817
rect 1553 3783 1586 3817
rect 1598 3783 1625 3817
rect 1625 3783 1650 3817
rect 1278 3774 1330 3783
rect 1342 3774 1394 3783
rect 1406 3774 1458 3783
rect 1470 3774 1522 3783
rect 1534 3774 1586 3783
rect 1598 3774 1650 3783
rect 1662 3817 1714 3826
rect 1662 3783 1663 3817
rect 1663 3783 1697 3817
rect 1697 3783 1714 3817
rect 1662 3774 1714 3783
rect 1726 3817 1778 3826
rect 1726 3783 1735 3817
rect 1735 3783 1769 3817
rect 1769 3783 1778 3817
rect 1726 3774 1778 3783
rect 1790 3817 1842 3826
rect 1790 3783 1807 3817
rect 1807 3783 1841 3817
rect 1841 3783 1842 3817
rect 1790 3774 1842 3783
rect 1854 3817 1906 3826
rect 1918 3817 1970 3826
rect 1982 3817 2034 3826
rect 2046 3817 2098 3826
rect 2110 3817 2162 3826
rect 2174 3817 2226 3826
rect 1854 3783 1879 3817
rect 1879 3783 1906 3817
rect 1918 3783 1951 3817
rect 1951 3783 1970 3817
rect 1982 3783 1985 3817
rect 1985 3783 2023 3817
rect 2023 3783 2034 3817
rect 2046 3783 2057 3817
rect 2057 3783 2095 3817
rect 2095 3783 2098 3817
rect 2110 3783 2129 3817
rect 2129 3783 2162 3817
rect 2174 3783 2201 3817
rect 2201 3783 2226 3817
rect 1854 3774 1906 3783
rect 1918 3774 1970 3783
rect 1982 3774 2034 3783
rect 2046 3774 2098 3783
rect 2110 3774 2162 3783
rect 2174 3774 2226 3783
rect 2238 3817 2290 3826
rect 2238 3783 2239 3817
rect 2239 3783 2273 3817
rect 2273 3783 2290 3817
rect 2238 3774 2290 3783
rect 2302 3817 2354 3826
rect 2302 3783 2311 3817
rect 2311 3783 2345 3817
rect 2345 3783 2354 3817
rect 2302 3774 2354 3783
rect 2366 3817 2418 3826
rect 2366 3783 2383 3817
rect 2383 3783 2417 3817
rect 2417 3783 2418 3817
rect 2366 3774 2418 3783
rect 2430 3817 2482 3826
rect 2494 3817 2546 3826
rect 2558 3817 2610 3826
rect 2622 3817 2674 3826
rect 2686 3817 2738 3826
rect 2750 3817 2802 3826
rect 2430 3783 2455 3817
rect 2455 3783 2482 3817
rect 2494 3783 2527 3817
rect 2527 3783 2546 3817
rect 2558 3783 2561 3817
rect 2561 3783 2599 3817
rect 2599 3783 2610 3817
rect 2622 3783 2633 3817
rect 2633 3783 2671 3817
rect 2671 3783 2674 3817
rect 2686 3783 2705 3817
rect 2705 3783 2738 3817
rect 2750 3783 2777 3817
rect 2777 3783 2802 3817
rect 2430 3774 2482 3783
rect 2494 3774 2546 3783
rect 2558 3774 2610 3783
rect 2622 3774 2674 3783
rect 2686 3774 2738 3783
rect 2750 3774 2802 3783
rect 2814 3817 2866 3826
rect 2814 3783 2815 3817
rect 2815 3783 2849 3817
rect 2849 3783 2866 3817
rect 2814 3774 2866 3783
rect 2878 3817 2930 3826
rect 2878 3783 2887 3817
rect 2887 3783 2921 3817
rect 2921 3783 2930 3817
rect 2878 3774 2930 3783
rect 2942 3817 2994 3826
rect 2942 3783 2959 3817
rect 2959 3783 2993 3817
rect 2993 3783 2994 3817
rect 2942 3774 2994 3783
rect 3006 3817 3058 3826
rect 3070 3817 3122 3826
rect 3134 3817 3186 3826
rect 3198 3817 3250 3826
rect 3262 3817 3314 3826
rect 3326 3817 3378 3826
rect 3006 3783 3031 3817
rect 3031 3783 3058 3817
rect 3070 3783 3103 3817
rect 3103 3783 3122 3817
rect 3134 3783 3137 3817
rect 3137 3783 3175 3817
rect 3175 3783 3186 3817
rect 3198 3783 3209 3817
rect 3209 3783 3247 3817
rect 3247 3783 3250 3817
rect 3262 3783 3281 3817
rect 3281 3783 3314 3817
rect 3326 3783 3353 3817
rect 3353 3783 3378 3817
rect 3006 3774 3058 3783
rect 3070 3774 3122 3783
rect 3134 3774 3186 3783
rect 3198 3774 3250 3783
rect 3262 3774 3314 3783
rect 3326 3774 3378 3783
rect 3390 3817 3442 3826
rect 3390 3783 3391 3817
rect 3391 3783 3425 3817
rect 3425 3783 3442 3817
rect 3390 3774 3442 3783
rect 3454 3817 3506 3826
rect 3454 3783 3463 3817
rect 3463 3783 3497 3817
rect 3497 3783 3506 3817
rect 3454 3774 3506 3783
rect 3518 3817 3570 3826
rect 3518 3783 3535 3817
rect 3535 3783 3569 3817
rect 3569 3783 3570 3817
rect 3518 3774 3570 3783
rect 3582 3817 3634 3826
rect 3646 3817 3698 3826
rect 3710 3817 3762 3826
rect 3774 3817 3826 3826
rect 3838 3817 3890 3826
rect 3902 3817 3954 3826
rect 3582 3783 3607 3817
rect 3607 3783 3634 3817
rect 3646 3783 3679 3817
rect 3679 3783 3698 3817
rect 3710 3783 3713 3817
rect 3713 3783 3751 3817
rect 3751 3783 3762 3817
rect 3774 3783 3785 3817
rect 3785 3783 3823 3817
rect 3823 3783 3826 3817
rect 3838 3783 3857 3817
rect 3857 3783 3890 3817
rect 3902 3783 3929 3817
rect 3929 3783 3954 3817
rect 3582 3774 3634 3783
rect 3646 3774 3698 3783
rect 3710 3774 3762 3783
rect 3774 3774 3826 3783
rect 3838 3774 3890 3783
rect 3902 3774 3954 3783
rect 3966 3817 4018 3826
rect 3966 3783 3967 3817
rect 3967 3783 4001 3817
rect 4001 3783 4018 3817
rect 3966 3774 4018 3783
rect -146 3454 -94 3506
rect 62 3497 114 3506
rect 62 3463 79 3497
rect 79 3463 113 3497
rect 113 3463 114 3497
rect 62 3454 114 3463
rect 126 3497 178 3506
rect 190 3497 242 3506
rect 254 3497 306 3506
rect 318 3497 370 3506
rect 382 3497 434 3506
rect 446 3497 498 3506
rect 126 3463 151 3497
rect 151 3463 178 3497
rect 190 3463 223 3497
rect 223 3463 242 3497
rect 254 3463 257 3497
rect 257 3463 295 3497
rect 295 3463 306 3497
rect 318 3463 329 3497
rect 329 3463 367 3497
rect 367 3463 370 3497
rect 382 3463 401 3497
rect 401 3463 434 3497
rect 446 3463 473 3497
rect 473 3463 498 3497
rect 126 3454 178 3463
rect 190 3454 242 3463
rect 254 3454 306 3463
rect 318 3454 370 3463
rect 382 3454 434 3463
rect 446 3454 498 3463
rect 510 3497 562 3506
rect 510 3463 511 3497
rect 511 3463 545 3497
rect 545 3463 562 3497
rect 510 3454 562 3463
rect 574 3497 626 3506
rect 574 3463 583 3497
rect 583 3463 617 3497
rect 617 3463 626 3497
rect 574 3454 626 3463
rect 638 3497 690 3506
rect 638 3463 655 3497
rect 655 3463 689 3497
rect 689 3463 690 3497
rect 638 3454 690 3463
rect 702 3497 754 3506
rect 766 3497 818 3506
rect 830 3497 882 3506
rect 894 3497 946 3506
rect 958 3497 1010 3506
rect 1022 3497 1074 3506
rect 702 3463 727 3497
rect 727 3463 754 3497
rect 766 3463 799 3497
rect 799 3463 818 3497
rect 830 3463 833 3497
rect 833 3463 871 3497
rect 871 3463 882 3497
rect 894 3463 905 3497
rect 905 3463 943 3497
rect 943 3463 946 3497
rect 958 3463 977 3497
rect 977 3463 1010 3497
rect 1022 3463 1049 3497
rect 1049 3463 1074 3497
rect 702 3454 754 3463
rect 766 3454 818 3463
rect 830 3454 882 3463
rect 894 3454 946 3463
rect 958 3454 1010 3463
rect 1022 3454 1074 3463
rect 1086 3497 1138 3506
rect 1086 3463 1087 3497
rect 1087 3463 1121 3497
rect 1121 3463 1138 3497
rect 1086 3454 1138 3463
rect 1150 3497 1202 3506
rect 1150 3463 1159 3497
rect 1159 3463 1193 3497
rect 1193 3463 1202 3497
rect 1150 3454 1202 3463
rect 1214 3497 1266 3506
rect 1214 3463 1231 3497
rect 1231 3463 1265 3497
rect 1265 3463 1266 3497
rect 1214 3454 1266 3463
rect 1278 3497 1330 3506
rect 1342 3497 1394 3506
rect 1406 3497 1458 3506
rect 1470 3497 1522 3506
rect 1534 3497 1586 3506
rect 1598 3497 1650 3506
rect 1278 3463 1303 3497
rect 1303 3463 1330 3497
rect 1342 3463 1375 3497
rect 1375 3463 1394 3497
rect 1406 3463 1409 3497
rect 1409 3463 1447 3497
rect 1447 3463 1458 3497
rect 1470 3463 1481 3497
rect 1481 3463 1519 3497
rect 1519 3463 1522 3497
rect 1534 3463 1553 3497
rect 1553 3463 1586 3497
rect 1598 3463 1625 3497
rect 1625 3463 1650 3497
rect 1278 3454 1330 3463
rect 1342 3454 1394 3463
rect 1406 3454 1458 3463
rect 1470 3454 1522 3463
rect 1534 3454 1586 3463
rect 1598 3454 1650 3463
rect 1662 3497 1714 3506
rect 1662 3463 1663 3497
rect 1663 3463 1697 3497
rect 1697 3463 1714 3497
rect 1662 3454 1714 3463
rect 1726 3497 1778 3506
rect 1726 3463 1735 3497
rect 1735 3463 1769 3497
rect 1769 3463 1778 3497
rect 1726 3454 1778 3463
rect 1790 3497 1842 3506
rect 1790 3463 1807 3497
rect 1807 3463 1841 3497
rect 1841 3463 1842 3497
rect 1790 3454 1842 3463
rect 1854 3497 1906 3506
rect 1918 3497 1970 3506
rect 1982 3497 2034 3506
rect 2046 3497 2098 3506
rect 2110 3497 2162 3506
rect 2174 3497 2226 3506
rect 1854 3463 1879 3497
rect 1879 3463 1906 3497
rect 1918 3463 1951 3497
rect 1951 3463 1970 3497
rect 1982 3463 1985 3497
rect 1985 3463 2023 3497
rect 2023 3463 2034 3497
rect 2046 3463 2057 3497
rect 2057 3463 2095 3497
rect 2095 3463 2098 3497
rect 2110 3463 2129 3497
rect 2129 3463 2162 3497
rect 2174 3463 2201 3497
rect 2201 3463 2226 3497
rect 1854 3454 1906 3463
rect 1918 3454 1970 3463
rect 1982 3454 2034 3463
rect 2046 3454 2098 3463
rect 2110 3454 2162 3463
rect 2174 3454 2226 3463
rect 2238 3497 2290 3506
rect 2238 3463 2239 3497
rect 2239 3463 2273 3497
rect 2273 3463 2290 3497
rect 2238 3454 2290 3463
rect 2302 3497 2354 3506
rect 2302 3463 2311 3497
rect 2311 3463 2345 3497
rect 2345 3463 2354 3497
rect 2302 3454 2354 3463
rect 2366 3497 2418 3506
rect 2366 3463 2383 3497
rect 2383 3463 2417 3497
rect 2417 3463 2418 3497
rect 2366 3454 2418 3463
rect 2430 3497 2482 3506
rect 2494 3497 2546 3506
rect 2558 3497 2610 3506
rect 2622 3497 2674 3506
rect 2686 3497 2738 3506
rect 2750 3497 2802 3506
rect 2430 3463 2455 3497
rect 2455 3463 2482 3497
rect 2494 3463 2527 3497
rect 2527 3463 2546 3497
rect 2558 3463 2561 3497
rect 2561 3463 2599 3497
rect 2599 3463 2610 3497
rect 2622 3463 2633 3497
rect 2633 3463 2671 3497
rect 2671 3463 2674 3497
rect 2686 3463 2705 3497
rect 2705 3463 2738 3497
rect 2750 3463 2777 3497
rect 2777 3463 2802 3497
rect 2430 3454 2482 3463
rect 2494 3454 2546 3463
rect 2558 3454 2610 3463
rect 2622 3454 2674 3463
rect 2686 3454 2738 3463
rect 2750 3454 2802 3463
rect 2814 3497 2866 3506
rect 2814 3463 2815 3497
rect 2815 3463 2849 3497
rect 2849 3463 2866 3497
rect 2814 3454 2866 3463
rect 2878 3497 2930 3506
rect 2878 3463 2887 3497
rect 2887 3463 2921 3497
rect 2921 3463 2930 3497
rect 2878 3454 2930 3463
rect 2942 3497 2994 3506
rect 2942 3463 2959 3497
rect 2959 3463 2993 3497
rect 2993 3463 2994 3497
rect 2942 3454 2994 3463
rect 3006 3497 3058 3506
rect 3070 3497 3122 3506
rect 3134 3497 3186 3506
rect 3198 3497 3250 3506
rect 3262 3497 3314 3506
rect 3326 3497 3378 3506
rect 3006 3463 3031 3497
rect 3031 3463 3058 3497
rect 3070 3463 3103 3497
rect 3103 3463 3122 3497
rect 3134 3463 3137 3497
rect 3137 3463 3175 3497
rect 3175 3463 3186 3497
rect 3198 3463 3209 3497
rect 3209 3463 3247 3497
rect 3247 3463 3250 3497
rect 3262 3463 3281 3497
rect 3281 3463 3314 3497
rect 3326 3463 3353 3497
rect 3353 3463 3378 3497
rect 3006 3454 3058 3463
rect 3070 3454 3122 3463
rect 3134 3454 3186 3463
rect 3198 3454 3250 3463
rect 3262 3454 3314 3463
rect 3326 3454 3378 3463
rect 3390 3497 3442 3506
rect 3390 3463 3391 3497
rect 3391 3463 3425 3497
rect 3425 3463 3442 3497
rect 3390 3454 3442 3463
rect 3454 3497 3506 3506
rect 3454 3463 3463 3497
rect 3463 3463 3497 3497
rect 3497 3463 3506 3497
rect 3454 3454 3506 3463
rect 3518 3497 3570 3506
rect 3518 3463 3535 3497
rect 3535 3463 3569 3497
rect 3569 3463 3570 3497
rect 3518 3454 3570 3463
rect 3582 3497 3634 3506
rect 3646 3497 3698 3506
rect 3710 3497 3762 3506
rect 3774 3497 3826 3506
rect 3838 3497 3890 3506
rect 3902 3497 3954 3506
rect 3582 3463 3607 3497
rect 3607 3463 3634 3497
rect 3646 3463 3679 3497
rect 3679 3463 3698 3497
rect 3710 3463 3713 3497
rect 3713 3463 3751 3497
rect 3751 3463 3762 3497
rect 3774 3463 3785 3497
rect 3785 3463 3823 3497
rect 3823 3463 3826 3497
rect 3838 3463 3857 3497
rect 3857 3463 3890 3497
rect 3902 3463 3929 3497
rect 3929 3463 3954 3497
rect 3582 3454 3634 3463
rect 3646 3454 3698 3463
rect 3710 3454 3762 3463
rect 3774 3454 3826 3463
rect 3838 3454 3890 3463
rect 3902 3454 3954 3463
rect 3966 3497 4018 3506
rect 3966 3463 3967 3497
rect 3967 3463 4001 3497
rect 4001 3463 4018 3497
rect 3966 3454 4018 3463
rect 62 2697 114 2706
rect 62 2663 79 2697
rect 79 2663 113 2697
rect 113 2663 114 2697
rect 62 2654 114 2663
rect 126 2697 178 2706
rect 190 2697 242 2706
rect 254 2697 306 2706
rect 318 2697 370 2706
rect 382 2697 434 2706
rect 446 2697 498 2706
rect 126 2663 151 2697
rect 151 2663 178 2697
rect 190 2663 223 2697
rect 223 2663 242 2697
rect 254 2663 257 2697
rect 257 2663 295 2697
rect 295 2663 306 2697
rect 318 2663 329 2697
rect 329 2663 367 2697
rect 367 2663 370 2697
rect 382 2663 401 2697
rect 401 2663 434 2697
rect 446 2663 473 2697
rect 473 2663 498 2697
rect 126 2654 178 2663
rect 190 2654 242 2663
rect 254 2654 306 2663
rect 318 2654 370 2663
rect 382 2654 434 2663
rect 446 2654 498 2663
rect 510 2697 562 2706
rect 510 2663 511 2697
rect 511 2663 545 2697
rect 545 2663 562 2697
rect 510 2654 562 2663
rect 574 2697 626 2706
rect 574 2663 583 2697
rect 583 2663 617 2697
rect 617 2663 626 2697
rect 574 2654 626 2663
rect 638 2697 690 2706
rect 638 2663 655 2697
rect 655 2663 689 2697
rect 689 2663 690 2697
rect 638 2654 690 2663
rect 702 2697 754 2706
rect 766 2697 818 2706
rect 830 2697 882 2706
rect 894 2697 946 2706
rect 958 2697 1010 2706
rect 1022 2697 1074 2706
rect 702 2663 727 2697
rect 727 2663 754 2697
rect 766 2663 799 2697
rect 799 2663 818 2697
rect 830 2663 833 2697
rect 833 2663 871 2697
rect 871 2663 882 2697
rect 894 2663 905 2697
rect 905 2663 943 2697
rect 943 2663 946 2697
rect 958 2663 977 2697
rect 977 2663 1010 2697
rect 1022 2663 1049 2697
rect 1049 2663 1074 2697
rect 702 2654 754 2663
rect 766 2654 818 2663
rect 830 2654 882 2663
rect 894 2654 946 2663
rect 958 2654 1010 2663
rect 1022 2654 1074 2663
rect 1086 2697 1138 2706
rect 1086 2663 1087 2697
rect 1087 2663 1121 2697
rect 1121 2663 1138 2697
rect 1086 2654 1138 2663
rect 1150 2697 1202 2706
rect 1150 2663 1159 2697
rect 1159 2663 1193 2697
rect 1193 2663 1202 2697
rect 1150 2654 1202 2663
rect 1214 2697 1266 2706
rect 1214 2663 1231 2697
rect 1231 2663 1265 2697
rect 1265 2663 1266 2697
rect 1214 2654 1266 2663
rect 1278 2697 1330 2706
rect 1342 2697 1394 2706
rect 1406 2697 1458 2706
rect 1470 2697 1522 2706
rect 1534 2697 1586 2706
rect 1598 2697 1650 2706
rect 1278 2663 1303 2697
rect 1303 2663 1330 2697
rect 1342 2663 1375 2697
rect 1375 2663 1394 2697
rect 1406 2663 1409 2697
rect 1409 2663 1447 2697
rect 1447 2663 1458 2697
rect 1470 2663 1481 2697
rect 1481 2663 1519 2697
rect 1519 2663 1522 2697
rect 1534 2663 1553 2697
rect 1553 2663 1586 2697
rect 1598 2663 1625 2697
rect 1625 2663 1650 2697
rect 1278 2654 1330 2663
rect 1342 2654 1394 2663
rect 1406 2654 1458 2663
rect 1470 2654 1522 2663
rect 1534 2654 1586 2663
rect 1598 2654 1650 2663
rect 1662 2697 1714 2706
rect 1662 2663 1663 2697
rect 1663 2663 1697 2697
rect 1697 2663 1714 2697
rect 1662 2654 1714 2663
rect 1726 2697 1778 2706
rect 1726 2663 1735 2697
rect 1735 2663 1769 2697
rect 1769 2663 1778 2697
rect 1726 2654 1778 2663
rect 1790 2697 1842 2706
rect 1790 2663 1807 2697
rect 1807 2663 1841 2697
rect 1841 2663 1842 2697
rect 1790 2654 1842 2663
rect 1854 2697 1906 2706
rect 1918 2697 1970 2706
rect 1982 2697 2034 2706
rect 2046 2697 2098 2706
rect 2110 2697 2162 2706
rect 2174 2697 2226 2706
rect 1854 2663 1879 2697
rect 1879 2663 1906 2697
rect 1918 2663 1951 2697
rect 1951 2663 1970 2697
rect 1982 2663 1985 2697
rect 1985 2663 2023 2697
rect 2023 2663 2034 2697
rect 2046 2663 2057 2697
rect 2057 2663 2095 2697
rect 2095 2663 2098 2697
rect 2110 2663 2129 2697
rect 2129 2663 2162 2697
rect 2174 2663 2201 2697
rect 2201 2663 2226 2697
rect 1854 2654 1906 2663
rect 1918 2654 1970 2663
rect 1982 2654 2034 2663
rect 2046 2654 2098 2663
rect 2110 2654 2162 2663
rect 2174 2654 2226 2663
rect 2238 2697 2290 2706
rect 2238 2663 2239 2697
rect 2239 2663 2273 2697
rect 2273 2663 2290 2697
rect 2238 2654 2290 2663
rect 2302 2697 2354 2706
rect 2302 2663 2311 2697
rect 2311 2663 2345 2697
rect 2345 2663 2354 2697
rect 2302 2654 2354 2663
rect 2366 2697 2418 2706
rect 2366 2663 2383 2697
rect 2383 2663 2417 2697
rect 2417 2663 2418 2697
rect 2366 2654 2418 2663
rect 2430 2697 2482 2706
rect 2494 2697 2546 2706
rect 2558 2697 2610 2706
rect 2622 2697 2674 2706
rect 2686 2697 2738 2706
rect 2750 2697 2802 2706
rect 2430 2663 2455 2697
rect 2455 2663 2482 2697
rect 2494 2663 2527 2697
rect 2527 2663 2546 2697
rect 2558 2663 2561 2697
rect 2561 2663 2599 2697
rect 2599 2663 2610 2697
rect 2622 2663 2633 2697
rect 2633 2663 2671 2697
rect 2671 2663 2674 2697
rect 2686 2663 2705 2697
rect 2705 2663 2738 2697
rect 2750 2663 2777 2697
rect 2777 2663 2802 2697
rect 2430 2654 2482 2663
rect 2494 2654 2546 2663
rect 2558 2654 2610 2663
rect 2622 2654 2674 2663
rect 2686 2654 2738 2663
rect 2750 2654 2802 2663
rect 2814 2697 2866 2706
rect 2814 2663 2815 2697
rect 2815 2663 2849 2697
rect 2849 2663 2866 2697
rect 2814 2654 2866 2663
rect 2878 2697 2930 2706
rect 2878 2663 2887 2697
rect 2887 2663 2921 2697
rect 2921 2663 2930 2697
rect 2878 2654 2930 2663
rect 2942 2697 2994 2706
rect 2942 2663 2959 2697
rect 2959 2663 2993 2697
rect 2993 2663 2994 2697
rect 2942 2654 2994 2663
rect 3006 2697 3058 2706
rect 3070 2697 3122 2706
rect 3134 2697 3186 2706
rect 3198 2697 3250 2706
rect 3262 2697 3314 2706
rect 3326 2697 3378 2706
rect 3006 2663 3031 2697
rect 3031 2663 3058 2697
rect 3070 2663 3103 2697
rect 3103 2663 3122 2697
rect 3134 2663 3137 2697
rect 3137 2663 3175 2697
rect 3175 2663 3186 2697
rect 3198 2663 3209 2697
rect 3209 2663 3247 2697
rect 3247 2663 3250 2697
rect 3262 2663 3281 2697
rect 3281 2663 3314 2697
rect 3326 2663 3353 2697
rect 3353 2663 3378 2697
rect 3006 2654 3058 2663
rect 3070 2654 3122 2663
rect 3134 2654 3186 2663
rect 3198 2654 3250 2663
rect 3262 2654 3314 2663
rect 3326 2654 3378 2663
rect 3390 2697 3442 2706
rect 3390 2663 3391 2697
rect 3391 2663 3425 2697
rect 3425 2663 3442 2697
rect 3390 2654 3442 2663
rect 3454 2697 3506 2706
rect 3454 2663 3463 2697
rect 3463 2663 3497 2697
rect 3497 2663 3506 2697
rect 3454 2654 3506 2663
rect 3518 2697 3570 2706
rect 3518 2663 3535 2697
rect 3535 2663 3569 2697
rect 3569 2663 3570 2697
rect 3518 2654 3570 2663
rect 3582 2697 3634 2706
rect 3646 2697 3698 2706
rect 3710 2697 3762 2706
rect 3774 2697 3826 2706
rect 3838 2697 3890 2706
rect 3902 2697 3954 2706
rect 3582 2663 3607 2697
rect 3607 2663 3634 2697
rect 3646 2663 3679 2697
rect 3679 2663 3698 2697
rect 3710 2663 3713 2697
rect 3713 2663 3751 2697
rect 3751 2663 3762 2697
rect 3774 2663 3785 2697
rect 3785 2663 3823 2697
rect 3823 2663 3826 2697
rect 3838 2663 3857 2697
rect 3857 2663 3890 2697
rect 3902 2663 3929 2697
rect 3929 2663 3954 2697
rect 3582 2654 3634 2663
rect 3646 2654 3698 2663
rect 3710 2654 3762 2663
rect 3774 2654 3826 2663
rect 3838 2654 3890 2663
rect 3902 2654 3954 2663
rect 3966 2697 4018 2706
rect 3966 2663 3967 2697
rect 3967 2663 4001 2697
rect 4001 2663 4018 2697
rect 3966 2654 4018 2663
rect 4174 2654 4226 2706
rect 62 2377 114 2386
rect 62 2343 79 2377
rect 79 2343 113 2377
rect 113 2343 114 2377
rect 62 2334 114 2343
rect 126 2377 178 2386
rect 190 2377 242 2386
rect 254 2377 306 2386
rect 318 2377 370 2386
rect 382 2377 434 2386
rect 446 2377 498 2386
rect 126 2343 151 2377
rect 151 2343 178 2377
rect 190 2343 223 2377
rect 223 2343 242 2377
rect 254 2343 257 2377
rect 257 2343 295 2377
rect 295 2343 306 2377
rect 318 2343 329 2377
rect 329 2343 367 2377
rect 367 2343 370 2377
rect 382 2343 401 2377
rect 401 2343 434 2377
rect 446 2343 473 2377
rect 473 2343 498 2377
rect 126 2334 178 2343
rect 190 2334 242 2343
rect 254 2334 306 2343
rect 318 2334 370 2343
rect 382 2334 434 2343
rect 446 2334 498 2343
rect 510 2377 562 2386
rect 510 2343 511 2377
rect 511 2343 545 2377
rect 545 2343 562 2377
rect 510 2334 562 2343
rect 574 2377 626 2386
rect 574 2343 583 2377
rect 583 2343 617 2377
rect 617 2343 626 2377
rect 574 2334 626 2343
rect 638 2377 690 2386
rect 638 2343 655 2377
rect 655 2343 689 2377
rect 689 2343 690 2377
rect 638 2334 690 2343
rect 702 2377 754 2386
rect 766 2377 818 2386
rect 830 2377 882 2386
rect 894 2377 946 2386
rect 958 2377 1010 2386
rect 1022 2377 1074 2386
rect 702 2343 727 2377
rect 727 2343 754 2377
rect 766 2343 799 2377
rect 799 2343 818 2377
rect 830 2343 833 2377
rect 833 2343 871 2377
rect 871 2343 882 2377
rect 894 2343 905 2377
rect 905 2343 943 2377
rect 943 2343 946 2377
rect 958 2343 977 2377
rect 977 2343 1010 2377
rect 1022 2343 1049 2377
rect 1049 2343 1074 2377
rect 702 2334 754 2343
rect 766 2334 818 2343
rect 830 2334 882 2343
rect 894 2334 946 2343
rect 958 2334 1010 2343
rect 1022 2334 1074 2343
rect 1086 2377 1138 2386
rect 1086 2343 1087 2377
rect 1087 2343 1121 2377
rect 1121 2343 1138 2377
rect 1086 2334 1138 2343
rect 1150 2377 1202 2386
rect 1150 2343 1159 2377
rect 1159 2343 1193 2377
rect 1193 2343 1202 2377
rect 1150 2334 1202 2343
rect 1214 2377 1266 2386
rect 1214 2343 1231 2377
rect 1231 2343 1265 2377
rect 1265 2343 1266 2377
rect 1214 2334 1266 2343
rect 1278 2377 1330 2386
rect 1342 2377 1394 2386
rect 1406 2377 1458 2386
rect 1470 2377 1522 2386
rect 1534 2377 1586 2386
rect 1598 2377 1650 2386
rect 1278 2343 1303 2377
rect 1303 2343 1330 2377
rect 1342 2343 1375 2377
rect 1375 2343 1394 2377
rect 1406 2343 1409 2377
rect 1409 2343 1447 2377
rect 1447 2343 1458 2377
rect 1470 2343 1481 2377
rect 1481 2343 1519 2377
rect 1519 2343 1522 2377
rect 1534 2343 1553 2377
rect 1553 2343 1586 2377
rect 1598 2343 1625 2377
rect 1625 2343 1650 2377
rect 1278 2334 1330 2343
rect 1342 2334 1394 2343
rect 1406 2334 1458 2343
rect 1470 2334 1522 2343
rect 1534 2334 1586 2343
rect 1598 2334 1650 2343
rect 1662 2377 1714 2386
rect 1662 2343 1663 2377
rect 1663 2343 1697 2377
rect 1697 2343 1714 2377
rect 1662 2334 1714 2343
rect 1726 2377 1778 2386
rect 1726 2343 1735 2377
rect 1735 2343 1769 2377
rect 1769 2343 1778 2377
rect 1726 2334 1778 2343
rect 1790 2377 1842 2386
rect 1790 2343 1807 2377
rect 1807 2343 1841 2377
rect 1841 2343 1842 2377
rect 1790 2334 1842 2343
rect 1854 2377 1906 2386
rect 1918 2377 1970 2386
rect 1982 2377 2034 2386
rect 2046 2377 2098 2386
rect 2110 2377 2162 2386
rect 2174 2377 2226 2386
rect 1854 2343 1879 2377
rect 1879 2343 1906 2377
rect 1918 2343 1951 2377
rect 1951 2343 1970 2377
rect 1982 2343 1985 2377
rect 1985 2343 2023 2377
rect 2023 2343 2034 2377
rect 2046 2343 2057 2377
rect 2057 2343 2095 2377
rect 2095 2343 2098 2377
rect 2110 2343 2129 2377
rect 2129 2343 2162 2377
rect 2174 2343 2201 2377
rect 2201 2343 2226 2377
rect 1854 2334 1906 2343
rect 1918 2334 1970 2343
rect 1982 2334 2034 2343
rect 2046 2334 2098 2343
rect 2110 2334 2162 2343
rect 2174 2334 2226 2343
rect 2238 2377 2290 2386
rect 2238 2343 2239 2377
rect 2239 2343 2273 2377
rect 2273 2343 2290 2377
rect 2238 2334 2290 2343
rect 2302 2377 2354 2386
rect 2302 2343 2311 2377
rect 2311 2343 2345 2377
rect 2345 2343 2354 2377
rect 2302 2334 2354 2343
rect 2366 2377 2418 2386
rect 2366 2343 2383 2377
rect 2383 2343 2417 2377
rect 2417 2343 2418 2377
rect 2366 2334 2418 2343
rect 2430 2377 2482 2386
rect 2494 2377 2546 2386
rect 2558 2377 2610 2386
rect 2622 2377 2674 2386
rect 2686 2377 2738 2386
rect 2750 2377 2802 2386
rect 2430 2343 2455 2377
rect 2455 2343 2482 2377
rect 2494 2343 2527 2377
rect 2527 2343 2546 2377
rect 2558 2343 2561 2377
rect 2561 2343 2599 2377
rect 2599 2343 2610 2377
rect 2622 2343 2633 2377
rect 2633 2343 2671 2377
rect 2671 2343 2674 2377
rect 2686 2343 2705 2377
rect 2705 2343 2738 2377
rect 2750 2343 2777 2377
rect 2777 2343 2802 2377
rect 2430 2334 2482 2343
rect 2494 2334 2546 2343
rect 2558 2334 2610 2343
rect 2622 2334 2674 2343
rect 2686 2334 2738 2343
rect 2750 2334 2802 2343
rect 2814 2377 2866 2386
rect 2814 2343 2815 2377
rect 2815 2343 2849 2377
rect 2849 2343 2866 2377
rect 2814 2334 2866 2343
rect 2878 2377 2930 2386
rect 2878 2343 2887 2377
rect 2887 2343 2921 2377
rect 2921 2343 2930 2377
rect 2878 2334 2930 2343
rect 2942 2377 2994 2386
rect 2942 2343 2959 2377
rect 2959 2343 2993 2377
rect 2993 2343 2994 2377
rect 2942 2334 2994 2343
rect 3006 2377 3058 2386
rect 3070 2377 3122 2386
rect 3134 2377 3186 2386
rect 3198 2377 3250 2386
rect 3262 2377 3314 2386
rect 3326 2377 3378 2386
rect 3006 2343 3031 2377
rect 3031 2343 3058 2377
rect 3070 2343 3103 2377
rect 3103 2343 3122 2377
rect 3134 2343 3137 2377
rect 3137 2343 3175 2377
rect 3175 2343 3186 2377
rect 3198 2343 3209 2377
rect 3209 2343 3247 2377
rect 3247 2343 3250 2377
rect 3262 2343 3281 2377
rect 3281 2343 3314 2377
rect 3326 2343 3353 2377
rect 3353 2343 3378 2377
rect 3006 2334 3058 2343
rect 3070 2334 3122 2343
rect 3134 2334 3186 2343
rect 3198 2334 3250 2343
rect 3262 2334 3314 2343
rect 3326 2334 3378 2343
rect 3390 2377 3442 2386
rect 3390 2343 3391 2377
rect 3391 2343 3425 2377
rect 3425 2343 3442 2377
rect 3390 2334 3442 2343
rect 3454 2377 3506 2386
rect 3454 2343 3463 2377
rect 3463 2343 3497 2377
rect 3497 2343 3506 2377
rect 3454 2334 3506 2343
rect 3518 2377 3570 2386
rect 3518 2343 3535 2377
rect 3535 2343 3569 2377
rect 3569 2343 3570 2377
rect 3518 2334 3570 2343
rect 3582 2377 3634 2386
rect 3646 2377 3698 2386
rect 3710 2377 3762 2386
rect 3774 2377 3826 2386
rect 3838 2377 3890 2386
rect 3902 2377 3954 2386
rect 3582 2343 3607 2377
rect 3607 2343 3634 2377
rect 3646 2343 3679 2377
rect 3679 2343 3698 2377
rect 3710 2343 3713 2377
rect 3713 2343 3751 2377
rect 3751 2343 3762 2377
rect 3774 2343 3785 2377
rect 3785 2343 3823 2377
rect 3823 2343 3826 2377
rect 3838 2343 3857 2377
rect 3857 2343 3890 2377
rect 3902 2343 3929 2377
rect 3929 2343 3954 2377
rect 3582 2334 3634 2343
rect 3646 2334 3698 2343
rect 3710 2334 3762 2343
rect 3774 2334 3826 2343
rect 3838 2334 3890 2343
rect 3902 2334 3954 2343
rect 3966 2377 4018 2386
rect 3966 2343 3967 2377
rect 3967 2343 4001 2377
rect 4001 2343 4018 2377
rect 3966 2334 4018 2343
rect 8542 3817 8594 3826
rect 8542 3783 8559 3817
rect 8559 3783 8593 3817
rect 8593 3783 8594 3817
rect 8542 3774 8594 3783
rect 8606 3817 8658 3826
rect 8670 3817 8722 3826
rect 8734 3817 8786 3826
rect 8798 3817 8850 3826
rect 8862 3817 8914 3826
rect 8926 3817 8978 3826
rect 8606 3783 8631 3817
rect 8631 3783 8658 3817
rect 8670 3783 8703 3817
rect 8703 3783 8722 3817
rect 8734 3783 8737 3817
rect 8737 3783 8775 3817
rect 8775 3783 8786 3817
rect 8798 3783 8809 3817
rect 8809 3783 8847 3817
rect 8847 3783 8850 3817
rect 8862 3783 8881 3817
rect 8881 3783 8914 3817
rect 8926 3783 8953 3817
rect 8953 3783 8978 3817
rect 8606 3774 8658 3783
rect 8670 3774 8722 3783
rect 8734 3774 8786 3783
rect 8798 3774 8850 3783
rect 8862 3774 8914 3783
rect 8926 3774 8978 3783
rect 8990 3817 9042 3826
rect 8990 3783 8991 3817
rect 8991 3783 9025 3817
rect 9025 3783 9042 3817
rect 8990 3774 9042 3783
rect 9054 3817 9106 3826
rect 9054 3783 9063 3817
rect 9063 3783 9097 3817
rect 9097 3783 9106 3817
rect 9054 3774 9106 3783
rect 9118 3817 9170 3826
rect 9118 3783 9135 3817
rect 9135 3783 9169 3817
rect 9169 3783 9170 3817
rect 9118 3774 9170 3783
rect 9182 3817 9234 3826
rect 9246 3817 9298 3826
rect 9310 3817 9362 3826
rect 9374 3817 9426 3826
rect 9438 3817 9490 3826
rect 9502 3817 9554 3826
rect 9182 3783 9207 3817
rect 9207 3783 9234 3817
rect 9246 3783 9279 3817
rect 9279 3783 9298 3817
rect 9310 3783 9313 3817
rect 9313 3783 9351 3817
rect 9351 3783 9362 3817
rect 9374 3783 9385 3817
rect 9385 3783 9423 3817
rect 9423 3783 9426 3817
rect 9438 3783 9457 3817
rect 9457 3783 9490 3817
rect 9502 3783 9529 3817
rect 9529 3783 9554 3817
rect 9182 3774 9234 3783
rect 9246 3774 9298 3783
rect 9310 3774 9362 3783
rect 9374 3774 9426 3783
rect 9438 3774 9490 3783
rect 9502 3774 9554 3783
rect 9566 3817 9618 3826
rect 9566 3783 9567 3817
rect 9567 3783 9601 3817
rect 9601 3783 9618 3817
rect 9566 3774 9618 3783
rect 9630 3817 9682 3826
rect 9630 3783 9639 3817
rect 9639 3783 9673 3817
rect 9673 3783 9682 3817
rect 9630 3774 9682 3783
rect 9694 3817 9746 3826
rect 9694 3783 9711 3817
rect 9711 3783 9745 3817
rect 9745 3783 9746 3817
rect 9694 3774 9746 3783
rect 9758 3817 9810 3826
rect 9822 3817 9874 3826
rect 9886 3817 9938 3826
rect 9950 3817 10002 3826
rect 10014 3817 10066 3826
rect 10078 3817 10130 3826
rect 9758 3783 9783 3817
rect 9783 3783 9810 3817
rect 9822 3783 9855 3817
rect 9855 3783 9874 3817
rect 9886 3783 9889 3817
rect 9889 3783 9927 3817
rect 9927 3783 9938 3817
rect 9950 3783 9961 3817
rect 9961 3783 9999 3817
rect 9999 3783 10002 3817
rect 10014 3783 10033 3817
rect 10033 3783 10066 3817
rect 10078 3783 10105 3817
rect 10105 3783 10130 3817
rect 9758 3774 9810 3783
rect 9822 3774 9874 3783
rect 9886 3774 9938 3783
rect 9950 3774 10002 3783
rect 10014 3774 10066 3783
rect 10078 3774 10130 3783
rect 10142 3817 10194 3826
rect 10142 3783 10143 3817
rect 10143 3783 10177 3817
rect 10177 3783 10194 3817
rect 10142 3774 10194 3783
rect 10206 3817 10258 3826
rect 10206 3783 10215 3817
rect 10215 3783 10249 3817
rect 10249 3783 10258 3817
rect 10206 3774 10258 3783
rect 10270 3817 10322 3826
rect 10270 3783 10287 3817
rect 10287 3783 10321 3817
rect 10321 3783 10322 3817
rect 10270 3774 10322 3783
rect 10334 3817 10386 3826
rect 10398 3817 10450 3826
rect 10462 3817 10514 3826
rect 10526 3817 10578 3826
rect 10590 3817 10642 3826
rect 10654 3817 10706 3826
rect 10334 3783 10359 3817
rect 10359 3783 10386 3817
rect 10398 3783 10431 3817
rect 10431 3783 10450 3817
rect 10462 3783 10465 3817
rect 10465 3783 10503 3817
rect 10503 3783 10514 3817
rect 10526 3783 10537 3817
rect 10537 3783 10575 3817
rect 10575 3783 10578 3817
rect 10590 3783 10609 3817
rect 10609 3783 10642 3817
rect 10654 3783 10681 3817
rect 10681 3783 10706 3817
rect 10334 3774 10386 3783
rect 10398 3774 10450 3783
rect 10462 3774 10514 3783
rect 10526 3774 10578 3783
rect 10590 3774 10642 3783
rect 10654 3774 10706 3783
rect 10718 3817 10770 3826
rect 10718 3783 10719 3817
rect 10719 3783 10753 3817
rect 10753 3783 10770 3817
rect 10718 3774 10770 3783
rect 10782 3817 10834 3826
rect 10782 3783 10791 3817
rect 10791 3783 10825 3817
rect 10825 3783 10834 3817
rect 10782 3774 10834 3783
rect 10846 3817 10898 3826
rect 10846 3783 10863 3817
rect 10863 3783 10897 3817
rect 10897 3783 10898 3817
rect 10846 3774 10898 3783
rect 10910 3817 10962 3826
rect 10974 3817 11026 3826
rect 11038 3817 11090 3826
rect 11102 3817 11154 3826
rect 11166 3817 11218 3826
rect 11230 3817 11282 3826
rect 10910 3783 10935 3817
rect 10935 3783 10962 3817
rect 10974 3783 11007 3817
rect 11007 3783 11026 3817
rect 11038 3783 11041 3817
rect 11041 3783 11079 3817
rect 11079 3783 11090 3817
rect 11102 3783 11113 3817
rect 11113 3783 11151 3817
rect 11151 3783 11154 3817
rect 11166 3783 11185 3817
rect 11185 3783 11218 3817
rect 11230 3783 11257 3817
rect 11257 3783 11282 3817
rect 10910 3774 10962 3783
rect 10974 3774 11026 3783
rect 11038 3774 11090 3783
rect 11102 3774 11154 3783
rect 11166 3774 11218 3783
rect 11230 3774 11282 3783
rect 11294 3817 11346 3826
rect 11294 3783 11295 3817
rect 11295 3783 11329 3817
rect 11329 3783 11346 3817
rect 11294 3774 11346 3783
rect 11358 3817 11410 3826
rect 11358 3783 11367 3817
rect 11367 3783 11401 3817
rect 11401 3783 11410 3817
rect 11358 3774 11410 3783
rect 11422 3817 11474 3826
rect 11422 3783 11439 3817
rect 11439 3783 11473 3817
rect 11473 3783 11474 3817
rect 11422 3774 11474 3783
rect 11486 3817 11538 3826
rect 11550 3817 11602 3826
rect 11614 3817 11666 3826
rect 11678 3817 11730 3826
rect 11742 3817 11794 3826
rect 11806 3817 11858 3826
rect 11486 3783 11511 3817
rect 11511 3783 11538 3817
rect 11550 3783 11583 3817
rect 11583 3783 11602 3817
rect 11614 3783 11617 3817
rect 11617 3783 11655 3817
rect 11655 3783 11666 3817
rect 11678 3783 11689 3817
rect 11689 3783 11727 3817
rect 11727 3783 11730 3817
rect 11742 3783 11761 3817
rect 11761 3783 11794 3817
rect 11806 3783 11833 3817
rect 11833 3783 11858 3817
rect 11486 3774 11538 3783
rect 11550 3774 11602 3783
rect 11614 3774 11666 3783
rect 11678 3774 11730 3783
rect 11742 3774 11794 3783
rect 11806 3774 11858 3783
rect 11870 3817 11922 3826
rect 11870 3783 11871 3817
rect 11871 3783 11905 3817
rect 11905 3783 11922 3817
rect 11870 3774 11922 3783
rect 11934 3817 11986 3826
rect 11934 3783 11943 3817
rect 11943 3783 11977 3817
rect 11977 3783 11986 3817
rect 11934 3774 11986 3783
rect 11998 3817 12050 3826
rect 11998 3783 12015 3817
rect 12015 3783 12049 3817
rect 12049 3783 12050 3817
rect 11998 3774 12050 3783
rect 12062 3817 12114 3826
rect 12126 3817 12178 3826
rect 12190 3817 12242 3826
rect 12254 3817 12306 3826
rect 12318 3817 12370 3826
rect 12382 3817 12434 3826
rect 12062 3783 12087 3817
rect 12087 3783 12114 3817
rect 12126 3783 12159 3817
rect 12159 3783 12178 3817
rect 12190 3783 12193 3817
rect 12193 3783 12231 3817
rect 12231 3783 12242 3817
rect 12254 3783 12265 3817
rect 12265 3783 12303 3817
rect 12303 3783 12306 3817
rect 12318 3783 12337 3817
rect 12337 3783 12370 3817
rect 12382 3783 12409 3817
rect 12409 3783 12434 3817
rect 12062 3774 12114 3783
rect 12126 3774 12178 3783
rect 12190 3774 12242 3783
rect 12254 3774 12306 3783
rect 12318 3774 12370 3783
rect 12382 3774 12434 3783
rect 12446 3817 12498 3826
rect 12446 3783 12447 3817
rect 12447 3783 12481 3817
rect 12481 3783 12498 3817
rect 12446 3774 12498 3783
rect 8542 3497 8594 3506
rect 8542 3463 8559 3497
rect 8559 3463 8593 3497
rect 8593 3463 8594 3497
rect 8542 3454 8594 3463
rect 8606 3497 8658 3506
rect 8670 3497 8722 3506
rect 8734 3497 8786 3506
rect 8798 3497 8850 3506
rect 8862 3497 8914 3506
rect 8926 3497 8978 3506
rect 8606 3463 8631 3497
rect 8631 3463 8658 3497
rect 8670 3463 8703 3497
rect 8703 3463 8722 3497
rect 8734 3463 8737 3497
rect 8737 3463 8775 3497
rect 8775 3463 8786 3497
rect 8798 3463 8809 3497
rect 8809 3463 8847 3497
rect 8847 3463 8850 3497
rect 8862 3463 8881 3497
rect 8881 3463 8914 3497
rect 8926 3463 8953 3497
rect 8953 3463 8978 3497
rect 8606 3454 8658 3463
rect 8670 3454 8722 3463
rect 8734 3454 8786 3463
rect 8798 3454 8850 3463
rect 8862 3454 8914 3463
rect 8926 3454 8978 3463
rect 8990 3497 9042 3506
rect 8990 3463 8991 3497
rect 8991 3463 9025 3497
rect 9025 3463 9042 3497
rect 8990 3454 9042 3463
rect 9054 3497 9106 3506
rect 9054 3463 9063 3497
rect 9063 3463 9097 3497
rect 9097 3463 9106 3497
rect 9054 3454 9106 3463
rect 9118 3497 9170 3506
rect 9118 3463 9135 3497
rect 9135 3463 9169 3497
rect 9169 3463 9170 3497
rect 9118 3454 9170 3463
rect 9182 3497 9234 3506
rect 9246 3497 9298 3506
rect 9310 3497 9362 3506
rect 9374 3497 9426 3506
rect 9438 3497 9490 3506
rect 9502 3497 9554 3506
rect 9182 3463 9207 3497
rect 9207 3463 9234 3497
rect 9246 3463 9279 3497
rect 9279 3463 9298 3497
rect 9310 3463 9313 3497
rect 9313 3463 9351 3497
rect 9351 3463 9362 3497
rect 9374 3463 9385 3497
rect 9385 3463 9423 3497
rect 9423 3463 9426 3497
rect 9438 3463 9457 3497
rect 9457 3463 9490 3497
rect 9502 3463 9529 3497
rect 9529 3463 9554 3497
rect 9182 3454 9234 3463
rect 9246 3454 9298 3463
rect 9310 3454 9362 3463
rect 9374 3454 9426 3463
rect 9438 3454 9490 3463
rect 9502 3454 9554 3463
rect 9566 3497 9618 3506
rect 9566 3463 9567 3497
rect 9567 3463 9601 3497
rect 9601 3463 9618 3497
rect 9566 3454 9618 3463
rect 9630 3497 9682 3506
rect 9630 3463 9639 3497
rect 9639 3463 9673 3497
rect 9673 3463 9682 3497
rect 9630 3454 9682 3463
rect 9694 3497 9746 3506
rect 9694 3463 9711 3497
rect 9711 3463 9745 3497
rect 9745 3463 9746 3497
rect 9694 3454 9746 3463
rect 9758 3497 9810 3506
rect 9822 3497 9874 3506
rect 9886 3497 9938 3506
rect 9950 3497 10002 3506
rect 10014 3497 10066 3506
rect 10078 3497 10130 3506
rect 9758 3463 9783 3497
rect 9783 3463 9810 3497
rect 9822 3463 9855 3497
rect 9855 3463 9874 3497
rect 9886 3463 9889 3497
rect 9889 3463 9927 3497
rect 9927 3463 9938 3497
rect 9950 3463 9961 3497
rect 9961 3463 9999 3497
rect 9999 3463 10002 3497
rect 10014 3463 10033 3497
rect 10033 3463 10066 3497
rect 10078 3463 10105 3497
rect 10105 3463 10130 3497
rect 9758 3454 9810 3463
rect 9822 3454 9874 3463
rect 9886 3454 9938 3463
rect 9950 3454 10002 3463
rect 10014 3454 10066 3463
rect 10078 3454 10130 3463
rect 10142 3497 10194 3506
rect 10142 3463 10143 3497
rect 10143 3463 10177 3497
rect 10177 3463 10194 3497
rect 10142 3454 10194 3463
rect 10206 3497 10258 3506
rect 10206 3463 10215 3497
rect 10215 3463 10249 3497
rect 10249 3463 10258 3497
rect 10206 3454 10258 3463
rect 10270 3497 10322 3506
rect 10270 3463 10287 3497
rect 10287 3463 10321 3497
rect 10321 3463 10322 3497
rect 10270 3454 10322 3463
rect 10334 3497 10386 3506
rect 10398 3497 10450 3506
rect 10462 3497 10514 3506
rect 10526 3497 10578 3506
rect 10590 3497 10642 3506
rect 10654 3497 10706 3506
rect 10334 3463 10359 3497
rect 10359 3463 10386 3497
rect 10398 3463 10431 3497
rect 10431 3463 10450 3497
rect 10462 3463 10465 3497
rect 10465 3463 10503 3497
rect 10503 3463 10514 3497
rect 10526 3463 10537 3497
rect 10537 3463 10575 3497
rect 10575 3463 10578 3497
rect 10590 3463 10609 3497
rect 10609 3463 10642 3497
rect 10654 3463 10681 3497
rect 10681 3463 10706 3497
rect 10334 3454 10386 3463
rect 10398 3454 10450 3463
rect 10462 3454 10514 3463
rect 10526 3454 10578 3463
rect 10590 3454 10642 3463
rect 10654 3454 10706 3463
rect 10718 3497 10770 3506
rect 10718 3463 10719 3497
rect 10719 3463 10753 3497
rect 10753 3463 10770 3497
rect 10718 3454 10770 3463
rect 10782 3497 10834 3506
rect 10782 3463 10791 3497
rect 10791 3463 10825 3497
rect 10825 3463 10834 3497
rect 10782 3454 10834 3463
rect 10846 3497 10898 3506
rect 10846 3463 10863 3497
rect 10863 3463 10897 3497
rect 10897 3463 10898 3497
rect 10846 3454 10898 3463
rect 10910 3497 10962 3506
rect 10974 3497 11026 3506
rect 11038 3497 11090 3506
rect 11102 3497 11154 3506
rect 11166 3497 11218 3506
rect 11230 3497 11282 3506
rect 10910 3463 10935 3497
rect 10935 3463 10962 3497
rect 10974 3463 11007 3497
rect 11007 3463 11026 3497
rect 11038 3463 11041 3497
rect 11041 3463 11079 3497
rect 11079 3463 11090 3497
rect 11102 3463 11113 3497
rect 11113 3463 11151 3497
rect 11151 3463 11154 3497
rect 11166 3463 11185 3497
rect 11185 3463 11218 3497
rect 11230 3463 11257 3497
rect 11257 3463 11282 3497
rect 10910 3454 10962 3463
rect 10974 3454 11026 3463
rect 11038 3454 11090 3463
rect 11102 3454 11154 3463
rect 11166 3454 11218 3463
rect 11230 3454 11282 3463
rect 11294 3497 11346 3506
rect 11294 3463 11295 3497
rect 11295 3463 11329 3497
rect 11329 3463 11346 3497
rect 11294 3454 11346 3463
rect 11358 3497 11410 3506
rect 11358 3463 11367 3497
rect 11367 3463 11401 3497
rect 11401 3463 11410 3497
rect 11358 3454 11410 3463
rect 11422 3497 11474 3506
rect 11422 3463 11439 3497
rect 11439 3463 11473 3497
rect 11473 3463 11474 3497
rect 11422 3454 11474 3463
rect 11486 3497 11538 3506
rect 11550 3497 11602 3506
rect 11614 3497 11666 3506
rect 11678 3497 11730 3506
rect 11742 3497 11794 3506
rect 11806 3497 11858 3506
rect 11486 3463 11511 3497
rect 11511 3463 11538 3497
rect 11550 3463 11583 3497
rect 11583 3463 11602 3497
rect 11614 3463 11617 3497
rect 11617 3463 11655 3497
rect 11655 3463 11666 3497
rect 11678 3463 11689 3497
rect 11689 3463 11727 3497
rect 11727 3463 11730 3497
rect 11742 3463 11761 3497
rect 11761 3463 11794 3497
rect 11806 3463 11833 3497
rect 11833 3463 11858 3497
rect 11486 3454 11538 3463
rect 11550 3454 11602 3463
rect 11614 3454 11666 3463
rect 11678 3454 11730 3463
rect 11742 3454 11794 3463
rect 11806 3454 11858 3463
rect 11870 3497 11922 3506
rect 11870 3463 11871 3497
rect 11871 3463 11905 3497
rect 11905 3463 11922 3497
rect 11870 3454 11922 3463
rect 11934 3497 11986 3506
rect 11934 3463 11943 3497
rect 11943 3463 11977 3497
rect 11977 3463 11986 3497
rect 11934 3454 11986 3463
rect 11998 3497 12050 3506
rect 11998 3463 12015 3497
rect 12015 3463 12049 3497
rect 12049 3463 12050 3497
rect 11998 3454 12050 3463
rect 12062 3497 12114 3506
rect 12126 3497 12178 3506
rect 12190 3497 12242 3506
rect 12254 3497 12306 3506
rect 12318 3497 12370 3506
rect 12382 3497 12434 3506
rect 12062 3463 12087 3497
rect 12087 3463 12114 3497
rect 12126 3463 12159 3497
rect 12159 3463 12178 3497
rect 12190 3463 12193 3497
rect 12193 3463 12231 3497
rect 12231 3463 12242 3497
rect 12254 3463 12265 3497
rect 12265 3463 12303 3497
rect 12303 3463 12306 3497
rect 12318 3463 12337 3497
rect 12337 3463 12370 3497
rect 12382 3463 12409 3497
rect 12409 3463 12434 3497
rect 12062 3454 12114 3463
rect 12126 3454 12178 3463
rect 12190 3454 12242 3463
rect 12254 3454 12306 3463
rect 12318 3454 12370 3463
rect 12382 3454 12434 3463
rect 12446 3497 12498 3506
rect 12446 3463 12447 3497
rect 12447 3463 12481 3497
rect 12481 3463 12498 3497
rect 12446 3454 12498 3463
rect 12654 3454 12706 3506
rect 8334 2654 8386 2706
rect 8542 2697 8594 2706
rect 8542 2663 8559 2697
rect 8559 2663 8593 2697
rect 8593 2663 8594 2697
rect 8542 2654 8594 2663
rect 8606 2697 8658 2706
rect 8670 2697 8722 2706
rect 8734 2697 8786 2706
rect 8798 2697 8850 2706
rect 8862 2697 8914 2706
rect 8926 2697 8978 2706
rect 8606 2663 8631 2697
rect 8631 2663 8658 2697
rect 8670 2663 8703 2697
rect 8703 2663 8722 2697
rect 8734 2663 8737 2697
rect 8737 2663 8775 2697
rect 8775 2663 8786 2697
rect 8798 2663 8809 2697
rect 8809 2663 8847 2697
rect 8847 2663 8850 2697
rect 8862 2663 8881 2697
rect 8881 2663 8914 2697
rect 8926 2663 8953 2697
rect 8953 2663 8978 2697
rect 8606 2654 8658 2663
rect 8670 2654 8722 2663
rect 8734 2654 8786 2663
rect 8798 2654 8850 2663
rect 8862 2654 8914 2663
rect 8926 2654 8978 2663
rect 8990 2697 9042 2706
rect 8990 2663 8991 2697
rect 8991 2663 9025 2697
rect 9025 2663 9042 2697
rect 8990 2654 9042 2663
rect 9054 2697 9106 2706
rect 9054 2663 9063 2697
rect 9063 2663 9097 2697
rect 9097 2663 9106 2697
rect 9054 2654 9106 2663
rect 9118 2697 9170 2706
rect 9118 2663 9135 2697
rect 9135 2663 9169 2697
rect 9169 2663 9170 2697
rect 9118 2654 9170 2663
rect 9182 2697 9234 2706
rect 9246 2697 9298 2706
rect 9310 2697 9362 2706
rect 9374 2697 9426 2706
rect 9438 2697 9490 2706
rect 9502 2697 9554 2706
rect 9182 2663 9207 2697
rect 9207 2663 9234 2697
rect 9246 2663 9279 2697
rect 9279 2663 9298 2697
rect 9310 2663 9313 2697
rect 9313 2663 9351 2697
rect 9351 2663 9362 2697
rect 9374 2663 9385 2697
rect 9385 2663 9423 2697
rect 9423 2663 9426 2697
rect 9438 2663 9457 2697
rect 9457 2663 9490 2697
rect 9502 2663 9529 2697
rect 9529 2663 9554 2697
rect 9182 2654 9234 2663
rect 9246 2654 9298 2663
rect 9310 2654 9362 2663
rect 9374 2654 9426 2663
rect 9438 2654 9490 2663
rect 9502 2654 9554 2663
rect 9566 2697 9618 2706
rect 9566 2663 9567 2697
rect 9567 2663 9601 2697
rect 9601 2663 9618 2697
rect 9566 2654 9618 2663
rect 9630 2697 9682 2706
rect 9630 2663 9639 2697
rect 9639 2663 9673 2697
rect 9673 2663 9682 2697
rect 9630 2654 9682 2663
rect 9694 2697 9746 2706
rect 9694 2663 9711 2697
rect 9711 2663 9745 2697
rect 9745 2663 9746 2697
rect 9694 2654 9746 2663
rect 9758 2697 9810 2706
rect 9822 2697 9874 2706
rect 9886 2697 9938 2706
rect 9950 2697 10002 2706
rect 10014 2697 10066 2706
rect 10078 2697 10130 2706
rect 9758 2663 9783 2697
rect 9783 2663 9810 2697
rect 9822 2663 9855 2697
rect 9855 2663 9874 2697
rect 9886 2663 9889 2697
rect 9889 2663 9927 2697
rect 9927 2663 9938 2697
rect 9950 2663 9961 2697
rect 9961 2663 9999 2697
rect 9999 2663 10002 2697
rect 10014 2663 10033 2697
rect 10033 2663 10066 2697
rect 10078 2663 10105 2697
rect 10105 2663 10130 2697
rect 9758 2654 9810 2663
rect 9822 2654 9874 2663
rect 9886 2654 9938 2663
rect 9950 2654 10002 2663
rect 10014 2654 10066 2663
rect 10078 2654 10130 2663
rect 10142 2697 10194 2706
rect 10142 2663 10143 2697
rect 10143 2663 10177 2697
rect 10177 2663 10194 2697
rect 10142 2654 10194 2663
rect 10206 2697 10258 2706
rect 10206 2663 10215 2697
rect 10215 2663 10249 2697
rect 10249 2663 10258 2697
rect 10206 2654 10258 2663
rect 10270 2697 10322 2706
rect 10270 2663 10287 2697
rect 10287 2663 10321 2697
rect 10321 2663 10322 2697
rect 10270 2654 10322 2663
rect 10334 2697 10386 2706
rect 10398 2697 10450 2706
rect 10462 2697 10514 2706
rect 10526 2697 10578 2706
rect 10590 2697 10642 2706
rect 10654 2697 10706 2706
rect 10334 2663 10359 2697
rect 10359 2663 10386 2697
rect 10398 2663 10431 2697
rect 10431 2663 10450 2697
rect 10462 2663 10465 2697
rect 10465 2663 10503 2697
rect 10503 2663 10514 2697
rect 10526 2663 10537 2697
rect 10537 2663 10575 2697
rect 10575 2663 10578 2697
rect 10590 2663 10609 2697
rect 10609 2663 10642 2697
rect 10654 2663 10681 2697
rect 10681 2663 10706 2697
rect 10334 2654 10386 2663
rect 10398 2654 10450 2663
rect 10462 2654 10514 2663
rect 10526 2654 10578 2663
rect 10590 2654 10642 2663
rect 10654 2654 10706 2663
rect 10718 2697 10770 2706
rect 10718 2663 10719 2697
rect 10719 2663 10753 2697
rect 10753 2663 10770 2697
rect 10718 2654 10770 2663
rect 10782 2697 10834 2706
rect 10782 2663 10791 2697
rect 10791 2663 10825 2697
rect 10825 2663 10834 2697
rect 10782 2654 10834 2663
rect 10846 2697 10898 2706
rect 10846 2663 10863 2697
rect 10863 2663 10897 2697
rect 10897 2663 10898 2697
rect 10846 2654 10898 2663
rect 10910 2697 10962 2706
rect 10974 2697 11026 2706
rect 11038 2697 11090 2706
rect 11102 2697 11154 2706
rect 11166 2697 11218 2706
rect 11230 2697 11282 2706
rect 10910 2663 10935 2697
rect 10935 2663 10962 2697
rect 10974 2663 11007 2697
rect 11007 2663 11026 2697
rect 11038 2663 11041 2697
rect 11041 2663 11079 2697
rect 11079 2663 11090 2697
rect 11102 2663 11113 2697
rect 11113 2663 11151 2697
rect 11151 2663 11154 2697
rect 11166 2663 11185 2697
rect 11185 2663 11218 2697
rect 11230 2663 11257 2697
rect 11257 2663 11282 2697
rect 10910 2654 10962 2663
rect 10974 2654 11026 2663
rect 11038 2654 11090 2663
rect 11102 2654 11154 2663
rect 11166 2654 11218 2663
rect 11230 2654 11282 2663
rect 11294 2697 11346 2706
rect 11294 2663 11295 2697
rect 11295 2663 11329 2697
rect 11329 2663 11346 2697
rect 11294 2654 11346 2663
rect 11358 2697 11410 2706
rect 11358 2663 11367 2697
rect 11367 2663 11401 2697
rect 11401 2663 11410 2697
rect 11358 2654 11410 2663
rect 11422 2697 11474 2706
rect 11422 2663 11439 2697
rect 11439 2663 11473 2697
rect 11473 2663 11474 2697
rect 11422 2654 11474 2663
rect 11486 2697 11538 2706
rect 11550 2697 11602 2706
rect 11614 2697 11666 2706
rect 11678 2697 11730 2706
rect 11742 2697 11794 2706
rect 11806 2697 11858 2706
rect 11486 2663 11511 2697
rect 11511 2663 11538 2697
rect 11550 2663 11583 2697
rect 11583 2663 11602 2697
rect 11614 2663 11617 2697
rect 11617 2663 11655 2697
rect 11655 2663 11666 2697
rect 11678 2663 11689 2697
rect 11689 2663 11727 2697
rect 11727 2663 11730 2697
rect 11742 2663 11761 2697
rect 11761 2663 11794 2697
rect 11806 2663 11833 2697
rect 11833 2663 11858 2697
rect 11486 2654 11538 2663
rect 11550 2654 11602 2663
rect 11614 2654 11666 2663
rect 11678 2654 11730 2663
rect 11742 2654 11794 2663
rect 11806 2654 11858 2663
rect 11870 2697 11922 2706
rect 11870 2663 11871 2697
rect 11871 2663 11905 2697
rect 11905 2663 11922 2697
rect 11870 2654 11922 2663
rect 11934 2697 11986 2706
rect 11934 2663 11943 2697
rect 11943 2663 11977 2697
rect 11977 2663 11986 2697
rect 11934 2654 11986 2663
rect 11998 2697 12050 2706
rect 11998 2663 12015 2697
rect 12015 2663 12049 2697
rect 12049 2663 12050 2697
rect 11998 2654 12050 2663
rect 12062 2697 12114 2706
rect 12126 2697 12178 2706
rect 12190 2697 12242 2706
rect 12254 2697 12306 2706
rect 12318 2697 12370 2706
rect 12382 2697 12434 2706
rect 12062 2663 12087 2697
rect 12087 2663 12114 2697
rect 12126 2663 12159 2697
rect 12159 2663 12178 2697
rect 12190 2663 12193 2697
rect 12193 2663 12231 2697
rect 12231 2663 12242 2697
rect 12254 2663 12265 2697
rect 12265 2663 12303 2697
rect 12303 2663 12306 2697
rect 12318 2663 12337 2697
rect 12337 2663 12370 2697
rect 12382 2663 12409 2697
rect 12409 2663 12434 2697
rect 12062 2654 12114 2663
rect 12126 2654 12178 2663
rect 12190 2654 12242 2663
rect 12254 2654 12306 2663
rect 12318 2654 12370 2663
rect 12382 2654 12434 2663
rect 12446 2697 12498 2706
rect 12446 2663 12447 2697
rect 12447 2663 12481 2697
rect 12481 2663 12498 2697
rect 12446 2654 12498 2663
rect 8542 2377 8594 2386
rect 8542 2343 8559 2377
rect 8559 2343 8593 2377
rect 8593 2343 8594 2377
rect 8542 2334 8594 2343
rect 8606 2377 8658 2386
rect 8670 2377 8722 2386
rect 8734 2377 8786 2386
rect 8798 2377 8850 2386
rect 8862 2377 8914 2386
rect 8926 2377 8978 2386
rect 8606 2343 8631 2377
rect 8631 2343 8658 2377
rect 8670 2343 8703 2377
rect 8703 2343 8722 2377
rect 8734 2343 8737 2377
rect 8737 2343 8775 2377
rect 8775 2343 8786 2377
rect 8798 2343 8809 2377
rect 8809 2343 8847 2377
rect 8847 2343 8850 2377
rect 8862 2343 8881 2377
rect 8881 2343 8914 2377
rect 8926 2343 8953 2377
rect 8953 2343 8978 2377
rect 8606 2334 8658 2343
rect 8670 2334 8722 2343
rect 8734 2334 8786 2343
rect 8798 2334 8850 2343
rect 8862 2334 8914 2343
rect 8926 2334 8978 2343
rect 8990 2377 9042 2386
rect 8990 2343 8991 2377
rect 8991 2343 9025 2377
rect 9025 2343 9042 2377
rect 8990 2334 9042 2343
rect 9054 2377 9106 2386
rect 9054 2343 9063 2377
rect 9063 2343 9097 2377
rect 9097 2343 9106 2377
rect 9054 2334 9106 2343
rect 9118 2377 9170 2386
rect 9118 2343 9135 2377
rect 9135 2343 9169 2377
rect 9169 2343 9170 2377
rect 9118 2334 9170 2343
rect 9182 2377 9234 2386
rect 9246 2377 9298 2386
rect 9310 2377 9362 2386
rect 9374 2377 9426 2386
rect 9438 2377 9490 2386
rect 9502 2377 9554 2386
rect 9182 2343 9207 2377
rect 9207 2343 9234 2377
rect 9246 2343 9279 2377
rect 9279 2343 9298 2377
rect 9310 2343 9313 2377
rect 9313 2343 9351 2377
rect 9351 2343 9362 2377
rect 9374 2343 9385 2377
rect 9385 2343 9423 2377
rect 9423 2343 9426 2377
rect 9438 2343 9457 2377
rect 9457 2343 9490 2377
rect 9502 2343 9529 2377
rect 9529 2343 9554 2377
rect 9182 2334 9234 2343
rect 9246 2334 9298 2343
rect 9310 2334 9362 2343
rect 9374 2334 9426 2343
rect 9438 2334 9490 2343
rect 9502 2334 9554 2343
rect 9566 2377 9618 2386
rect 9566 2343 9567 2377
rect 9567 2343 9601 2377
rect 9601 2343 9618 2377
rect 9566 2334 9618 2343
rect 9630 2377 9682 2386
rect 9630 2343 9639 2377
rect 9639 2343 9673 2377
rect 9673 2343 9682 2377
rect 9630 2334 9682 2343
rect 9694 2377 9746 2386
rect 9694 2343 9711 2377
rect 9711 2343 9745 2377
rect 9745 2343 9746 2377
rect 9694 2334 9746 2343
rect 9758 2377 9810 2386
rect 9822 2377 9874 2386
rect 9886 2377 9938 2386
rect 9950 2377 10002 2386
rect 10014 2377 10066 2386
rect 10078 2377 10130 2386
rect 9758 2343 9783 2377
rect 9783 2343 9810 2377
rect 9822 2343 9855 2377
rect 9855 2343 9874 2377
rect 9886 2343 9889 2377
rect 9889 2343 9927 2377
rect 9927 2343 9938 2377
rect 9950 2343 9961 2377
rect 9961 2343 9999 2377
rect 9999 2343 10002 2377
rect 10014 2343 10033 2377
rect 10033 2343 10066 2377
rect 10078 2343 10105 2377
rect 10105 2343 10130 2377
rect 9758 2334 9810 2343
rect 9822 2334 9874 2343
rect 9886 2334 9938 2343
rect 9950 2334 10002 2343
rect 10014 2334 10066 2343
rect 10078 2334 10130 2343
rect 10142 2377 10194 2386
rect 10142 2343 10143 2377
rect 10143 2343 10177 2377
rect 10177 2343 10194 2377
rect 10142 2334 10194 2343
rect 10206 2377 10258 2386
rect 10206 2343 10215 2377
rect 10215 2343 10249 2377
rect 10249 2343 10258 2377
rect 10206 2334 10258 2343
rect 10270 2377 10322 2386
rect 10270 2343 10287 2377
rect 10287 2343 10321 2377
rect 10321 2343 10322 2377
rect 10270 2334 10322 2343
rect 10334 2377 10386 2386
rect 10398 2377 10450 2386
rect 10462 2377 10514 2386
rect 10526 2377 10578 2386
rect 10590 2377 10642 2386
rect 10654 2377 10706 2386
rect 10334 2343 10359 2377
rect 10359 2343 10386 2377
rect 10398 2343 10431 2377
rect 10431 2343 10450 2377
rect 10462 2343 10465 2377
rect 10465 2343 10503 2377
rect 10503 2343 10514 2377
rect 10526 2343 10537 2377
rect 10537 2343 10575 2377
rect 10575 2343 10578 2377
rect 10590 2343 10609 2377
rect 10609 2343 10642 2377
rect 10654 2343 10681 2377
rect 10681 2343 10706 2377
rect 10334 2334 10386 2343
rect 10398 2334 10450 2343
rect 10462 2334 10514 2343
rect 10526 2334 10578 2343
rect 10590 2334 10642 2343
rect 10654 2334 10706 2343
rect 10718 2377 10770 2386
rect 10718 2343 10719 2377
rect 10719 2343 10753 2377
rect 10753 2343 10770 2377
rect 10718 2334 10770 2343
rect 10782 2377 10834 2386
rect 10782 2343 10791 2377
rect 10791 2343 10825 2377
rect 10825 2343 10834 2377
rect 10782 2334 10834 2343
rect 10846 2377 10898 2386
rect 10846 2343 10863 2377
rect 10863 2343 10897 2377
rect 10897 2343 10898 2377
rect 10846 2334 10898 2343
rect 10910 2377 10962 2386
rect 10974 2377 11026 2386
rect 11038 2377 11090 2386
rect 11102 2377 11154 2386
rect 11166 2377 11218 2386
rect 11230 2377 11282 2386
rect 10910 2343 10935 2377
rect 10935 2343 10962 2377
rect 10974 2343 11007 2377
rect 11007 2343 11026 2377
rect 11038 2343 11041 2377
rect 11041 2343 11079 2377
rect 11079 2343 11090 2377
rect 11102 2343 11113 2377
rect 11113 2343 11151 2377
rect 11151 2343 11154 2377
rect 11166 2343 11185 2377
rect 11185 2343 11218 2377
rect 11230 2343 11257 2377
rect 11257 2343 11282 2377
rect 10910 2334 10962 2343
rect 10974 2334 11026 2343
rect 11038 2334 11090 2343
rect 11102 2334 11154 2343
rect 11166 2334 11218 2343
rect 11230 2334 11282 2343
rect 11294 2377 11346 2386
rect 11294 2343 11295 2377
rect 11295 2343 11329 2377
rect 11329 2343 11346 2377
rect 11294 2334 11346 2343
rect 11358 2377 11410 2386
rect 11358 2343 11367 2377
rect 11367 2343 11401 2377
rect 11401 2343 11410 2377
rect 11358 2334 11410 2343
rect 11422 2377 11474 2386
rect 11422 2343 11439 2377
rect 11439 2343 11473 2377
rect 11473 2343 11474 2377
rect 11422 2334 11474 2343
rect 11486 2377 11538 2386
rect 11550 2377 11602 2386
rect 11614 2377 11666 2386
rect 11678 2377 11730 2386
rect 11742 2377 11794 2386
rect 11806 2377 11858 2386
rect 11486 2343 11511 2377
rect 11511 2343 11538 2377
rect 11550 2343 11583 2377
rect 11583 2343 11602 2377
rect 11614 2343 11617 2377
rect 11617 2343 11655 2377
rect 11655 2343 11666 2377
rect 11678 2343 11689 2377
rect 11689 2343 11727 2377
rect 11727 2343 11730 2377
rect 11742 2343 11761 2377
rect 11761 2343 11794 2377
rect 11806 2343 11833 2377
rect 11833 2343 11858 2377
rect 11486 2334 11538 2343
rect 11550 2334 11602 2343
rect 11614 2334 11666 2343
rect 11678 2334 11730 2343
rect 11742 2334 11794 2343
rect 11806 2334 11858 2343
rect 11870 2377 11922 2386
rect 11870 2343 11871 2377
rect 11871 2343 11905 2377
rect 11905 2343 11922 2377
rect 11870 2334 11922 2343
rect 11934 2377 11986 2386
rect 11934 2343 11943 2377
rect 11943 2343 11977 2377
rect 11977 2343 11986 2377
rect 11934 2334 11986 2343
rect 11998 2377 12050 2386
rect 11998 2343 12015 2377
rect 12015 2343 12049 2377
rect 12049 2343 12050 2377
rect 11998 2334 12050 2343
rect 12062 2377 12114 2386
rect 12126 2377 12178 2386
rect 12190 2377 12242 2386
rect 12254 2377 12306 2386
rect 12318 2377 12370 2386
rect 12382 2377 12434 2386
rect 12062 2343 12087 2377
rect 12087 2343 12114 2377
rect 12126 2343 12159 2377
rect 12159 2343 12178 2377
rect 12190 2343 12193 2377
rect 12193 2343 12231 2377
rect 12231 2343 12242 2377
rect 12254 2343 12265 2377
rect 12265 2343 12303 2377
rect 12303 2343 12306 2377
rect 12318 2343 12337 2377
rect 12337 2343 12370 2377
rect 12382 2343 12409 2377
rect 12409 2343 12434 2377
rect 12062 2334 12114 2343
rect 12126 2334 12178 2343
rect 12190 2334 12242 2343
rect 12254 2334 12306 2343
rect 12318 2334 12370 2343
rect 12382 2334 12434 2343
rect 12446 2377 12498 2386
rect 12446 2343 12447 2377
rect 12447 2343 12481 2377
rect 12481 2343 12498 2377
rect 12446 2334 12498 2343
rect -306 1817 -254 1826
rect -306 1783 -297 1817
rect -297 1783 -263 1817
rect -263 1783 -254 1817
rect -306 1774 -254 1783
rect 12814 1817 12866 1826
rect 12814 1783 12823 1817
rect 12823 1783 12857 1817
rect 12857 1783 12866 1817
rect 12814 1774 12866 1783
rect 62 1257 114 1266
rect 62 1223 79 1257
rect 79 1223 113 1257
rect 113 1223 114 1257
rect 62 1214 114 1223
rect 126 1257 178 1266
rect 190 1257 242 1266
rect 254 1257 306 1266
rect 318 1257 370 1266
rect 382 1257 434 1266
rect 446 1257 498 1266
rect 126 1223 151 1257
rect 151 1223 178 1257
rect 190 1223 223 1257
rect 223 1223 242 1257
rect 254 1223 257 1257
rect 257 1223 295 1257
rect 295 1223 306 1257
rect 318 1223 329 1257
rect 329 1223 367 1257
rect 367 1223 370 1257
rect 382 1223 401 1257
rect 401 1223 434 1257
rect 446 1223 473 1257
rect 473 1223 498 1257
rect 126 1214 178 1223
rect 190 1214 242 1223
rect 254 1214 306 1223
rect 318 1214 370 1223
rect 382 1214 434 1223
rect 446 1214 498 1223
rect 510 1257 562 1266
rect 510 1223 511 1257
rect 511 1223 545 1257
rect 545 1223 562 1257
rect 510 1214 562 1223
rect 574 1257 626 1266
rect 574 1223 583 1257
rect 583 1223 617 1257
rect 617 1223 626 1257
rect 574 1214 626 1223
rect 638 1257 690 1266
rect 638 1223 655 1257
rect 655 1223 689 1257
rect 689 1223 690 1257
rect 638 1214 690 1223
rect 702 1257 754 1266
rect 766 1257 818 1266
rect 830 1257 882 1266
rect 894 1257 946 1266
rect 958 1257 1010 1266
rect 1022 1257 1074 1266
rect 702 1223 727 1257
rect 727 1223 754 1257
rect 766 1223 799 1257
rect 799 1223 818 1257
rect 830 1223 833 1257
rect 833 1223 871 1257
rect 871 1223 882 1257
rect 894 1223 905 1257
rect 905 1223 943 1257
rect 943 1223 946 1257
rect 958 1223 977 1257
rect 977 1223 1010 1257
rect 1022 1223 1049 1257
rect 1049 1223 1074 1257
rect 702 1214 754 1223
rect 766 1214 818 1223
rect 830 1214 882 1223
rect 894 1214 946 1223
rect 958 1214 1010 1223
rect 1022 1214 1074 1223
rect 1086 1257 1138 1266
rect 1086 1223 1087 1257
rect 1087 1223 1121 1257
rect 1121 1223 1138 1257
rect 1086 1214 1138 1223
rect 1150 1257 1202 1266
rect 1150 1223 1159 1257
rect 1159 1223 1193 1257
rect 1193 1223 1202 1257
rect 1150 1214 1202 1223
rect 1214 1257 1266 1266
rect 1214 1223 1231 1257
rect 1231 1223 1265 1257
rect 1265 1223 1266 1257
rect 1214 1214 1266 1223
rect 1278 1257 1330 1266
rect 1342 1257 1394 1266
rect 1406 1257 1458 1266
rect 1470 1257 1522 1266
rect 1534 1257 1586 1266
rect 1598 1257 1650 1266
rect 1278 1223 1303 1257
rect 1303 1223 1330 1257
rect 1342 1223 1375 1257
rect 1375 1223 1394 1257
rect 1406 1223 1409 1257
rect 1409 1223 1447 1257
rect 1447 1223 1458 1257
rect 1470 1223 1481 1257
rect 1481 1223 1519 1257
rect 1519 1223 1522 1257
rect 1534 1223 1553 1257
rect 1553 1223 1586 1257
rect 1598 1223 1625 1257
rect 1625 1223 1650 1257
rect 1278 1214 1330 1223
rect 1342 1214 1394 1223
rect 1406 1214 1458 1223
rect 1470 1214 1522 1223
rect 1534 1214 1586 1223
rect 1598 1214 1650 1223
rect 1662 1257 1714 1266
rect 1662 1223 1663 1257
rect 1663 1223 1697 1257
rect 1697 1223 1714 1257
rect 1662 1214 1714 1223
rect 1726 1257 1778 1266
rect 1726 1223 1735 1257
rect 1735 1223 1769 1257
rect 1769 1223 1778 1257
rect 1726 1214 1778 1223
rect 1790 1257 1842 1266
rect 1790 1223 1807 1257
rect 1807 1223 1841 1257
rect 1841 1223 1842 1257
rect 1790 1214 1842 1223
rect 1854 1257 1906 1266
rect 1918 1257 1970 1266
rect 1982 1257 2034 1266
rect 2046 1257 2098 1266
rect 2110 1257 2162 1266
rect 2174 1257 2226 1266
rect 1854 1223 1879 1257
rect 1879 1223 1906 1257
rect 1918 1223 1951 1257
rect 1951 1223 1970 1257
rect 1982 1223 1985 1257
rect 1985 1223 2023 1257
rect 2023 1223 2034 1257
rect 2046 1223 2057 1257
rect 2057 1223 2095 1257
rect 2095 1223 2098 1257
rect 2110 1223 2129 1257
rect 2129 1223 2162 1257
rect 2174 1223 2201 1257
rect 2201 1223 2226 1257
rect 1854 1214 1906 1223
rect 1918 1214 1970 1223
rect 1982 1214 2034 1223
rect 2046 1214 2098 1223
rect 2110 1214 2162 1223
rect 2174 1214 2226 1223
rect 2238 1257 2290 1266
rect 2238 1223 2239 1257
rect 2239 1223 2273 1257
rect 2273 1223 2290 1257
rect 2238 1214 2290 1223
rect 2302 1257 2354 1266
rect 2302 1223 2311 1257
rect 2311 1223 2345 1257
rect 2345 1223 2354 1257
rect 2302 1214 2354 1223
rect 2366 1257 2418 1266
rect 2366 1223 2383 1257
rect 2383 1223 2417 1257
rect 2417 1223 2418 1257
rect 2366 1214 2418 1223
rect 2430 1257 2482 1266
rect 2494 1257 2546 1266
rect 2558 1257 2610 1266
rect 2622 1257 2674 1266
rect 2686 1257 2738 1266
rect 2750 1257 2802 1266
rect 2430 1223 2455 1257
rect 2455 1223 2482 1257
rect 2494 1223 2527 1257
rect 2527 1223 2546 1257
rect 2558 1223 2561 1257
rect 2561 1223 2599 1257
rect 2599 1223 2610 1257
rect 2622 1223 2633 1257
rect 2633 1223 2671 1257
rect 2671 1223 2674 1257
rect 2686 1223 2705 1257
rect 2705 1223 2738 1257
rect 2750 1223 2777 1257
rect 2777 1223 2802 1257
rect 2430 1214 2482 1223
rect 2494 1214 2546 1223
rect 2558 1214 2610 1223
rect 2622 1214 2674 1223
rect 2686 1214 2738 1223
rect 2750 1214 2802 1223
rect 2814 1257 2866 1266
rect 2814 1223 2815 1257
rect 2815 1223 2849 1257
rect 2849 1223 2866 1257
rect 2814 1214 2866 1223
rect 2878 1257 2930 1266
rect 2878 1223 2887 1257
rect 2887 1223 2921 1257
rect 2921 1223 2930 1257
rect 2878 1214 2930 1223
rect 2942 1257 2994 1266
rect 2942 1223 2959 1257
rect 2959 1223 2993 1257
rect 2993 1223 2994 1257
rect 2942 1214 2994 1223
rect 3006 1257 3058 1266
rect 3070 1257 3122 1266
rect 3134 1257 3186 1266
rect 3198 1257 3250 1266
rect 3262 1257 3314 1266
rect 3326 1257 3378 1266
rect 3006 1223 3031 1257
rect 3031 1223 3058 1257
rect 3070 1223 3103 1257
rect 3103 1223 3122 1257
rect 3134 1223 3137 1257
rect 3137 1223 3175 1257
rect 3175 1223 3186 1257
rect 3198 1223 3209 1257
rect 3209 1223 3247 1257
rect 3247 1223 3250 1257
rect 3262 1223 3281 1257
rect 3281 1223 3314 1257
rect 3326 1223 3353 1257
rect 3353 1223 3378 1257
rect 3006 1214 3058 1223
rect 3070 1214 3122 1223
rect 3134 1214 3186 1223
rect 3198 1214 3250 1223
rect 3262 1214 3314 1223
rect 3326 1214 3378 1223
rect 3390 1257 3442 1266
rect 3390 1223 3391 1257
rect 3391 1223 3425 1257
rect 3425 1223 3442 1257
rect 3390 1214 3442 1223
rect 3454 1257 3506 1266
rect 3454 1223 3463 1257
rect 3463 1223 3497 1257
rect 3497 1223 3506 1257
rect 3454 1214 3506 1223
rect 3518 1257 3570 1266
rect 3518 1223 3535 1257
rect 3535 1223 3569 1257
rect 3569 1223 3570 1257
rect 3518 1214 3570 1223
rect 3582 1257 3634 1266
rect 3646 1257 3698 1266
rect 3710 1257 3762 1266
rect 3774 1257 3826 1266
rect 3838 1257 3890 1266
rect 3902 1257 3954 1266
rect 3582 1223 3607 1257
rect 3607 1223 3634 1257
rect 3646 1223 3679 1257
rect 3679 1223 3698 1257
rect 3710 1223 3713 1257
rect 3713 1223 3751 1257
rect 3751 1223 3762 1257
rect 3774 1223 3785 1257
rect 3785 1223 3823 1257
rect 3823 1223 3826 1257
rect 3838 1223 3857 1257
rect 3857 1223 3890 1257
rect 3902 1223 3929 1257
rect 3929 1223 3954 1257
rect 3582 1214 3634 1223
rect 3646 1214 3698 1223
rect 3710 1214 3762 1223
rect 3774 1214 3826 1223
rect 3838 1214 3890 1223
rect 3902 1214 3954 1223
rect 3966 1257 4018 1266
rect 3966 1223 3967 1257
rect 3967 1223 4001 1257
rect 4001 1223 4018 1257
rect 3966 1214 4018 1223
rect 62 937 114 946
rect 62 903 79 937
rect 79 903 113 937
rect 113 903 114 937
rect 62 894 114 903
rect 126 937 178 946
rect 190 937 242 946
rect 254 937 306 946
rect 318 937 370 946
rect 382 937 434 946
rect 446 937 498 946
rect 126 903 151 937
rect 151 903 178 937
rect 190 903 223 937
rect 223 903 242 937
rect 254 903 257 937
rect 257 903 295 937
rect 295 903 306 937
rect 318 903 329 937
rect 329 903 367 937
rect 367 903 370 937
rect 382 903 401 937
rect 401 903 434 937
rect 446 903 473 937
rect 473 903 498 937
rect 126 894 178 903
rect 190 894 242 903
rect 254 894 306 903
rect 318 894 370 903
rect 382 894 434 903
rect 446 894 498 903
rect 510 937 562 946
rect 510 903 511 937
rect 511 903 545 937
rect 545 903 562 937
rect 510 894 562 903
rect 574 937 626 946
rect 574 903 583 937
rect 583 903 617 937
rect 617 903 626 937
rect 574 894 626 903
rect 638 937 690 946
rect 638 903 655 937
rect 655 903 689 937
rect 689 903 690 937
rect 638 894 690 903
rect 702 937 754 946
rect 766 937 818 946
rect 830 937 882 946
rect 894 937 946 946
rect 958 937 1010 946
rect 1022 937 1074 946
rect 702 903 727 937
rect 727 903 754 937
rect 766 903 799 937
rect 799 903 818 937
rect 830 903 833 937
rect 833 903 871 937
rect 871 903 882 937
rect 894 903 905 937
rect 905 903 943 937
rect 943 903 946 937
rect 958 903 977 937
rect 977 903 1010 937
rect 1022 903 1049 937
rect 1049 903 1074 937
rect 702 894 754 903
rect 766 894 818 903
rect 830 894 882 903
rect 894 894 946 903
rect 958 894 1010 903
rect 1022 894 1074 903
rect 1086 937 1138 946
rect 1086 903 1087 937
rect 1087 903 1121 937
rect 1121 903 1138 937
rect 1086 894 1138 903
rect 1150 937 1202 946
rect 1150 903 1159 937
rect 1159 903 1193 937
rect 1193 903 1202 937
rect 1150 894 1202 903
rect 1214 937 1266 946
rect 1214 903 1231 937
rect 1231 903 1265 937
rect 1265 903 1266 937
rect 1214 894 1266 903
rect 1278 937 1330 946
rect 1342 937 1394 946
rect 1406 937 1458 946
rect 1470 937 1522 946
rect 1534 937 1586 946
rect 1598 937 1650 946
rect 1278 903 1303 937
rect 1303 903 1330 937
rect 1342 903 1375 937
rect 1375 903 1394 937
rect 1406 903 1409 937
rect 1409 903 1447 937
rect 1447 903 1458 937
rect 1470 903 1481 937
rect 1481 903 1519 937
rect 1519 903 1522 937
rect 1534 903 1553 937
rect 1553 903 1586 937
rect 1598 903 1625 937
rect 1625 903 1650 937
rect 1278 894 1330 903
rect 1342 894 1394 903
rect 1406 894 1458 903
rect 1470 894 1522 903
rect 1534 894 1586 903
rect 1598 894 1650 903
rect 1662 937 1714 946
rect 1662 903 1663 937
rect 1663 903 1697 937
rect 1697 903 1714 937
rect 1662 894 1714 903
rect 1726 937 1778 946
rect 1726 903 1735 937
rect 1735 903 1769 937
rect 1769 903 1778 937
rect 1726 894 1778 903
rect 1790 937 1842 946
rect 1790 903 1807 937
rect 1807 903 1841 937
rect 1841 903 1842 937
rect 1790 894 1842 903
rect 1854 937 1906 946
rect 1918 937 1970 946
rect 1982 937 2034 946
rect 2046 937 2098 946
rect 2110 937 2162 946
rect 2174 937 2226 946
rect 1854 903 1879 937
rect 1879 903 1906 937
rect 1918 903 1951 937
rect 1951 903 1970 937
rect 1982 903 1985 937
rect 1985 903 2023 937
rect 2023 903 2034 937
rect 2046 903 2057 937
rect 2057 903 2095 937
rect 2095 903 2098 937
rect 2110 903 2129 937
rect 2129 903 2162 937
rect 2174 903 2201 937
rect 2201 903 2226 937
rect 1854 894 1906 903
rect 1918 894 1970 903
rect 1982 894 2034 903
rect 2046 894 2098 903
rect 2110 894 2162 903
rect 2174 894 2226 903
rect 2238 937 2290 946
rect 2238 903 2239 937
rect 2239 903 2273 937
rect 2273 903 2290 937
rect 2238 894 2290 903
rect 2302 937 2354 946
rect 2302 903 2311 937
rect 2311 903 2345 937
rect 2345 903 2354 937
rect 2302 894 2354 903
rect 2366 937 2418 946
rect 2366 903 2383 937
rect 2383 903 2417 937
rect 2417 903 2418 937
rect 2366 894 2418 903
rect 2430 937 2482 946
rect 2494 937 2546 946
rect 2558 937 2610 946
rect 2622 937 2674 946
rect 2686 937 2738 946
rect 2750 937 2802 946
rect 2430 903 2455 937
rect 2455 903 2482 937
rect 2494 903 2527 937
rect 2527 903 2546 937
rect 2558 903 2561 937
rect 2561 903 2599 937
rect 2599 903 2610 937
rect 2622 903 2633 937
rect 2633 903 2671 937
rect 2671 903 2674 937
rect 2686 903 2705 937
rect 2705 903 2738 937
rect 2750 903 2777 937
rect 2777 903 2802 937
rect 2430 894 2482 903
rect 2494 894 2546 903
rect 2558 894 2610 903
rect 2622 894 2674 903
rect 2686 894 2738 903
rect 2750 894 2802 903
rect 2814 937 2866 946
rect 2814 903 2815 937
rect 2815 903 2849 937
rect 2849 903 2866 937
rect 2814 894 2866 903
rect 2878 937 2930 946
rect 2878 903 2887 937
rect 2887 903 2921 937
rect 2921 903 2930 937
rect 2878 894 2930 903
rect 2942 937 2994 946
rect 2942 903 2959 937
rect 2959 903 2993 937
rect 2993 903 2994 937
rect 2942 894 2994 903
rect 3006 937 3058 946
rect 3070 937 3122 946
rect 3134 937 3186 946
rect 3198 937 3250 946
rect 3262 937 3314 946
rect 3326 937 3378 946
rect 3006 903 3031 937
rect 3031 903 3058 937
rect 3070 903 3103 937
rect 3103 903 3122 937
rect 3134 903 3137 937
rect 3137 903 3175 937
rect 3175 903 3186 937
rect 3198 903 3209 937
rect 3209 903 3247 937
rect 3247 903 3250 937
rect 3262 903 3281 937
rect 3281 903 3314 937
rect 3326 903 3353 937
rect 3353 903 3378 937
rect 3006 894 3058 903
rect 3070 894 3122 903
rect 3134 894 3186 903
rect 3198 894 3250 903
rect 3262 894 3314 903
rect 3326 894 3378 903
rect 3390 937 3442 946
rect 3390 903 3391 937
rect 3391 903 3425 937
rect 3425 903 3442 937
rect 3390 894 3442 903
rect 3454 937 3506 946
rect 3454 903 3463 937
rect 3463 903 3497 937
rect 3497 903 3506 937
rect 3454 894 3506 903
rect 3518 937 3570 946
rect 3518 903 3535 937
rect 3535 903 3569 937
rect 3569 903 3570 937
rect 3518 894 3570 903
rect 3582 937 3634 946
rect 3646 937 3698 946
rect 3710 937 3762 946
rect 3774 937 3826 946
rect 3838 937 3890 946
rect 3902 937 3954 946
rect 3582 903 3607 937
rect 3607 903 3634 937
rect 3646 903 3679 937
rect 3679 903 3698 937
rect 3710 903 3713 937
rect 3713 903 3751 937
rect 3751 903 3762 937
rect 3774 903 3785 937
rect 3785 903 3823 937
rect 3823 903 3826 937
rect 3838 903 3857 937
rect 3857 903 3890 937
rect 3902 903 3929 937
rect 3929 903 3954 937
rect 3582 894 3634 903
rect 3646 894 3698 903
rect 3710 894 3762 903
rect 3774 894 3826 903
rect 3838 894 3890 903
rect 3902 894 3954 903
rect 3966 937 4018 946
rect 3966 903 3967 937
rect 3967 903 4001 937
rect 4001 903 4018 937
rect 3966 894 4018 903
rect 4174 894 4226 946
rect -146 94 -94 146
rect 62 137 114 146
rect 62 103 79 137
rect 79 103 113 137
rect 113 103 114 137
rect 62 94 114 103
rect 126 137 178 146
rect 190 137 242 146
rect 254 137 306 146
rect 318 137 370 146
rect 382 137 434 146
rect 446 137 498 146
rect 126 103 151 137
rect 151 103 178 137
rect 190 103 223 137
rect 223 103 242 137
rect 254 103 257 137
rect 257 103 295 137
rect 295 103 306 137
rect 318 103 329 137
rect 329 103 367 137
rect 367 103 370 137
rect 382 103 401 137
rect 401 103 434 137
rect 446 103 473 137
rect 473 103 498 137
rect 126 94 178 103
rect 190 94 242 103
rect 254 94 306 103
rect 318 94 370 103
rect 382 94 434 103
rect 446 94 498 103
rect 510 137 562 146
rect 510 103 511 137
rect 511 103 545 137
rect 545 103 562 137
rect 510 94 562 103
rect 574 137 626 146
rect 574 103 583 137
rect 583 103 617 137
rect 617 103 626 137
rect 574 94 626 103
rect 638 137 690 146
rect 638 103 655 137
rect 655 103 689 137
rect 689 103 690 137
rect 638 94 690 103
rect 702 137 754 146
rect 766 137 818 146
rect 830 137 882 146
rect 894 137 946 146
rect 958 137 1010 146
rect 1022 137 1074 146
rect 702 103 727 137
rect 727 103 754 137
rect 766 103 799 137
rect 799 103 818 137
rect 830 103 833 137
rect 833 103 871 137
rect 871 103 882 137
rect 894 103 905 137
rect 905 103 943 137
rect 943 103 946 137
rect 958 103 977 137
rect 977 103 1010 137
rect 1022 103 1049 137
rect 1049 103 1074 137
rect 702 94 754 103
rect 766 94 818 103
rect 830 94 882 103
rect 894 94 946 103
rect 958 94 1010 103
rect 1022 94 1074 103
rect 1086 137 1138 146
rect 1086 103 1087 137
rect 1087 103 1121 137
rect 1121 103 1138 137
rect 1086 94 1138 103
rect 1150 137 1202 146
rect 1150 103 1159 137
rect 1159 103 1193 137
rect 1193 103 1202 137
rect 1150 94 1202 103
rect 1214 137 1266 146
rect 1214 103 1231 137
rect 1231 103 1265 137
rect 1265 103 1266 137
rect 1214 94 1266 103
rect 1278 137 1330 146
rect 1342 137 1394 146
rect 1406 137 1458 146
rect 1470 137 1522 146
rect 1534 137 1586 146
rect 1598 137 1650 146
rect 1278 103 1303 137
rect 1303 103 1330 137
rect 1342 103 1375 137
rect 1375 103 1394 137
rect 1406 103 1409 137
rect 1409 103 1447 137
rect 1447 103 1458 137
rect 1470 103 1481 137
rect 1481 103 1519 137
rect 1519 103 1522 137
rect 1534 103 1553 137
rect 1553 103 1586 137
rect 1598 103 1625 137
rect 1625 103 1650 137
rect 1278 94 1330 103
rect 1342 94 1394 103
rect 1406 94 1458 103
rect 1470 94 1522 103
rect 1534 94 1586 103
rect 1598 94 1650 103
rect 1662 137 1714 146
rect 1662 103 1663 137
rect 1663 103 1697 137
rect 1697 103 1714 137
rect 1662 94 1714 103
rect 1726 137 1778 146
rect 1726 103 1735 137
rect 1735 103 1769 137
rect 1769 103 1778 137
rect 1726 94 1778 103
rect 1790 137 1842 146
rect 1790 103 1807 137
rect 1807 103 1841 137
rect 1841 103 1842 137
rect 1790 94 1842 103
rect 1854 137 1906 146
rect 1918 137 1970 146
rect 1982 137 2034 146
rect 2046 137 2098 146
rect 2110 137 2162 146
rect 2174 137 2226 146
rect 1854 103 1879 137
rect 1879 103 1906 137
rect 1918 103 1951 137
rect 1951 103 1970 137
rect 1982 103 1985 137
rect 1985 103 2023 137
rect 2023 103 2034 137
rect 2046 103 2057 137
rect 2057 103 2095 137
rect 2095 103 2098 137
rect 2110 103 2129 137
rect 2129 103 2162 137
rect 2174 103 2201 137
rect 2201 103 2226 137
rect 1854 94 1906 103
rect 1918 94 1970 103
rect 1982 94 2034 103
rect 2046 94 2098 103
rect 2110 94 2162 103
rect 2174 94 2226 103
rect 2238 137 2290 146
rect 2238 103 2239 137
rect 2239 103 2273 137
rect 2273 103 2290 137
rect 2238 94 2290 103
rect 2302 137 2354 146
rect 2302 103 2311 137
rect 2311 103 2345 137
rect 2345 103 2354 137
rect 2302 94 2354 103
rect 2366 137 2418 146
rect 2366 103 2383 137
rect 2383 103 2417 137
rect 2417 103 2418 137
rect 2366 94 2418 103
rect 2430 137 2482 146
rect 2494 137 2546 146
rect 2558 137 2610 146
rect 2622 137 2674 146
rect 2686 137 2738 146
rect 2750 137 2802 146
rect 2430 103 2455 137
rect 2455 103 2482 137
rect 2494 103 2527 137
rect 2527 103 2546 137
rect 2558 103 2561 137
rect 2561 103 2599 137
rect 2599 103 2610 137
rect 2622 103 2633 137
rect 2633 103 2671 137
rect 2671 103 2674 137
rect 2686 103 2705 137
rect 2705 103 2738 137
rect 2750 103 2777 137
rect 2777 103 2802 137
rect 2430 94 2482 103
rect 2494 94 2546 103
rect 2558 94 2610 103
rect 2622 94 2674 103
rect 2686 94 2738 103
rect 2750 94 2802 103
rect 2814 137 2866 146
rect 2814 103 2815 137
rect 2815 103 2849 137
rect 2849 103 2866 137
rect 2814 94 2866 103
rect 2878 137 2930 146
rect 2878 103 2887 137
rect 2887 103 2921 137
rect 2921 103 2930 137
rect 2878 94 2930 103
rect 2942 137 2994 146
rect 2942 103 2959 137
rect 2959 103 2993 137
rect 2993 103 2994 137
rect 2942 94 2994 103
rect 3006 137 3058 146
rect 3070 137 3122 146
rect 3134 137 3186 146
rect 3198 137 3250 146
rect 3262 137 3314 146
rect 3326 137 3378 146
rect 3006 103 3031 137
rect 3031 103 3058 137
rect 3070 103 3103 137
rect 3103 103 3122 137
rect 3134 103 3137 137
rect 3137 103 3175 137
rect 3175 103 3186 137
rect 3198 103 3209 137
rect 3209 103 3247 137
rect 3247 103 3250 137
rect 3262 103 3281 137
rect 3281 103 3314 137
rect 3326 103 3353 137
rect 3353 103 3378 137
rect 3006 94 3058 103
rect 3070 94 3122 103
rect 3134 94 3186 103
rect 3198 94 3250 103
rect 3262 94 3314 103
rect 3326 94 3378 103
rect 3390 137 3442 146
rect 3390 103 3391 137
rect 3391 103 3425 137
rect 3425 103 3442 137
rect 3390 94 3442 103
rect 3454 137 3506 146
rect 3454 103 3463 137
rect 3463 103 3497 137
rect 3497 103 3506 137
rect 3454 94 3506 103
rect 3518 137 3570 146
rect 3518 103 3535 137
rect 3535 103 3569 137
rect 3569 103 3570 137
rect 3518 94 3570 103
rect 3582 137 3634 146
rect 3646 137 3698 146
rect 3710 137 3762 146
rect 3774 137 3826 146
rect 3838 137 3890 146
rect 3902 137 3954 146
rect 3582 103 3607 137
rect 3607 103 3634 137
rect 3646 103 3679 137
rect 3679 103 3698 137
rect 3710 103 3713 137
rect 3713 103 3751 137
rect 3751 103 3762 137
rect 3774 103 3785 137
rect 3785 103 3823 137
rect 3823 103 3826 137
rect 3838 103 3857 137
rect 3857 103 3890 137
rect 3902 103 3929 137
rect 3929 103 3954 137
rect 3582 94 3634 103
rect 3646 94 3698 103
rect 3710 94 3762 103
rect 3774 94 3826 103
rect 3838 94 3890 103
rect 3902 94 3954 103
rect 3966 137 4018 146
rect 3966 103 3967 137
rect 3967 103 4001 137
rect 4001 103 4018 137
rect 3966 94 4018 103
rect 62 -183 114 -174
rect 62 -217 79 -183
rect 79 -217 113 -183
rect 113 -217 114 -183
rect 62 -226 114 -217
rect 126 -183 178 -174
rect 190 -183 242 -174
rect 254 -183 306 -174
rect 318 -183 370 -174
rect 382 -183 434 -174
rect 446 -183 498 -174
rect 126 -217 151 -183
rect 151 -217 178 -183
rect 190 -217 223 -183
rect 223 -217 242 -183
rect 254 -217 257 -183
rect 257 -217 295 -183
rect 295 -217 306 -183
rect 318 -217 329 -183
rect 329 -217 367 -183
rect 367 -217 370 -183
rect 382 -217 401 -183
rect 401 -217 434 -183
rect 446 -217 473 -183
rect 473 -217 498 -183
rect 126 -226 178 -217
rect 190 -226 242 -217
rect 254 -226 306 -217
rect 318 -226 370 -217
rect 382 -226 434 -217
rect 446 -226 498 -217
rect 510 -183 562 -174
rect 510 -217 511 -183
rect 511 -217 545 -183
rect 545 -217 562 -183
rect 510 -226 562 -217
rect 574 -183 626 -174
rect 574 -217 583 -183
rect 583 -217 617 -183
rect 617 -217 626 -183
rect 574 -226 626 -217
rect 638 -183 690 -174
rect 638 -217 655 -183
rect 655 -217 689 -183
rect 689 -217 690 -183
rect 638 -226 690 -217
rect 702 -183 754 -174
rect 766 -183 818 -174
rect 830 -183 882 -174
rect 894 -183 946 -174
rect 958 -183 1010 -174
rect 1022 -183 1074 -174
rect 702 -217 727 -183
rect 727 -217 754 -183
rect 766 -217 799 -183
rect 799 -217 818 -183
rect 830 -217 833 -183
rect 833 -217 871 -183
rect 871 -217 882 -183
rect 894 -217 905 -183
rect 905 -217 943 -183
rect 943 -217 946 -183
rect 958 -217 977 -183
rect 977 -217 1010 -183
rect 1022 -217 1049 -183
rect 1049 -217 1074 -183
rect 702 -226 754 -217
rect 766 -226 818 -217
rect 830 -226 882 -217
rect 894 -226 946 -217
rect 958 -226 1010 -217
rect 1022 -226 1074 -217
rect 1086 -183 1138 -174
rect 1086 -217 1087 -183
rect 1087 -217 1121 -183
rect 1121 -217 1138 -183
rect 1086 -226 1138 -217
rect 1150 -183 1202 -174
rect 1150 -217 1159 -183
rect 1159 -217 1193 -183
rect 1193 -217 1202 -183
rect 1150 -226 1202 -217
rect 1214 -183 1266 -174
rect 1214 -217 1231 -183
rect 1231 -217 1265 -183
rect 1265 -217 1266 -183
rect 1214 -226 1266 -217
rect 1278 -183 1330 -174
rect 1342 -183 1394 -174
rect 1406 -183 1458 -174
rect 1470 -183 1522 -174
rect 1534 -183 1586 -174
rect 1598 -183 1650 -174
rect 1278 -217 1303 -183
rect 1303 -217 1330 -183
rect 1342 -217 1375 -183
rect 1375 -217 1394 -183
rect 1406 -217 1409 -183
rect 1409 -217 1447 -183
rect 1447 -217 1458 -183
rect 1470 -217 1481 -183
rect 1481 -217 1519 -183
rect 1519 -217 1522 -183
rect 1534 -217 1553 -183
rect 1553 -217 1586 -183
rect 1598 -217 1625 -183
rect 1625 -217 1650 -183
rect 1278 -226 1330 -217
rect 1342 -226 1394 -217
rect 1406 -226 1458 -217
rect 1470 -226 1522 -217
rect 1534 -226 1586 -217
rect 1598 -226 1650 -217
rect 1662 -183 1714 -174
rect 1662 -217 1663 -183
rect 1663 -217 1697 -183
rect 1697 -217 1714 -183
rect 1662 -226 1714 -217
rect 1726 -183 1778 -174
rect 1726 -217 1735 -183
rect 1735 -217 1769 -183
rect 1769 -217 1778 -183
rect 1726 -226 1778 -217
rect 1790 -183 1842 -174
rect 1790 -217 1807 -183
rect 1807 -217 1841 -183
rect 1841 -217 1842 -183
rect 1790 -226 1842 -217
rect 1854 -183 1906 -174
rect 1918 -183 1970 -174
rect 1982 -183 2034 -174
rect 2046 -183 2098 -174
rect 2110 -183 2162 -174
rect 2174 -183 2226 -174
rect 1854 -217 1879 -183
rect 1879 -217 1906 -183
rect 1918 -217 1951 -183
rect 1951 -217 1970 -183
rect 1982 -217 1985 -183
rect 1985 -217 2023 -183
rect 2023 -217 2034 -183
rect 2046 -217 2057 -183
rect 2057 -217 2095 -183
rect 2095 -217 2098 -183
rect 2110 -217 2129 -183
rect 2129 -217 2162 -183
rect 2174 -217 2201 -183
rect 2201 -217 2226 -183
rect 1854 -226 1906 -217
rect 1918 -226 1970 -217
rect 1982 -226 2034 -217
rect 2046 -226 2098 -217
rect 2110 -226 2162 -217
rect 2174 -226 2226 -217
rect 2238 -183 2290 -174
rect 2238 -217 2239 -183
rect 2239 -217 2273 -183
rect 2273 -217 2290 -183
rect 2238 -226 2290 -217
rect 2302 -183 2354 -174
rect 2302 -217 2311 -183
rect 2311 -217 2345 -183
rect 2345 -217 2354 -183
rect 2302 -226 2354 -217
rect 2366 -183 2418 -174
rect 2366 -217 2383 -183
rect 2383 -217 2417 -183
rect 2417 -217 2418 -183
rect 2366 -226 2418 -217
rect 2430 -183 2482 -174
rect 2494 -183 2546 -174
rect 2558 -183 2610 -174
rect 2622 -183 2674 -174
rect 2686 -183 2738 -174
rect 2750 -183 2802 -174
rect 2430 -217 2455 -183
rect 2455 -217 2482 -183
rect 2494 -217 2527 -183
rect 2527 -217 2546 -183
rect 2558 -217 2561 -183
rect 2561 -217 2599 -183
rect 2599 -217 2610 -183
rect 2622 -217 2633 -183
rect 2633 -217 2671 -183
rect 2671 -217 2674 -183
rect 2686 -217 2705 -183
rect 2705 -217 2738 -183
rect 2750 -217 2777 -183
rect 2777 -217 2802 -183
rect 2430 -226 2482 -217
rect 2494 -226 2546 -217
rect 2558 -226 2610 -217
rect 2622 -226 2674 -217
rect 2686 -226 2738 -217
rect 2750 -226 2802 -217
rect 2814 -183 2866 -174
rect 2814 -217 2815 -183
rect 2815 -217 2849 -183
rect 2849 -217 2866 -183
rect 2814 -226 2866 -217
rect 2878 -183 2930 -174
rect 2878 -217 2887 -183
rect 2887 -217 2921 -183
rect 2921 -217 2930 -183
rect 2878 -226 2930 -217
rect 2942 -183 2994 -174
rect 2942 -217 2959 -183
rect 2959 -217 2993 -183
rect 2993 -217 2994 -183
rect 2942 -226 2994 -217
rect 3006 -183 3058 -174
rect 3070 -183 3122 -174
rect 3134 -183 3186 -174
rect 3198 -183 3250 -174
rect 3262 -183 3314 -174
rect 3326 -183 3378 -174
rect 3006 -217 3031 -183
rect 3031 -217 3058 -183
rect 3070 -217 3103 -183
rect 3103 -217 3122 -183
rect 3134 -217 3137 -183
rect 3137 -217 3175 -183
rect 3175 -217 3186 -183
rect 3198 -217 3209 -183
rect 3209 -217 3247 -183
rect 3247 -217 3250 -183
rect 3262 -217 3281 -183
rect 3281 -217 3314 -183
rect 3326 -217 3353 -183
rect 3353 -217 3378 -183
rect 3006 -226 3058 -217
rect 3070 -226 3122 -217
rect 3134 -226 3186 -217
rect 3198 -226 3250 -217
rect 3262 -226 3314 -217
rect 3326 -226 3378 -217
rect 3390 -183 3442 -174
rect 3390 -217 3391 -183
rect 3391 -217 3425 -183
rect 3425 -217 3442 -183
rect 3390 -226 3442 -217
rect 3454 -183 3506 -174
rect 3454 -217 3463 -183
rect 3463 -217 3497 -183
rect 3497 -217 3506 -183
rect 3454 -226 3506 -217
rect 3518 -183 3570 -174
rect 3518 -217 3535 -183
rect 3535 -217 3569 -183
rect 3569 -217 3570 -183
rect 3518 -226 3570 -217
rect 3582 -183 3634 -174
rect 3646 -183 3698 -174
rect 3710 -183 3762 -174
rect 3774 -183 3826 -174
rect 3838 -183 3890 -174
rect 3902 -183 3954 -174
rect 3582 -217 3607 -183
rect 3607 -217 3634 -183
rect 3646 -217 3679 -183
rect 3679 -217 3698 -183
rect 3710 -217 3713 -183
rect 3713 -217 3751 -183
rect 3751 -217 3762 -183
rect 3774 -217 3785 -183
rect 3785 -217 3823 -183
rect 3823 -217 3826 -183
rect 3838 -217 3857 -183
rect 3857 -217 3890 -183
rect 3902 -217 3929 -183
rect 3929 -217 3954 -183
rect 3582 -226 3634 -217
rect 3646 -226 3698 -217
rect 3710 -226 3762 -217
rect 3774 -226 3826 -217
rect 3838 -226 3890 -217
rect 3902 -226 3954 -217
rect 3966 -183 4018 -174
rect 3966 -217 3967 -183
rect 3967 -217 4001 -183
rect 4001 -217 4018 -183
rect 3966 -226 4018 -217
rect 8542 1257 8594 1266
rect 8542 1223 8559 1257
rect 8559 1223 8593 1257
rect 8593 1223 8594 1257
rect 8542 1214 8594 1223
rect 8606 1257 8658 1266
rect 8670 1257 8722 1266
rect 8734 1257 8786 1266
rect 8798 1257 8850 1266
rect 8862 1257 8914 1266
rect 8926 1257 8978 1266
rect 8606 1223 8631 1257
rect 8631 1223 8658 1257
rect 8670 1223 8703 1257
rect 8703 1223 8722 1257
rect 8734 1223 8737 1257
rect 8737 1223 8775 1257
rect 8775 1223 8786 1257
rect 8798 1223 8809 1257
rect 8809 1223 8847 1257
rect 8847 1223 8850 1257
rect 8862 1223 8881 1257
rect 8881 1223 8914 1257
rect 8926 1223 8953 1257
rect 8953 1223 8978 1257
rect 8606 1214 8658 1223
rect 8670 1214 8722 1223
rect 8734 1214 8786 1223
rect 8798 1214 8850 1223
rect 8862 1214 8914 1223
rect 8926 1214 8978 1223
rect 8990 1257 9042 1266
rect 8990 1223 8991 1257
rect 8991 1223 9025 1257
rect 9025 1223 9042 1257
rect 8990 1214 9042 1223
rect 9054 1257 9106 1266
rect 9054 1223 9063 1257
rect 9063 1223 9097 1257
rect 9097 1223 9106 1257
rect 9054 1214 9106 1223
rect 9118 1257 9170 1266
rect 9118 1223 9135 1257
rect 9135 1223 9169 1257
rect 9169 1223 9170 1257
rect 9118 1214 9170 1223
rect 9182 1257 9234 1266
rect 9246 1257 9298 1266
rect 9310 1257 9362 1266
rect 9374 1257 9426 1266
rect 9438 1257 9490 1266
rect 9502 1257 9554 1266
rect 9182 1223 9207 1257
rect 9207 1223 9234 1257
rect 9246 1223 9279 1257
rect 9279 1223 9298 1257
rect 9310 1223 9313 1257
rect 9313 1223 9351 1257
rect 9351 1223 9362 1257
rect 9374 1223 9385 1257
rect 9385 1223 9423 1257
rect 9423 1223 9426 1257
rect 9438 1223 9457 1257
rect 9457 1223 9490 1257
rect 9502 1223 9529 1257
rect 9529 1223 9554 1257
rect 9182 1214 9234 1223
rect 9246 1214 9298 1223
rect 9310 1214 9362 1223
rect 9374 1214 9426 1223
rect 9438 1214 9490 1223
rect 9502 1214 9554 1223
rect 9566 1257 9618 1266
rect 9566 1223 9567 1257
rect 9567 1223 9601 1257
rect 9601 1223 9618 1257
rect 9566 1214 9618 1223
rect 9630 1257 9682 1266
rect 9630 1223 9639 1257
rect 9639 1223 9673 1257
rect 9673 1223 9682 1257
rect 9630 1214 9682 1223
rect 9694 1257 9746 1266
rect 9694 1223 9711 1257
rect 9711 1223 9745 1257
rect 9745 1223 9746 1257
rect 9694 1214 9746 1223
rect 9758 1257 9810 1266
rect 9822 1257 9874 1266
rect 9886 1257 9938 1266
rect 9950 1257 10002 1266
rect 10014 1257 10066 1266
rect 10078 1257 10130 1266
rect 9758 1223 9783 1257
rect 9783 1223 9810 1257
rect 9822 1223 9855 1257
rect 9855 1223 9874 1257
rect 9886 1223 9889 1257
rect 9889 1223 9927 1257
rect 9927 1223 9938 1257
rect 9950 1223 9961 1257
rect 9961 1223 9999 1257
rect 9999 1223 10002 1257
rect 10014 1223 10033 1257
rect 10033 1223 10066 1257
rect 10078 1223 10105 1257
rect 10105 1223 10130 1257
rect 9758 1214 9810 1223
rect 9822 1214 9874 1223
rect 9886 1214 9938 1223
rect 9950 1214 10002 1223
rect 10014 1214 10066 1223
rect 10078 1214 10130 1223
rect 10142 1257 10194 1266
rect 10142 1223 10143 1257
rect 10143 1223 10177 1257
rect 10177 1223 10194 1257
rect 10142 1214 10194 1223
rect 10206 1257 10258 1266
rect 10206 1223 10215 1257
rect 10215 1223 10249 1257
rect 10249 1223 10258 1257
rect 10206 1214 10258 1223
rect 10270 1257 10322 1266
rect 10270 1223 10287 1257
rect 10287 1223 10321 1257
rect 10321 1223 10322 1257
rect 10270 1214 10322 1223
rect 10334 1257 10386 1266
rect 10398 1257 10450 1266
rect 10462 1257 10514 1266
rect 10526 1257 10578 1266
rect 10590 1257 10642 1266
rect 10654 1257 10706 1266
rect 10334 1223 10359 1257
rect 10359 1223 10386 1257
rect 10398 1223 10431 1257
rect 10431 1223 10450 1257
rect 10462 1223 10465 1257
rect 10465 1223 10503 1257
rect 10503 1223 10514 1257
rect 10526 1223 10537 1257
rect 10537 1223 10575 1257
rect 10575 1223 10578 1257
rect 10590 1223 10609 1257
rect 10609 1223 10642 1257
rect 10654 1223 10681 1257
rect 10681 1223 10706 1257
rect 10334 1214 10386 1223
rect 10398 1214 10450 1223
rect 10462 1214 10514 1223
rect 10526 1214 10578 1223
rect 10590 1214 10642 1223
rect 10654 1214 10706 1223
rect 10718 1257 10770 1266
rect 10718 1223 10719 1257
rect 10719 1223 10753 1257
rect 10753 1223 10770 1257
rect 10718 1214 10770 1223
rect 10782 1257 10834 1266
rect 10782 1223 10791 1257
rect 10791 1223 10825 1257
rect 10825 1223 10834 1257
rect 10782 1214 10834 1223
rect 10846 1257 10898 1266
rect 10846 1223 10863 1257
rect 10863 1223 10897 1257
rect 10897 1223 10898 1257
rect 10846 1214 10898 1223
rect 10910 1257 10962 1266
rect 10974 1257 11026 1266
rect 11038 1257 11090 1266
rect 11102 1257 11154 1266
rect 11166 1257 11218 1266
rect 11230 1257 11282 1266
rect 10910 1223 10935 1257
rect 10935 1223 10962 1257
rect 10974 1223 11007 1257
rect 11007 1223 11026 1257
rect 11038 1223 11041 1257
rect 11041 1223 11079 1257
rect 11079 1223 11090 1257
rect 11102 1223 11113 1257
rect 11113 1223 11151 1257
rect 11151 1223 11154 1257
rect 11166 1223 11185 1257
rect 11185 1223 11218 1257
rect 11230 1223 11257 1257
rect 11257 1223 11282 1257
rect 10910 1214 10962 1223
rect 10974 1214 11026 1223
rect 11038 1214 11090 1223
rect 11102 1214 11154 1223
rect 11166 1214 11218 1223
rect 11230 1214 11282 1223
rect 11294 1257 11346 1266
rect 11294 1223 11295 1257
rect 11295 1223 11329 1257
rect 11329 1223 11346 1257
rect 11294 1214 11346 1223
rect 11358 1257 11410 1266
rect 11358 1223 11367 1257
rect 11367 1223 11401 1257
rect 11401 1223 11410 1257
rect 11358 1214 11410 1223
rect 11422 1257 11474 1266
rect 11422 1223 11439 1257
rect 11439 1223 11473 1257
rect 11473 1223 11474 1257
rect 11422 1214 11474 1223
rect 11486 1257 11538 1266
rect 11550 1257 11602 1266
rect 11614 1257 11666 1266
rect 11678 1257 11730 1266
rect 11742 1257 11794 1266
rect 11806 1257 11858 1266
rect 11486 1223 11511 1257
rect 11511 1223 11538 1257
rect 11550 1223 11583 1257
rect 11583 1223 11602 1257
rect 11614 1223 11617 1257
rect 11617 1223 11655 1257
rect 11655 1223 11666 1257
rect 11678 1223 11689 1257
rect 11689 1223 11727 1257
rect 11727 1223 11730 1257
rect 11742 1223 11761 1257
rect 11761 1223 11794 1257
rect 11806 1223 11833 1257
rect 11833 1223 11858 1257
rect 11486 1214 11538 1223
rect 11550 1214 11602 1223
rect 11614 1214 11666 1223
rect 11678 1214 11730 1223
rect 11742 1214 11794 1223
rect 11806 1214 11858 1223
rect 11870 1257 11922 1266
rect 11870 1223 11871 1257
rect 11871 1223 11905 1257
rect 11905 1223 11922 1257
rect 11870 1214 11922 1223
rect 11934 1257 11986 1266
rect 11934 1223 11943 1257
rect 11943 1223 11977 1257
rect 11977 1223 11986 1257
rect 11934 1214 11986 1223
rect 11998 1257 12050 1266
rect 11998 1223 12015 1257
rect 12015 1223 12049 1257
rect 12049 1223 12050 1257
rect 11998 1214 12050 1223
rect 12062 1257 12114 1266
rect 12126 1257 12178 1266
rect 12190 1257 12242 1266
rect 12254 1257 12306 1266
rect 12318 1257 12370 1266
rect 12382 1257 12434 1266
rect 12062 1223 12087 1257
rect 12087 1223 12114 1257
rect 12126 1223 12159 1257
rect 12159 1223 12178 1257
rect 12190 1223 12193 1257
rect 12193 1223 12231 1257
rect 12231 1223 12242 1257
rect 12254 1223 12265 1257
rect 12265 1223 12303 1257
rect 12303 1223 12306 1257
rect 12318 1223 12337 1257
rect 12337 1223 12370 1257
rect 12382 1223 12409 1257
rect 12409 1223 12434 1257
rect 12062 1214 12114 1223
rect 12126 1214 12178 1223
rect 12190 1214 12242 1223
rect 12254 1214 12306 1223
rect 12318 1214 12370 1223
rect 12382 1214 12434 1223
rect 12446 1257 12498 1266
rect 12446 1223 12447 1257
rect 12447 1223 12481 1257
rect 12481 1223 12498 1257
rect 12446 1214 12498 1223
rect 8334 894 8386 946
rect 8542 937 8594 946
rect 8542 903 8559 937
rect 8559 903 8593 937
rect 8593 903 8594 937
rect 8542 894 8594 903
rect 8606 937 8658 946
rect 8670 937 8722 946
rect 8734 937 8786 946
rect 8798 937 8850 946
rect 8862 937 8914 946
rect 8926 937 8978 946
rect 8606 903 8631 937
rect 8631 903 8658 937
rect 8670 903 8703 937
rect 8703 903 8722 937
rect 8734 903 8737 937
rect 8737 903 8775 937
rect 8775 903 8786 937
rect 8798 903 8809 937
rect 8809 903 8847 937
rect 8847 903 8850 937
rect 8862 903 8881 937
rect 8881 903 8914 937
rect 8926 903 8953 937
rect 8953 903 8978 937
rect 8606 894 8658 903
rect 8670 894 8722 903
rect 8734 894 8786 903
rect 8798 894 8850 903
rect 8862 894 8914 903
rect 8926 894 8978 903
rect 8990 937 9042 946
rect 8990 903 8991 937
rect 8991 903 9025 937
rect 9025 903 9042 937
rect 8990 894 9042 903
rect 9054 937 9106 946
rect 9054 903 9063 937
rect 9063 903 9097 937
rect 9097 903 9106 937
rect 9054 894 9106 903
rect 9118 937 9170 946
rect 9118 903 9135 937
rect 9135 903 9169 937
rect 9169 903 9170 937
rect 9118 894 9170 903
rect 9182 937 9234 946
rect 9246 937 9298 946
rect 9310 937 9362 946
rect 9374 937 9426 946
rect 9438 937 9490 946
rect 9502 937 9554 946
rect 9182 903 9207 937
rect 9207 903 9234 937
rect 9246 903 9279 937
rect 9279 903 9298 937
rect 9310 903 9313 937
rect 9313 903 9351 937
rect 9351 903 9362 937
rect 9374 903 9385 937
rect 9385 903 9423 937
rect 9423 903 9426 937
rect 9438 903 9457 937
rect 9457 903 9490 937
rect 9502 903 9529 937
rect 9529 903 9554 937
rect 9182 894 9234 903
rect 9246 894 9298 903
rect 9310 894 9362 903
rect 9374 894 9426 903
rect 9438 894 9490 903
rect 9502 894 9554 903
rect 9566 937 9618 946
rect 9566 903 9567 937
rect 9567 903 9601 937
rect 9601 903 9618 937
rect 9566 894 9618 903
rect 9630 937 9682 946
rect 9630 903 9639 937
rect 9639 903 9673 937
rect 9673 903 9682 937
rect 9630 894 9682 903
rect 9694 937 9746 946
rect 9694 903 9711 937
rect 9711 903 9745 937
rect 9745 903 9746 937
rect 9694 894 9746 903
rect 9758 937 9810 946
rect 9822 937 9874 946
rect 9886 937 9938 946
rect 9950 937 10002 946
rect 10014 937 10066 946
rect 10078 937 10130 946
rect 9758 903 9783 937
rect 9783 903 9810 937
rect 9822 903 9855 937
rect 9855 903 9874 937
rect 9886 903 9889 937
rect 9889 903 9927 937
rect 9927 903 9938 937
rect 9950 903 9961 937
rect 9961 903 9999 937
rect 9999 903 10002 937
rect 10014 903 10033 937
rect 10033 903 10066 937
rect 10078 903 10105 937
rect 10105 903 10130 937
rect 9758 894 9810 903
rect 9822 894 9874 903
rect 9886 894 9938 903
rect 9950 894 10002 903
rect 10014 894 10066 903
rect 10078 894 10130 903
rect 10142 937 10194 946
rect 10142 903 10143 937
rect 10143 903 10177 937
rect 10177 903 10194 937
rect 10142 894 10194 903
rect 10206 937 10258 946
rect 10206 903 10215 937
rect 10215 903 10249 937
rect 10249 903 10258 937
rect 10206 894 10258 903
rect 10270 937 10322 946
rect 10270 903 10287 937
rect 10287 903 10321 937
rect 10321 903 10322 937
rect 10270 894 10322 903
rect 10334 937 10386 946
rect 10398 937 10450 946
rect 10462 937 10514 946
rect 10526 937 10578 946
rect 10590 937 10642 946
rect 10654 937 10706 946
rect 10334 903 10359 937
rect 10359 903 10386 937
rect 10398 903 10431 937
rect 10431 903 10450 937
rect 10462 903 10465 937
rect 10465 903 10503 937
rect 10503 903 10514 937
rect 10526 903 10537 937
rect 10537 903 10575 937
rect 10575 903 10578 937
rect 10590 903 10609 937
rect 10609 903 10642 937
rect 10654 903 10681 937
rect 10681 903 10706 937
rect 10334 894 10386 903
rect 10398 894 10450 903
rect 10462 894 10514 903
rect 10526 894 10578 903
rect 10590 894 10642 903
rect 10654 894 10706 903
rect 10718 937 10770 946
rect 10718 903 10719 937
rect 10719 903 10753 937
rect 10753 903 10770 937
rect 10718 894 10770 903
rect 10782 937 10834 946
rect 10782 903 10791 937
rect 10791 903 10825 937
rect 10825 903 10834 937
rect 10782 894 10834 903
rect 10846 937 10898 946
rect 10846 903 10863 937
rect 10863 903 10897 937
rect 10897 903 10898 937
rect 10846 894 10898 903
rect 10910 937 10962 946
rect 10974 937 11026 946
rect 11038 937 11090 946
rect 11102 937 11154 946
rect 11166 937 11218 946
rect 11230 937 11282 946
rect 10910 903 10935 937
rect 10935 903 10962 937
rect 10974 903 11007 937
rect 11007 903 11026 937
rect 11038 903 11041 937
rect 11041 903 11079 937
rect 11079 903 11090 937
rect 11102 903 11113 937
rect 11113 903 11151 937
rect 11151 903 11154 937
rect 11166 903 11185 937
rect 11185 903 11218 937
rect 11230 903 11257 937
rect 11257 903 11282 937
rect 10910 894 10962 903
rect 10974 894 11026 903
rect 11038 894 11090 903
rect 11102 894 11154 903
rect 11166 894 11218 903
rect 11230 894 11282 903
rect 11294 937 11346 946
rect 11294 903 11295 937
rect 11295 903 11329 937
rect 11329 903 11346 937
rect 11294 894 11346 903
rect 11358 937 11410 946
rect 11358 903 11367 937
rect 11367 903 11401 937
rect 11401 903 11410 937
rect 11358 894 11410 903
rect 11422 937 11474 946
rect 11422 903 11439 937
rect 11439 903 11473 937
rect 11473 903 11474 937
rect 11422 894 11474 903
rect 11486 937 11538 946
rect 11550 937 11602 946
rect 11614 937 11666 946
rect 11678 937 11730 946
rect 11742 937 11794 946
rect 11806 937 11858 946
rect 11486 903 11511 937
rect 11511 903 11538 937
rect 11550 903 11583 937
rect 11583 903 11602 937
rect 11614 903 11617 937
rect 11617 903 11655 937
rect 11655 903 11666 937
rect 11678 903 11689 937
rect 11689 903 11727 937
rect 11727 903 11730 937
rect 11742 903 11761 937
rect 11761 903 11794 937
rect 11806 903 11833 937
rect 11833 903 11858 937
rect 11486 894 11538 903
rect 11550 894 11602 903
rect 11614 894 11666 903
rect 11678 894 11730 903
rect 11742 894 11794 903
rect 11806 894 11858 903
rect 11870 937 11922 946
rect 11870 903 11871 937
rect 11871 903 11905 937
rect 11905 903 11922 937
rect 11870 894 11922 903
rect 11934 937 11986 946
rect 11934 903 11943 937
rect 11943 903 11977 937
rect 11977 903 11986 937
rect 11934 894 11986 903
rect 11998 937 12050 946
rect 11998 903 12015 937
rect 12015 903 12049 937
rect 12049 903 12050 937
rect 11998 894 12050 903
rect 12062 937 12114 946
rect 12126 937 12178 946
rect 12190 937 12242 946
rect 12254 937 12306 946
rect 12318 937 12370 946
rect 12382 937 12434 946
rect 12062 903 12087 937
rect 12087 903 12114 937
rect 12126 903 12159 937
rect 12159 903 12178 937
rect 12190 903 12193 937
rect 12193 903 12231 937
rect 12231 903 12242 937
rect 12254 903 12265 937
rect 12265 903 12303 937
rect 12303 903 12306 937
rect 12318 903 12337 937
rect 12337 903 12370 937
rect 12382 903 12409 937
rect 12409 903 12434 937
rect 12062 894 12114 903
rect 12126 894 12178 903
rect 12190 894 12242 903
rect 12254 894 12306 903
rect 12318 894 12370 903
rect 12382 894 12434 903
rect 12446 937 12498 946
rect 12446 903 12447 937
rect 12447 903 12481 937
rect 12481 903 12498 937
rect 12446 894 12498 903
rect 8542 137 8594 146
rect 8542 103 8559 137
rect 8559 103 8593 137
rect 8593 103 8594 137
rect 8542 94 8594 103
rect 8606 137 8658 146
rect 8670 137 8722 146
rect 8734 137 8786 146
rect 8798 137 8850 146
rect 8862 137 8914 146
rect 8926 137 8978 146
rect 8606 103 8631 137
rect 8631 103 8658 137
rect 8670 103 8703 137
rect 8703 103 8722 137
rect 8734 103 8737 137
rect 8737 103 8775 137
rect 8775 103 8786 137
rect 8798 103 8809 137
rect 8809 103 8847 137
rect 8847 103 8850 137
rect 8862 103 8881 137
rect 8881 103 8914 137
rect 8926 103 8953 137
rect 8953 103 8978 137
rect 8606 94 8658 103
rect 8670 94 8722 103
rect 8734 94 8786 103
rect 8798 94 8850 103
rect 8862 94 8914 103
rect 8926 94 8978 103
rect 8990 137 9042 146
rect 8990 103 8991 137
rect 8991 103 9025 137
rect 9025 103 9042 137
rect 8990 94 9042 103
rect 9054 137 9106 146
rect 9054 103 9063 137
rect 9063 103 9097 137
rect 9097 103 9106 137
rect 9054 94 9106 103
rect 9118 137 9170 146
rect 9118 103 9135 137
rect 9135 103 9169 137
rect 9169 103 9170 137
rect 9118 94 9170 103
rect 9182 137 9234 146
rect 9246 137 9298 146
rect 9310 137 9362 146
rect 9374 137 9426 146
rect 9438 137 9490 146
rect 9502 137 9554 146
rect 9182 103 9207 137
rect 9207 103 9234 137
rect 9246 103 9279 137
rect 9279 103 9298 137
rect 9310 103 9313 137
rect 9313 103 9351 137
rect 9351 103 9362 137
rect 9374 103 9385 137
rect 9385 103 9423 137
rect 9423 103 9426 137
rect 9438 103 9457 137
rect 9457 103 9490 137
rect 9502 103 9529 137
rect 9529 103 9554 137
rect 9182 94 9234 103
rect 9246 94 9298 103
rect 9310 94 9362 103
rect 9374 94 9426 103
rect 9438 94 9490 103
rect 9502 94 9554 103
rect 9566 137 9618 146
rect 9566 103 9567 137
rect 9567 103 9601 137
rect 9601 103 9618 137
rect 9566 94 9618 103
rect 9630 137 9682 146
rect 9630 103 9639 137
rect 9639 103 9673 137
rect 9673 103 9682 137
rect 9630 94 9682 103
rect 9694 137 9746 146
rect 9694 103 9711 137
rect 9711 103 9745 137
rect 9745 103 9746 137
rect 9694 94 9746 103
rect 9758 137 9810 146
rect 9822 137 9874 146
rect 9886 137 9938 146
rect 9950 137 10002 146
rect 10014 137 10066 146
rect 10078 137 10130 146
rect 9758 103 9783 137
rect 9783 103 9810 137
rect 9822 103 9855 137
rect 9855 103 9874 137
rect 9886 103 9889 137
rect 9889 103 9927 137
rect 9927 103 9938 137
rect 9950 103 9961 137
rect 9961 103 9999 137
rect 9999 103 10002 137
rect 10014 103 10033 137
rect 10033 103 10066 137
rect 10078 103 10105 137
rect 10105 103 10130 137
rect 9758 94 9810 103
rect 9822 94 9874 103
rect 9886 94 9938 103
rect 9950 94 10002 103
rect 10014 94 10066 103
rect 10078 94 10130 103
rect 10142 137 10194 146
rect 10142 103 10143 137
rect 10143 103 10177 137
rect 10177 103 10194 137
rect 10142 94 10194 103
rect 10206 137 10258 146
rect 10206 103 10215 137
rect 10215 103 10249 137
rect 10249 103 10258 137
rect 10206 94 10258 103
rect 10270 137 10322 146
rect 10270 103 10287 137
rect 10287 103 10321 137
rect 10321 103 10322 137
rect 10270 94 10322 103
rect 10334 137 10386 146
rect 10398 137 10450 146
rect 10462 137 10514 146
rect 10526 137 10578 146
rect 10590 137 10642 146
rect 10654 137 10706 146
rect 10334 103 10359 137
rect 10359 103 10386 137
rect 10398 103 10431 137
rect 10431 103 10450 137
rect 10462 103 10465 137
rect 10465 103 10503 137
rect 10503 103 10514 137
rect 10526 103 10537 137
rect 10537 103 10575 137
rect 10575 103 10578 137
rect 10590 103 10609 137
rect 10609 103 10642 137
rect 10654 103 10681 137
rect 10681 103 10706 137
rect 10334 94 10386 103
rect 10398 94 10450 103
rect 10462 94 10514 103
rect 10526 94 10578 103
rect 10590 94 10642 103
rect 10654 94 10706 103
rect 10718 137 10770 146
rect 10718 103 10719 137
rect 10719 103 10753 137
rect 10753 103 10770 137
rect 10718 94 10770 103
rect 10782 137 10834 146
rect 10782 103 10791 137
rect 10791 103 10825 137
rect 10825 103 10834 137
rect 10782 94 10834 103
rect 10846 137 10898 146
rect 10846 103 10863 137
rect 10863 103 10897 137
rect 10897 103 10898 137
rect 10846 94 10898 103
rect 10910 137 10962 146
rect 10974 137 11026 146
rect 11038 137 11090 146
rect 11102 137 11154 146
rect 11166 137 11218 146
rect 11230 137 11282 146
rect 10910 103 10935 137
rect 10935 103 10962 137
rect 10974 103 11007 137
rect 11007 103 11026 137
rect 11038 103 11041 137
rect 11041 103 11079 137
rect 11079 103 11090 137
rect 11102 103 11113 137
rect 11113 103 11151 137
rect 11151 103 11154 137
rect 11166 103 11185 137
rect 11185 103 11218 137
rect 11230 103 11257 137
rect 11257 103 11282 137
rect 10910 94 10962 103
rect 10974 94 11026 103
rect 11038 94 11090 103
rect 11102 94 11154 103
rect 11166 94 11218 103
rect 11230 94 11282 103
rect 11294 137 11346 146
rect 11294 103 11295 137
rect 11295 103 11329 137
rect 11329 103 11346 137
rect 11294 94 11346 103
rect 11358 137 11410 146
rect 11358 103 11367 137
rect 11367 103 11401 137
rect 11401 103 11410 137
rect 11358 94 11410 103
rect 11422 137 11474 146
rect 11422 103 11439 137
rect 11439 103 11473 137
rect 11473 103 11474 137
rect 11422 94 11474 103
rect 11486 137 11538 146
rect 11550 137 11602 146
rect 11614 137 11666 146
rect 11678 137 11730 146
rect 11742 137 11794 146
rect 11806 137 11858 146
rect 11486 103 11511 137
rect 11511 103 11538 137
rect 11550 103 11583 137
rect 11583 103 11602 137
rect 11614 103 11617 137
rect 11617 103 11655 137
rect 11655 103 11666 137
rect 11678 103 11689 137
rect 11689 103 11727 137
rect 11727 103 11730 137
rect 11742 103 11761 137
rect 11761 103 11794 137
rect 11806 103 11833 137
rect 11833 103 11858 137
rect 11486 94 11538 103
rect 11550 94 11602 103
rect 11614 94 11666 103
rect 11678 94 11730 103
rect 11742 94 11794 103
rect 11806 94 11858 103
rect 11870 137 11922 146
rect 11870 103 11871 137
rect 11871 103 11905 137
rect 11905 103 11922 137
rect 11870 94 11922 103
rect 11934 137 11986 146
rect 11934 103 11943 137
rect 11943 103 11977 137
rect 11977 103 11986 137
rect 11934 94 11986 103
rect 11998 137 12050 146
rect 11998 103 12015 137
rect 12015 103 12049 137
rect 12049 103 12050 137
rect 11998 94 12050 103
rect 12062 137 12114 146
rect 12126 137 12178 146
rect 12190 137 12242 146
rect 12254 137 12306 146
rect 12318 137 12370 146
rect 12382 137 12434 146
rect 12062 103 12087 137
rect 12087 103 12114 137
rect 12126 103 12159 137
rect 12159 103 12178 137
rect 12190 103 12193 137
rect 12193 103 12231 137
rect 12231 103 12242 137
rect 12254 103 12265 137
rect 12265 103 12303 137
rect 12303 103 12306 137
rect 12318 103 12337 137
rect 12337 103 12370 137
rect 12382 103 12409 137
rect 12409 103 12434 137
rect 12062 94 12114 103
rect 12126 94 12178 103
rect 12190 94 12242 103
rect 12254 94 12306 103
rect 12318 94 12370 103
rect 12382 94 12434 103
rect 12446 137 12498 146
rect 12446 103 12447 137
rect 12447 103 12481 137
rect 12481 103 12498 137
rect 12446 94 12498 103
rect 12654 94 12706 146
rect 8542 -183 8594 -174
rect 8542 -217 8559 -183
rect 8559 -217 8593 -183
rect 8593 -217 8594 -183
rect 8542 -226 8594 -217
rect 8606 -183 8658 -174
rect 8670 -183 8722 -174
rect 8734 -183 8786 -174
rect 8798 -183 8850 -174
rect 8862 -183 8914 -174
rect 8926 -183 8978 -174
rect 8606 -217 8631 -183
rect 8631 -217 8658 -183
rect 8670 -217 8703 -183
rect 8703 -217 8722 -183
rect 8734 -217 8737 -183
rect 8737 -217 8775 -183
rect 8775 -217 8786 -183
rect 8798 -217 8809 -183
rect 8809 -217 8847 -183
rect 8847 -217 8850 -183
rect 8862 -217 8881 -183
rect 8881 -217 8914 -183
rect 8926 -217 8953 -183
rect 8953 -217 8978 -183
rect 8606 -226 8658 -217
rect 8670 -226 8722 -217
rect 8734 -226 8786 -217
rect 8798 -226 8850 -217
rect 8862 -226 8914 -217
rect 8926 -226 8978 -217
rect 8990 -183 9042 -174
rect 8990 -217 8991 -183
rect 8991 -217 9025 -183
rect 9025 -217 9042 -183
rect 8990 -226 9042 -217
rect 9054 -183 9106 -174
rect 9054 -217 9063 -183
rect 9063 -217 9097 -183
rect 9097 -217 9106 -183
rect 9054 -226 9106 -217
rect 9118 -183 9170 -174
rect 9118 -217 9135 -183
rect 9135 -217 9169 -183
rect 9169 -217 9170 -183
rect 9118 -226 9170 -217
rect 9182 -183 9234 -174
rect 9246 -183 9298 -174
rect 9310 -183 9362 -174
rect 9374 -183 9426 -174
rect 9438 -183 9490 -174
rect 9502 -183 9554 -174
rect 9182 -217 9207 -183
rect 9207 -217 9234 -183
rect 9246 -217 9279 -183
rect 9279 -217 9298 -183
rect 9310 -217 9313 -183
rect 9313 -217 9351 -183
rect 9351 -217 9362 -183
rect 9374 -217 9385 -183
rect 9385 -217 9423 -183
rect 9423 -217 9426 -183
rect 9438 -217 9457 -183
rect 9457 -217 9490 -183
rect 9502 -217 9529 -183
rect 9529 -217 9554 -183
rect 9182 -226 9234 -217
rect 9246 -226 9298 -217
rect 9310 -226 9362 -217
rect 9374 -226 9426 -217
rect 9438 -226 9490 -217
rect 9502 -226 9554 -217
rect 9566 -183 9618 -174
rect 9566 -217 9567 -183
rect 9567 -217 9601 -183
rect 9601 -217 9618 -183
rect 9566 -226 9618 -217
rect 9630 -183 9682 -174
rect 9630 -217 9639 -183
rect 9639 -217 9673 -183
rect 9673 -217 9682 -183
rect 9630 -226 9682 -217
rect 9694 -183 9746 -174
rect 9694 -217 9711 -183
rect 9711 -217 9745 -183
rect 9745 -217 9746 -183
rect 9694 -226 9746 -217
rect 9758 -183 9810 -174
rect 9822 -183 9874 -174
rect 9886 -183 9938 -174
rect 9950 -183 10002 -174
rect 10014 -183 10066 -174
rect 10078 -183 10130 -174
rect 9758 -217 9783 -183
rect 9783 -217 9810 -183
rect 9822 -217 9855 -183
rect 9855 -217 9874 -183
rect 9886 -217 9889 -183
rect 9889 -217 9927 -183
rect 9927 -217 9938 -183
rect 9950 -217 9961 -183
rect 9961 -217 9999 -183
rect 9999 -217 10002 -183
rect 10014 -217 10033 -183
rect 10033 -217 10066 -183
rect 10078 -217 10105 -183
rect 10105 -217 10130 -183
rect 9758 -226 9810 -217
rect 9822 -226 9874 -217
rect 9886 -226 9938 -217
rect 9950 -226 10002 -217
rect 10014 -226 10066 -217
rect 10078 -226 10130 -217
rect 10142 -183 10194 -174
rect 10142 -217 10143 -183
rect 10143 -217 10177 -183
rect 10177 -217 10194 -183
rect 10142 -226 10194 -217
rect 10206 -183 10258 -174
rect 10206 -217 10215 -183
rect 10215 -217 10249 -183
rect 10249 -217 10258 -183
rect 10206 -226 10258 -217
rect 10270 -183 10322 -174
rect 10270 -217 10287 -183
rect 10287 -217 10321 -183
rect 10321 -217 10322 -183
rect 10270 -226 10322 -217
rect 10334 -183 10386 -174
rect 10398 -183 10450 -174
rect 10462 -183 10514 -174
rect 10526 -183 10578 -174
rect 10590 -183 10642 -174
rect 10654 -183 10706 -174
rect 10334 -217 10359 -183
rect 10359 -217 10386 -183
rect 10398 -217 10431 -183
rect 10431 -217 10450 -183
rect 10462 -217 10465 -183
rect 10465 -217 10503 -183
rect 10503 -217 10514 -183
rect 10526 -217 10537 -183
rect 10537 -217 10575 -183
rect 10575 -217 10578 -183
rect 10590 -217 10609 -183
rect 10609 -217 10642 -183
rect 10654 -217 10681 -183
rect 10681 -217 10706 -183
rect 10334 -226 10386 -217
rect 10398 -226 10450 -217
rect 10462 -226 10514 -217
rect 10526 -226 10578 -217
rect 10590 -226 10642 -217
rect 10654 -226 10706 -217
rect 10718 -183 10770 -174
rect 10718 -217 10719 -183
rect 10719 -217 10753 -183
rect 10753 -217 10770 -183
rect 10718 -226 10770 -217
rect 10782 -183 10834 -174
rect 10782 -217 10791 -183
rect 10791 -217 10825 -183
rect 10825 -217 10834 -183
rect 10782 -226 10834 -217
rect 10846 -183 10898 -174
rect 10846 -217 10863 -183
rect 10863 -217 10897 -183
rect 10897 -217 10898 -183
rect 10846 -226 10898 -217
rect 10910 -183 10962 -174
rect 10974 -183 11026 -174
rect 11038 -183 11090 -174
rect 11102 -183 11154 -174
rect 11166 -183 11218 -174
rect 11230 -183 11282 -174
rect 10910 -217 10935 -183
rect 10935 -217 10962 -183
rect 10974 -217 11007 -183
rect 11007 -217 11026 -183
rect 11038 -217 11041 -183
rect 11041 -217 11079 -183
rect 11079 -217 11090 -183
rect 11102 -217 11113 -183
rect 11113 -217 11151 -183
rect 11151 -217 11154 -183
rect 11166 -217 11185 -183
rect 11185 -217 11218 -183
rect 11230 -217 11257 -183
rect 11257 -217 11282 -183
rect 10910 -226 10962 -217
rect 10974 -226 11026 -217
rect 11038 -226 11090 -217
rect 11102 -226 11154 -217
rect 11166 -226 11218 -217
rect 11230 -226 11282 -217
rect 11294 -183 11346 -174
rect 11294 -217 11295 -183
rect 11295 -217 11329 -183
rect 11329 -217 11346 -183
rect 11294 -226 11346 -217
rect 11358 -183 11410 -174
rect 11358 -217 11367 -183
rect 11367 -217 11401 -183
rect 11401 -217 11410 -183
rect 11358 -226 11410 -217
rect 11422 -183 11474 -174
rect 11422 -217 11439 -183
rect 11439 -217 11473 -183
rect 11473 -217 11474 -183
rect 11422 -226 11474 -217
rect 11486 -183 11538 -174
rect 11550 -183 11602 -174
rect 11614 -183 11666 -174
rect 11678 -183 11730 -174
rect 11742 -183 11794 -174
rect 11806 -183 11858 -174
rect 11486 -217 11511 -183
rect 11511 -217 11538 -183
rect 11550 -217 11583 -183
rect 11583 -217 11602 -183
rect 11614 -217 11617 -183
rect 11617 -217 11655 -183
rect 11655 -217 11666 -183
rect 11678 -217 11689 -183
rect 11689 -217 11727 -183
rect 11727 -217 11730 -183
rect 11742 -217 11761 -183
rect 11761 -217 11794 -183
rect 11806 -217 11833 -183
rect 11833 -217 11858 -183
rect 11486 -226 11538 -217
rect 11550 -226 11602 -217
rect 11614 -226 11666 -217
rect 11678 -226 11730 -217
rect 11742 -226 11794 -217
rect 11806 -226 11858 -217
rect 11870 -183 11922 -174
rect 11870 -217 11871 -183
rect 11871 -217 11905 -183
rect 11905 -217 11922 -183
rect 11870 -226 11922 -217
rect 11934 -183 11986 -174
rect 11934 -217 11943 -183
rect 11943 -217 11977 -183
rect 11977 -217 11986 -183
rect 11934 -226 11986 -217
rect 11998 -183 12050 -174
rect 11998 -217 12015 -183
rect 12015 -217 12049 -183
rect 12049 -217 12050 -183
rect 11998 -226 12050 -217
rect 12062 -183 12114 -174
rect 12126 -183 12178 -174
rect 12190 -183 12242 -174
rect 12254 -183 12306 -174
rect 12318 -183 12370 -174
rect 12382 -183 12434 -174
rect 12062 -217 12087 -183
rect 12087 -217 12114 -183
rect 12126 -217 12159 -183
rect 12159 -217 12178 -183
rect 12190 -217 12193 -183
rect 12193 -217 12231 -183
rect 12231 -217 12242 -183
rect 12254 -217 12265 -183
rect 12265 -217 12303 -183
rect 12303 -217 12306 -183
rect 12318 -217 12337 -183
rect 12337 -217 12370 -183
rect 12382 -217 12409 -183
rect 12409 -217 12434 -183
rect 12062 -226 12114 -217
rect 12126 -226 12178 -217
rect 12190 -226 12242 -217
rect 12254 -226 12306 -217
rect 12318 -226 12370 -217
rect 12382 -226 12434 -217
rect 12446 -183 12498 -174
rect 12446 -217 12447 -183
rect 12447 -217 12481 -183
rect 12481 -217 12498 -183
rect 12446 -226 12498 -217
rect -306 -503 -254 -494
rect -306 -537 -297 -503
rect -297 -537 -263 -503
rect -263 -537 -254 -503
rect -306 -546 -254 -537
rect 12814 -503 12866 -494
rect 12814 -537 12823 -503
rect 12823 -537 12857 -503
rect 12857 -537 12866 -503
rect 12814 -546 12866 -537
<< metal2 >>
rect 4640 4308 7920 4320
rect 4640 4252 4652 4308
rect 4708 4252 4972 4308
rect 5028 4252 5292 4308
rect 5348 4252 5612 4308
rect 5668 4252 5932 4308
rect 5988 4252 6252 4308
rect 6308 4252 6572 4308
rect 6628 4252 6892 4308
rect 6948 4252 7212 4308
rect 7268 4252 7532 4308
rect 7588 4252 7852 4308
rect 7908 4252 7920 4308
rect 4640 4240 7920 4252
rect -480 4148 13040 4160
rect -480 4146 6412 4148
rect -480 4094 -306 4146
rect -254 4094 6412 4146
rect -480 4092 6412 4094
rect 6468 4146 13040 4148
rect 6468 4094 12814 4146
rect 12866 4094 13040 4146
rect 6468 4092 13040 4094
rect -480 4080 13040 4092
rect 4640 3988 7920 4000
rect 4640 3932 4652 3988
rect 4708 3932 4972 3988
rect 5028 3932 5292 3988
rect 5348 3932 5612 3988
rect 5668 3932 5932 3988
rect 5988 3932 6252 3988
rect 6308 3932 6572 3988
rect 6628 3932 6892 3988
rect 6948 3932 7212 3988
rect 7268 3932 7532 3988
rect 7588 3932 7852 3988
rect 7908 3932 7920 3988
rect 4640 3920 7920 3932
rect -480 3828 13040 3840
rect -480 3826 6092 3828
rect -480 3774 62 3826
rect 114 3774 126 3826
rect 178 3774 190 3826
rect 242 3774 254 3826
rect 306 3774 318 3826
rect 370 3774 382 3826
rect 434 3774 446 3826
rect 498 3774 510 3826
rect 562 3774 574 3826
rect 626 3774 638 3826
rect 690 3774 702 3826
rect 754 3774 766 3826
rect 818 3774 830 3826
rect 882 3774 894 3826
rect 946 3774 958 3826
rect 1010 3774 1022 3826
rect 1074 3774 1086 3826
rect 1138 3774 1150 3826
rect 1202 3774 1214 3826
rect 1266 3774 1278 3826
rect 1330 3774 1342 3826
rect 1394 3774 1406 3826
rect 1458 3774 1470 3826
rect 1522 3774 1534 3826
rect 1586 3774 1598 3826
rect 1650 3774 1662 3826
rect 1714 3774 1726 3826
rect 1778 3774 1790 3826
rect 1842 3774 1854 3826
rect 1906 3774 1918 3826
rect 1970 3774 1982 3826
rect 2034 3774 2046 3826
rect 2098 3774 2110 3826
rect 2162 3774 2174 3826
rect 2226 3774 2238 3826
rect 2290 3774 2302 3826
rect 2354 3774 2366 3826
rect 2418 3774 2430 3826
rect 2482 3774 2494 3826
rect 2546 3774 2558 3826
rect 2610 3774 2622 3826
rect 2674 3774 2686 3826
rect 2738 3774 2750 3826
rect 2802 3774 2814 3826
rect 2866 3774 2878 3826
rect 2930 3774 2942 3826
rect 2994 3774 3006 3826
rect 3058 3774 3070 3826
rect 3122 3774 3134 3826
rect 3186 3774 3198 3826
rect 3250 3774 3262 3826
rect 3314 3774 3326 3826
rect 3378 3774 3390 3826
rect 3442 3774 3454 3826
rect 3506 3774 3518 3826
rect 3570 3774 3582 3826
rect 3634 3774 3646 3826
rect 3698 3774 3710 3826
rect 3762 3774 3774 3826
rect 3826 3774 3838 3826
rect 3890 3774 3902 3826
rect 3954 3774 3966 3826
rect 4018 3774 6092 3826
rect -480 3772 6092 3774
rect 6148 3826 13040 3828
rect 6148 3774 8542 3826
rect 8594 3774 8606 3826
rect 8658 3774 8670 3826
rect 8722 3774 8734 3826
rect 8786 3774 8798 3826
rect 8850 3774 8862 3826
rect 8914 3774 8926 3826
rect 8978 3774 8990 3826
rect 9042 3774 9054 3826
rect 9106 3774 9118 3826
rect 9170 3774 9182 3826
rect 9234 3774 9246 3826
rect 9298 3774 9310 3826
rect 9362 3774 9374 3826
rect 9426 3774 9438 3826
rect 9490 3774 9502 3826
rect 9554 3774 9566 3826
rect 9618 3774 9630 3826
rect 9682 3774 9694 3826
rect 9746 3774 9758 3826
rect 9810 3774 9822 3826
rect 9874 3774 9886 3826
rect 9938 3774 9950 3826
rect 10002 3774 10014 3826
rect 10066 3774 10078 3826
rect 10130 3774 10142 3826
rect 10194 3774 10206 3826
rect 10258 3774 10270 3826
rect 10322 3774 10334 3826
rect 10386 3774 10398 3826
rect 10450 3774 10462 3826
rect 10514 3774 10526 3826
rect 10578 3774 10590 3826
rect 10642 3774 10654 3826
rect 10706 3774 10718 3826
rect 10770 3774 10782 3826
rect 10834 3774 10846 3826
rect 10898 3774 10910 3826
rect 10962 3774 10974 3826
rect 11026 3774 11038 3826
rect 11090 3774 11102 3826
rect 11154 3774 11166 3826
rect 11218 3774 11230 3826
rect 11282 3774 11294 3826
rect 11346 3774 11358 3826
rect 11410 3774 11422 3826
rect 11474 3774 11486 3826
rect 11538 3774 11550 3826
rect 11602 3774 11614 3826
rect 11666 3774 11678 3826
rect 11730 3774 11742 3826
rect 11794 3774 11806 3826
rect 11858 3774 11870 3826
rect 11922 3774 11934 3826
rect 11986 3774 11998 3826
rect 12050 3774 12062 3826
rect 12114 3774 12126 3826
rect 12178 3774 12190 3826
rect 12242 3774 12254 3826
rect 12306 3774 12318 3826
rect 12370 3774 12382 3826
rect 12434 3774 12446 3826
rect 12498 3774 13040 3826
rect 6148 3772 13040 3774
rect -480 3760 13040 3772
rect 4640 3668 7920 3680
rect 4640 3612 4652 3668
rect 4708 3612 4972 3668
rect 5028 3612 5292 3668
rect 5348 3612 5612 3668
rect 5668 3612 5932 3668
rect 5988 3612 6252 3668
rect 6308 3612 6572 3668
rect 6628 3612 6892 3668
rect 6948 3612 7212 3668
rect 7268 3612 7532 3668
rect 7588 3612 7852 3668
rect 7908 3612 7920 3668
rect 4640 3600 7920 3612
rect -480 3508 5840 3520
rect -480 3506 5452 3508
rect -480 3454 -146 3506
rect -94 3454 62 3506
rect 114 3454 126 3506
rect 178 3454 190 3506
rect 242 3454 254 3506
rect 306 3454 318 3506
rect 370 3454 382 3506
rect 434 3454 446 3506
rect 498 3454 510 3506
rect 562 3454 574 3506
rect 626 3454 638 3506
rect 690 3454 702 3506
rect 754 3454 766 3506
rect 818 3454 830 3506
rect 882 3454 894 3506
rect 946 3454 958 3506
rect 1010 3454 1022 3506
rect 1074 3454 1086 3506
rect 1138 3454 1150 3506
rect 1202 3454 1214 3506
rect 1266 3454 1278 3506
rect 1330 3454 1342 3506
rect 1394 3454 1406 3506
rect 1458 3454 1470 3506
rect 1522 3454 1534 3506
rect 1586 3454 1598 3506
rect 1650 3454 1662 3506
rect 1714 3454 1726 3506
rect 1778 3454 1790 3506
rect 1842 3454 1854 3506
rect 1906 3454 1918 3506
rect 1970 3454 1982 3506
rect 2034 3454 2046 3506
rect 2098 3454 2110 3506
rect 2162 3454 2174 3506
rect 2226 3454 2238 3506
rect 2290 3454 2302 3506
rect 2354 3454 2366 3506
rect 2418 3454 2430 3506
rect 2482 3454 2494 3506
rect 2546 3454 2558 3506
rect 2610 3454 2622 3506
rect 2674 3454 2686 3506
rect 2738 3454 2750 3506
rect 2802 3454 2814 3506
rect 2866 3454 2878 3506
rect 2930 3454 2942 3506
rect 2994 3454 3006 3506
rect 3058 3454 3070 3506
rect 3122 3454 3134 3506
rect 3186 3454 3198 3506
rect 3250 3454 3262 3506
rect 3314 3454 3326 3506
rect 3378 3454 3390 3506
rect 3442 3454 3454 3506
rect 3506 3454 3518 3506
rect 3570 3454 3582 3506
rect 3634 3454 3646 3506
rect 3698 3454 3710 3506
rect 3762 3454 3774 3506
rect 3826 3454 3838 3506
rect 3890 3454 3902 3506
rect 3954 3454 3966 3506
rect 4018 3454 5452 3506
rect -480 3452 5452 3454
rect 5508 3452 5840 3508
rect -480 3440 5840 3452
rect 5920 3508 6640 3520
rect 5920 3452 5932 3508
rect 5988 3452 6252 3508
rect 6308 3452 6572 3508
rect 6628 3452 6640 3508
rect 5920 3440 6640 3452
rect 6720 3508 13040 3520
rect 6720 3452 7692 3508
rect 7748 3506 13040 3508
rect 7748 3454 8542 3506
rect 8594 3454 8606 3506
rect 8658 3454 8670 3506
rect 8722 3454 8734 3506
rect 8786 3454 8798 3506
rect 8850 3454 8862 3506
rect 8914 3454 8926 3506
rect 8978 3454 8990 3506
rect 9042 3454 9054 3506
rect 9106 3454 9118 3506
rect 9170 3454 9182 3506
rect 9234 3454 9246 3506
rect 9298 3454 9310 3506
rect 9362 3454 9374 3506
rect 9426 3454 9438 3506
rect 9490 3454 9502 3506
rect 9554 3454 9566 3506
rect 9618 3454 9630 3506
rect 9682 3454 9694 3506
rect 9746 3454 9758 3506
rect 9810 3454 9822 3506
rect 9874 3454 9886 3506
rect 9938 3454 9950 3506
rect 10002 3454 10014 3506
rect 10066 3454 10078 3506
rect 10130 3454 10142 3506
rect 10194 3454 10206 3506
rect 10258 3454 10270 3506
rect 10322 3454 10334 3506
rect 10386 3454 10398 3506
rect 10450 3454 10462 3506
rect 10514 3454 10526 3506
rect 10578 3454 10590 3506
rect 10642 3454 10654 3506
rect 10706 3454 10718 3506
rect 10770 3454 10782 3506
rect 10834 3454 10846 3506
rect 10898 3454 10910 3506
rect 10962 3454 10974 3506
rect 11026 3454 11038 3506
rect 11090 3454 11102 3506
rect 11154 3454 11166 3506
rect 11218 3454 11230 3506
rect 11282 3454 11294 3506
rect 11346 3454 11358 3506
rect 11410 3454 11422 3506
rect 11474 3454 11486 3506
rect 11538 3454 11550 3506
rect 11602 3454 11614 3506
rect 11666 3454 11678 3506
rect 11730 3454 11742 3506
rect 11794 3454 11806 3506
rect 11858 3454 11870 3506
rect 11922 3454 11934 3506
rect 11986 3454 11998 3506
rect 12050 3454 12062 3506
rect 12114 3454 12126 3506
rect 12178 3454 12190 3506
rect 12242 3454 12254 3506
rect 12306 3454 12318 3506
rect 12370 3454 12382 3506
rect 12434 3454 12446 3506
rect 12498 3454 12654 3506
rect 12706 3454 13040 3506
rect 7748 3452 13040 3454
rect 6720 3440 13040 3452
rect 4640 3348 7920 3360
rect 4640 3292 4652 3348
rect 4708 3292 4972 3348
rect 5028 3292 5292 3348
rect 5348 3292 5612 3348
rect 5668 3292 5932 3348
rect 5988 3292 6252 3348
rect 6308 3292 6572 3348
rect 6628 3292 6892 3348
rect 6948 3292 7212 3348
rect 7268 3292 7532 3348
rect 7588 3292 7852 3348
rect 7908 3292 7920 3348
rect 4640 3280 7920 3292
rect 4640 3188 7920 3200
rect 4640 3132 4652 3188
rect 4708 3132 4972 3188
rect 5028 3132 5292 3188
rect 5348 3132 5612 3188
rect 5668 3132 5932 3188
rect 5988 3132 6252 3188
rect 6308 3132 6572 3188
rect 6628 3132 6892 3188
rect 6948 3132 7212 3188
rect 7268 3132 7532 3188
rect 7588 3132 7852 3188
rect 7908 3132 7920 3188
rect 4640 3120 7920 3132
rect 4640 3028 7920 3040
rect 4640 2972 5772 3028
rect 5828 2972 6732 3028
rect 6788 2972 7920 3028
rect 4640 2960 7920 2972
rect 4640 2868 7920 2880
rect 4640 2812 4652 2868
rect 4708 2812 4972 2868
rect 5028 2812 5292 2868
rect 5348 2812 5612 2868
rect 5668 2812 5932 2868
rect 5988 2812 6252 2868
rect 6308 2812 6572 2868
rect 6628 2812 6892 2868
rect 6948 2812 7212 2868
rect 7268 2812 7532 2868
rect 7588 2812 7852 2868
rect 7908 2812 7920 2868
rect 4640 2800 7920 2812
rect -480 2708 5840 2720
rect -480 2706 5772 2708
rect -480 2654 62 2706
rect 114 2654 126 2706
rect 178 2654 190 2706
rect 242 2654 254 2706
rect 306 2654 318 2706
rect 370 2654 382 2706
rect 434 2654 446 2706
rect 498 2654 510 2706
rect 562 2654 574 2706
rect 626 2654 638 2706
rect 690 2654 702 2706
rect 754 2654 766 2706
rect 818 2654 830 2706
rect 882 2654 894 2706
rect 946 2654 958 2706
rect 1010 2654 1022 2706
rect 1074 2654 1086 2706
rect 1138 2654 1150 2706
rect 1202 2654 1214 2706
rect 1266 2654 1278 2706
rect 1330 2654 1342 2706
rect 1394 2654 1406 2706
rect 1458 2654 1470 2706
rect 1522 2654 1534 2706
rect 1586 2654 1598 2706
rect 1650 2654 1662 2706
rect 1714 2654 1726 2706
rect 1778 2654 1790 2706
rect 1842 2654 1854 2706
rect 1906 2654 1918 2706
rect 1970 2654 1982 2706
rect 2034 2654 2046 2706
rect 2098 2654 2110 2706
rect 2162 2654 2174 2706
rect 2226 2654 2238 2706
rect 2290 2654 2302 2706
rect 2354 2654 2366 2706
rect 2418 2654 2430 2706
rect 2482 2654 2494 2706
rect 2546 2654 2558 2706
rect 2610 2654 2622 2706
rect 2674 2654 2686 2706
rect 2738 2654 2750 2706
rect 2802 2654 2814 2706
rect 2866 2654 2878 2706
rect 2930 2654 2942 2706
rect 2994 2654 3006 2706
rect 3058 2654 3070 2706
rect 3122 2654 3134 2706
rect 3186 2654 3198 2706
rect 3250 2654 3262 2706
rect 3314 2654 3326 2706
rect 3378 2654 3390 2706
rect 3442 2654 3454 2706
rect 3506 2654 3518 2706
rect 3570 2654 3582 2706
rect 3634 2654 3646 2706
rect 3698 2654 3710 2706
rect 3762 2654 3774 2706
rect 3826 2654 3838 2706
rect 3890 2654 3902 2706
rect 3954 2654 3966 2706
rect 4018 2654 4174 2706
rect 4226 2654 5772 2706
rect -480 2652 5772 2654
rect 5828 2652 5840 2708
rect -480 2640 5840 2652
rect 5920 2708 6640 2720
rect 5920 2652 5932 2708
rect 5988 2652 6252 2708
rect 6308 2652 6572 2708
rect 6628 2652 6640 2708
rect 5920 2640 6640 2652
rect 6720 2708 13040 2720
rect 6720 2652 7372 2708
rect 7428 2706 13040 2708
rect 7428 2654 8334 2706
rect 8386 2654 8542 2706
rect 8594 2654 8606 2706
rect 8658 2654 8670 2706
rect 8722 2654 8734 2706
rect 8786 2654 8798 2706
rect 8850 2654 8862 2706
rect 8914 2654 8926 2706
rect 8978 2654 8990 2706
rect 9042 2654 9054 2706
rect 9106 2654 9118 2706
rect 9170 2654 9182 2706
rect 9234 2654 9246 2706
rect 9298 2654 9310 2706
rect 9362 2654 9374 2706
rect 9426 2654 9438 2706
rect 9490 2654 9502 2706
rect 9554 2654 9566 2706
rect 9618 2654 9630 2706
rect 9682 2654 9694 2706
rect 9746 2654 9758 2706
rect 9810 2654 9822 2706
rect 9874 2654 9886 2706
rect 9938 2654 9950 2706
rect 10002 2654 10014 2706
rect 10066 2654 10078 2706
rect 10130 2654 10142 2706
rect 10194 2654 10206 2706
rect 10258 2654 10270 2706
rect 10322 2654 10334 2706
rect 10386 2654 10398 2706
rect 10450 2654 10462 2706
rect 10514 2654 10526 2706
rect 10578 2654 10590 2706
rect 10642 2654 10654 2706
rect 10706 2654 10718 2706
rect 10770 2654 10782 2706
rect 10834 2654 10846 2706
rect 10898 2654 10910 2706
rect 10962 2654 10974 2706
rect 11026 2654 11038 2706
rect 11090 2654 11102 2706
rect 11154 2654 11166 2706
rect 11218 2654 11230 2706
rect 11282 2654 11294 2706
rect 11346 2654 11358 2706
rect 11410 2654 11422 2706
rect 11474 2654 11486 2706
rect 11538 2654 11550 2706
rect 11602 2654 11614 2706
rect 11666 2654 11678 2706
rect 11730 2654 11742 2706
rect 11794 2654 11806 2706
rect 11858 2654 11870 2706
rect 11922 2654 11934 2706
rect 11986 2654 11998 2706
rect 12050 2654 12062 2706
rect 12114 2654 12126 2706
rect 12178 2654 12190 2706
rect 12242 2654 12254 2706
rect 12306 2654 12318 2706
rect 12370 2654 12382 2706
rect 12434 2654 12446 2706
rect 12498 2654 13040 2706
rect 7428 2652 13040 2654
rect 6720 2640 13040 2652
rect 4640 2548 7920 2560
rect 4640 2492 4652 2548
rect 4708 2492 4972 2548
rect 5028 2492 5292 2548
rect 5348 2492 5612 2548
rect 5668 2492 5932 2548
rect 5988 2492 6252 2548
rect 6308 2492 6572 2548
rect 6628 2492 6892 2548
rect 6948 2492 7212 2548
rect 7268 2492 7532 2548
rect 7588 2492 7852 2548
rect 7908 2492 7920 2548
rect 4640 2480 7920 2492
rect -480 2388 13040 2400
rect -480 2386 6092 2388
rect -480 2334 62 2386
rect 114 2334 126 2386
rect 178 2334 190 2386
rect 242 2334 254 2386
rect 306 2334 318 2386
rect 370 2334 382 2386
rect 434 2334 446 2386
rect 498 2334 510 2386
rect 562 2334 574 2386
rect 626 2334 638 2386
rect 690 2334 702 2386
rect 754 2334 766 2386
rect 818 2334 830 2386
rect 882 2334 894 2386
rect 946 2334 958 2386
rect 1010 2334 1022 2386
rect 1074 2334 1086 2386
rect 1138 2334 1150 2386
rect 1202 2334 1214 2386
rect 1266 2334 1278 2386
rect 1330 2334 1342 2386
rect 1394 2334 1406 2386
rect 1458 2334 1470 2386
rect 1522 2334 1534 2386
rect 1586 2334 1598 2386
rect 1650 2334 1662 2386
rect 1714 2334 1726 2386
rect 1778 2334 1790 2386
rect 1842 2334 1854 2386
rect 1906 2334 1918 2386
rect 1970 2334 1982 2386
rect 2034 2334 2046 2386
rect 2098 2334 2110 2386
rect 2162 2334 2174 2386
rect 2226 2334 2238 2386
rect 2290 2334 2302 2386
rect 2354 2334 2366 2386
rect 2418 2334 2430 2386
rect 2482 2334 2494 2386
rect 2546 2334 2558 2386
rect 2610 2334 2622 2386
rect 2674 2334 2686 2386
rect 2738 2334 2750 2386
rect 2802 2334 2814 2386
rect 2866 2334 2878 2386
rect 2930 2334 2942 2386
rect 2994 2334 3006 2386
rect 3058 2334 3070 2386
rect 3122 2334 3134 2386
rect 3186 2334 3198 2386
rect 3250 2334 3262 2386
rect 3314 2334 3326 2386
rect 3378 2334 3390 2386
rect 3442 2334 3454 2386
rect 3506 2334 3518 2386
rect 3570 2334 3582 2386
rect 3634 2334 3646 2386
rect 3698 2334 3710 2386
rect 3762 2334 3774 2386
rect 3826 2334 3838 2386
rect 3890 2334 3902 2386
rect 3954 2334 3966 2386
rect 4018 2334 6092 2386
rect -480 2332 6092 2334
rect 6148 2386 13040 2388
rect 6148 2334 8542 2386
rect 8594 2334 8606 2386
rect 8658 2334 8670 2386
rect 8722 2334 8734 2386
rect 8786 2334 8798 2386
rect 8850 2334 8862 2386
rect 8914 2334 8926 2386
rect 8978 2334 8990 2386
rect 9042 2334 9054 2386
rect 9106 2334 9118 2386
rect 9170 2334 9182 2386
rect 9234 2334 9246 2386
rect 9298 2334 9310 2386
rect 9362 2334 9374 2386
rect 9426 2334 9438 2386
rect 9490 2334 9502 2386
rect 9554 2334 9566 2386
rect 9618 2334 9630 2386
rect 9682 2334 9694 2386
rect 9746 2334 9758 2386
rect 9810 2334 9822 2386
rect 9874 2334 9886 2386
rect 9938 2334 9950 2386
rect 10002 2334 10014 2386
rect 10066 2334 10078 2386
rect 10130 2334 10142 2386
rect 10194 2334 10206 2386
rect 10258 2334 10270 2386
rect 10322 2334 10334 2386
rect 10386 2334 10398 2386
rect 10450 2334 10462 2386
rect 10514 2334 10526 2386
rect 10578 2334 10590 2386
rect 10642 2334 10654 2386
rect 10706 2334 10718 2386
rect 10770 2334 10782 2386
rect 10834 2334 10846 2386
rect 10898 2334 10910 2386
rect 10962 2334 10974 2386
rect 11026 2334 11038 2386
rect 11090 2334 11102 2386
rect 11154 2334 11166 2386
rect 11218 2334 11230 2386
rect 11282 2334 11294 2386
rect 11346 2334 11358 2386
rect 11410 2334 11422 2386
rect 11474 2334 11486 2386
rect 11538 2334 11550 2386
rect 11602 2334 11614 2386
rect 11666 2334 11678 2386
rect 11730 2334 11742 2386
rect 11794 2334 11806 2386
rect 11858 2334 11870 2386
rect 11922 2334 11934 2386
rect 11986 2334 11998 2386
rect 12050 2334 12062 2386
rect 12114 2334 12126 2386
rect 12178 2334 12190 2386
rect 12242 2334 12254 2386
rect 12306 2334 12318 2386
rect 12370 2334 12382 2386
rect 12434 2334 12446 2386
rect 12498 2334 13040 2386
rect 6148 2332 13040 2334
rect -480 2320 13040 2332
rect 4640 2228 7920 2240
rect 4640 2172 4652 2228
rect 4708 2172 4972 2228
rect 5028 2172 5292 2228
rect 5348 2172 5612 2228
rect 5668 2172 5932 2228
rect 5988 2172 6252 2228
rect 6308 2172 6572 2228
rect 6628 2172 6892 2228
rect 6948 2172 7212 2228
rect 7268 2172 7532 2228
rect 7588 2172 7852 2228
rect 7908 2172 7920 2228
rect 4640 2160 7920 2172
rect -480 2000 4560 2080
rect 4640 2068 7920 2080
rect 4640 2012 5452 2068
rect 5508 2012 7052 2068
rect 7108 2012 7920 2068
rect 4640 2000 7920 2012
rect 8000 2000 13040 2080
rect -400 1828 -160 1920
rect 4640 1908 7920 1920
rect 4640 1852 4652 1908
rect 4708 1852 4972 1908
rect 5028 1852 5292 1908
rect 5348 1852 5612 1908
rect 5668 1852 5932 1908
rect 5988 1852 6252 1908
rect 6308 1852 6572 1908
rect 6628 1852 6892 1908
rect 6948 1852 7212 1908
rect 7268 1852 7532 1908
rect 7588 1852 7852 1908
rect 7908 1852 7920 1908
rect 4640 1840 7920 1852
rect -400 1772 -308 1828
rect -252 1772 -160 1828
rect -400 1680 -160 1772
rect 12720 1828 12960 1920
rect 12720 1772 12812 1828
rect 12868 1772 12960 1828
rect 4640 1748 7920 1760
rect 4640 1692 4652 1748
rect 4708 1692 4972 1748
rect 5028 1692 5292 1748
rect 5348 1692 5612 1748
rect 5668 1692 5932 1748
rect 5988 1692 6252 1748
rect 6308 1692 6572 1748
rect 6628 1692 6892 1748
rect 6948 1692 7212 1748
rect 7268 1692 7532 1748
rect 7588 1692 7852 1748
rect 7908 1692 7920 1748
rect 4640 1680 7920 1692
rect 12720 1680 12960 1772
rect -480 1520 4560 1600
rect 4640 1588 7920 1600
rect 4640 1532 4812 1588
rect 4868 1532 7692 1588
rect 7748 1532 7920 1588
rect 4640 1520 7920 1532
rect 8000 1520 13040 1600
rect 4640 1428 7920 1440
rect 4640 1372 4652 1428
rect 4708 1372 4972 1428
rect 5028 1372 5292 1428
rect 5348 1372 5612 1428
rect 5668 1372 5932 1428
rect 5988 1372 6252 1428
rect 6308 1372 6572 1428
rect 6628 1372 6892 1428
rect 6948 1372 7212 1428
rect 7268 1372 7532 1428
rect 7588 1372 7852 1428
rect 7908 1372 7920 1428
rect 4640 1360 7920 1372
rect -480 1268 13040 1280
rect -480 1266 6092 1268
rect -480 1214 62 1266
rect 114 1214 126 1266
rect 178 1214 190 1266
rect 242 1214 254 1266
rect 306 1214 318 1266
rect 370 1214 382 1266
rect 434 1214 446 1266
rect 498 1214 510 1266
rect 562 1214 574 1266
rect 626 1214 638 1266
rect 690 1214 702 1266
rect 754 1214 766 1266
rect 818 1214 830 1266
rect 882 1214 894 1266
rect 946 1214 958 1266
rect 1010 1214 1022 1266
rect 1074 1214 1086 1266
rect 1138 1214 1150 1266
rect 1202 1214 1214 1266
rect 1266 1214 1278 1266
rect 1330 1214 1342 1266
rect 1394 1214 1406 1266
rect 1458 1214 1470 1266
rect 1522 1214 1534 1266
rect 1586 1214 1598 1266
rect 1650 1214 1662 1266
rect 1714 1214 1726 1266
rect 1778 1214 1790 1266
rect 1842 1214 1854 1266
rect 1906 1214 1918 1266
rect 1970 1214 1982 1266
rect 2034 1214 2046 1266
rect 2098 1214 2110 1266
rect 2162 1214 2174 1266
rect 2226 1214 2238 1266
rect 2290 1214 2302 1266
rect 2354 1214 2366 1266
rect 2418 1214 2430 1266
rect 2482 1214 2494 1266
rect 2546 1214 2558 1266
rect 2610 1214 2622 1266
rect 2674 1214 2686 1266
rect 2738 1214 2750 1266
rect 2802 1214 2814 1266
rect 2866 1214 2878 1266
rect 2930 1214 2942 1266
rect 2994 1214 3006 1266
rect 3058 1214 3070 1266
rect 3122 1214 3134 1266
rect 3186 1214 3198 1266
rect 3250 1214 3262 1266
rect 3314 1214 3326 1266
rect 3378 1214 3390 1266
rect 3442 1214 3454 1266
rect 3506 1214 3518 1266
rect 3570 1214 3582 1266
rect 3634 1214 3646 1266
rect 3698 1214 3710 1266
rect 3762 1214 3774 1266
rect 3826 1214 3838 1266
rect 3890 1214 3902 1266
rect 3954 1214 3966 1266
rect 4018 1214 6092 1266
rect -480 1212 6092 1214
rect 6148 1266 13040 1268
rect 6148 1214 8542 1266
rect 8594 1214 8606 1266
rect 8658 1214 8670 1266
rect 8722 1214 8734 1266
rect 8786 1214 8798 1266
rect 8850 1214 8862 1266
rect 8914 1214 8926 1266
rect 8978 1214 8990 1266
rect 9042 1214 9054 1266
rect 9106 1214 9118 1266
rect 9170 1214 9182 1266
rect 9234 1214 9246 1266
rect 9298 1214 9310 1266
rect 9362 1214 9374 1266
rect 9426 1214 9438 1266
rect 9490 1214 9502 1266
rect 9554 1214 9566 1266
rect 9618 1214 9630 1266
rect 9682 1214 9694 1266
rect 9746 1214 9758 1266
rect 9810 1214 9822 1266
rect 9874 1214 9886 1266
rect 9938 1214 9950 1266
rect 10002 1214 10014 1266
rect 10066 1214 10078 1266
rect 10130 1214 10142 1266
rect 10194 1214 10206 1266
rect 10258 1214 10270 1266
rect 10322 1214 10334 1266
rect 10386 1214 10398 1266
rect 10450 1214 10462 1266
rect 10514 1214 10526 1266
rect 10578 1214 10590 1266
rect 10642 1214 10654 1266
rect 10706 1214 10718 1266
rect 10770 1214 10782 1266
rect 10834 1214 10846 1266
rect 10898 1214 10910 1266
rect 10962 1214 10974 1266
rect 11026 1214 11038 1266
rect 11090 1214 11102 1266
rect 11154 1214 11166 1266
rect 11218 1214 11230 1266
rect 11282 1214 11294 1266
rect 11346 1214 11358 1266
rect 11410 1214 11422 1266
rect 11474 1214 11486 1266
rect 11538 1214 11550 1266
rect 11602 1214 11614 1266
rect 11666 1214 11678 1266
rect 11730 1214 11742 1266
rect 11794 1214 11806 1266
rect 11858 1214 11870 1266
rect 11922 1214 11934 1266
rect 11986 1214 11998 1266
rect 12050 1214 12062 1266
rect 12114 1214 12126 1266
rect 12178 1214 12190 1266
rect 12242 1214 12254 1266
rect 12306 1214 12318 1266
rect 12370 1214 12382 1266
rect 12434 1214 12446 1266
rect 12498 1214 13040 1266
rect 6148 1212 13040 1214
rect -480 1200 13040 1212
rect 4640 1108 7920 1120
rect 4640 1052 4652 1108
rect 4708 1052 4972 1108
rect 5028 1052 5292 1108
rect 5348 1052 5612 1108
rect 5668 1052 5932 1108
rect 5988 1052 6252 1108
rect 6308 1052 6572 1108
rect 6628 1052 6892 1108
rect 6948 1052 7212 1108
rect 7268 1052 7532 1108
rect 7588 1052 7852 1108
rect 7908 1052 7920 1108
rect 4640 1040 7920 1052
rect -480 948 5840 960
rect -480 946 5132 948
rect -480 894 62 946
rect 114 894 126 946
rect 178 894 190 946
rect 242 894 254 946
rect 306 894 318 946
rect 370 894 382 946
rect 434 894 446 946
rect 498 894 510 946
rect 562 894 574 946
rect 626 894 638 946
rect 690 894 702 946
rect 754 894 766 946
rect 818 894 830 946
rect 882 894 894 946
rect 946 894 958 946
rect 1010 894 1022 946
rect 1074 894 1086 946
rect 1138 894 1150 946
rect 1202 894 1214 946
rect 1266 894 1278 946
rect 1330 894 1342 946
rect 1394 894 1406 946
rect 1458 894 1470 946
rect 1522 894 1534 946
rect 1586 894 1598 946
rect 1650 894 1662 946
rect 1714 894 1726 946
rect 1778 894 1790 946
rect 1842 894 1854 946
rect 1906 894 1918 946
rect 1970 894 1982 946
rect 2034 894 2046 946
rect 2098 894 2110 946
rect 2162 894 2174 946
rect 2226 894 2238 946
rect 2290 894 2302 946
rect 2354 894 2366 946
rect 2418 894 2430 946
rect 2482 894 2494 946
rect 2546 894 2558 946
rect 2610 894 2622 946
rect 2674 894 2686 946
rect 2738 894 2750 946
rect 2802 894 2814 946
rect 2866 894 2878 946
rect 2930 894 2942 946
rect 2994 894 3006 946
rect 3058 894 3070 946
rect 3122 894 3134 946
rect 3186 894 3198 946
rect 3250 894 3262 946
rect 3314 894 3326 946
rect 3378 894 3390 946
rect 3442 894 3454 946
rect 3506 894 3518 946
rect 3570 894 3582 946
rect 3634 894 3646 946
rect 3698 894 3710 946
rect 3762 894 3774 946
rect 3826 894 3838 946
rect 3890 894 3902 946
rect 3954 894 3966 946
rect 4018 894 4174 946
rect 4226 894 5132 946
rect -480 892 5132 894
rect 5188 892 5840 948
rect -480 880 5840 892
rect 5920 948 6640 960
rect 5920 892 5932 948
rect 5988 892 6252 948
rect 6308 892 6572 948
rect 6628 892 6640 948
rect 5920 880 6640 892
rect 6720 948 13040 960
rect 6720 892 6732 948
rect 6788 946 13040 948
rect 6788 894 8334 946
rect 8386 894 8542 946
rect 8594 894 8606 946
rect 8658 894 8670 946
rect 8722 894 8734 946
rect 8786 894 8798 946
rect 8850 894 8862 946
rect 8914 894 8926 946
rect 8978 894 8990 946
rect 9042 894 9054 946
rect 9106 894 9118 946
rect 9170 894 9182 946
rect 9234 894 9246 946
rect 9298 894 9310 946
rect 9362 894 9374 946
rect 9426 894 9438 946
rect 9490 894 9502 946
rect 9554 894 9566 946
rect 9618 894 9630 946
rect 9682 894 9694 946
rect 9746 894 9758 946
rect 9810 894 9822 946
rect 9874 894 9886 946
rect 9938 894 9950 946
rect 10002 894 10014 946
rect 10066 894 10078 946
rect 10130 894 10142 946
rect 10194 894 10206 946
rect 10258 894 10270 946
rect 10322 894 10334 946
rect 10386 894 10398 946
rect 10450 894 10462 946
rect 10514 894 10526 946
rect 10578 894 10590 946
rect 10642 894 10654 946
rect 10706 894 10718 946
rect 10770 894 10782 946
rect 10834 894 10846 946
rect 10898 894 10910 946
rect 10962 894 10974 946
rect 11026 894 11038 946
rect 11090 894 11102 946
rect 11154 894 11166 946
rect 11218 894 11230 946
rect 11282 894 11294 946
rect 11346 894 11358 946
rect 11410 894 11422 946
rect 11474 894 11486 946
rect 11538 894 11550 946
rect 11602 894 11614 946
rect 11666 894 11678 946
rect 11730 894 11742 946
rect 11794 894 11806 946
rect 11858 894 11870 946
rect 11922 894 11934 946
rect 11986 894 11998 946
rect 12050 894 12062 946
rect 12114 894 12126 946
rect 12178 894 12190 946
rect 12242 894 12254 946
rect 12306 894 12318 946
rect 12370 894 12382 946
rect 12434 894 12446 946
rect 12498 894 13040 946
rect 6788 892 13040 894
rect 6720 880 13040 892
rect 4640 788 7920 800
rect 4640 732 4652 788
rect 4708 732 4972 788
rect 5028 732 5292 788
rect 5348 732 5612 788
rect 5668 732 5932 788
rect 5988 732 6252 788
rect 6308 732 6572 788
rect 6628 732 6892 788
rect 6948 732 7212 788
rect 7268 732 7532 788
rect 7588 732 7852 788
rect 7908 732 7920 788
rect 4640 720 7920 732
rect 4640 628 7920 640
rect 4640 572 5132 628
rect 5188 572 7372 628
rect 7428 572 7920 628
rect 4640 560 7920 572
rect 4640 468 7920 480
rect 4640 412 4652 468
rect 4708 412 4972 468
rect 5028 412 5292 468
rect 5348 412 5612 468
rect 5668 412 5932 468
rect 5988 412 6252 468
rect 6308 412 6572 468
rect 6628 412 6892 468
rect 6948 412 7212 468
rect 7268 412 7532 468
rect 7588 412 7852 468
rect 7908 412 7920 468
rect 4640 400 7920 412
rect 4640 308 7920 320
rect 4640 252 4652 308
rect 4708 252 4972 308
rect 5028 252 5292 308
rect 5348 252 5612 308
rect 5668 252 5932 308
rect 5988 252 6252 308
rect 6308 252 6572 308
rect 6628 252 6892 308
rect 6948 252 7212 308
rect 7268 252 7532 308
rect 7588 252 7852 308
rect 7908 252 7920 308
rect 4640 240 7920 252
rect -480 148 5840 160
rect -480 146 4812 148
rect -480 94 -146 146
rect -94 94 62 146
rect 114 94 126 146
rect 178 94 190 146
rect 242 94 254 146
rect 306 94 318 146
rect 370 94 382 146
rect 434 94 446 146
rect 498 94 510 146
rect 562 94 574 146
rect 626 94 638 146
rect 690 94 702 146
rect 754 94 766 146
rect 818 94 830 146
rect 882 94 894 146
rect 946 94 958 146
rect 1010 94 1022 146
rect 1074 94 1086 146
rect 1138 94 1150 146
rect 1202 94 1214 146
rect 1266 94 1278 146
rect 1330 94 1342 146
rect 1394 94 1406 146
rect 1458 94 1470 146
rect 1522 94 1534 146
rect 1586 94 1598 146
rect 1650 94 1662 146
rect 1714 94 1726 146
rect 1778 94 1790 146
rect 1842 94 1854 146
rect 1906 94 1918 146
rect 1970 94 1982 146
rect 2034 94 2046 146
rect 2098 94 2110 146
rect 2162 94 2174 146
rect 2226 94 2238 146
rect 2290 94 2302 146
rect 2354 94 2366 146
rect 2418 94 2430 146
rect 2482 94 2494 146
rect 2546 94 2558 146
rect 2610 94 2622 146
rect 2674 94 2686 146
rect 2738 94 2750 146
rect 2802 94 2814 146
rect 2866 94 2878 146
rect 2930 94 2942 146
rect 2994 94 3006 146
rect 3058 94 3070 146
rect 3122 94 3134 146
rect 3186 94 3198 146
rect 3250 94 3262 146
rect 3314 94 3326 146
rect 3378 94 3390 146
rect 3442 94 3454 146
rect 3506 94 3518 146
rect 3570 94 3582 146
rect 3634 94 3646 146
rect 3698 94 3710 146
rect 3762 94 3774 146
rect 3826 94 3838 146
rect 3890 94 3902 146
rect 3954 94 3966 146
rect 4018 94 4812 146
rect -480 92 4812 94
rect 4868 92 5840 148
rect -480 80 5840 92
rect 5920 148 6640 160
rect 5920 92 5932 148
rect 5988 92 6252 148
rect 6308 92 6572 148
rect 6628 92 6640 148
rect 5920 80 6640 92
rect 6720 148 13040 160
rect 6720 92 7052 148
rect 7108 146 13040 148
rect 7108 94 8542 146
rect 8594 94 8606 146
rect 8658 94 8670 146
rect 8722 94 8734 146
rect 8786 94 8798 146
rect 8850 94 8862 146
rect 8914 94 8926 146
rect 8978 94 8990 146
rect 9042 94 9054 146
rect 9106 94 9118 146
rect 9170 94 9182 146
rect 9234 94 9246 146
rect 9298 94 9310 146
rect 9362 94 9374 146
rect 9426 94 9438 146
rect 9490 94 9502 146
rect 9554 94 9566 146
rect 9618 94 9630 146
rect 9682 94 9694 146
rect 9746 94 9758 146
rect 9810 94 9822 146
rect 9874 94 9886 146
rect 9938 94 9950 146
rect 10002 94 10014 146
rect 10066 94 10078 146
rect 10130 94 10142 146
rect 10194 94 10206 146
rect 10258 94 10270 146
rect 10322 94 10334 146
rect 10386 94 10398 146
rect 10450 94 10462 146
rect 10514 94 10526 146
rect 10578 94 10590 146
rect 10642 94 10654 146
rect 10706 94 10718 146
rect 10770 94 10782 146
rect 10834 94 10846 146
rect 10898 94 10910 146
rect 10962 94 10974 146
rect 11026 94 11038 146
rect 11090 94 11102 146
rect 11154 94 11166 146
rect 11218 94 11230 146
rect 11282 94 11294 146
rect 11346 94 11358 146
rect 11410 94 11422 146
rect 11474 94 11486 146
rect 11538 94 11550 146
rect 11602 94 11614 146
rect 11666 94 11678 146
rect 11730 94 11742 146
rect 11794 94 11806 146
rect 11858 94 11870 146
rect 11922 94 11934 146
rect 11986 94 11998 146
rect 12050 94 12062 146
rect 12114 94 12126 146
rect 12178 94 12190 146
rect 12242 94 12254 146
rect 12306 94 12318 146
rect 12370 94 12382 146
rect 12434 94 12446 146
rect 12498 94 12654 146
rect 12706 94 13040 146
rect 7108 92 13040 94
rect 6720 80 13040 92
rect 4640 -12 7920 0
rect 4640 -68 4652 -12
rect 4708 -68 4972 -12
rect 5028 -68 5292 -12
rect 5348 -68 5612 -12
rect 5668 -68 5932 -12
rect 5988 -68 6252 -12
rect 6308 -68 6572 -12
rect 6628 -68 6892 -12
rect 6948 -68 7212 -12
rect 7268 -68 7532 -12
rect 7588 -68 7852 -12
rect 7908 -68 7920 -12
rect 4640 -80 7920 -68
rect -480 -172 13040 -160
rect -480 -174 6092 -172
rect -480 -226 62 -174
rect 114 -226 126 -174
rect 178 -226 190 -174
rect 242 -226 254 -174
rect 306 -226 318 -174
rect 370 -226 382 -174
rect 434 -226 446 -174
rect 498 -226 510 -174
rect 562 -226 574 -174
rect 626 -226 638 -174
rect 690 -226 702 -174
rect 754 -226 766 -174
rect 818 -226 830 -174
rect 882 -226 894 -174
rect 946 -226 958 -174
rect 1010 -226 1022 -174
rect 1074 -226 1086 -174
rect 1138 -226 1150 -174
rect 1202 -226 1214 -174
rect 1266 -226 1278 -174
rect 1330 -226 1342 -174
rect 1394 -226 1406 -174
rect 1458 -226 1470 -174
rect 1522 -226 1534 -174
rect 1586 -226 1598 -174
rect 1650 -226 1662 -174
rect 1714 -226 1726 -174
rect 1778 -226 1790 -174
rect 1842 -226 1854 -174
rect 1906 -226 1918 -174
rect 1970 -226 1982 -174
rect 2034 -226 2046 -174
rect 2098 -226 2110 -174
rect 2162 -226 2174 -174
rect 2226 -226 2238 -174
rect 2290 -226 2302 -174
rect 2354 -226 2366 -174
rect 2418 -226 2430 -174
rect 2482 -226 2494 -174
rect 2546 -226 2558 -174
rect 2610 -226 2622 -174
rect 2674 -226 2686 -174
rect 2738 -226 2750 -174
rect 2802 -226 2814 -174
rect 2866 -226 2878 -174
rect 2930 -226 2942 -174
rect 2994 -226 3006 -174
rect 3058 -226 3070 -174
rect 3122 -226 3134 -174
rect 3186 -226 3198 -174
rect 3250 -226 3262 -174
rect 3314 -226 3326 -174
rect 3378 -226 3390 -174
rect 3442 -226 3454 -174
rect 3506 -226 3518 -174
rect 3570 -226 3582 -174
rect 3634 -226 3646 -174
rect 3698 -226 3710 -174
rect 3762 -226 3774 -174
rect 3826 -226 3838 -174
rect 3890 -226 3902 -174
rect 3954 -226 3966 -174
rect 4018 -226 6092 -174
rect -480 -228 6092 -226
rect 6148 -174 13040 -172
rect 6148 -226 8542 -174
rect 8594 -226 8606 -174
rect 8658 -226 8670 -174
rect 8722 -226 8734 -174
rect 8786 -226 8798 -174
rect 8850 -226 8862 -174
rect 8914 -226 8926 -174
rect 8978 -226 8990 -174
rect 9042 -226 9054 -174
rect 9106 -226 9118 -174
rect 9170 -226 9182 -174
rect 9234 -226 9246 -174
rect 9298 -226 9310 -174
rect 9362 -226 9374 -174
rect 9426 -226 9438 -174
rect 9490 -226 9502 -174
rect 9554 -226 9566 -174
rect 9618 -226 9630 -174
rect 9682 -226 9694 -174
rect 9746 -226 9758 -174
rect 9810 -226 9822 -174
rect 9874 -226 9886 -174
rect 9938 -226 9950 -174
rect 10002 -226 10014 -174
rect 10066 -226 10078 -174
rect 10130 -226 10142 -174
rect 10194 -226 10206 -174
rect 10258 -226 10270 -174
rect 10322 -226 10334 -174
rect 10386 -226 10398 -174
rect 10450 -226 10462 -174
rect 10514 -226 10526 -174
rect 10578 -226 10590 -174
rect 10642 -226 10654 -174
rect 10706 -226 10718 -174
rect 10770 -226 10782 -174
rect 10834 -226 10846 -174
rect 10898 -226 10910 -174
rect 10962 -226 10974 -174
rect 11026 -226 11038 -174
rect 11090 -226 11102 -174
rect 11154 -226 11166 -174
rect 11218 -226 11230 -174
rect 11282 -226 11294 -174
rect 11346 -226 11358 -174
rect 11410 -226 11422 -174
rect 11474 -226 11486 -174
rect 11538 -226 11550 -174
rect 11602 -226 11614 -174
rect 11666 -226 11678 -174
rect 11730 -226 11742 -174
rect 11794 -226 11806 -174
rect 11858 -226 11870 -174
rect 11922 -226 11934 -174
rect 11986 -226 11998 -174
rect 12050 -226 12062 -174
rect 12114 -226 12126 -174
rect 12178 -226 12190 -174
rect 12242 -226 12254 -174
rect 12306 -226 12318 -174
rect 12370 -226 12382 -174
rect 12434 -226 12446 -174
rect 12498 -226 13040 -174
rect 6148 -228 13040 -226
rect -480 -240 13040 -228
rect 4640 -332 7920 -320
rect 4640 -388 4652 -332
rect 4708 -388 4972 -332
rect 5028 -388 5292 -332
rect 5348 -388 5612 -332
rect 5668 -388 5932 -332
rect 5988 -388 6252 -332
rect 6308 -388 6572 -332
rect 6628 -388 6892 -332
rect 6948 -388 7212 -332
rect 7268 -388 7532 -332
rect 7588 -388 7852 -332
rect 7908 -388 7920 -332
rect 4640 -400 7920 -388
rect -480 -492 13040 -480
rect -480 -494 6412 -492
rect -480 -546 -306 -494
rect -254 -546 6412 -494
rect -480 -548 6412 -546
rect 6468 -494 13040 -492
rect 6468 -546 12814 -494
rect 12866 -546 13040 -494
rect 6468 -548 13040 -546
rect -480 -560 13040 -548
rect 4640 -652 7920 -640
rect 4640 -708 4652 -652
rect 4708 -708 4972 -652
rect 5028 -708 5292 -652
rect 5348 -708 5612 -652
rect 5668 -708 5932 -652
rect 5988 -708 6252 -652
rect 6308 -708 6572 -652
rect 6628 -708 6892 -652
rect 6948 -708 7212 -652
rect 7268 -708 7532 -652
rect 7588 -708 7852 -652
rect 7908 -708 7920 -652
rect 4640 -720 7920 -708
<< via2 >>
rect 4652 4252 4708 4308
rect 4972 4252 5028 4308
rect 5292 4252 5348 4308
rect 5612 4252 5668 4308
rect 5932 4252 5988 4308
rect 6252 4252 6308 4308
rect 6572 4252 6628 4308
rect 6892 4252 6948 4308
rect 7212 4252 7268 4308
rect 7532 4252 7588 4308
rect 7852 4252 7908 4308
rect 6412 4092 6468 4148
rect 4652 3932 4708 3988
rect 4972 3932 5028 3988
rect 5292 3932 5348 3988
rect 5612 3932 5668 3988
rect 5932 3932 5988 3988
rect 6252 3932 6308 3988
rect 6572 3932 6628 3988
rect 6892 3932 6948 3988
rect 7212 3932 7268 3988
rect 7532 3932 7588 3988
rect 7852 3932 7908 3988
rect 6092 3772 6148 3828
rect 4652 3612 4708 3668
rect 4972 3612 5028 3668
rect 5292 3612 5348 3668
rect 5612 3612 5668 3668
rect 5932 3612 5988 3668
rect 6252 3612 6308 3668
rect 6572 3612 6628 3668
rect 6892 3612 6948 3668
rect 7212 3612 7268 3668
rect 7532 3612 7588 3668
rect 7852 3612 7908 3668
rect 5452 3452 5508 3508
rect 5932 3452 5988 3508
rect 6252 3452 6308 3508
rect 6572 3452 6628 3508
rect 7692 3452 7748 3508
rect 4652 3292 4708 3348
rect 4972 3292 5028 3348
rect 5292 3292 5348 3348
rect 5612 3292 5668 3348
rect 5932 3292 5988 3348
rect 6252 3292 6308 3348
rect 6572 3292 6628 3348
rect 6892 3292 6948 3348
rect 7212 3292 7268 3348
rect 7532 3292 7588 3348
rect 7852 3292 7908 3348
rect 4652 3132 4708 3188
rect 4972 3132 5028 3188
rect 5292 3132 5348 3188
rect 5612 3132 5668 3188
rect 5932 3132 5988 3188
rect 6252 3132 6308 3188
rect 6572 3132 6628 3188
rect 6892 3132 6948 3188
rect 7212 3132 7268 3188
rect 7532 3132 7588 3188
rect 7852 3132 7908 3188
rect 5772 2972 5828 3028
rect 6732 2972 6788 3028
rect 4652 2812 4708 2868
rect 4972 2812 5028 2868
rect 5292 2812 5348 2868
rect 5612 2812 5668 2868
rect 5932 2812 5988 2868
rect 6252 2812 6308 2868
rect 6572 2812 6628 2868
rect 6892 2812 6948 2868
rect 7212 2812 7268 2868
rect 7532 2812 7588 2868
rect 7852 2812 7908 2868
rect 5772 2652 5828 2708
rect 5932 2652 5988 2708
rect 6252 2652 6308 2708
rect 6572 2652 6628 2708
rect 7372 2652 7428 2708
rect 4652 2492 4708 2548
rect 4972 2492 5028 2548
rect 5292 2492 5348 2548
rect 5612 2492 5668 2548
rect 5932 2492 5988 2548
rect 6252 2492 6308 2548
rect 6572 2492 6628 2548
rect 6892 2492 6948 2548
rect 7212 2492 7268 2548
rect 7532 2492 7588 2548
rect 7852 2492 7908 2548
rect 6092 2332 6148 2388
rect 4652 2172 4708 2228
rect 4972 2172 5028 2228
rect 5292 2172 5348 2228
rect 5612 2172 5668 2228
rect 5932 2172 5988 2228
rect 6252 2172 6308 2228
rect 6572 2172 6628 2228
rect 6892 2172 6948 2228
rect 7212 2172 7268 2228
rect 7532 2172 7588 2228
rect 7852 2172 7908 2228
rect 5452 2012 5508 2068
rect 7052 2012 7108 2068
rect 4652 1852 4708 1908
rect 4972 1852 5028 1908
rect 5292 1852 5348 1908
rect 5612 1852 5668 1908
rect 5932 1852 5988 1908
rect 6252 1852 6308 1908
rect 6572 1852 6628 1908
rect 6892 1852 6948 1908
rect 7212 1852 7268 1908
rect 7532 1852 7588 1908
rect 7852 1852 7908 1908
rect -308 1826 -252 1828
rect -308 1774 -306 1826
rect -306 1774 -254 1826
rect -254 1774 -252 1826
rect -308 1772 -252 1774
rect 12812 1826 12868 1828
rect 12812 1774 12814 1826
rect 12814 1774 12866 1826
rect 12866 1774 12868 1826
rect 12812 1772 12868 1774
rect 4652 1692 4708 1748
rect 4972 1692 5028 1748
rect 5292 1692 5348 1748
rect 5612 1692 5668 1748
rect 5932 1692 5988 1748
rect 6252 1692 6308 1748
rect 6572 1692 6628 1748
rect 6892 1692 6948 1748
rect 7212 1692 7268 1748
rect 7532 1692 7588 1748
rect 7852 1692 7908 1748
rect 4812 1532 4868 1588
rect 7692 1532 7748 1588
rect 4652 1372 4708 1428
rect 4972 1372 5028 1428
rect 5292 1372 5348 1428
rect 5612 1372 5668 1428
rect 5932 1372 5988 1428
rect 6252 1372 6308 1428
rect 6572 1372 6628 1428
rect 6892 1372 6948 1428
rect 7212 1372 7268 1428
rect 7532 1372 7588 1428
rect 7852 1372 7908 1428
rect 6092 1212 6148 1268
rect 4652 1052 4708 1108
rect 4972 1052 5028 1108
rect 5292 1052 5348 1108
rect 5612 1052 5668 1108
rect 5932 1052 5988 1108
rect 6252 1052 6308 1108
rect 6572 1052 6628 1108
rect 6892 1052 6948 1108
rect 7212 1052 7268 1108
rect 7532 1052 7588 1108
rect 7852 1052 7908 1108
rect 5132 892 5188 948
rect 5932 892 5988 948
rect 6252 892 6308 948
rect 6572 892 6628 948
rect 6732 892 6788 948
rect 4652 732 4708 788
rect 4972 732 5028 788
rect 5292 732 5348 788
rect 5612 732 5668 788
rect 5932 732 5988 788
rect 6252 732 6308 788
rect 6572 732 6628 788
rect 6892 732 6948 788
rect 7212 732 7268 788
rect 7532 732 7588 788
rect 7852 732 7908 788
rect 5132 572 5188 628
rect 7372 572 7428 628
rect 4652 412 4708 468
rect 4972 412 5028 468
rect 5292 412 5348 468
rect 5612 412 5668 468
rect 5932 412 5988 468
rect 6252 412 6308 468
rect 6572 412 6628 468
rect 6892 412 6948 468
rect 7212 412 7268 468
rect 7532 412 7588 468
rect 7852 412 7908 468
rect 4652 252 4708 308
rect 4972 252 5028 308
rect 5292 252 5348 308
rect 5612 252 5668 308
rect 5932 252 5988 308
rect 6252 252 6308 308
rect 6572 252 6628 308
rect 6892 252 6948 308
rect 7212 252 7268 308
rect 7532 252 7588 308
rect 7852 252 7908 308
rect 4812 92 4868 148
rect 5932 92 5988 148
rect 6252 92 6308 148
rect 6572 92 6628 148
rect 7052 92 7108 148
rect 4652 -68 4708 -12
rect 4972 -68 5028 -12
rect 5292 -68 5348 -12
rect 5612 -68 5668 -12
rect 5932 -68 5988 -12
rect 6252 -68 6308 -12
rect 6572 -68 6628 -12
rect 6892 -68 6948 -12
rect 7212 -68 7268 -12
rect 7532 -68 7588 -12
rect 7852 -68 7908 -12
rect 6092 -228 6148 -172
rect 4652 -388 4708 -332
rect 4972 -388 5028 -332
rect 5292 -388 5348 -332
rect 5612 -388 5668 -332
rect 5932 -388 5988 -332
rect 6252 -388 6308 -332
rect 6572 -388 6628 -332
rect 6892 -388 6948 -332
rect 7212 -388 7268 -332
rect 7532 -388 7588 -332
rect 7852 -388 7908 -332
rect 6412 -548 6468 -492
rect 4652 -708 4708 -652
rect 4972 -708 5028 -652
rect 5292 -708 5348 -652
rect 5612 -708 5668 -652
rect 5932 -708 5988 -652
rect 6252 -708 6308 -652
rect 6572 -708 6628 -652
rect 6892 -708 6948 -652
rect 7212 -708 7268 -652
rect 7532 -708 7588 -652
rect 7852 -708 7908 -652
<< metal3 >>
rect 4640 4312 4720 4320
rect 4640 4248 4648 4312
rect 4712 4248 4720 4312
rect 4640 3992 4720 4248
rect 4640 3928 4648 3992
rect 4712 3928 4720 3992
rect 4640 3672 4720 3928
rect 4640 3608 4648 3672
rect 4712 3608 4720 3672
rect 4640 3352 4720 3608
rect 4640 3288 4648 3352
rect 4712 3288 4720 3352
rect 4640 3192 4720 3288
rect 4640 3128 4648 3192
rect 4712 3128 4720 3192
rect 4640 2872 4720 3128
rect 4640 2808 4648 2872
rect 4712 2808 4720 2872
rect 4640 2552 4720 2808
rect 4640 2488 4648 2552
rect 4712 2488 4720 2552
rect 4640 2232 4720 2488
rect 4640 2168 4648 2232
rect 4712 2168 4720 2232
rect -400 1832 -160 1920
rect -400 1768 -312 1832
rect -248 1768 -160 1832
rect -400 1680 -160 1768
rect 4640 1912 4720 2168
rect 4640 1848 4648 1912
rect 4712 1848 4720 1912
rect 4640 1752 4720 1848
rect 4640 1688 4648 1752
rect 4712 1688 4720 1752
rect 4640 1432 4720 1688
rect 4640 1368 4648 1432
rect 4712 1368 4720 1432
rect 4640 1112 4720 1368
rect 4640 1048 4648 1112
rect 4712 1048 4720 1112
rect 4640 792 4720 1048
rect 4640 728 4648 792
rect 4712 728 4720 792
rect 4640 472 4720 728
rect 4640 408 4648 472
rect 4712 408 4720 472
rect 4640 312 4720 408
rect 4640 248 4648 312
rect 4712 248 4720 312
rect 4640 -8 4720 248
rect 4640 -72 4648 -8
rect 4712 -72 4720 -8
rect 4640 -328 4720 -72
rect 4640 -392 4648 -328
rect 4712 -392 4720 -328
rect 4640 -648 4720 -392
rect 4640 -712 4648 -648
rect 4712 -712 4720 -648
rect 4640 -720 4720 -712
rect 4800 1588 4880 4320
rect 4800 1532 4812 1588
rect 4868 1532 4880 1588
rect 4800 148 4880 1532
rect 4800 92 4812 148
rect 4868 92 4880 148
rect 4800 -720 4880 92
rect 4960 4312 5040 4320
rect 4960 4248 4968 4312
rect 5032 4248 5040 4312
rect 4960 3992 5040 4248
rect 4960 3928 4968 3992
rect 5032 3928 5040 3992
rect 4960 3672 5040 3928
rect 4960 3608 4968 3672
rect 5032 3608 5040 3672
rect 4960 3352 5040 3608
rect 4960 3288 4968 3352
rect 5032 3288 5040 3352
rect 4960 3192 5040 3288
rect 4960 3128 4968 3192
rect 5032 3128 5040 3192
rect 4960 2872 5040 3128
rect 4960 2808 4968 2872
rect 5032 2808 5040 2872
rect 4960 2552 5040 2808
rect 4960 2488 4968 2552
rect 5032 2488 5040 2552
rect 4960 2232 5040 2488
rect 4960 2168 4968 2232
rect 5032 2168 5040 2232
rect 4960 1912 5040 2168
rect 4960 1848 4968 1912
rect 5032 1848 5040 1912
rect 4960 1752 5040 1848
rect 4960 1688 4968 1752
rect 5032 1688 5040 1752
rect 4960 1432 5040 1688
rect 4960 1368 4968 1432
rect 5032 1368 5040 1432
rect 4960 1112 5040 1368
rect 4960 1048 4968 1112
rect 5032 1048 5040 1112
rect 4960 792 5040 1048
rect 4960 728 4968 792
rect 5032 728 5040 792
rect 4960 472 5040 728
rect 4960 408 4968 472
rect 5032 408 5040 472
rect 4960 312 5040 408
rect 4960 248 4968 312
rect 5032 248 5040 312
rect 4960 -8 5040 248
rect 4960 -72 4968 -8
rect 5032 -72 5040 -8
rect 4960 -328 5040 -72
rect 4960 -392 4968 -328
rect 5032 -392 5040 -328
rect 4960 -648 5040 -392
rect 4960 -712 4968 -648
rect 5032 -712 5040 -648
rect 4960 -720 5040 -712
rect 5120 948 5200 4320
rect 5120 892 5132 948
rect 5188 892 5200 948
rect 5120 628 5200 892
rect 5120 572 5132 628
rect 5188 572 5200 628
rect 5120 -720 5200 572
rect 5280 4312 5360 4320
rect 5280 4248 5288 4312
rect 5352 4248 5360 4312
rect 5280 3992 5360 4248
rect 5280 3928 5288 3992
rect 5352 3928 5360 3992
rect 5280 3672 5360 3928
rect 5280 3608 5288 3672
rect 5352 3608 5360 3672
rect 5280 3352 5360 3608
rect 5280 3288 5288 3352
rect 5352 3288 5360 3352
rect 5280 3192 5360 3288
rect 5280 3128 5288 3192
rect 5352 3128 5360 3192
rect 5280 2872 5360 3128
rect 5280 2808 5288 2872
rect 5352 2808 5360 2872
rect 5280 2552 5360 2808
rect 5280 2488 5288 2552
rect 5352 2488 5360 2552
rect 5280 2232 5360 2488
rect 5280 2168 5288 2232
rect 5352 2168 5360 2232
rect 5280 1912 5360 2168
rect 5280 1848 5288 1912
rect 5352 1848 5360 1912
rect 5280 1752 5360 1848
rect 5280 1688 5288 1752
rect 5352 1688 5360 1752
rect 5280 1432 5360 1688
rect 5280 1368 5288 1432
rect 5352 1368 5360 1432
rect 5280 1112 5360 1368
rect 5280 1048 5288 1112
rect 5352 1048 5360 1112
rect 5280 792 5360 1048
rect 5280 728 5288 792
rect 5352 728 5360 792
rect 5280 472 5360 728
rect 5280 408 5288 472
rect 5352 408 5360 472
rect 5280 312 5360 408
rect 5280 248 5288 312
rect 5352 248 5360 312
rect 5280 -8 5360 248
rect 5280 -72 5288 -8
rect 5352 -72 5360 -8
rect 5280 -328 5360 -72
rect 5280 -392 5288 -328
rect 5352 -392 5360 -328
rect 5280 -648 5360 -392
rect 5280 -712 5288 -648
rect 5352 -712 5360 -648
rect 5280 -720 5360 -712
rect 5440 3508 5520 4320
rect 5440 3452 5452 3508
rect 5508 3452 5520 3508
rect 5440 2068 5520 3452
rect 5440 2012 5452 2068
rect 5508 2012 5520 2068
rect 5440 -720 5520 2012
rect 5600 4312 5680 4320
rect 5600 4248 5608 4312
rect 5672 4248 5680 4312
rect 5600 3992 5680 4248
rect 5600 3928 5608 3992
rect 5672 3928 5680 3992
rect 5600 3672 5680 3928
rect 5600 3608 5608 3672
rect 5672 3608 5680 3672
rect 5600 3352 5680 3608
rect 5600 3288 5608 3352
rect 5672 3288 5680 3352
rect 5600 3192 5680 3288
rect 5600 3128 5608 3192
rect 5672 3128 5680 3192
rect 5600 2872 5680 3128
rect 5600 2808 5608 2872
rect 5672 2808 5680 2872
rect 5600 2552 5680 2808
rect 5600 2488 5608 2552
rect 5672 2488 5680 2552
rect 5600 2232 5680 2488
rect 5600 2168 5608 2232
rect 5672 2168 5680 2232
rect 5600 1912 5680 2168
rect 5600 1848 5608 1912
rect 5672 1848 5680 1912
rect 5600 1752 5680 1848
rect 5600 1688 5608 1752
rect 5672 1688 5680 1752
rect 5600 1432 5680 1688
rect 5600 1368 5608 1432
rect 5672 1368 5680 1432
rect 5600 1112 5680 1368
rect 5600 1048 5608 1112
rect 5672 1048 5680 1112
rect 5600 792 5680 1048
rect 5600 728 5608 792
rect 5672 728 5680 792
rect 5600 472 5680 728
rect 5600 408 5608 472
rect 5672 408 5680 472
rect 5600 312 5680 408
rect 5600 248 5608 312
rect 5672 248 5680 312
rect 5600 -8 5680 248
rect 5600 -72 5608 -8
rect 5672 -72 5680 -8
rect 5600 -328 5680 -72
rect 5600 -392 5608 -328
rect 5672 -392 5680 -328
rect 5600 -648 5680 -392
rect 5600 -712 5608 -648
rect 5672 -712 5680 -648
rect 5600 -720 5680 -712
rect 5760 3028 5840 4320
rect 5760 2972 5772 3028
rect 5828 2972 5840 3028
rect 5760 2708 5840 2972
rect 5760 2652 5772 2708
rect 5828 2652 5840 2708
rect 5760 -720 5840 2652
rect 5920 4312 6000 4320
rect 5920 4248 5928 4312
rect 5992 4248 6000 4312
rect 5920 3992 6000 4248
rect 5920 3928 5928 3992
rect 5992 3928 6000 3992
rect 5920 3672 6000 3928
rect 5920 3608 5928 3672
rect 5992 3608 6000 3672
rect 5920 3512 6000 3608
rect 5920 3448 5928 3512
rect 5992 3448 6000 3512
rect 5920 3352 6000 3448
rect 5920 3288 5928 3352
rect 5992 3288 6000 3352
rect 5920 3192 6000 3288
rect 5920 3128 5928 3192
rect 5992 3128 6000 3192
rect 5920 2872 6000 3128
rect 5920 2808 5928 2872
rect 5992 2808 6000 2872
rect 5920 2712 6000 2808
rect 5920 2648 5928 2712
rect 5992 2648 6000 2712
rect 5920 2552 6000 2648
rect 5920 2488 5928 2552
rect 5992 2488 6000 2552
rect 5920 2232 6000 2488
rect 5920 2168 5928 2232
rect 5992 2168 6000 2232
rect 5920 1912 6000 2168
rect 5920 1848 5928 1912
rect 5992 1848 6000 1912
rect 5920 1752 6000 1848
rect 5920 1688 5928 1752
rect 5992 1688 6000 1752
rect 5920 1432 6000 1688
rect 5920 1368 5928 1432
rect 5992 1368 6000 1432
rect 5920 1112 6000 1368
rect 5920 1048 5928 1112
rect 5992 1048 6000 1112
rect 5920 952 6000 1048
rect 5920 888 5928 952
rect 5992 888 6000 952
rect 5920 792 6000 888
rect 5920 728 5928 792
rect 5992 728 6000 792
rect 5920 472 6000 728
rect 5920 408 5928 472
rect 5992 408 6000 472
rect 5920 312 6000 408
rect 5920 248 5928 312
rect 5992 248 6000 312
rect 5920 152 6000 248
rect 5920 88 5928 152
rect 5992 88 6000 152
rect 5920 -8 6000 88
rect 5920 -72 5928 -8
rect 5992 -72 6000 -8
rect 5920 -328 6000 -72
rect 5920 -392 5928 -328
rect 5992 -392 6000 -328
rect 5920 -648 6000 -392
rect 5920 -712 5928 -648
rect 5992 -712 6000 -648
rect 5920 -720 6000 -712
rect 6080 3828 6160 4320
rect 6080 3772 6092 3828
rect 6148 3772 6160 3828
rect 6080 2388 6160 3772
rect 6080 2332 6092 2388
rect 6148 2332 6160 2388
rect 6080 1268 6160 2332
rect 6080 1212 6092 1268
rect 6148 1212 6160 1268
rect 6080 -172 6160 1212
rect 6080 -228 6092 -172
rect 6148 -228 6160 -172
rect 6080 -720 6160 -228
rect 6240 4312 6320 4320
rect 6240 4248 6248 4312
rect 6312 4248 6320 4312
rect 6240 3992 6320 4248
rect 6240 3928 6248 3992
rect 6312 3928 6320 3992
rect 6240 3672 6320 3928
rect 6240 3608 6248 3672
rect 6312 3608 6320 3672
rect 6240 3512 6320 3608
rect 6240 3448 6248 3512
rect 6312 3448 6320 3512
rect 6240 3352 6320 3448
rect 6240 3288 6248 3352
rect 6312 3288 6320 3352
rect 6240 3192 6320 3288
rect 6240 3128 6248 3192
rect 6312 3128 6320 3192
rect 6240 2872 6320 3128
rect 6240 2808 6248 2872
rect 6312 2808 6320 2872
rect 6240 2712 6320 2808
rect 6240 2648 6248 2712
rect 6312 2648 6320 2712
rect 6240 2552 6320 2648
rect 6240 2488 6248 2552
rect 6312 2488 6320 2552
rect 6240 2232 6320 2488
rect 6240 2168 6248 2232
rect 6312 2168 6320 2232
rect 6240 1912 6320 2168
rect 6240 1848 6248 1912
rect 6312 1848 6320 1912
rect 6240 1752 6320 1848
rect 6240 1688 6248 1752
rect 6312 1688 6320 1752
rect 6240 1432 6320 1688
rect 6240 1368 6248 1432
rect 6312 1368 6320 1432
rect 6240 1112 6320 1368
rect 6240 1048 6248 1112
rect 6312 1048 6320 1112
rect 6240 952 6320 1048
rect 6240 888 6248 952
rect 6312 888 6320 952
rect 6240 792 6320 888
rect 6240 728 6248 792
rect 6312 728 6320 792
rect 6240 472 6320 728
rect 6240 408 6248 472
rect 6312 408 6320 472
rect 6240 312 6320 408
rect 6240 248 6248 312
rect 6312 248 6320 312
rect 6240 152 6320 248
rect 6240 88 6248 152
rect 6312 88 6320 152
rect 6240 -8 6320 88
rect 6240 -72 6248 -8
rect 6312 -72 6320 -8
rect 6240 -328 6320 -72
rect 6240 -392 6248 -328
rect 6312 -392 6320 -328
rect 6240 -648 6320 -392
rect 6240 -712 6248 -648
rect 6312 -712 6320 -648
rect 6240 -720 6320 -712
rect 6400 4148 6480 4320
rect 6400 4092 6412 4148
rect 6468 4092 6480 4148
rect 6400 -492 6480 4092
rect 6400 -548 6412 -492
rect 6468 -548 6480 -492
rect 6400 -720 6480 -548
rect 6560 4312 6640 4320
rect 6560 4248 6568 4312
rect 6632 4248 6640 4312
rect 6560 3992 6640 4248
rect 6560 3928 6568 3992
rect 6632 3928 6640 3992
rect 6560 3672 6640 3928
rect 6560 3608 6568 3672
rect 6632 3608 6640 3672
rect 6560 3512 6640 3608
rect 6560 3448 6568 3512
rect 6632 3448 6640 3512
rect 6560 3352 6640 3448
rect 6560 3288 6568 3352
rect 6632 3288 6640 3352
rect 6560 3192 6640 3288
rect 6560 3128 6568 3192
rect 6632 3128 6640 3192
rect 6560 2872 6640 3128
rect 6560 2808 6568 2872
rect 6632 2808 6640 2872
rect 6560 2712 6640 2808
rect 6560 2648 6568 2712
rect 6632 2648 6640 2712
rect 6560 2552 6640 2648
rect 6560 2488 6568 2552
rect 6632 2488 6640 2552
rect 6560 2232 6640 2488
rect 6560 2168 6568 2232
rect 6632 2168 6640 2232
rect 6560 1912 6640 2168
rect 6560 1848 6568 1912
rect 6632 1848 6640 1912
rect 6560 1752 6640 1848
rect 6560 1688 6568 1752
rect 6632 1688 6640 1752
rect 6560 1432 6640 1688
rect 6560 1368 6568 1432
rect 6632 1368 6640 1432
rect 6560 1112 6640 1368
rect 6560 1048 6568 1112
rect 6632 1048 6640 1112
rect 6560 952 6640 1048
rect 6560 888 6568 952
rect 6632 888 6640 952
rect 6560 792 6640 888
rect 6560 728 6568 792
rect 6632 728 6640 792
rect 6560 472 6640 728
rect 6560 408 6568 472
rect 6632 408 6640 472
rect 6560 312 6640 408
rect 6560 248 6568 312
rect 6632 248 6640 312
rect 6560 152 6640 248
rect 6560 88 6568 152
rect 6632 88 6640 152
rect 6560 -8 6640 88
rect 6560 -72 6568 -8
rect 6632 -72 6640 -8
rect 6560 -328 6640 -72
rect 6560 -392 6568 -328
rect 6632 -392 6640 -328
rect 6560 -648 6640 -392
rect 6560 -712 6568 -648
rect 6632 -712 6640 -648
rect 6560 -720 6640 -712
rect 6720 3028 6800 4320
rect 6720 2972 6732 3028
rect 6788 2972 6800 3028
rect 6720 948 6800 2972
rect 6720 892 6732 948
rect 6788 892 6800 948
rect 6720 -720 6800 892
rect 6880 4312 6960 4320
rect 6880 4248 6888 4312
rect 6952 4248 6960 4312
rect 6880 3992 6960 4248
rect 6880 3928 6888 3992
rect 6952 3928 6960 3992
rect 6880 3672 6960 3928
rect 6880 3608 6888 3672
rect 6952 3608 6960 3672
rect 6880 3352 6960 3608
rect 6880 3288 6888 3352
rect 6952 3288 6960 3352
rect 6880 3192 6960 3288
rect 6880 3128 6888 3192
rect 6952 3128 6960 3192
rect 6880 2872 6960 3128
rect 6880 2808 6888 2872
rect 6952 2808 6960 2872
rect 6880 2552 6960 2808
rect 6880 2488 6888 2552
rect 6952 2488 6960 2552
rect 6880 2232 6960 2488
rect 6880 2168 6888 2232
rect 6952 2168 6960 2232
rect 6880 1912 6960 2168
rect 6880 1848 6888 1912
rect 6952 1848 6960 1912
rect 6880 1752 6960 1848
rect 6880 1688 6888 1752
rect 6952 1688 6960 1752
rect 6880 1432 6960 1688
rect 6880 1368 6888 1432
rect 6952 1368 6960 1432
rect 6880 1112 6960 1368
rect 6880 1048 6888 1112
rect 6952 1048 6960 1112
rect 6880 792 6960 1048
rect 6880 728 6888 792
rect 6952 728 6960 792
rect 6880 472 6960 728
rect 6880 408 6888 472
rect 6952 408 6960 472
rect 6880 312 6960 408
rect 6880 248 6888 312
rect 6952 248 6960 312
rect 6880 -8 6960 248
rect 6880 -72 6888 -8
rect 6952 -72 6960 -8
rect 6880 -328 6960 -72
rect 6880 -392 6888 -328
rect 6952 -392 6960 -328
rect 6880 -648 6960 -392
rect 6880 -712 6888 -648
rect 6952 -712 6960 -648
rect 6880 -720 6960 -712
rect 7040 2068 7120 4320
rect 7040 2012 7052 2068
rect 7108 2012 7120 2068
rect 7040 148 7120 2012
rect 7040 92 7052 148
rect 7108 92 7120 148
rect 7040 -720 7120 92
rect 7200 4312 7280 4320
rect 7200 4248 7208 4312
rect 7272 4248 7280 4312
rect 7200 3992 7280 4248
rect 7200 3928 7208 3992
rect 7272 3928 7280 3992
rect 7200 3672 7280 3928
rect 7200 3608 7208 3672
rect 7272 3608 7280 3672
rect 7200 3352 7280 3608
rect 7200 3288 7208 3352
rect 7272 3288 7280 3352
rect 7200 3192 7280 3288
rect 7200 3128 7208 3192
rect 7272 3128 7280 3192
rect 7200 2872 7280 3128
rect 7200 2808 7208 2872
rect 7272 2808 7280 2872
rect 7200 2552 7280 2808
rect 7200 2488 7208 2552
rect 7272 2488 7280 2552
rect 7200 2232 7280 2488
rect 7200 2168 7208 2232
rect 7272 2168 7280 2232
rect 7200 1912 7280 2168
rect 7200 1848 7208 1912
rect 7272 1848 7280 1912
rect 7200 1752 7280 1848
rect 7200 1688 7208 1752
rect 7272 1688 7280 1752
rect 7200 1432 7280 1688
rect 7200 1368 7208 1432
rect 7272 1368 7280 1432
rect 7200 1112 7280 1368
rect 7200 1048 7208 1112
rect 7272 1048 7280 1112
rect 7200 792 7280 1048
rect 7200 728 7208 792
rect 7272 728 7280 792
rect 7200 472 7280 728
rect 7200 408 7208 472
rect 7272 408 7280 472
rect 7200 312 7280 408
rect 7200 248 7208 312
rect 7272 248 7280 312
rect 7200 -8 7280 248
rect 7200 -72 7208 -8
rect 7272 -72 7280 -8
rect 7200 -328 7280 -72
rect 7200 -392 7208 -328
rect 7272 -392 7280 -328
rect 7200 -648 7280 -392
rect 7200 -712 7208 -648
rect 7272 -712 7280 -648
rect 7200 -720 7280 -712
rect 7360 2708 7440 4320
rect 7360 2652 7372 2708
rect 7428 2652 7440 2708
rect 7360 628 7440 2652
rect 7360 572 7372 628
rect 7428 572 7440 628
rect 7360 -720 7440 572
rect 7520 4312 7600 4320
rect 7520 4248 7528 4312
rect 7592 4248 7600 4312
rect 7520 3992 7600 4248
rect 7520 3928 7528 3992
rect 7592 3928 7600 3992
rect 7520 3672 7600 3928
rect 7520 3608 7528 3672
rect 7592 3608 7600 3672
rect 7520 3352 7600 3608
rect 7520 3288 7528 3352
rect 7592 3288 7600 3352
rect 7520 3192 7600 3288
rect 7520 3128 7528 3192
rect 7592 3128 7600 3192
rect 7520 2872 7600 3128
rect 7520 2808 7528 2872
rect 7592 2808 7600 2872
rect 7520 2552 7600 2808
rect 7520 2488 7528 2552
rect 7592 2488 7600 2552
rect 7520 2232 7600 2488
rect 7520 2168 7528 2232
rect 7592 2168 7600 2232
rect 7520 1912 7600 2168
rect 7520 1848 7528 1912
rect 7592 1848 7600 1912
rect 7520 1752 7600 1848
rect 7520 1688 7528 1752
rect 7592 1688 7600 1752
rect 7520 1432 7600 1688
rect 7520 1368 7528 1432
rect 7592 1368 7600 1432
rect 7520 1112 7600 1368
rect 7520 1048 7528 1112
rect 7592 1048 7600 1112
rect 7520 792 7600 1048
rect 7520 728 7528 792
rect 7592 728 7600 792
rect 7520 472 7600 728
rect 7520 408 7528 472
rect 7592 408 7600 472
rect 7520 312 7600 408
rect 7520 248 7528 312
rect 7592 248 7600 312
rect 7520 -8 7600 248
rect 7520 -72 7528 -8
rect 7592 -72 7600 -8
rect 7520 -328 7600 -72
rect 7520 -392 7528 -328
rect 7592 -392 7600 -328
rect 7520 -648 7600 -392
rect 7520 -712 7528 -648
rect 7592 -712 7600 -648
rect 7520 -720 7600 -712
rect 7680 3508 7760 4320
rect 7680 3452 7692 3508
rect 7748 3452 7760 3508
rect 7680 1588 7760 3452
rect 7680 1532 7692 1588
rect 7748 1532 7760 1588
rect 7680 -720 7760 1532
rect 7840 4312 7920 4320
rect 7840 4248 7848 4312
rect 7912 4248 7920 4312
rect 7840 3992 7920 4248
rect 7840 3928 7848 3992
rect 7912 3928 7920 3992
rect 7840 3672 7920 3928
rect 7840 3608 7848 3672
rect 7912 3608 7920 3672
rect 7840 3352 7920 3608
rect 7840 3288 7848 3352
rect 7912 3288 7920 3352
rect 7840 3192 7920 3288
rect 7840 3128 7848 3192
rect 7912 3128 7920 3192
rect 7840 2872 7920 3128
rect 7840 2808 7848 2872
rect 7912 2808 7920 2872
rect 7840 2552 7920 2808
rect 7840 2488 7848 2552
rect 7912 2488 7920 2552
rect 7840 2232 7920 2488
rect 7840 2168 7848 2232
rect 7912 2168 7920 2232
rect 7840 1912 7920 2168
rect 7840 1848 7848 1912
rect 7912 1848 7920 1912
rect 7840 1752 7920 1848
rect 7840 1688 7848 1752
rect 7912 1688 7920 1752
rect 7840 1432 7920 1688
rect 12720 1832 12960 1920
rect 12720 1768 12808 1832
rect 12872 1768 12960 1832
rect 12720 1680 12960 1768
rect 7840 1368 7848 1432
rect 7912 1368 7920 1432
rect 7840 1112 7920 1368
rect 7840 1048 7848 1112
rect 7912 1048 7920 1112
rect 7840 792 7920 1048
rect 7840 728 7848 792
rect 7912 728 7920 792
rect 7840 472 7920 728
rect 7840 408 7848 472
rect 7912 408 7920 472
rect 7840 312 7920 408
rect 7840 248 7848 312
rect 7912 248 7920 312
rect 7840 -8 7920 248
rect 7840 -72 7848 -8
rect 7912 -72 7920 -8
rect 7840 -328 7920 -72
rect 7840 -392 7848 -328
rect 7912 -392 7920 -328
rect 7840 -648 7920 -392
rect 7840 -712 7848 -648
rect 7912 -712 7920 -648
rect 7840 -720 7920 -712
<< via3 >>
rect 4648 4308 4712 4312
rect 4648 4252 4652 4308
rect 4652 4252 4708 4308
rect 4708 4252 4712 4308
rect 4648 4248 4712 4252
rect 4648 3988 4712 3992
rect 4648 3932 4652 3988
rect 4652 3932 4708 3988
rect 4708 3932 4712 3988
rect 4648 3928 4712 3932
rect 4648 3668 4712 3672
rect 4648 3612 4652 3668
rect 4652 3612 4708 3668
rect 4708 3612 4712 3668
rect 4648 3608 4712 3612
rect 4648 3348 4712 3352
rect 4648 3292 4652 3348
rect 4652 3292 4708 3348
rect 4708 3292 4712 3348
rect 4648 3288 4712 3292
rect 4648 3188 4712 3192
rect 4648 3132 4652 3188
rect 4652 3132 4708 3188
rect 4708 3132 4712 3188
rect 4648 3128 4712 3132
rect 4648 2868 4712 2872
rect 4648 2812 4652 2868
rect 4652 2812 4708 2868
rect 4708 2812 4712 2868
rect 4648 2808 4712 2812
rect 4648 2548 4712 2552
rect 4648 2492 4652 2548
rect 4652 2492 4708 2548
rect 4708 2492 4712 2548
rect 4648 2488 4712 2492
rect 4648 2228 4712 2232
rect 4648 2172 4652 2228
rect 4652 2172 4708 2228
rect 4708 2172 4712 2228
rect 4648 2168 4712 2172
rect -312 1828 -248 1832
rect -312 1772 -308 1828
rect -308 1772 -252 1828
rect -252 1772 -248 1828
rect -312 1768 -248 1772
rect 4648 1908 4712 1912
rect 4648 1852 4652 1908
rect 4652 1852 4708 1908
rect 4708 1852 4712 1908
rect 4648 1848 4712 1852
rect 4648 1748 4712 1752
rect 4648 1692 4652 1748
rect 4652 1692 4708 1748
rect 4708 1692 4712 1748
rect 4648 1688 4712 1692
rect 4648 1428 4712 1432
rect 4648 1372 4652 1428
rect 4652 1372 4708 1428
rect 4708 1372 4712 1428
rect 4648 1368 4712 1372
rect 4648 1108 4712 1112
rect 4648 1052 4652 1108
rect 4652 1052 4708 1108
rect 4708 1052 4712 1108
rect 4648 1048 4712 1052
rect 4648 788 4712 792
rect 4648 732 4652 788
rect 4652 732 4708 788
rect 4708 732 4712 788
rect 4648 728 4712 732
rect 4648 468 4712 472
rect 4648 412 4652 468
rect 4652 412 4708 468
rect 4708 412 4712 468
rect 4648 408 4712 412
rect 4648 308 4712 312
rect 4648 252 4652 308
rect 4652 252 4708 308
rect 4708 252 4712 308
rect 4648 248 4712 252
rect 4648 -12 4712 -8
rect 4648 -68 4652 -12
rect 4652 -68 4708 -12
rect 4708 -68 4712 -12
rect 4648 -72 4712 -68
rect 4648 -332 4712 -328
rect 4648 -388 4652 -332
rect 4652 -388 4708 -332
rect 4708 -388 4712 -332
rect 4648 -392 4712 -388
rect 4648 -652 4712 -648
rect 4648 -708 4652 -652
rect 4652 -708 4708 -652
rect 4708 -708 4712 -652
rect 4648 -712 4712 -708
rect 4968 4308 5032 4312
rect 4968 4252 4972 4308
rect 4972 4252 5028 4308
rect 5028 4252 5032 4308
rect 4968 4248 5032 4252
rect 4968 3988 5032 3992
rect 4968 3932 4972 3988
rect 4972 3932 5028 3988
rect 5028 3932 5032 3988
rect 4968 3928 5032 3932
rect 4968 3668 5032 3672
rect 4968 3612 4972 3668
rect 4972 3612 5028 3668
rect 5028 3612 5032 3668
rect 4968 3608 5032 3612
rect 4968 3348 5032 3352
rect 4968 3292 4972 3348
rect 4972 3292 5028 3348
rect 5028 3292 5032 3348
rect 4968 3288 5032 3292
rect 4968 3188 5032 3192
rect 4968 3132 4972 3188
rect 4972 3132 5028 3188
rect 5028 3132 5032 3188
rect 4968 3128 5032 3132
rect 4968 2868 5032 2872
rect 4968 2812 4972 2868
rect 4972 2812 5028 2868
rect 5028 2812 5032 2868
rect 4968 2808 5032 2812
rect 4968 2548 5032 2552
rect 4968 2492 4972 2548
rect 4972 2492 5028 2548
rect 5028 2492 5032 2548
rect 4968 2488 5032 2492
rect 4968 2228 5032 2232
rect 4968 2172 4972 2228
rect 4972 2172 5028 2228
rect 5028 2172 5032 2228
rect 4968 2168 5032 2172
rect 4968 1908 5032 1912
rect 4968 1852 4972 1908
rect 4972 1852 5028 1908
rect 5028 1852 5032 1908
rect 4968 1848 5032 1852
rect 4968 1748 5032 1752
rect 4968 1692 4972 1748
rect 4972 1692 5028 1748
rect 5028 1692 5032 1748
rect 4968 1688 5032 1692
rect 4968 1428 5032 1432
rect 4968 1372 4972 1428
rect 4972 1372 5028 1428
rect 5028 1372 5032 1428
rect 4968 1368 5032 1372
rect 4968 1108 5032 1112
rect 4968 1052 4972 1108
rect 4972 1052 5028 1108
rect 5028 1052 5032 1108
rect 4968 1048 5032 1052
rect 4968 788 5032 792
rect 4968 732 4972 788
rect 4972 732 5028 788
rect 5028 732 5032 788
rect 4968 728 5032 732
rect 4968 468 5032 472
rect 4968 412 4972 468
rect 4972 412 5028 468
rect 5028 412 5032 468
rect 4968 408 5032 412
rect 4968 308 5032 312
rect 4968 252 4972 308
rect 4972 252 5028 308
rect 5028 252 5032 308
rect 4968 248 5032 252
rect 4968 -12 5032 -8
rect 4968 -68 4972 -12
rect 4972 -68 5028 -12
rect 5028 -68 5032 -12
rect 4968 -72 5032 -68
rect 4968 -332 5032 -328
rect 4968 -388 4972 -332
rect 4972 -388 5028 -332
rect 5028 -388 5032 -332
rect 4968 -392 5032 -388
rect 4968 -652 5032 -648
rect 4968 -708 4972 -652
rect 4972 -708 5028 -652
rect 5028 -708 5032 -652
rect 4968 -712 5032 -708
rect 5288 4308 5352 4312
rect 5288 4252 5292 4308
rect 5292 4252 5348 4308
rect 5348 4252 5352 4308
rect 5288 4248 5352 4252
rect 5288 3988 5352 3992
rect 5288 3932 5292 3988
rect 5292 3932 5348 3988
rect 5348 3932 5352 3988
rect 5288 3928 5352 3932
rect 5288 3668 5352 3672
rect 5288 3612 5292 3668
rect 5292 3612 5348 3668
rect 5348 3612 5352 3668
rect 5288 3608 5352 3612
rect 5288 3348 5352 3352
rect 5288 3292 5292 3348
rect 5292 3292 5348 3348
rect 5348 3292 5352 3348
rect 5288 3288 5352 3292
rect 5288 3188 5352 3192
rect 5288 3132 5292 3188
rect 5292 3132 5348 3188
rect 5348 3132 5352 3188
rect 5288 3128 5352 3132
rect 5288 2868 5352 2872
rect 5288 2812 5292 2868
rect 5292 2812 5348 2868
rect 5348 2812 5352 2868
rect 5288 2808 5352 2812
rect 5288 2548 5352 2552
rect 5288 2492 5292 2548
rect 5292 2492 5348 2548
rect 5348 2492 5352 2548
rect 5288 2488 5352 2492
rect 5288 2228 5352 2232
rect 5288 2172 5292 2228
rect 5292 2172 5348 2228
rect 5348 2172 5352 2228
rect 5288 2168 5352 2172
rect 5288 1908 5352 1912
rect 5288 1852 5292 1908
rect 5292 1852 5348 1908
rect 5348 1852 5352 1908
rect 5288 1848 5352 1852
rect 5288 1748 5352 1752
rect 5288 1692 5292 1748
rect 5292 1692 5348 1748
rect 5348 1692 5352 1748
rect 5288 1688 5352 1692
rect 5288 1428 5352 1432
rect 5288 1372 5292 1428
rect 5292 1372 5348 1428
rect 5348 1372 5352 1428
rect 5288 1368 5352 1372
rect 5288 1108 5352 1112
rect 5288 1052 5292 1108
rect 5292 1052 5348 1108
rect 5348 1052 5352 1108
rect 5288 1048 5352 1052
rect 5288 788 5352 792
rect 5288 732 5292 788
rect 5292 732 5348 788
rect 5348 732 5352 788
rect 5288 728 5352 732
rect 5288 468 5352 472
rect 5288 412 5292 468
rect 5292 412 5348 468
rect 5348 412 5352 468
rect 5288 408 5352 412
rect 5288 308 5352 312
rect 5288 252 5292 308
rect 5292 252 5348 308
rect 5348 252 5352 308
rect 5288 248 5352 252
rect 5288 -12 5352 -8
rect 5288 -68 5292 -12
rect 5292 -68 5348 -12
rect 5348 -68 5352 -12
rect 5288 -72 5352 -68
rect 5288 -332 5352 -328
rect 5288 -388 5292 -332
rect 5292 -388 5348 -332
rect 5348 -388 5352 -332
rect 5288 -392 5352 -388
rect 5288 -652 5352 -648
rect 5288 -708 5292 -652
rect 5292 -708 5348 -652
rect 5348 -708 5352 -652
rect 5288 -712 5352 -708
rect 5608 4308 5672 4312
rect 5608 4252 5612 4308
rect 5612 4252 5668 4308
rect 5668 4252 5672 4308
rect 5608 4248 5672 4252
rect 5608 3988 5672 3992
rect 5608 3932 5612 3988
rect 5612 3932 5668 3988
rect 5668 3932 5672 3988
rect 5608 3928 5672 3932
rect 5608 3668 5672 3672
rect 5608 3612 5612 3668
rect 5612 3612 5668 3668
rect 5668 3612 5672 3668
rect 5608 3608 5672 3612
rect 5608 3348 5672 3352
rect 5608 3292 5612 3348
rect 5612 3292 5668 3348
rect 5668 3292 5672 3348
rect 5608 3288 5672 3292
rect 5608 3188 5672 3192
rect 5608 3132 5612 3188
rect 5612 3132 5668 3188
rect 5668 3132 5672 3188
rect 5608 3128 5672 3132
rect 5608 2868 5672 2872
rect 5608 2812 5612 2868
rect 5612 2812 5668 2868
rect 5668 2812 5672 2868
rect 5608 2808 5672 2812
rect 5608 2548 5672 2552
rect 5608 2492 5612 2548
rect 5612 2492 5668 2548
rect 5668 2492 5672 2548
rect 5608 2488 5672 2492
rect 5608 2228 5672 2232
rect 5608 2172 5612 2228
rect 5612 2172 5668 2228
rect 5668 2172 5672 2228
rect 5608 2168 5672 2172
rect 5608 1908 5672 1912
rect 5608 1852 5612 1908
rect 5612 1852 5668 1908
rect 5668 1852 5672 1908
rect 5608 1848 5672 1852
rect 5608 1748 5672 1752
rect 5608 1692 5612 1748
rect 5612 1692 5668 1748
rect 5668 1692 5672 1748
rect 5608 1688 5672 1692
rect 5608 1428 5672 1432
rect 5608 1372 5612 1428
rect 5612 1372 5668 1428
rect 5668 1372 5672 1428
rect 5608 1368 5672 1372
rect 5608 1108 5672 1112
rect 5608 1052 5612 1108
rect 5612 1052 5668 1108
rect 5668 1052 5672 1108
rect 5608 1048 5672 1052
rect 5608 788 5672 792
rect 5608 732 5612 788
rect 5612 732 5668 788
rect 5668 732 5672 788
rect 5608 728 5672 732
rect 5608 468 5672 472
rect 5608 412 5612 468
rect 5612 412 5668 468
rect 5668 412 5672 468
rect 5608 408 5672 412
rect 5608 308 5672 312
rect 5608 252 5612 308
rect 5612 252 5668 308
rect 5668 252 5672 308
rect 5608 248 5672 252
rect 5608 -12 5672 -8
rect 5608 -68 5612 -12
rect 5612 -68 5668 -12
rect 5668 -68 5672 -12
rect 5608 -72 5672 -68
rect 5608 -332 5672 -328
rect 5608 -388 5612 -332
rect 5612 -388 5668 -332
rect 5668 -388 5672 -332
rect 5608 -392 5672 -388
rect 5608 -652 5672 -648
rect 5608 -708 5612 -652
rect 5612 -708 5668 -652
rect 5668 -708 5672 -652
rect 5608 -712 5672 -708
rect 5928 4308 5992 4312
rect 5928 4252 5932 4308
rect 5932 4252 5988 4308
rect 5988 4252 5992 4308
rect 5928 4248 5992 4252
rect 5928 3988 5992 3992
rect 5928 3932 5932 3988
rect 5932 3932 5988 3988
rect 5988 3932 5992 3988
rect 5928 3928 5992 3932
rect 5928 3668 5992 3672
rect 5928 3612 5932 3668
rect 5932 3612 5988 3668
rect 5988 3612 5992 3668
rect 5928 3608 5992 3612
rect 5928 3508 5992 3512
rect 5928 3452 5932 3508
rect 5932 3452 5988 3508
rect 5988 3452 5992 3508
rect 5928 3448 5992 3452
rect 5928 3348 5992 3352
rect 5928 3292 5932 3348
rect 5932 3292 5988 3348
rect 5988 3292 5992 3348
rect 5928 3288 5992 3292
rect 5928 3188 5992 3192
rect 5928 3132 5932 3188
rect 5932 3132 5988 3188
rect 5988 3132 5992 3188
rect 5928 3128 5992 3132
rect 5928 2868 5992 2872
rect 5928 2812 5932 2868
rect 5932 2812 5988 2868
rect 5988 2812 5992 2868
rect 5928 2808 5992 2812
rect 5928 2708 5992 2712
rect 5928 2652 5932 2708
rect 5932 2652 5988 2708
rect 5988 2652 5992 2708
rect 5928 2648 5992 2652
rect 5928 2548 5992 2552
rect 5928 2492 5932 2548
rect 5932 2492 5988 2548
rect 5988 2492 5992 2548
rect 5928 2488 5992 2492
rect 5928 2228 5992 2232
rect 5928 2172 5932 2228
rect 5932 2172 5988 2228
rect 5988 2172 5992 2228
rect 5928 2168 5992 2172
rect 5928 1908 5992 1912
rect 5928 1852 5932 1908
rect 5932 1852 5988 1908
rect 5988 1852 5992 1908
rect 5928 1848 5992 1852
rect 5928 1748 5992 1752
rect 5928 1692 5932 1748
rect 5932 1692 5988 1748
rect 5988 1692 5992 1748
rect 5928 1688 5992 1692
rect 5928 1428 5992 1432
rect 5928 1372 5932 1428
rect 5932 1372 5988 1428
rect 5988 1372 5992 1428
rect 5928 1368 5992 1372
rect 5928 1108 5992 1112
rect 5928 1052 5932 1108
rect 5932 1052 5988 1108
rect 5988 1052 5992 1108
rect 5928 1048 5992 1052
rect 5928 948 5992 952
rect 5928 892 5932 948
rect 5932 892 5988 948
rect 5988 892 5992 948
rect 5928 888 5992 892
rect 5928 788 5992 792
rect 5928 732 5932 788
rect 5932 732 5988 788
rect 5988 732 5992 788
rect 5928 728 5992 732
rect 5928 468 5992 472
rect 5928 412 5932 468
rect 5932 412 5988 468
rect 5988 412 5992 468
rect 5928 408 5992 412
rect 5928 308 5992 312
rect 5928 252 5932 308
rect 5932 252 5988 308
rect 5988 252 5992 308
rect 5928 248 5992 252
rect 5928 148 5992 152
rect 5928 92 5932 148
rect 5932 92 5988 148
rect 5988 92 5992 148
rect 5928 88 5992 92
rect 5928 -12 5992 -8
rect 5928 -68 5932 -12
rect 5932 -68 5988 -12
rect 5988 -68 5992 -12
rect 5928 -72 5992 -68
rect 5928 -332 5992 -328
rect 5928 -388 5932 -332
rect 5932 -388 5988 -332
rect 5988 -388 5992 -332
rect 5928 -392 5992 -388
rect 5928 -652 5992 -648
rect 5928 -708 5932 -652
rect 5932 -708 5988 -652
rect 5988 -708 5992 -652
rect 5928 -712 5992 -708
rect 6248 4308 6312 4312
rect 6248 4252 6252 4308
rect 6252 4252 6308 4308
rect 6308 4252 6312 4308
rect 6248 4248 6312 4252
rect 6248 3988 6312 3992
rect 6248 3932 6252 3988
rect 6252 3932 6308 3988
rect 6308 3932 6312 3988
rect 6248 3928 6312 3932
rect 6248 3668 6312 3672
rect 6248 3612 6252 3668
rect 6252 3612 6308 3668
rect 6308 3612 6312 3668
rect 6248 3608 6312 3612
rect 6248 3508 6312 3512
rect 6248 3452 6252 3508
rect 6252 3452 6308 3508
rect 6308 3452 6312 3508
rect 6248 3448 6312 3452
rect 6248 3348 6312 3352
rect 6248 3292 6252 3348
rect 6252 3292 6308 3348
rect 6308 3292 6312 3348
rect 6248 3288 6312 3292
rect 6248 3188 6312 3192
rect 6248 3132 6252 3188
rect 6252 3132 6308 3188
rect 6308 3132 6312 3188
rect 6248 3128 6312 3132
rect 6248 2868 6312 2872
rect 6248 2812 6252 2868
rect 6252 2812 6308 2868
rect 6308 2812 6312 2868
rect 6248 2808 6312 2812
rect 6248 2708 6312 2712
rect 6248 2652 6252 2708
rect 6252 2652 6308 2708
rect 6308 2652 6312 2708
rect 6248 2648 6312 2652
rect 6248 2548 6312 2552
rect 6248 2492 6252 2548
rect 6252 2492 6308 2548
rect 6308 2492 6312 2548
rect 6248 2488 6312 2492
rect 6248 2228 6312 2232
rect 6248 2172 6252 2228
rect 6252 2172 6308 2228
rect 6308 2172 6312 2228
rect 6248 2168 6312 2172
rect 6248 1908 6312 1912
rect 6248 1852 6252 1908
rect 6252 1852 6308 1908
rect 6308 1852 6312 1908
rect 6248 1848 6312 1852
rect 6248 1748 6312 1752
rect 6248 1692 6252 1748
rect 6252 1692 6308 1748
rect 6308 1692 6312 1748
rect 6248 1688 6312 1692
rect 6248 1428 6312 1432
rect 6248 1372 6252 1428
rect 6252 1372 6308 1428
rect 6308 1372 6312 1428
rect 6248 1368 6312 1372
rect 6248 1108 6312 1112
rect 6248 1052 6252 1108
rect 6252 1052 6308 1108
rect 6308 1052 6312 1108
rect 6248 1048 6312 1052
rect 6248 948 6312 952
rect 6248 892 6252 948
rect 6252 892 6308 948
rect 6308 892 6312 948
rect 6248 888 6312 892
rect 6248 788 6312 792
rect 6248 732 6252 788
rect 6252 732 6308 788
rect 6308 732 6312 788
rect 6248 728 6312 732
rect 6248 468 6312 472
rect 6248 412 6252 468
rect 6252 412 6308 468
rect 6308 412 6312 468
rect 6248 408 6312 412
rect 6248 308 6312 312
rect 6248 252 6252 308
rect 6252 252 6308 308
rect 6308 252 6312 308
rect 6248 248 6312 252
rect 6248 148 6312 152
rect 6248 92 6252 148
rect 6252 92 6308 148
rect 6308 92 6312 148
rect 6248 88 6312 92
rect 6248 -12 6312 -8
rect 6248 -68 6252 -12
rect 6252 -68 6308 -12
rect 6308 -68 6312 -12
rect 6248 -72 6312 -68
rect 6248 -332 6312 -328
rect 6248 -388 6252 -332
rect 6252 -388 6308 -332
rect 6308 -388 6312 -332
rect 6248 -392 6312 -388
rect 6248 -652 6312 -648
rect 6248 -708 6252 -652
rect 6252 -708 6308 -652
rect 6308 -708 6312 -652
rect 6248 -712 6312 -708
rect 6568 4308 6632 4312
rect 6568 4252 6572 4308
rect 6572 4252 6628 4308
rect 6628 4252 6632 4308
rect 6568 4248 6632 4252
rect 6568 3988 6632 3992
rect 6568 3932 6572 3988
rect 6572 3932 6628 3988
rect 6628 3932 6632 3988
rect 6568 3928 6632 3932
rect 6568 3668 6632 3672
rect 6568 3612 6572 3668
rect 6572 3612 6628 3668
rect 6628 3612 6632 3668
rect 6568 3608 6632 3612
rect 6568 3508 6632 3512
rect 6568 3452 6572 3508
rect 6572 3452 6628 3508
rect 6628 3452 6632 3508
rect 6568 3448 6632 3452
rect 6568 3348 6632 3352
rect 6568 3292 6572 3348
rect 6572 3292 6628 3348
rect 6628 3292 6632 3348
rect 6568 3288 6632 3292
rect 6568 3188 6632 3192
rect 6568 3132 6572 3188
rect 6572 3132 6628 3188
rect 6628 3132 6632 3188
rect 6568 3128 6632 3132
rect 6568 2868 6632 2872
rect 6568 2812 6572 2868
rect 6572 2812 6628 2868
rect 6628 2812 6632 2868
rect 6568 2808 6632 2812
rect 6568 2708 6632 2712
rect 6568 2652 6572 2708
rect 6572 2652 6628 2708
rect 6628 2652 6632 2708
rect 6568 2648 6632 2652
rect 6568 2548 6632 2552
rect 6568 2492 6572 2548
rect 6572 2492 6628 2548
rect 6628 2492 6632 2548
rect 6568 2488 6632 2492
rect 6568 2228 6632 2232
rect 6568 2172 6572 2228
rect 6572 2172 6628 2228
rect 6628 2172 6632 2228
rect 6568 2168 6632 2172
rect 6568 1908 6632 1912
rect 6568 1852 6572 1908
rect 6572 1852 6628 1908
rect 6628 1852 6632 1908
rect 6568 1848 6632 1852
rect 6568 1748 6632 1752
rect 6568 1692 6572 1748
rect 6572 1692 6628 1748
rect 6628 1692 6632 1748
rect 6568 1688 6632 1692
rect 6568 1428 6632 1432
rect 6568 1372 6572 1428
rect 6572 1372 6628 1428
rect 6628 1372 6632 1428
rect 6568 1368 6632 1372
rect 6568 1108 6632 1112
rect 6568 1052 6572 1108
rect 6572 1052 6628 1108
rect 6628 1052 6632 1108
rect 6568 1048 6632 1052
rect 6568 948 6632 952
rect 6568 892 6572 948
rect 6572 892 6628 948
rect 6628 892 6632 948
rect 6568 888 6632 892
rect 6568 788 6632 792
rect 6568 732 6572 788
rect 6572 732 6628 788
rect 6628 732 6632 788
rect 6568 728 6632 732
rect 6568 468 6632 472
rect 6568 412 6572 468
rect 6572 412 6628 468
rect 6628 412 6632 468
rect 6568 408 6632 412
rect 6568 308 6632 312
rect 6568 252 6572 308
rect 6572 252 6628 308
rect 6628 252 6632 308
rect 6568 248 6632 252
rect 6568 148 6632 152
rect 6568 92 6572 148
rect 6572 92 6628 148
rect 6628 92 6632 148
rect 6568 88 6632 92
rect 6568 -12 6632 -8
rect 6568 -68 6572 -12
rect 6572 -68 6628 -12
rect 6628 -68 6632 -12
rect 6568 -72 6632 -68
rect 6568 -332 6632 -328
rect 6568 -388 6572 -332
rect 6572 -388 6628 -332
rect 6628 -388 6632 -332
rect 6568 -392 6632 -388
rect 6568 -652 6632 -648
rect 6568 -708 6572 -652
rect 6572 -708 6628 -652
rect 6628 -708 6632 -652
rect 6568 -712 6632 -708
rect 6888 4308 6952 4312
rect 6888 4252 6892 4308
rect 6892 4252 6948 4308
rect 6948 4252 6952 4308
rect 6888 4248 6952 4252
rect 6888 3988 6952 3992
rect 6888 3932 6892 3988
rect 6892 3932 6948 3988
rect 6948 3932 6952 3988
rect 6888 3928 6952 3932
rect 6888 3668 6952 3672
rect 6888 3612 6892 3668
rect 6892 3612 6948 3668
rect 6948 3612 6952 3668
rect 6888 3608 6952 3612
rect 6888 3348 6952 3352
rect 6888 3292 6892 3348
rect 6892 3292 6948 3348
rect 6948 3292 6952 3348
rect 6888 3288 6952 3292
rect 6888 3188 6952 3192
rect 6888 3132 6892 3188
rect 6892 3132 6948 3188
rect 6948 3132 6952 3188
rect 6888 3128 6952 3132
rect 6888 2868 6952 2872
rect 6888 2812 6892 2868
rect 6892 2812 6948 2868
rect 6948 2812 6952 2868
rect 6888 2808 6952 2812
rect 6888 2548 6952 2552
rect 6888 2492 6892 2548
rect 6892 2492 6948 2548
rect 6948 2492 6952 2548
rect 6888 2488 6952 2492
rect 6888 2228 6952 2232
rect 6888 2172 6892 2228
rect 6892 2172 6948 2228
rect 6948 2172 6952 2228
rect 6888 2168 6952 2172
rect 6888 1908 6952 1912
rect 6888 1852 6892 1908
rect 6892 1852 6948 1908
rect 6948 1852 6952 1908
rect 6888 1848 6952 1852
rect 6888 1748 6952 1752
rect 6888 1692 6892 1748
rect 6892 1692 6948 1748
rect 6948 1692 6952 1748
rect 6888 1688 6952 1692
rect 6888 1428 6952 1432
rect 6888 1372 6892 1428
rect 6892 1372 6948 1428
rect 6948 1372 6952 1428
rect 6888 1368 6952 1372
rect 6888 1108 6952 1112
rect 6888 1052 6892 1108
rect 6892 1052 6948 1108
rect 6948 1052 6952 1108
rect 6888 1048 6952 1052
rect 6888 788 6952 792
rect 6888 732 6892 788
rect 6892 732 6948 788
rect 6948 732 6952 788
rect 6888 728 6952 732
rect 6888 468 6952 472
rect 6888 412 6892 468
rect 6892 412 6948 468
rect 6948 412 6952 468
rect 6888 408 6952 412
rect 6888 308 6952 312
rect 6888 252 6892 308
rect 6892 252 6948 308
rect 6948 252 6952 308
rect 6888 248 6952 252
rect 6888 -12 6952 -8
rect 6888 -68 6892 -12
rect 6892 -68 6948 -12
rect 6948 -68 6952 -12
rect 6888 -72 6952 -68
rect 6888 -332 6952 -328
rect 6888 -388 6892 -332
rect 6892 -388 6948 -332
rect 6948 -388 6952 -332
rect 6888 -392 6952 -388
rect 6888 -652 6952 -648
rect 6888 -708 6892 -652
rect 6892 -708 6948 -652
rect 6948 -708 6952 -652
rect 6888 -712 6952 -708
rect 7208 4308 7272 4312
rect 7208 4252 7212 4308
rect 7212 4252 7268 4308
rect 7268 4252 7272 4308
rect 7208 4248 7272 4252
rect 7208 3988 7272 3992
rect 7208 3932 7212 3988
rect 7212 3932 7268 3988
rect 7268 3932 7272 3988
rect 7208 3928 7272 3932
rect 7208 3668 7272 3672
rect 7208 3612 7212 3668
rect 7212 3612 7268 3668
rect 7268 3612 7272 3668
rect 7208 3608 7272 3612
rect 7208 3348 7272 3352
rect 7208 3292 7212 3348
rect 7212 3292 7268 3348
rect 7268 3292 7272 3348
rect 7208 3288 7272 3292
rect 7208 3188 7272 3192
rect 7208 3132 7212 3188
rect 7212 3132 7268 3188
rect 7268 3132 7272 3188
rect 7208 3128 7272 3132
rect 7208 2868 7272 2872
rect 7208 2812 7212 2868
rect 7212 2812 7268 2868
rect 7268 2812 7272 2868
rect 7208 2808 7272 2812
rect 7208 2548 7272 2552
rect 7208 2492 7212 2548
rect 7212 2492 7268 2548
rect 7268 2492 7272 2548
rect 7208 2488 7272 2492
rect 7208 2228 7272 2232
rect 7208 2172 7212 2228
rect 7212 2172 7268 2228
rect 7268 2172 7272 2228
rect 7208 2168 7272 2172
rect 7208 1908 7272 1912
rect 7208 1852 7212 1908
rect 7212 1852 7268 1908
rect 7268 1852 7272 1908
rect 7208 1848 7272 1852
rect 7208 1748 7272 1752
rect 7208 1692 7212 1748
rect 7212 1692 7268 1748
rect 7268 1692 7272 1748
rect 7208 1688 7272 1692
rect 7208 1428 7272 1432
rect 7208 1372 7212 1428
rect 7212 1372 7268 1428
rect 7268 1372 7272 1428
rect 7208 1368 7272 1372
rect 7208 1108 7272 1112
rect 7208 1052 7212 1108
rect 7212 1052 7268 1108
rect 7268 1052 7272 1108
rect 7208 1048 7272 1052
rect 7208 788 7272 792
rect 7208 732 7212 788
rect 7212 732 7268 788
rect 7268 732 7272 788
rect 7208 728 7272 732
rect 7208 468 7272 472
rect 7208 412 7212 468
rect 7212 412 7268 468
rect 7268 412 7272 468
rect 7208 408 7272 412
rect 7208 308 7272 312
rect 7208 252 7212 308
rect 7212 252 7268 308
rect 7268 252 7272 308
rect 7208 248 7272 252
rect 7208 -12 7272 -8
rect 7208 -68 7212 -12
rect 7212 -68 7268 -12
rect 7268 -68 7272 -12
rect 7208 -72 7272 -68
rect 7208 -332 7272 -328
rect 7208 -388 7212 -332
rect 7212 -388 7268 -332
rect 7268 -388 7272 -332
rect 7208 -392 7272 -388
rect 7208 -652 7272 -648
rect 7208 -708 7212 -652
rect 7212 -708 7268 -652
rect 7268 -708 7272 -652
rect 7208 -712 7272 -708
rect 7528 4308 7592 4312
rect 7528 4252 7532 4308
rect 7532 4252 7588 4308
rect 7588 4252 7592 4308
rect 7528 4248 7592 4252
rect 7528 3988 7592 3992
rect 7528 3932 7532 3988
rect 7532 3932 7588 3988
rect 7588 3932 7592 3988
rect 7528 3928 7592 3932
rect 7528 3668 7592 3672
rect 7528 3612 7532 3668
rect 7532 3612 7588 3668
rect 7588 3612 7592 3668
rect 7528 3608 7592 3612
rect 7528 3348 7592 3352
rect 7528 3292 7532 3348
rect 7532 3292 7588 3348
rect 7588 3292 7592 3348
rect 7528 3288 7592 3292
rect 7528 3188 7592 3192
rect 7528 3132 7532 3188
rect 7532 3132 7588 3188
rect 7588 3132 7592 3188
rect 7528 3128 7592 3132
rect 7528 2868 7592 2872
rect 7528 2812 7532 2868
rect 7532 2812 7588 2868
rect 7588 2812 7592 2868
rect 7528 2808 7592 2812
rect 7528 2548 7592 2552
rect 7528 2492 7532 2548
rect 7532 2492 7588 2548
rect 7588 2492 7592 2548
rect 7528 2488 7592 2492
rect 7528 2228 7592 2232
rect 7528 2172 7532 2228
rect 7532 2172 7588 2228
rect 7588 2172 7592 2228
rect 7528 2168 7592 2172
rect 7528 1908 7592 1912
rect 7528 1852 7532 1908
rect 7532 1852 7588 1908
rect 7588 1852 7592 1908
rect 7528 1848 7592 1852
rect 7528 1748 7592 1752
rect 7528 1692 7532 1748
rect 7532 1692 7588 1748
rect 7588 1692 7592 1748
rect 7528 1688 7592 1692
rect 7528 1428 7592 1432
rect 7528 1372 7532 1428
rect 7532 1372 7588 1428
rect 7588 1372 7592 1428
rect 7528 1368 7592 1372
rect 7528 1108 7592 1112
rect 7528 1052 7532 1108
rect 7532 1052 7588 1108
rect 7588 1052 7592 1108
rect 7528 1048 7592 1052
rect 7528 788 7592 792
rect 7528 732 7532 788
rect 7532 732 7588 788
rect 7588 732 7592 788
rect 7528 728 7592 732
rect 7528 468 7592 472
rect 7528 412 7532 468
rect 7532 412 7588 468
rect 7588 412 7592 468
rect 7528 408 7592 412
rect 7528 308 7592 312
rect 7528 252 7532 308
rect 7532 252 7588 308
rect 7588 252 7592 308
rect 7528 248 7592 252
rect 7528 -12 7592 -8
rect 7528 -68 7532 -12
rect 7532 -68 7588 -12
rect 7588 -68 7592 -12
rect 7528 -72 7592 -68
rect 7528 -332 7592 -328
rect 7528 -388 7532 -332
rect 7532 -388 7588 -332
rect 7588 -388 7592 -332
rect 7528 -392 7592 -388
rect 7528 -652 7592 -648
rect 7528 -708 7532 -652
rect 7532 -708 7588 -652
rect 7588 -708 7592 -652
rect 7528 -712 7592 -708
rect 7848 4308 7912 4312
rect 7848 4252 7852 4308
rect 7852 4252 7908 4308
rect 7908 4252 7912 4308
rect 7848 4248 7912 4252
rect 7848 3988 7912 3992
rect 7848 3932 7852 3988
rect 7852 3932 7908 3988
rect 7908 3932 7912 3988
rect 7848 3928 7912 3932
rect 7848 3668 7912 3672
rect 7848 3612 7852 3668
rect 7852 3612 7908 3668
rect 7908 3612 7912 3668
rect 7848 3608 7912 3612
rect 7848 3348 7912 3352
rect 7848 3292 7852 3348
rect 7852 3292 7908 3348
rect 7908 3292 7912 3348
rect 7848 3288 7912 3292
rect 7848 3188 7912 3192
rect 7848 3132 7852 3188
rect 7852 3132 7908 3188
rect 7908 3132 7912 3188
rect 7848 3128 7912 3132
rect 7848 2868 7912 2872
rect 7848 2812 7852 2868
rect 7852 2812 7908 2868
rect 7908 2812 7912 2868
rect 7848 2808 7912 2812
rect 7848 2548 7912 2552
rect 7848 2492 7852 2548
rect 7852 2492 7908 2548
rect 7908 2492 7912 2548
rect 7848 2488 7912 2492
rect 7848 2228 7912 2232
rect 7848 2172 7852 2228
rect 7852 2172 7908 2228
rect 7908 2172 7912 2228
rect 7848 2168 7912 2172
rect 7848 1908 7912 1912
rect 7848 1852 7852 1908
rect 7852 1852 7908 1908
rect 7908 1852 7912 1908
rect 7848 1848 7912 1852
rect 7848 1748 7912 1752
rect 7848 1692 7852 1748
rect 7852 1692 7908 1748
rect 7908 1692 7912 1748
rect 7848 1688 7912 1692
rect 12808 1828 12872 1832
rect 12808 1772 12812 1828
rect 12812 1772 12868 1828
rect 12868 1772 12872 1828
rect 12808 1768 12872 1772
rect 7848 1428 7912 1432
rect 7848 1372 7852 1428
rect 7852 1372 7908 1428
rect 7908 1372 7912 1428
rect 7848 1368 7912 1372
rect 7848 1108 7912 1112
rect 7848 1052 7852 1108
rect 7852 1052 7908 1108
rect 7908 1052 7912 1108
rect 7848 1048 7912 1052
rect 7848 788 7912 792
rect 7848 732 7852 788
rect 7852 732 7908 788
rect 7908 732 7912 788
rect 7848 728 7912 732
rect 7848 468 7912 472
rect 7848 412 7852 468
rect 7852 412 7908 468
rect 7908 412 7912 468
rect 7848 408 7912 412
rect 7848 308 7912 312
rect 7848 252 7852 308
rect 7852 252 7908 308
rect 7908 252 7912 308
rect 7848 248 7912 252
rect 7848 -12 7912 -8
rect 7848 -68 7852 -12
rect 7852 -68 7908 -12
rect 7908 -68 7912 -12
rect 7848 -72 7912 -68
rect 7848 -332 7912 -328
rect 7848 -388 7852 -332
rect 7852 -388 7908 -332
rect 7908 -388 7912 -332
rect 7848 -392 7912 -388
rect 7848 -652 7912 -648
rect 7848 -708 7852 -652
rect 7852 -708 7908 -652
rect 7908 -708 7912 -652
rect 7848 -712 7912 -708
<< metal4 >>
rect 4640 4312 7920 4320
rect 4640 4248 4648 4312
rect 4712 4248 4968 4312
rect 5032 4248 5288 4312
rect 5352 4248 5608 4312
rect 5672 4248 5928 4312
rect 5992 4248 6248 4312
rect 6312 4248 6568 4312
rect 6632 4248 6888 4312
rect 6952 4248 7208 4312
rect 7272 4248 7528 4312
rect 7592 4248 7848 4312
rect 7912 4248 7920 4312
rect 4640 4240 7920 4248
rect 4640 3992 7920 4000
rect 4640 3928 4648 3992
rect 4712 3928 4968 3992
rect 5032 3928 5288 3992
rect 5352 3928 5608 3992
rect 5672 3928 5928 3992
rect 5992 3928 6248 3992
rect 6312 3928 6568 3992
rect 6632 3928 6888 3992
rect 6952 3928 7208 3992
rect 7272 3928 7528 3992
rect 7592 3928 7848 3992
rect 7912 3928 7920 3992
rect 4640 3920 7920 3928
rect 4640 3672 7920 3680
rect 4640 3608 4648 3672
rect 4712 3608 4968 3672
rect 5032 3608 5288 3672
rect 5352 3608 5608 3672
rect 5672 3608 5928 3672
rect 5992 3608 6248 3672
rect 6312 3608 6568 3672
rect 6632 3608 6888 3672
rect 6952 3608 7208 3672
rect 7272 3608 7528 3672
rect 7592 3608 7848 3672
rect 7912 3608 7920 3672
rect 4640 3600 7920 3608
rect 5920 3512 6640 3520
rect 5920 3448 5928 3512
rect 5992 3448 6248 3512
rect 6312 3448 6568 3512
rect 6632 3448 6640 3512
rect 5920 3440 6640 3448
rect 4640 3352 7920 3360
rect 4640 3288 4648 3352
rect 4712 3288 4968 3352
rect 5032 3288 5288 3352
rect 5352 3288 5608 3352
rect 5672 3288 5928 3352
rect 5992 3288 6248 3352
rect 6312 3288 6568 3352
rect 6632 3288 6888 3352
rect 6952 3288 7208 3352
rect 7272 3288 7528 3352
rect 7592 3288 7848 3352
rect 7912 3288 7920 3352
rect 4640 3280 7920 3288
rect 4640 3192 7920 3200
rect 4640 3128 4648 3192
rect 4712 3128 4968 3192
rect 5032 3128 5288 3192
rect 5352 3128 5608 3192
rect 5672 3128 5928 3192
rect 5992 3128 6248 3192
rect 6312 3128 6568 3192
rect 6632 3128 6888 3192
rect 6952 3128 7208 3192
rect 7272 3128 7528 3192
rect 7592 3128 7848 3192
rect 7912 3128 7920 3192
rect 4640 3120 7920 3128
rect 4640 2872 7920 2880
rect 4640 2808 4648 2872
rect 4712 2808 4968 2872
rect 5032 2808 5288 2872
rect 5352 2808 5608 2872
rect 5672 2808 5928 2872
rect 5992 2808 6248 2872
rect 6312 2808 6568 2872
rect 6632 2808 6888 2872
rect 6952 2808 7208 2872
rect 7272 2808 7528 2872
rect 7592 2808 7848 2872
rect 7912 2808 7920 2872
rect 4640 2800 7920 2808
rect 5920 2712 6640 2720
rect 5920 2648 5928 2712
rect 5992 2648 6248 2712
rect 6312 2648 6568 2712
rect 6632 2648 6640 2712
rect 5920 2640 6640 2648
rect 4640 2552 7920 2560
rect 4640 2488 4648 2552
rect 4712 2488 4968 2552
rect 5032 2488 5288 2552
rect 5352 2488 5608 2552
rect 5672 2488 5928 2552
rect 5992 2488 6248 2552
rect 6312 2488 6568 2552
rect 6632 2488 6888 2552
rect 6952 2488 7208 2552
rect 7272 2488 7528 2552
rect 7592 2488 7848 2552
rect 7912 2488 7920 2552
rect 4640 2480 7920 2488
rect 4640 2232 7920 2240
rect 4640 2168 4648 2232
rect 4712 2168 4968 2232
rect 5032 2168 5288 2232
rect 5352 2168 5608 2232
rect 5672 2168 5928 2232
rect 5992 2168 6248 2232
rect 6312 2168 6568 2232
rect 6632 2168 6888 2232
rect 6952 2168 7208 2232
rect 7272 2168 7528 2232
rect 7592 2168 7848 2232
rect 7912 2168 7920 2232
rect 4640 2160 7920 2168
rect -480 1918 -80 2000
rect -480 1682 -398 1918
rect -162 1682 -80 1918
rect 4640 1912 7920 1920
rect 4640 1848 4648 1912
rect 4712 1848 4968 1912
rect 5032 1848 5288 1912
rect 5352 1848 5608 1912
rect 5672 1848 5928 1912
rect 5992 1848 6248 1912
rect 6312 1848 6568 1912
rect 6632 1848 6888 1912
rect 6952 1848 7208 1912
rect 7272 1848 7528 1912
rect 7592 1848 7848 1912
rect 7912 1848 7920 1912
rect 4640 1840 7920 1848
rect 12640 1918 13040 2000
rect -480 1600 -80 1682
rect 4640 1752 7920 1760
rect 4640 1688 4648 1752
rect 4712 1688 4968 1752
rect 5032 1688 5288 1752
rect 5352 1688 5608 1752
rect 5672 1688 5928 1752
rect 5992 1688 6248 1752
rect 6312 1688 6568 1752
rect 6632 1688 6888 1752
rect 6952 1688 7208 1752
rect 7272 1688 7528 1752
rect 7592 1688 7848 1752
rect 7912 1688 7920 1752
rect 4640 1680 7920 1688
rect 12640 1682 12722 1918
rect 12958 1682 13040 1918
rect 12640 1600 13040 1682
rect 4640 1432 7920 1440
rect 4640 1368 4648 1432
rect 4712 1368 4968 1432
rect 5032 1368 5288 1432
rect 5352 1368 5608 1432
rect 5672 1368 5928 1432
rect 5992 1368 6248 1432
rect 6312 1368 6568 1432
rect 6632 1368 6888 1432
rect 6952 1368 7208 1432
rect 7272 1368 7528 1432
rect 7592 1368 7848 1432
rect 7912 1368 7920 1432
rect 4640 1360 7920 1368
rect 4640 1112 7920 1120
rect 4640 1048 4648 1112
rect 4712 1048 4968 1112
rect 5032 1048 5288 1112
rect 5352 1048 5608 1112
rect 5672 1048 5928 1112
rect 5992 1048 6248 1112
rect 6312 1048 6568 1112
rect 6632 1048 6888 1112
rect 6952 1048 7208 1112
rect 7272 1048 7528 1112
rect 7592 1048 7848 1112
rect 7912 1048 7920 1112
rect 4640 1040 7920 1048
rect 5920 952 6640 960
rect 5920 888 5928 952
rect 5992 888 6248 952
rect 6312 888 6568 952
rect 6632 888 6640 952
rect 5920 880 6640 888
rect 4640 792 7920 800
rect 4640 728 4648 792
rect 4712 728 4968 792
rect 5032 728 5288 792
rect 5352 728 5608 792
rect 5672 728 5928 792
rect 5992 728 6248 792
rect 6312 728 6568 792
rect 6632 728 6888 792
rect 6952 728 7208 792
rect 7272 728 7528 792
rect 7592 728 7848 792
rect 7912 728 7920 792
rect 4640 720 7920 728
rect 4640 472 7920 480
rect 4640 408 4648 472
rect 4712 408 4968 472
rect 5032 408 5288 472
rect 5352 408 5608 472
rect 5672 408 5928 472
rect 5992 408 6248 472
rect 6312 408 6568 472
rect 6632 408 6888 472
rect 6952 408 7208 472
rect 7272 408 7528 472
rect 7592 408 7848 472
rect 7912 408 7920 472
rect 4640 400 7920 408
rect 4640 312 7920 320
rect 4640 248 4648 312
rect 4712 248 4968 312
rect 5032 248 5288 312
rect 5352 248 5608 312
rect 5672 248 5928 312
rect 5992 248 6248 312
rect 6312 248 6568 312
rect 6632 248 6888 312
rect 6952 248 7208 312
rect 7272 248 7528 312
rect 7592 248 7848 312
rect 7912 248 7920 312
rect 4640 240 7920 248
rect 5920 152 6640 160
rect 5920 88 5928 152
rect 5992 88 6248 152
rect 6312 88 6568 152
rect 6632 88 6640 152
rect 5920 80 6640 88
rect 4640 -8 7920 0
rect 4640 -72 4648 -8
rect 4712 -72 4968 -8
rect 5032 -72 5288 -8
rect 5352 -72 5608 -8
rect 5672 -72 5928 -8
rect 5992 -72 6248 -8
rect 6312 -72 6568 -8
rect 6632 -72 6888 -8
rect 6952 -72 7208 -8
rect 7272 -72 7528 -8
rect 7592 -72 7848 -8
rect 7912 -72 7920 -8
rect 4640 -80 7920 -72
rect 4640 -328 7920 -320
rect 4640 -392 4648 -328
rect 4712 -392 4968 -328
rect 5032 -392 5288 -328
rect 5352 -392 5608 -328
rect 5672 -392 5928 -328
rect 5992 -392 6248 -328
rect 6312 -392 6568 -328
rect 6632 -392 6888 -328
rect 6952 -392 7208 -328
rect 7272 -392 7528 -328
rect 7592 -392 7848 -328
rect 7912 -392 7920 -328
rect 4640 -400 7920 -392
rect 4640 -648 7920 -640
rect 4640 -712 4648 -648
rect 4712 -712 4968 -648
rect 5032 -712 5288 -648
rect 5352 -712 5608 -648
rect 5672 -712 5928 -648
rect 5992 -712 6248 -648
rect 6312 -712 6568 -648
rect 6632 -712 6888 -648
rect 6952 -712 7208 -648
rect 7272 -712 7528 -648
rect 7592 -712 7848 -648
rect 7912 -712 7920 -648
rect 4640 -720 7920 -712
<< via4 >>
rect -398 1832 -162 1918
rect -398 1768 -312 1832
rect -312 1768 -248 1832
rect -248 1768 -162 1832
rect -398 1682 -162 1768
rect 12722 1832 12958 1918
rect 12722 1768 12808 1832
rect 12808 1768 12872 1832
rect 12872 1768 12958 1832
rect 12722 1682 12958 1768
<< metal5 >>
rect -480 1918 -80 4320
rect -480 1682 -398 1918
rect -162 1682 -80 1918
rect -480 -720 -80 1682
rect 12640 1918 13040 4320
rect 12640 1682 12722 1918
rect 12958 1682 13040 1918
rect 12640 -720 13040 1682
<< labels >>
rlabel metal3 s 4800 -720 4880 4320 4 xp
port 1 nsew
rlabel metal3 s 5120 -720 5200 4320 4 om
port 2 nsew
rlabel metal3 s 5440 -720 5520 4320 4 xm
port 3 nsew
rlabel metal3 s 5760 -720 5840 4320 4 op
port 4 nsew
rlabel metal3 s 6080 -720 6160 4320 4 fsb
port 5 nsew
rlabel metal3 s 6400 -720 6480 4320 4 q
port 6 nsew
rlabel metal3 s 4640 -640 4720 -560 4 gnda
port 7 nsew
rlabel metal5 s -480 -720 -80 -640 4 vssa
port 8 nsew
<< end >>
