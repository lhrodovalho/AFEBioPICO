magic
tech sky130A
timestamp 1634665005
<< nwell >>
rect 0 70 940 2900
<< pwell >>
rect 0 2900 940 2970
<< pmoslvt >>
rect 70 2520 870 2820
rect 70 2190 870 2490
rect 70 1860 870 2160
rect 70 1530 870 1830
rect 70 1200 870 1500
rect 70 870 870 1170
rect 70 540 870 840
rect 70 210 870 510
<< pdiff >>
rect 20 2810 70 2820
rect 20 2530 30 2810
rect 60 2530 70 2810
rect 20 2520 70 2530
rect 870 2810 920 2820
rect 870 2530 880 2810
rect 910 2530 920 2810
rect 870 2520 920 2530
rect 20 2480 70 2490
rect 20 2200 30 2480
rect 60 2200 70 2480
rect 20 2190 70 2200
rect 870 2480 920 2490
rect 870 2200 880 2480
rect 910 2200 920 2480
rect 870 2190 920 2200
rect 20 2150 70 2160
rect 20 1870 30 2150
rect 60 1870 70 2150
rect 20 1860 70 1870
rect 870 2150 920 2160
rect 870 1870 880 2150
rect 910 1870 920 2150
rect 870 1860 920 1870
rect 20 1820 70 1830
rect 20 1540 30 1820
rect 60 1540 70 1820
rect 20 1530 70 1540
rect 870 1820 920 1830
rect 870 1540 880 1820
rect 910 1540 920 1820
rect 870 1530 920 1540
rect 20 1490 70 1500
rect 20 1210 30 1490
rect 60 1210 70 1490
rect 20 1200 70 1210
rect 870 1490 920 1500
rect 870 1210 880 1490
rect 910 1210 920 1490
rect 870 1200 920 1210
rect 20 1160 70 1170
rect 20 880 30 1160
rect 60 880 70 1160
rect 20 870 70 880
rect 870 1160 920 1170
rect 870 880 880 1160
rect 910 880 920 1160
rect 870 870 920 880
rect 20 830 70 840
rect 20 550 30 830
rect 60 550 70 830
rect 20 540 70 550
rect 870 830 920 840
rect 870 550 880 830
rect 910 550 920 830
rect 870 540 920 550
rect 20 500 70 510
rect 20 220 30 500
rect 60 220 70 500
rect 20 210 70 220
rect 870 500 920 510
rect 870 220 880 500
rect 910 220 920 500
rect 870 210 920 220
<< pdiffc >>
rect 30 2530 60 2810
rect 880 2530 910 2810
rect 30 2200 60 2480
rect 880 2200 910 2480
rect 30 1870 60 2150
rect 880 1870 910 2150
rect 30 1540 60 1820
rect 880 1540 910 1820
rect 30 1210 60 1490
rect 880 1210 910 1490
rect 30 880 60 1160
rect 880 880 910 1160
rect 30 550 60 830
rect 880 550 910 830
rect 30 220 60 500
rect 880 220 910 500
<< psubdiff >>
rect 0 2920 70 2950
rect 870 2920 940 2950
<< nsubdiff >>
rect 20 2850 70 2880
rect 870 2850 920 2880
rect 20 90 70 120
rect 870 90 920 120
<< psubdiffcont >>
rect 70 2920 870 2950
<< nsubdiffcont >>
rect 70 2850 870 2880
rect 70 90 870 120
<< poly >>
rect 70 2820 870 2840
rect 70 2490 870 2520
rect 70 2160 870 2190
rect 70 1830 870 1860
rect 70 1500 870 1530
rect 70 1170 870 1200
rect 70 840 870 870
rect 70 510 870 540
rect 70 180 870 210
rect 70 150 90 180
rect 850 150 870 180
rect 70 140 870 150
<< polycont >>
rect 90 150 850 180
<< locali >>
rect 0 2920 70 2950
rect 870 2920 940 2950
rect 0 2850 70 2880
rect 870 2850 940 2880
rect 30 2810 60 2820
rect 30 2480 60 2530
rect 30 2150 60 2200
rect 30 1820 60 1870
rect 30 1490 60 1540
rect 880 2810 910 2820
rect 880 2480 910 2530
rect 880 2150 910 2200
rect 880 1820 910 1870
rect 880 1530 910 1540
rect 30 1160 60 1210
rect 30 830 60 880
rect 30 500 60 550
rect 30 210 60 220
rect 880 1490 910 1500
rect 880 1160 910 1210
rect 880 830 910 880
rect 880 500 910 550
rect 880 210 910 220
rect 80 150 90 180
rect 850 150 860 180
rect 0 90 70 120
rect 870 90 940 120
<< viali >>
rect 880 2530 910 2810
rect 880 220 910 500
rect 150 150 180 180
<< metal1 >>
rect 880 2820 910 2970
rect 870 2810 920 2820
rect 870 2530 880 2810
rect 910 2530 920 2810
rect 870 2520 920 2530
rect 870 500 920 510
rect 870 220 880 500
rect 910 220 920 500
rect 870 210 920 220
rect 140 180 190 190
rect 140 150 150 180
rect 180 150 190 180
rect 140 140 190 150
rect 150 0 180 140
rect 880 0 910 210
<< labels >>
rlabel metal1 880 0 910 10 1 D
port 1 n
rlabel metal1 150 0 180 10 1 G
port 2 n
rlabel metal1 880 2960 910 2970 5 S
port 3 s
rlabel locali 0 2850 10 2880 3 B
port 4 e
rlabel locali 0 2920 10 2950 3 SUB
port 5 e
rlabel locali 40 1510 50 1520 1 X
<< end >>
