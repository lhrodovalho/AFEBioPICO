magic
tech sky130A
timestamp 1634602342
<< pwell >>
rect -1970 -3360 -1880 -390
<< psubdiff >>
rect -1880 -3340 -1810 -3310
rect 10270 -3340 10340 -3310
rect -1880 -6310 10340 -6280
<< psubdiffcont >>
rect -1810 -3340 10270 -3310
<< locali >>
rect -1010 -480 -960 -470
rect -1010 -510 -1000 -480
rect -970 -510 -960 -480
rect -1010 -520 -960 -510
rect -1880 -3340 -1850 -3310
rect -1820 -3340 -1810 -3310
rect 10270 -3340 10340 -3310
rect -1880 -3490 10340 -3400
rect -1880 -3520 -1850 -3490
rect -1880 -3610 10340 -3520
rect -1880 -3640 -1850 -3610
rect -1880 -3730 10340 -3640
rect -1880 -3760 -1850 -3730
rect -1880 -3850 10340 -3760
rect -1880 -3880 -1850 -3850
rect -1880 -3970 10340 -3880
rect -1880 -4000 -1850 -3970
rect -1880 -4090 10340 -4000
rect -1880 -4120 -1850 -4090
rect -1880 -4150 10340 -4120
rect -1880 -4310 -1790 -4150
rect -1760 -4310 10340 -4150
rect -1880 -4340 10340 -4310
rect -1880 -4370 -1850 -4340
rect -1880 -4460 10340 -4370
rect -1880 -4490 -1850 -4460
rect -1880 -4580 10340 -4490
rect -1880 -4610 -1850 -4580
rect -1880 -4700 10340 -4610
rect -1880 -4730 -1850 -4700
rect -1880 -4820 10340 -4730
rect -1880 -4850 -1850 -4820
rect -1880 -4940 10340 -4850
rect -1880 -4970 -1850 -4940
rect -1880 -5060 10340 -4970
rect -1860 -6280 -1810 -6270
rect -1880 -6310 -1850 -6280
rect -1820 -6310 10340 -6280
rect -1860 -6320 -1810 -6310
<< viali >>
rect -1000 -510 -970 -480
rect -1850 -3340 -1820 -3310
rect -1790 -4310 -1760 -4150
rect -1850 -6310 -1820 -6280
<< metal1 >>
rect -1000 -230 -970 -220
rect -1000 -390 -970 -370
rect 880 -230 910 -220
rect 880 -450 910 -370
rect 1820 -230 1850 -220
rect 1820 -450 1850 -370
rect 3700 -230 3730 -220
rect 3700 -390 3730 -370
rect 5580 -230 5610 -220
rect 5580 -390 5610 -370
rect 7460 -230 7490 -220
rect 7460 -390 7490 -370
rect 10280 -230 10310 -220
rect 10280 -390 10310 -370
rect -1010 -480 -960 -470
rect -1010 -510 -1000 -480
rect -970 -510 -960 -480
rect -1010 -520 -960 -510
rect -1860 -3310 -1810 -3300
rect -1860 -3340 -1850 -3310
rect -1820 -3340 -1810 -3310
rect -1860 -3350 -1810 -3340
rect -1850 -6270 -1820 -3350
rect -1790 -3370 -1760 -3360
rect -1790 -3490 -1760 -3400
rect -1730 -3430 -1700 -3360
rect -1730 -3470 -1700 -3460
rect -1000 -3430 -970 -3360
rect -1000 -3470 -970 -3460
rect -1790 -3610 -1760 -3520
rect -910 -3550 -880 -3360
rect -910 -3590 -880 -3580
rect -790 -3550 -760 -3360
rect -60 -3430 -30 -3150
rect 1820 -3160 1850 -3150
rect -60 -3470 -30 -3460
rect 150 -3430 180 -3360
rect 150 -3470 180 -3460
rect -790 -3590 -760 -3580
rect -1790 -3730 -1760 -3640
rect -1790 -3850 -1760 -3760
rect -1790 -3970 -1760 -3880
rect -1790 -4090 -1760 -4000
rect -1790 -4140 -1760 -4120
rect -1800 -4150 -1750 -4140
rect -1800 -4310 -1790 -4150
rect -1760 -4310 -1750 -4150
rect -1800 -4320 -1750 -4310
rect -1790 -4340 -1760 -4320
rect -1790 -4460 -1760 -4370
rect -1790 -4580 -1760 -4490
rect -1790 -4700 -1760 -4610
rect -1790 -4820 -1760 -4730
rect -1790 -4940 -1760 -4850
rect -1790 -5060 -1760 -4970
rect 760 -4880 790 -4870
rect -1790 -5100 -1760 -5090
rect -1120 -5000 -1090 -4990
rect -1120 -5100 -1090 -5030
rect -910 -5000 -880 -4990
rect -910 -5100 -880 -5030
rect -180 -5000 -150 -4990
rect -180 -5100 -150 -5030
rect 30 -5000 60 -4990
rect 30 -5240 60 -5030
rect 760 -5100 790 -4910
rect 880 -4880 910 -3360
rect 1090 -3430 1120 -3360
rect 1090 -3470 1120 -3460
rect 1820 -3670 1850 -3360
rect 1820 -3710 1850 -3700
rect 1910 -3670 1940 -3360
rect 1910 -3710 1940 -3700
rect 2030 -3790 2060 -3360
rect 2030 -3830 2060 -3820
rect 880 -5100 910 -4910
rect 970 -4030 1000 -4020
rect 970 -5100 1000 -4060
rect 1910 -4030 1940 -4020
rect 1700 -4520 1730 -4510
rect 1700 -5100 1730 -4550
rect 1910 -5240 1940 -4060
rect 2760 -4030 2790 -3150
rect 2970 -3430 3000 -3360
rect 2970 -3470 3000 -3460
rect 3700 -3670 3730 -3360
rect 3700 -3710 3730 -3700
rect 3790 -3670 3820 -3360
rect 3790 -3710 3820 -3700
rect 3910 -3910 3940 -3350
rect 3910 -3950 3940 -3940
rect 2760 -4070 2790 -4060
rect 2850 -4400 2880 -4390
rect 2640 -4520 2670 -4510
rect 2640 -5100 2670 -4550
rect 2760 -4520 2790 -4510
rect 2760 -5100 2790 -4550
rect 2850 -5100 2880 -4430
rect 3790 -4400 3820 -4390
rect 3580 -4520 3610 -4510
rect 3580 -5100 3610 -4550
rect 3790 -5240 3820 -4430
rect 4640 -4400 4670 -3150
rect 4850 -3430 4880 -3360
rect 4850 -3470 4880 -3460
rect 4640 -4440 4670 -4430
rect 4730 -4400 4760 -4390
rect 4520 -4520 4550 -4510
rect 4520 -5100 4550 -4550
rect 4640 -4760 4670 -4750
rect 4640 -5100 4670 -4790
rect 4730 -5100 4760 -4430
rect 5460 -4520 5490 -4510
rect 5460 -5100 5490 -4550
rect 5580 -4520 5610 -3360
rect 5670 -3670 5700 -3360
rect 5670 -3710 5700 -3700
rect 5790 -3910 5820 -3360
rect 5790 -3950 5820 -3940
rect 5580 -4560 5610 -4550
rect 5670 -4400 5700 -4390
rect 5670 -5240 5700 -4430
rect 6520 -4400 6550 -3150
rect 6730 -3430 6760 -3360
rect 6730 -3470 6760 -3460
rect 6520 -4440 6550 -4430
rect 6610 -4030 6640 -4020
rect 6400 -4520 6430 -4510
rect 6400 -5100 6430 -4550
rect 6520 -4760 6550 -4750
rect 6520 -5100 6550 -4790
rect 6610 -5100 6640 -4060
rect 7340 -4520 7370 -4510
rect 7340 -5100 7370 -4550
rect 7460 -4640 7490 -3360
rect 7550 -3670 7580 -3360
rect 7550 -3710 7580 -3700
rect 7670 -3790 7700 -3360
rect 7670 -3830 7700 -3820
rect 7460 -4680 7490 -4670
rect 7550 -4030 7580 -4020
rect 7550 -5240 7580 -4060
rect 8400 -4030 8430 -3150
rect 8400 -4070 8430 -4060
rect 8280 -4520 8310 -4510
rect 8280 -5100 8310 -4550
rect 8400 -4520 8430 -4510
rect 8400 -5100 8430 -4550
rect 8490 -4640 8520 -3360
rect 8610 -3550 8640 -3360
rect 8610 -3590 8640 -3580
rect 8490 -5240 8520 -4670
rect 9340 -4760 9370 -3150
rect 9430 -4160 9460 -3360
rect 9430 -4310 9460 -4300
rect 9550 -4640 9580 -3360
rect 9550 -4680 9580 -4670
rect 10280 -4160 10310 -4150
rect 9220 -4880 9250 -4870
rect 9220 -5100 9250 -4910
rect 9340 -5100 9370 -4790
rect 10160 -4760 10190 -4750
rect 10160 -5100 10190 -4790
rect 10280 -5100 10310 -4300
rect -1860 -6280 -1810 -6270
rect -1860 -6310 -1850 -6280
rect -1820 -6310 -1810 -6280
rect -1860 -6320 -1810 -6310
rect -1850 -6350 -1820 -6320
rect -1850 -6500 -1820 -6490
rect -910 -6350 -880 -6330
rect -910 -6500 -880 -6490
rect 970 -6350 1000 -6330
rect 970 -6500 1000 -6490
rect 2850 -6350 2880 -6330
rect 2850 -6500 2880 -6490
rect 4730 -6350 4760 -6330
rect 4730 -6500 4760 -6490
rect 6610 -6350 6640 -6330
rect 6610 -6500 6640 -6490
rect 9430 -6350 9460 -6330
rect 9430 -6500 9460 -6490
<< via1 >>
rect -1000 -370 -970 -230
rect 880 -370 910 -230
rect 1820 -370 1850 -230
rect 3700 -370 3730 -230
rect 5580 -370 5610 -230
rect 7460 -370 7490 -230
rect 10280 -370 10310 -230
rect -1790 -3400 -1760 -3370
rect -1730 -3460 -1700 -3430
rect -1000 -3460 -970 -3430
rect -1790 -3520 -1760 -3490
rect -910 -3580 -880 -3550
rect -60 -3460 -30 -3430
rect 150 -3460 180 -3430
rect -790 -3580 -760 -3550
rect -1790 -3640 -1760 -3610
rect -1790 -3760 -1760 -3730
rect -1790 -3880 -1760 -3850
rect -1790 -4000 -1760 -3970
rect -1790 -4120 -1760 -4090
rect -1790 -4370 -1760 -4340
rect -1790 -4490 -1760 -4460
rect -1790 -4610 -1760 -4580
rect -1790 -4730 -1760 -4700
rect -1790 -4850 -1760 -4820
rect -1790 -4970 -1760 -4940
rect 760 -4910 790 -4880
rect -1790 -5090 -1760 -5060
rect -1120 -5030 -1090 -5000
rect -910 -5030 -880 -5000
rect -180 -5030 -150 -5000
rect 30 -5030 60 -5000
rect 1090 -3460 1120 -3430
rect 1820 -3700 1850 -3670
rect 1910 -3700 1940 -3670
rect 2030 -3820 2060 -3790
rect 880 -4910 910 -4880
rect 970 -4060 1000 -4030
rect 1910 -4060 1940 -4030
rect 1700 -4550 1730 -4520
rect 2970 -3460 3000 -3430
rect 3700 -3700 3730 -3670
rect 3790 -3700 3820 -3670
rect 3910 -3940 3940 -3910
rect 2760 -4060 2790 -4030
rect 2850 -4430 2880 -4400
rect 2640 -4550 2670 -4520
rect 2760 -4550 2790 -4520
rect 3790 -4430 3820 -4400
rect 3580 -4550 3610 -4520
rect 4850 -3460 4880 -3430
rect 4640 -4430 4670 -4400
rect 4730 -4430 4760 -4400
rect 4520 -4550 4550 -4520
rect 4640 -4790 4670 -4760
rect 5460 -4550 5490 -4520
rect 5670 -3700 5700 -3670
rect 5790 -3940 5820 -3910
rect 5580 -4550 5610 -4520
rect 5670 -4430 5700 -4400
rect 6730 -3460 6760 -3430
rect 6520 -4430 6550 -4400
rect 6610 -4060 6640 -4030
rect 6400 -4550 6430 -4520
rect 6520 -4790 6550 -4760
rect 7340 -4550 7370 -4520
rect 7550 -3700 7580 -3670
rect 7670 -3820 7700 -3790
rect 7460 -4670 7490 -4640
rect 7550 -4060 7580 -4030
rect 8400 -4060 8430 -4030
rect 8280 -4550 8310 -4520
rect 8400 -4550 8430 -4520
rect 8610 -3580 8640 -3550
rect 8490 -4670 8520 -4640
rect 9430 -4300 9460 -4160
rect 9550 -4670 9580 -4640
rect 10280 -4300 10310 -4160
rect 9340 -4790 9370 -4760
rect 9220 -4910 9250 -4880
rect 10160 -4790 10190 -4760
rect -1850 -6490 -1820 -6350
rect -910 -6490 -880 -6350
rect 970 -6490 1000 -6350
rect 2850 -6490 2880 -6350
rect 4730 -6490 4760 -6350
rect 6610 -6490 6640 -6350
rect 9430 -6490 9460 -6350
<< metal2 >>
rect -1880 -230 10340 -220
rect -1880 -370 -1000 -230
rect -970 -370 880 -230
rect 910 -370 1820 -230
rect 1850 -370 3700 -230
rect 3730 -370 5580 -230
rect 5610 -370 7460 -230
rect 7490 -370 10280 -230
rect 10310 -370 10340 -230
rect -1880 -380 10340 -370
rect -1880 -3400 -1790 -3370
rect -1760 -3400 10340 -3370
rect -1880 -3460 -1730 -3430
rect -1700 -3460 -1000 -3430
rect -970 -3460 -60 -3430
rect -30 -3460 150 -3430
rect 180 -3460 1090 -3430
rect 1120 -3460 2970 -3430
rect 3000 -3460 4850 -3430
rect 4880 -3460 6730 -3430
rect 6760 -3460 10340 -3430
rect -1880 -3520 -1790 -3490
rect -1760 -3520 10340 -3490
rect -1880 -3580 -910 -3550
rect -880 -3580 -790 -3550
rect -760 -3580 8610 -3550
rect 8640 -3580 10340 -3550
rect -1880 -3640 -1790 -3610
rect -1760 -3640 10340 -3610
rect -1880 -3700 1820 -3670
rect 1850 -3700 1910 -3670
rect 1940 -3700 3700 -3670
rect 3730 -3700 3790 -3670
rect 3820 -3700 5670 -3670
rect 5700 -3700 7550 -3670
rect 7580 -3700 10340 -3670
rect -1880 -3760 -1790 -3730
rect -1760 -3760 10340 -3730
rect -1880 -3820 2030 -3790
rect 2060 -3820 7670 -3790
rect 7700 -3820 10340 -3790
rect -1880 -3880 -1790 -3850
rect -1760 -3880 10340 -3850
rect -1880 -3940 3910 -3910
rect 3940 -3940 5790 -3910
rect 5820 -3940 10340 -3910
rect -1880 -4000 -1790 -3970
rect -1760 -4000 10340 -3970
rect -1880 -4060 970 -4030
rect 1000 -4060 1910 -4030
rect 1940 -4060 2760 -4030
rect 2790 -4060 6610 -4030
rect 6640 -4060 7550 -4030
rect 7580 -4060 8400 -4030
rect 8430 -4060 10340 -4030
rect -1880 -4120 -1790 -4090
rect -1760 -4120 10340 -4090
rect -1880 -4160 10340 -4150
rect -1880 -4300 9430 -4160
rect 9460 -4300 10280 -4160
rect 10310 -4300 10340 -4160
rect -1880 -4310 10340 -4300
rect -1880 -4370 -1790 -4340
rect -1760 -4370 10340 -4340
rect -1880 -4430 2850 -4400
rect 2880 -4430 3790 -4400
rect 3820 -4430 4640 -4400
rect 4670 -4430 4730 -4400
rect 4760 -4430 5670 -4400
rect 5700 -4430 6520 -4400
rect 6550 -4430 10340 -4400
rect -1880 -4490 -1790 -4460
rect -1760 -4490 10340 -4460
rect -1880 -4550 1700 -4520
rect 1730 -4550 2640 -4520
rect 2670 -4550 2760 -4520
rect 2790 -4550 3580 -4520
rect 3610 -4550 4520 -4520
rect 4550 -4550 5460 -4520
rect 5490 -4550 5580 -4520
rect 5610 -4550 6400 -4520
rect 6430 -4550 7340 -4520
rect 7370 -4550 8280 -4520
rect 8310 -4550 8400 -4520
rect 8430 -4550 10340 -4520
rect -1880 -4610 -1790 -4580
rect -1760 -4610 10340 -4580
rect -1880 -4670 7460 -4640
rect 7490 -4670 8490 -4640
rect 8520 -4670 9550 -4640
rect 9580 -4670 10340 -4640
rect -1880 -4730 -1790 -4700
rect -1760 -4730 10340 -4700
rect -1880 -4790 4640 -4760
rect 4670 -4790 6520 -4760
rect 6550 -4790 9340 -4760
rect 9370 -4790 10160 -4760
rect 10190 -4790 10340 -4760
rect -1880 -4850 -1790 -4820
rect -1760 -4850 10340 -4820
rect -1880 -4910 760 -4880
rect 790 -4910 880 -4880
rect 910 -4910 9220 -4880
rect 9250 -4910 10340 -4880
rect -1880 -4970 -1790 -4940
rect -1760 -4970 10340 -4940
rect -1880 -5030 -1120 -5000
rect -1090 -5030 -910 -5000
rect -880 -5030 -180 -5000
rect -150 -5030 30 -5000
rect 60 -5030 10340 -5000
rect -1880 -5090 -1790 -5060
rect -1760 -5090 10340 -5060
rect -1880 -6350 10340 -6340
rect -1880 -6490 -1850 -6350
rect -1820 -6490 -910 -6350
rect -880 -6490 970 -6350
rect 1000 -6490 2850 -6350
rect 2880 -6490 4730 -6350
rect 4760 -6490 6610 -6350
rect 6640 -6490 9430 -6350
rect 9460 -6490 10340 -6350
rect -1880 -6500 10340 -6490
use p8_1  pa2_1
timestamp 1634440961
transform 1 0 -940 0 1 -3360
box 0 0 940 2970
use p1_8  pa1_1
timestamp 1634440922
transform 1 0 -1880 0 1 -3360
box 0 0 940 2970
use n1_8  nb4_1
timestamp 1634337365
transform 1 0 -940 0 1 -6330
box 0 0 940 1230
use n1_8  na4_1
timestamp 1634337365
transform 1 0 -1880 0 1 -6330
box 0 0 940 1230
use p1_8  pb1_1
timestamp 1634440922
transform 1 0 0 0 1 -3360
box 0 0 940 2970
use n8_1  nb3_1
timestamp 1634429522
transform 1 0 0 0 1 -6330
box 0 0 940 1230
use p1_8  pc1_1
timestamp 1634440922
transform 1 0 940 0 1 -3360
box 0 0 940 2970
use n1_8  ne4_1
timestamp 1634337365
transform 1 0 940 0 1 -6330
box 0 0 940 1230
use p8_1  pc2_1
timestamp 1634440961
transform 1 0 1880 0 1 -3360
box 0 0 940 2970
use n8_1  ne3_1
timestamp 1634429522
transform 1 0 1880 0 1 -6330
box 0 0 940 1230
use p1_8  pd1_1
timestamp 1634440922
transform 1 0 2820 0 1 -3360
box 0 0 940 2970
use n1_8  nf4_1
timestamp 1634337365
transform 1 0 2820 0 1 -6330
box 0 0 940 1230
use p8_1  pd2_1
timestamp 1634440961
transform 1 0 3760 0 1 -3360
box 0 0 940 2970
use n8_1  nf3_1
timestamp 1634429522
transform 1 0 3760 0 1 -6330
box 0 0 940 1230
use p1_8  pe1_1
timestamp 1634440922
transform 1 0 4700 0 1 -3360
box 0 0 940 2970
use n1_8  nf4_2
timestamp 1634337365
transform 1 0 4700 0 1 -6330
box 0 0 940 1230
use p8_1  pd2_2
timestamp 1634440961
transform 1 0 5640 0 1 -3360
box 0 0 940 2970
use n8_1  nf3_2
timestamp 1634429522
transform 1 0 5640 0 1 -6330
box 0 0 940 1230
use p1_8  pf1_1
timestamp 1634440922
transform 1 0 6580 0 1 -3360
box 0 0 940 2970
use n1_8  ne4_2
timestamp 1634337365
transform 1 0 6580 0 1 -6330
box 0 0 940 1230
use p8_1  pc2_2
timestamp 1634440961
transform 1 0 7520 0 1 -3360
box 0 0 940 2970
use n8_1  ne3_2
timestamp 1634429522
transform 1 0 7520 0 1 -6330
box 0 0 940 1230
use p8_1  pf2_1
timestamp 1634440961
transform 1 0 8460 0 1 -3360
box 0 0 940 2970
use n8_1  nf2_1
timestamp 1634429522
transform 1 0 8460 0 1 -6330
box 0 0 940 1230
use p8_1  pg1_1
timestamp 1634440961
transform 1 0 9400 0 1 -3360
box 0 0 940 2970
use n8_1  ng4_1
timestamp 1634429522
transform 1 0 9400 0 1 -6330
box 0 0 940 1230
<< labels >>
rlabel metal2 -1880 -4550 -1870 -4520 3 a
rlabel metal2 -1880 -4670 -1870 -4640 3 b
rlabel metal2 -1880 -4790 -1870 -4760 3 c
rlabel metal2 -1880 -4910 -1870 -4880 3 n2
rlabel metal2 -1880 -5030 -1870 -5000 3 n1
rlabel metal2 -1880 -3700 -1870 -3670 3 x
rlabel metal2 -1880 -3460 -1870 -3430 3 p1
rlabel metal2 -1880 -3820 -1870 -3790 1 inm
port 4 n
rlabel metal2 -1880 -3940 -1870 -3910 1 inp
port 5 n
rlabel metal2 -1880 -4060 -1870 -4030 1 xm
rlabel metal2 -1880 -4430 -1870 -4400 1 xp
rlabel metal2 -1880 -4310 -1870 -4150 1 out
port 6 n
rlabel metal2 -1880 -3580 -1870 -3550 1 ib
port 7 n
rlabel metal2 -1880 -380 -1870 -220 1 vdda
port 8 n
rlabel locali -1880 -3420 -1870 -3410 1 gnda
port 9 n
rlabel metal2 -1880 -6500 -1870 -6340 1 vssa
port 10 n
<< end >>
