magic
tech sky130A
timestamp 1633696713
<< pwell >>
rect 5130 6720 6070 7950
<< nmoslvt >>
rect 5200 7710 6000 7810
rect 5200 7580 6000 7680
rect 5200 7450 6000 7550
rect 5200 7320 6000 7420
rect 5200 7190 6000 7290
rect 5200 7060 6000 7160
rect 5200 6930 6000 7030
rect 5200 6800 6000 6900
<< ndiff >>
rect 5150 7800 5200 7810
rect 5150 7720 5160 7800
rect 5190 7720 5200 7800
rect 5150 7710 5200 7720
rect 6000 7800 6050 7810
rect 6000 7720 6010 7800
rect 6040 7720 6050 7800
rect 6000 7710 6050 7720
rect 5150 7670 5200 7680
rect 5150 7590 5160 7670
rect 5190 7590 5200 7670
rect 5150 7580 5200 7590
rect 6000 7670 6050 7680
rect 6000 7590 6010 7670
rect 6040 7590 6050 7670
rect 6000 7580 6050 7590
rect 5150 7540 5200 7550
rect 5150 7460 5160 7540
rect 5190 7460 5200 7540
rect 5150 7450 5200 7460
rect 6000 7540 6050 7550
rect 6000 7460 6010 7540
rect 6040 7460 6050 7540
rect 6000 7450 6050 7460
rect 5150 7410 5200 7420
rect 5150 7330 5160 7410
rect 5190 7330 5200 7410
rect 5150 7320 5200 7330
rect 6000 7410 6050 7420
rect 6000 7330 6010 7410
rect 6040 7330 6050 7410
rect 6000 7320 6050 7330
rect 5150 7280 5200 7290
rect 5150 7200 5160 7280
rect 5190 7200 5200 7280
rect 5150 7190 5200 7200
rect 6000 7280 6050 7290
rect 6000 7200 6010 7280
rect 6040 7200 6050 7280
rect 6000 7190 6050 7200
rect 5150 7150 5200 7160
rect 5150 7070 5160 7150
rect 5190 7070 5200 7150
rect 5150 7060 5200 7070
rect 6000 7150 6050 7160
rect 6000 7070 6010 7150
rect 6040 7070 6050 7150
rect 6000 7060 6050 7070
rect 5150 7020 5200 7030
rect 5150 6940 5160 7020
rect 5190 6940 5200 7020
rect 5150 6930 5200 6940
rect 6000 7020 6050 7030
rect 6000 6940 6010 7020
rect 6040 6940 6050 7020
rect 6000 6930 6050 6940
rect 5150 6890 5200 6900
rect 5150 6810 5160 6890
rect 5190 6810 5200 6890
rect 5150 6800 5200 6810
rect 6000 6890 6050 6900
rect 6000 6810 6010 6890
rect 6040 6810 6050 6890
rect 6000 6800 6050 6810
<< ndiffc >>
rect 5160 7720 5190 7800
rect 6010 7720 6040 7800
rect 5160 7590 5190 7670
rect 6010 7590 6040 7670
rect 5160 7460 5190 7540
rect 6010 7460 6040 7540
rect 5160 7330 5190 7410
rect 6010 7330 6040 7410
rect 5160 7200 5190 7280
rect 6010 7200 6040 7280
rect 5160 7070 5190 7150
rect 6010 7070 6040 7150
rect 5160 6940 5190 7020
rect 6010 6940 6040 7020
rect 5160 6810 5190 6890
rect 6010 6810 6040 6890
<< psubdiff >>
rect 5150 6740 5200 6770
rect 6000 6740 6050 6770
<< psubdiffcont >>
rect 5200 6740 6000 6770
<< poly >>
rect 5200 7870 6000 7880
rect 5200 7840 5220 7870
rect 5980 7840 6000 7870
rect 5200 7810 6000 7840
rect 5200 7680 6000 7710
rect 5200 7550 6000 7580
rect 5200 7420 6000 7450
rect 5200 7290 6000 7320
rect 5200 7160 6000 7190
rect 5200 7030 6000 7060
rect 5200 6900 6000 6930
rect 5200 6780 6000 6800
<< polycont >>
rect 5220 7840 5980 7870
<< locali >>
rect 5210 7840 5220 7870
rect 5980 7840 5990 7870
rect 5160 7800 5190 7810
rect 5160 7710 5190 7720
rect 6010 7800 6040 7810
rect 5160 7670 5190 7680
rect 5160 7540 5190 7590
rect 6010 7670 6040 7720
rect 6010 7580 6040 7590
rect 5160 7450 5190 7460
rect 6010 7540 6040 7550
rect 5160 7410 5190 7420
rect 5160 7280 5190 7330
rect 6010 7410 6040 7460
rect 6010 7320 6040 7330
rect 5160 7190 5190 7200
rect 6010 7280 6040 7290
rect 5160 7150 5190 7160
rect 5160 7020 5190 7070
rect 6010 7150 6040 7200
rect 6010 7060 6040 7070
rect 5160 6930 5190 6940
rect 6010 7020 6040 7030
rect 5160 6890 5190 6900
rect 5160 6800 5190 6810
rect 6010 6890 6040 6940
rect 6010 6800 6040 6810
rect 5150 6740 5200 6770
rect 6000 6740 6050 6770
<< viali >>
rect 5950 7840 5980 7870
rect 5160 7720 5190 7800
rect 5160 6810 5190 6890
<< metal1 >>
rect 5160 7810 5190 7930
rect 5950 7880 5980 7930
rect 5940 7870 5990 7880
rect 5940 7840 5950 7870
rect 5980 7840 5990 7870
rect 5940 7830 5990 7840
rect 5150 7800 5200 7810
rect 5150 7720 5160 7800
rect 5190 7720 5200 7800
rect 5150 7710 5200 7720
rect 5150 6890 5200 6900
rect 5150 6810 5160 6890
rect 5190 6810 5200 6890
rect 5150 6800 5200 6810
rect 5160 6740 5190 6800
<< labels >>
rlabel metal1 5170 6750 5180 6760 1 S
port 3 n
rlabel pwell 6020 6750 6030 6760 1 B
port 4 n
rlabel metal1 5960 7910 5970 7920 1 G
port 2 n
rlabel metal1 5170 7910 5180 7920 1 D
port 1 n
rlabel locali 6020 6910 6030 6920 1 x1
rlabel locali 5170 7040 5180 7050 1 x2
rlabel locali 6020 7170 6030 7180 1 x3
rlabel locali 5170 7300 5180 7310 1 x4
rlabel locali 6020 7430 6030 7440 1 x5
rlabel locali 5170 7560 5180 7570 1 x6
rlabel locali 6020 7690 6030 7700 1 x7
<< end >>
