magic
tech sky130A
magscale 1 2
timestamp 1634089225
<< error_p >>
rect 48606 14486 48610 14934
rect 48640 14520 48644 14900
<< pwell >>
rect 48540 -1240 80424 15084
<< psubdiff >>
rect 48576 15014 48672 15048
rect 80292 15014 80388 15048
rect 48576 14952 48610 15014
rect 80354 14952 80388 15014
rect 48576 -1170 48610 -1108
rect 80354 -1170 80388 -1108
rect 48576 -1204 48672 -1170
rect 80292 -1204 80388 -1170
<< psubdiffcont >>
rect 48672 15014 80292 15048
rect 48576 -1108 48610 14952
rect 80354 -1108 80388 14952
rect 48672 -1204 80292 -1170
<< xpolycontact >>
rect 48706 14486 48776 14918
rect 48706 7054 48776 7486
rect 49024 14486 49094 14918
rect 49024 7054 49094 7486
rect 49342 14486 49412 14918
rect 49342 7054 49412 7486
rect 49660 14486 49730 14918
rect 49660 7054 49730 7486
rect 49978 14486 50048 14918
rect 49978 7054 50048 7486
rect 50296 14486 50366 14918
rect 50296 7054 50366 7486
rect 50614 14486 50684 14918
rect 50614 7054 50684 7486
rect 50932 14486 51002 14918
rect 50932 7054 51002 7486
rect 51250 14486 51320 14918
rect 51250 7054 51320 7486
rect 51568 14486 51638 14918
rect 51568 7054 51638 7486
rect 51886 14486 51956 14918
rect 51886 7054 51956 7486
rect 52204 14486 52274 14918
rect 52204 7054 52274 7486
rect 52522 14486 52592 14918
rect 52522 7054 52592 7486
rect 52840 14486 52910 14918
rect 52840 7054 52910 7486
rect 53158 14486 53228 14918
rect 53158 7054 53228 7486
rect 53476 14486 53546 14918
rect 53476 7054 53546 7486
rect 53794 14486 53864 14918
rect 53794 7054 53864 7486
rect 54112 14486 54182 14918
rect 54112 7054 54182 7486
rect 54430 14486 54500 14918
rect 54430 7054 54500 7486
rect 54748 14486 54818 14918
rect 54748 7054 54818 7486
rect 55066 14486 55136 14918
rect 55066 7054 55136 7486
rect 55384 14486 55454 14918
rect 55384 7054 55454 7486
rect 55702 14486 55772 14918
rect 55702 7054 55772 7486
rect 56020 14486 56090 14918
rect 56020 7054 56090 7486
rect 56338 14486 56408 14918
rect 56338 7054 56408 7486
rect 56656 14486 56726 14918
rect 56656 7054 56726 7486
rect 56974 14486 57044 14918
rect 56974 7054 57044 7486
rect 57292 14486 57362 14918
rect 57292 7054 57362 7486
rect 57610 14486 57680 14918
rect 57610 7054 57680 7486
rect 57928 14486 57998 14918
rect 57928 7054 57998 7486
rect 58246 14486 58316 14918
rect 58246 7054 58316 7486
rect 58564 14486 58634 14918
rect 58564 7054 58634 7486
rect 58882 14486 58952 14918
rect 58882 7054 58952 7486
rect 59200 14486 59270 14918
rect 59200 7054 59270 7486
rect 59518 14486 59588 14918
rect 59518 7054 59588 7486
rect 59836 14486 59906 14918
rect 59836 7054 59906 7486
rect 60154 14486 60224 14918
rect 60154 7054 60224 7486
rect 60472 14486 60542 14918
rect 60472 7054 60542 7486
rect 60790 14486 60860 14918
rect 60790 7054 60860 7486
rect 61108 14486 61178 14918
rect 61108 7054 61178 7486
rect 61426 14486 61496 14918
rect 61426 7054 61496 7486
rect 61744 14486 61814 14918
rect 61744 7054 61814 7486
rect 62062 14486 62132 14918
rect 62062 7054 62132 7486
rect 62380 14486 62450 14918
rect 62380 7054 62450 7486
rect 62698 14486 62768 14918
rect 62698 7054 62768 7486
rect 63016 14486 63086 14918
rect 63016 7054 63086 7486
rect 63334 14486 63404 14918
rect 63334 7054 63404 7486
rect 63652 14486 63722 14918
rect 63652 7054 63722 7486
rect 63970 14486 64040 14918
rect 63970 7054 64040 7486
rect 64288 14486 64358 14918
rect 64288 7054 64358 7486
rect 64606 14486 64676 14918
rect 64606 7054 64676 7486
rect 64924 14486 64994 14918
rect 64924 7054 64994 7486
rect 65242 14486 65312 14918
rect 65242 7054 65312 7486
rect 65560 14486 65630 14918
rect 65560 7054 65630 7486
rect 65878 14486 65948 14918
rect 65878 7054 65948 7486
rect 66196 14486 66266 14918
rect 66196 7054 66266 7486
rect 66514 14486 66584 14918
rect 66514 7054 66584 7486
rect 66832 14486 66902 14918
rect 66832 7054 66902 7486
rect 67150 14486 67220 14918
rect 67150 7054 67220 7486
rect 67468 14486 67538 14918
rect 67468 7054 67538 7486
rect 67786 14486 67856 14918
rect 67786 7054 67856 7486
rect 68104 14486 68174 14918
rect 68104 7054 68174 7486
rect 68422 14486 68492 14918
rect 68422 7054 68492 7486
rect 68740 14486 68810 14918
rect 68740 7054 68810 7486
rect 69058 14486 69128 14918
rect 69058 7054 69128 7486
rect 69376 14486 69446 14918
rect 69376 7054 69446 7486
rect 69694 14486 69764 14918
rect 69694 7054 69764 7486
rect 70012 14486 70082 14918
rect 70012 7054 70082 7486
rect 70330 14486 70400 14918
rect 70330 7054 70400 7486
rect 70648 14486 70718 14918
rect 70648 7054 70718 7486
rect 70966 14486 71036 14918
rect 70966 7054 71036 7486
rect 71284 14486 71354 14918
rect 71284 7054 71354 7486
rect 71602 14486 71672 14918
rect 71602 7054 71672 7486
rect 71920 14486 71990 14918
rect 71920 7054 71990 7486
rect 72238 14486 72308 14918
rect 72238 7054 72308 7486
rect 72556 14486 72626 14918
rect 72556 7054 72626 7486
rect 72874 14486 72944 14918
rect 72874 7054 72944 7486
rect 73192 14486 73262 14918
rect 73192 7054 73262 7486
rect 73510 14486 73580 14918
rect 73510 7054 73580 7486
rect 73828 14486 73898 14918
rect 73828 7054 73898 7486
rect 74146 14486 74216 14918
rect 74146 7054 74216 7486
rect 74464 14486 74534 14918
rect 74464 7054 74534 7486
rect 74782 14486 74852 14918
rect 74782 7054 74852 7486
rect 75100 14486 75170 14918
rect 75100 7054 75170 7486
rect 75418 14486 75488 14918
rect 75418 7054 75488 7486
rect 75736 14486 75806 14918
rect 75736 7054 75806 7486
rect 76054 14486 76124 14918
rect 76054 7054 76124 7486
rect 76372 14486 76442 14918
rect 76372 7054 76442 7486
rect 76690 14486 76760 14918
rect 76690 7054 76760 7486
rect 77008 14486 77078 14918
rect 77008 7054 77078 7486
rect 77326 14486 77396 14918
rect 77326 7054 77396 7486
rect 77644 14486 77714 14918
rect 77644 7054 77714 7486
rect 77962 14486 78032 14918
rect 77962 7054 78032 7486
rect 78280 14486 78350 14918
rect 78280 7054 78350 7486
rect 78598 14486 78668 14918
rect 78598 7054 78668 7486
rect 78916 14486 78986 14918
rect 78916 7054 78986 7486
rect 79234 14486 79304 14918
rect 79234 7054 79304 7486
rect 79552 14486 79622 14918
rect 79552 7054 79622 7486
rect 79870 14486 79940 14918
rect 79870 7054 79940 7486
rect 80188 14486 80258 14918
rect 80188 7054 80258 7486
rect 48706 6358 48776 6790
rect 48706 -1074 48776 -642
rect 49024 6358 49094 6790
rect 49024 -1074 49094 -642
rect 49342 6358 49412 6790
rect 49342 -1074 49412 -642
rect 49660 6358 49730 6790
rect 49660 -1074 49730 -642
rect 49978 6358 50048 6790
rect 49978 -1074 50048 -642
rect 50296 6358 50366 6790
rect 50296 -1074 50366 -642
rect 50614 6358 50684 6790
rect 50614 -1074 50684 -642
rect 50932 6358 51002 6790
rect 50932 -1074 51002 -642
rect 51250 6358 51320 6790
rect 51250 -1074 51320 -642
rect 51568 6358 51638 6790
rect 51568 -1074 51638 -642
rect 51886 6358 51956 6790
rect 51886 -1074 51956 -642
rect 52204 6358 52274 6790
rect 52204 -1074 52274 -642
rect 52522 6358 52592 6790
rect 52522 -1074 52592 -642
rect 52840 6358 52910 6790
rect 52840 -1074 52910 -642
rect 53158 6358 53228 6790
rect 53158 -1074 53228 -642
rect 53476 6358 53546 6790
rect 53476 -1074 53546 -642
rect 53794 6358 53864 6790
rect 53794 -1074 53864 -642
rect 54112 6358 54182 6790
rect 54112 -1074 54182 -642
rect 54430 6358 54500 6790
rect 54430 -1074 54500 -642
rect 54748 6358 54818 6790
rect 54748 -1074 54818 -642
rect 55066 6358 55136 6790
rect 55066 -1074 55136 -642
rect 55384 6358 55454 6790
rect 55384 -1074 55454 -642
rect 55702 6358 55772 6790
rect 55702 -1074 55772 -642
rect 56020 6358 56090 6790
rect 56020 -1074 56090 -642
rect 56338 6358 56408 6790
rect 56338 -1074 56408 -642
rect 56656 6358 56726 6790
rect 56656 -1074 56726 -642
rect 56974 6358 57044 6790
rect 56974 -1074 57044 -642
rect 57292 6358 57362 6790
rect 57292 -1074 57362 -642
rect 57610 6358 57680 6790
rect 57610 -1074 57680 -642
rect 57928 6358 57998 6790
rect 57928 -1074 57998 -642
rect 58246 6358 58316 6790
rect 58246 -1074 58316 -642
rect 58564 6358 58634 6790
rect 58564 -1074 58634 -642
rect 58882 6358 58952 6790
rect 58882 -1074 58952 -642
rect 59200 6358 59270 6790
rect 59200 -1074 59270 -642
rect 59518 6358 59588 6790
rect 59518 -1074 59588 -642
rect 59836 6358 59906 6790
rect 59836 -1074 59906 -642
rect 60154 6358 60224 6790
rect 60154 -1074 60224 -642
rect 60472 6358 60542 6790
rect 60472 -1074 60542 -642
rect 60790 6358 60860 6790
rect 60790 -1074 60860 -642
rect 61108 6358 61178 6790
rect 61108 -1074 61178 -642
rect 61426 6358 61496 6790
rect 61426 -1074 61496 -642
rect 61744 6358 61814 6790
rect 61744 -1074 61814 -642
rect 62062 6358 62132 6790
rect 62062 -1074 62132 -642
rect 62380 6358 62450 6790
rect 62380 -1074 62450 -642
rect 62698 6358 62768 6790
rect 62698 -1074 62768 -642
rect 63016 6358 63086 6790
rect 63016 -1074 63086 -642
rect 63334 6358 63404 6790
rect 63334 -1074 63404 -642
rect 63652 6358 63722 6790
rect 63652 -1074 63722 -642
rect 63970 6358 64040 6790
rect 63970 -1074 64040 -642
rect 64288 6358 64358 6790
rect 64288 -1074 64358 -642
rect 64606 6358 64676 6790
rect 64606 -1074 64676 -642
rect 64924 6358 64994 6790
rect 64924 -1074 64994 -642
rect 65242 6358 65312 6790
rect 65242 -1074 65312 -642
rect 65560 6358 65630 6790
rect 65560 -1074 65630 -642
rect 65878 6358 65948 6790
rect 65878 -1074 65948 -642
rect 66196 6358 66266 6790
rect 66196 -1074 66266 -642
rect 66514 6358 66584 6790
rect 66514 -1074 66584 -642
rect 66832 6358 66902 6790
rect 66832 -1074 66902 -642
rect 67150 6358 67220 6790
rect 67150 -1074 67220 -642
rect 67468 6358 67538 6790
rect 67468 -1074 67538 -642
rect 67786 6358 67856 6790
rect 67786 -1074 67856 -642
rect 68104 6358 68174 6790
rect 68104 -1074 68174 -642
rect 68422 6358 68492 6790
rect 68422 -1074 68492 -642
rect 68740 6358 68810 6790
rect 68740 -1074 68810 -642
rect 69058 6358 69128 6790
rect 69058 -1074 69128 -642
rect 69376 6358 69446 6790
rect 69376 -1074 69446 -642
rect 69694 6358 69764 6790
rect 69694 -1074 69764 -642
rect 70012 6358 70082 6790
rect 70012 -1074 70082 -642
rect 70330 6358 70400 6790
rect 70330 -1074 70400 -642
rect 70648 6358 70718 6790
rect 70648 -1074 70718 -642
rect 70966 6358 71036 6790
rect 70966 -1074 71036 -642
rect 71284 6358 71354 6790
rect 71284 -1074 71354 -642
rect 71602 6358 71672 6790
rect 71602 -1074 71672 -642
rect 71920 6358 71990 6790
rect 71920 -1074 71990 -642
rect 72238 6358 72308 6790
rect 72238 -1074 72308 -642
rect 72556 6358 72626 6790
rect 72556 -1074 72626 -642
rect 72874 6358 72944 6790
rect 72874 -1074 72944 -642
rect 73192 6358 73262 6790
rect 73192 -1074 73262 -642
rect 73510 6358 73580 6790
rect 73510 -1074 73580 -642
rect 73828 6358 73898 6790
rect 73828 -1074 73898 -642
rect 74146 6358 74216 6790
rect 74146 -1074 74216 -642
rect 74464 6358 74534 6790
rect 74464 -1074 74534 -642
rect 74782 6358 74852 6790
rect 74782 -1074 74852 -642
rect 75100 6358 75170 6790
rect 75100 -1074 75170 -642
rect 75418 6358 75488 6790
rect 75418 -1074 75488 -642
rect 75736 6358 75806 6790
rect 75736 -1074 75806 -642
rect 76054 6358 76124 6790
rect 76054 -1074 76124 -642
rect 76372 6358 76442 6790
rect 76372 -1074 76442 -642
rect 76690 6358 76760 6790
rect 76690 -1074 76760 -642
rect 77008 6358 77078 6790
rect 77008 -1074 77078 -642
rect 77326 6358 77396 6790
rect 77326 -1074 77396 -642
rect 77644 6358 77714 6790
rect 77644 -1074 77714 -642
rect 77962 6358 78032 6790
rect 77962 -1074 78032 -642
rect 78280 6358 78350 6790
rect 78280 -1074 78350 -642
rect 78598 6358 78668 6790
rect 78598 -1074 78668 -642
rect 78916 6358 78986 6790
rect 78916 -1074 78986 -642
rect 79234 6358 79304 6790
rect 79234 -1074 79304 -642
rect 79552 6358 79622 6790
rect 79552 -1074 79622 -642
rect 79870 6358 79940 6790
rect 79870 -1074 79940 -642
rect 80188 6358 80258 6790
rect 80188 -1074 80258 -642
<< xpolyres >>
rect 48706 7486 48776 14486
rect 49024 7486 49094 14486
rect 49342 7486 49412 14486
rect 49660 7486 49730 14486
rect 49978 7486 50048 14486
rect 50296 7486 50366 14486
rect 50614 7486 50684 14486
rect 50932 7486 51002 14486
rect 51250 7486 51320 14486
rect 51568 7486 51638 14486
rect 51886 7486 51956 14486
rect 52204 7486 52274 14486
rect 52522 7486 52592 14486
rect 52840 7486 52910 14486
rect 53158 7486 53228 14486
rect 53476 7486 53546 14486
rect 53794 7486 53864 14486
rect 54112 7486 54182 14486
rect 54430 7486 54500 14486
rect 54748 7486 54818 14486
rect 55066 7486 55136 14486
rect 55384 7486 55454 14486
rect 55702 7486 55772 14486
rect 56020 7486 56090 14486
rect 56338 7486 56408 14486
rect 56656 7486 56726 14486
rect 56974 7486 57044 14486
rect 57292 7486 57362 14486
rect 57610 7486 57680 14486
rect 57928 7486 57998 14486
rect 58246 7486 58316 14486
rect 58564 7486 58634 14486
rect 58882 7486 58952 14486
rect 59200 7486 59270 14486
rect 59518 7486 59588 14486
rect 59836 7486 59906 14486
rect 60154 7486 60224 14486
rect 60472 7486 60542 14486
rect 60790 7486 60860 14486
rect 61108 7486 61178 14486
rect 61426 7486 61496 14486
rect 61744 7486 61814 14486
rect 62062 7486 62132 14486
rect 62380 7486 62450 14486
rect 62698 7486 62768 14486
rect 63016 7486 63086 14486
rect 63334 7486 63404 14486
rect 63652 7486 63722 14486
rect 63970 7486 64040 14486
rect 64288 7486 64358 14486
rect 64606 7486 64676 14486
rect 64924 7486 64994 14486
rect 65242 7486 65312 14486
rect 65560 7486 65630 14486
rect 65878 7486 65948 14486
rect 66196 7486 66266 14486
rect 66514 7486 66584 14486
rect 66832 7486 66902 14486
rect 67150 7486 67220 14486
rect 67468 7486 67538 14486
rect 67786 7486 67856 14486
rect 68104 7486 68174 14486
rect 68422 7486 68492 14486
rect 68740 7486 68810 14486
rect 69058 7486 69128 14486
rect 69376 7486 69446 14486
rect 69694 7486 69764 14486
rect 70012 7486 70082 14486
rect 70330 7486 70400 14486
rect 70648 7486 70718 14486
rect 70966 7486 71036 14486
rect 71284 7486 71354 14486
rect 71602 7486 71672 14486
rect 71920 7486 71990 14486
rect 72238 7486 72308 14486
rect 72556 7486 72626 14486
rect 72874 7486 72944 14486
rect 73192 7486 73262 14486
rect 73510 7486 73580 14486
rect 73828 7486 73898 14486
rect 74146 7486 74216 14486
rect 74464 7486 74534 14486
rect 74782 7486 74852 14486
rect 75100 7486 75170 14486
rect 75418 7486 75488 14486
rect 75736 7486 75806 14486
rect 76054 7486 76124 14486
rect 76372 7486 76442 14486
rect 76690 7486 76760 14486
rect 77008 7486 77078 14486
rect 77326 7486 77396 14486
rect 77644 7486 77714 14486
rect 77962 7486 78032 14486
rect 78280 7486 78350 14486
rect 78598 7486 78668 14486
rect 78916 7486 78986 14486
rect 79234 7486 79304 14486
rect 79552 7486 79622 14486
rect 79870 7486 79940 14486
rect 80188 7486 80258 14486
rect 48706 -642 48776 6358
rect 49024 -642 49094 6358
rect 49342 -642 49412 6358
rect 49660 -642 49730 6358
rect 49978 -642 50048 6358
rect 50296 -642 50366 6358
rect 50614 -642 50684 6358
rect 50932 -642 51002 6358
rect 51250 -642 51320 6358
rect 51568 -642 51638 6358
rect 51886 -642 51956 6358
rect 52204 -642 52274 6358
rect 52522 -642 52592 6358
rect 52840 -642 52910 6358
rect 53158 -642 53228 6358
rect 53476 -642 53546 6358
rect 53794 -642 53864 6358
rect 54112 -642 54182 6358
rect 54430 -642 54500 6358
rect 54748 -642 54818 6358
rect 55066 -642 55136 6358
rect 55384 -642 55454 6358
rect 55702 -642 55772 6358
rect 56020 -642 56090 6358
rect 56338 -642 56408 6358
rect 56656 -642 56726 6358
rect 56974 -642 57044 6358
rect 57292 -642 57362 6358
rect 57610 -642 57680 6358
rect 57928 -642 57998 6358
rect 58246 -642 58316 6358
rect 58564 -642 58634 6358
rect 58882 -642 58952 6358
rect 59200 -642 59270 6358
rect 59518 -642 59588 6358
rect 59836 -642 59906 6358
rect 60154 -642 60224 6358
rect 60472 -642 60542 6358
rect 60790 -642 60860 6358
rect 61108 -642 61178 6358
rect 61426 -642 61496 6358
rect 61744 -642 61814 6358
rect 62062 -642 62132 6358
rect 62380 -642 62450 6358
rect 62698 -642 62768 6358
rect 63016 -642 63086 6358
rect 63334 -642 63404 6358
rect 63652 -642 63722 6358
rect 63970 -642 64040 6358
rect 64288 -642 64358 6358
rect 64606 -642 64676 6358
rect 64924 -642 64994 6358
rect 65242 -642 65312 6358
rect 65560 -642 65630 6358
rect 65878 -642 65948 6358
rect 66196 -642 66266 6358
rect 66514 -642 66584 6358
rect 66832 -642 66902 6358
rect 67150 -642 67220 6358
rect 67468 -642 67538 6358
rect 67786 -642 67856 6358
rect 68104 -642 68174 6358
rect 68422 -642 68492 6358
rect 68740 -642 68810 6358
rect 69058 -642 69128 6358
rect 69376 -642 69446 6358
rect 69694 -642 69764 6358
rect 70012 -642 70082 6358
rect 70330 -642 70400 6358
rect 70648 -642 70718 6358
rect 70966 -642 71036 6358
rect 71284 -642 71354 6358
rect 71602 -642 71672 6358
rect 71920 -642 71990 6358
rect 72238 -642 72308 6358
rect 72556 -642 72626 6358
rect 72874 -642 72944 6358
rect 73192 -642 73262 6358
rect 73510 -642 73580 6358
rect 73828 -642 73898 6358
rect 74146 -642 74216 6358
rect 74464 -642 74534 6358
rect 74782 -642 74852 6358
rect 75100 -642 75170 6358
rect 75418 -642 75488 6358
rect 75736 -642 75806 6358
rect 76054 -642 76124 6358
rect 76372 -642 76442 6358
rect 76690 -642 76760 6358
rect 77008 -642 77078 6358
rect 77326 -642 77396 6358
rect 77644 -642 77714 6358
rect 77962 -642 78032 6358
rect 78280 -642 78350 6358
rect 78598 -642 78668 6358
rect 78916 -642 78986 6358
rect 79234 -642 79304 6358
rect 79552 -642 79622 6358
rect 79870 -642 79940 6358
rect 80188 -642 80258 6358
<< locali >>
rect 48576 15014 48672 15048
rect 80292 15014 80388 15048
rect 48576 14952 48610 15014
rect 80354 14952 80388 15014
rect 48640 14520 48706 14900
rect 48776 14520 49024 14900
rect 49094 14520 49342 14900
rect 49412 14520 49660 14900
rect 49730 14520 49978 14900
rect 50048 14520 50296 14900
rect 50366 14520 50614 14900
rect 50684 14520 50932 14900
rect 51002 14520 51250 14900
rect 51320 14520 51568 14900
rect 51638 14520 51886 14900
rect 51956 14520 52204 14900
rect 52274 14520 52522 14900
rect 52592 14520 52840 14900
rect 52910 14520 53158 14900
rect 53228 14520 53476 14900
rect 53546 14520 53794 14900
rect 53864 14520 54112 14900
rect 54182 14520 54430 14900
rect 54500 14520 54748 14900
rect 54818 14520 55066 14900
rect 55136 14520 55384 14900
rect 55454 14520 55702 14900
rect 55772 14520 56020 14900
rect 56090 14520 56338 14900
rect 56408 14520 56656 14900
rect 56726 14520 56974 14900
rect 57044 14520 57292 14900
rect 57362 14520 57610 14900
rect 57680 14520 57928 14900
rect 57998 14520 58246 14900
rect 58316 14520 58564 14900
rect 58634 14520 58882 14900
rect 58952 14520 59200 14900
rect 59270 14520 59518 14900
rect 59588 14520 59836 14900
rect 59906 14520 60154 14900
rect 60224 14520 60472 14900
rect 60542 14520 60790 14900
rect 60860 14520 61108 14900
rect 61178 14520 61426 14900
rect 61496 14520 61744 14900
rect 61814 14520 62062 14900
rect 62132 14520 62380 14900
rect 62450 14520 62698 14900
rect 62768 14520 63016 14900
rect 63086 14520 63334 14900
rect 63404 14520 63652 14900
rect 63722 14520 63970 14900
rect 64040 14520 64288 14900
rect 64358 14520 64606 14900
rect 64676 14520 64924 14900
rect 64994 14520 65242 14900
rect 65312 14520 65560 14900
rect 65630 14520 65878 14900
rect 65948 14520 66196 14900
rect 66266 14520 66514 14900
rect 66584 14520 66832 14900
rect 66902 14520 67150 14900
rect 67220 14520 67468 14900
rect 67538 14520 67786 14900
rect 67856 14520 68104 14900
rect 68174 14520 68422 14900
rect 68492 14520 68740 14900
rect 68810 14520 69058 14900
rect 69128 14520 69376 14900
rect 69446 14520 69694 14900
rect 69764 14520 70012 14900
rect 70082 14520 70330 14900
rect 70400 14520 70648 14900
rect 70718 14520 70966 14900
rect 71036 14520 71284 14900
rect 71354 14520 71602 14900
rect 71672 14520 71920 14900
rect 71990 14520 72238 14900
rect 72308 14520 72556 14900
rect 72626 14520 72874 14900
rect 72944 14520 73192 14900
rect 73262 14520 73510 14900
rect 73580 14520 73828 14900
rect 73898 14520 74146 14900
rect 74216 14520 74464 14900
rect 74534 14520 74782 14900
rect 74852 14520 75100 14900
rect 75170 14520 75418 14900
rect 75488 14520 75736 14900
rect 75806 14520 76054 14900
rect 76124 14520 76372 14900
rect 76442 14520 76690 14900
rect 76760 14520 77008 14900
rect 77078 14520 77326 14900
rect 77396 14520 77644 14900
rect 77714 14520 77962 14900
rect 78032 14520 78280 14900
rect 78350 14520 78598 14900
rect 78668 14520 78916 14900
rect 78986 14520 79234 14900
rect 79304 14520 79552 14900
rect 79622 14520 79870 14900
rect 79940 14520 80188 14900
rect 80258 14520 80280 14900
rect 48680 7054 48706 7080
rect 48776 7054 49024 7080
rect 49094 7054 49342 7080
rect 49412 7054 49660 7080
rect 49730 7054 49978 7080
rect 50048 7054 50296 7080
rect 50366 7054 50614 7080
rect 50684 7054 50932 7080
rect 51002 7054 51250 7080
rect 51320 7054 51568 7080
rect 51638 7054 51886 7080
rect 51956 7054 52204 7080
rect 52274 7054 52522 7080
rect 52592 7054 52840 7080
rect 52910 7054 53158 7080
rect 53228 7054 53476 7080
rect 53546 7054 53794 7080
rect 53864 7054 54112 7080
rect 54182 7054 54430 7080
rect 54500 7054 54748 7080
rect 54818 7054 55066 7080
rect 55136 7054 55384 7080
rect 55454 7054 55702 7080
rect 55772 7054 56020 7080
rect 56090 7054 56338 7080
rect 56408 7054 56656 7080
rect 56726 7054 56974 7080
rect 57044 7054 57292 7080
rect 57362 7054 57610 7080
rect 57680 7054 57928 7080
rect 57998 7054 58246 7080
rect 58316 7054 58564 7080
rect 58634 7054 58882 7080
rect 58952 7054 59200 7080
rect 59270 7054 59518 7080
rect 59588 7054 59836 7080
rect 59906 7054 60154 7080
rect 60224 7054 60472 7080
rect 60542 7054 60790 7080
rect 60860 7054 61108 7080
rect 61178 7054 61426 7080
rect 61496 7054 61744 7080
rect 61814 7054 62062 7080
rect 62132 7054 62380 7080
rect 62450 7054 62698 7080
rect 62768 7054 63016 7080
rect 63086 7054 63334 7080
rect 63404 7054 63652 7080
rect 63722 7054 63970 7080
rect 64040 7054 64288 7080
rect 64358 7054 64606 7080
rect 64676 7054 64924 7080
rect 64994 7054 65242 7080
rect 65312 7054 65560 7080
rect 65630 7054 65878 7080
rect 65948 7054 66196 7080
rect 66266 7054 66514 7080
rect 66584 7054 66832 7080
rect 66902 7054 67150 7080
rect 67220 7054 67468 7080
rect 67538 7054 67786 7080
rect 67856 7054 68104 7080
rect 68174 7054 68422 7080
rect 68492 7054 68740 7080
rect 68810 7054 69058 7080
rect 69128 7054 69376 7080
rect 69446 7054 69694 7080
rect 69764 7054 70012 7080
rect 70082 7054 70330 7080
rect 70400 7054 70648 7080
rect 70718 7054 70966 7080
rect 71036 7054 71284 7080
rect 71354 7054 71602 7080
rect 71672 7054 71920 7080
rect 71990 7054 72238 7080
rect 72308 7054 72556 7080
rect 72626 7054 72874 7080
rect 72944 7054 73192 7080
rect 73262 7054 73510 7080
rect 73580 7054 73828 7080
rect 73898 7054 74146 7080
rect 74216 7054 74464 7080
rect 74534 7054 74782 7080
rect 74852 7054 75100 7080
rect 75170 7054 75418 7080
rect 75488 7054 75736 7080
rect 75806 7054 76054 7080
rect 76124 7054 76372 7080
rect 76442 7054 76690 7080
rect 76760 7054 77008 7080
rect 77078 7054 77326 7080
rect 77396 7054 77644 7080
rect 77714 7054 77962 7080
rect 78032 7054 78280 7080
rect 78350 7054 78598 7080
rect 78668 7054 78916 7080
rect 78986 7054 79234 7080
rect 79304 7054 79552 7080
rect 79622 7054 79870 7080
rect 79940 7054 80188 7080
rect 80258 7054 80320 7080
rect 48680 6790 80320 7054
rect 48680 6700 48706 6790
rect 48776 6700 49024 6790
rect 49094 6700 49342 6790
rect 49412 6700 49660 6790
rect 49730 6700 49978 6790
rect 50048 6700 50296 6790
rect 50366 6700 50614 6790
rect 50684 6700 50932 6790
rect 51002 6700 51250 6790
rect 51320 6700 51568 6790
rect 51638 6700 51886 6790
rect 51956 6700 52204 6790
rect 52274 6700 52522 6790
rect 52592 6700 52840 6790
rect 52910 6700 53158 6790
rect 53228 6700 53476 6790
rect 53546 6700 53794 6790
rect 53864 6700 54112 6790
rect 54182 6700 54430 6790
rect 54500 6700 54748 6790
rect 54818 6700 55066 6790
rect 55136 6700 55384 6790
rect 55454 6700 55702 6790
rect 55772 6700 56020 6790
rect 56090 6700 56338 6790
rect 56408 6700 56656 6790
rect 56726 6700 56974 6790
rect 57044 6700 57292 6790
rect 57362 6700 57610 6790
rect 57680 6700 57928 6790
rect 57998 6700 58246 6790
rect 58316 6700 58564 6790
rect 58634 6700 58882 6790
rect 58952 6700 59200 6790
rect 59270 6700 59518 6790
rect 59588 6700 59836 6790
rect 59906 6700 60154 6790
rect 60224 6700 60472 6790
rect 60542 6700 60790 6790
rect 60860 6700 61108 6790
rect 61178 6700 61426 6790
rect 61496 6700 61744 6790
rect 61814 6700 62062 6790
rect 62132 6700 62380 6790
rect 62450 6700 62698 6790
rect 62768 6700 63016 6790
rect 63086 6700 63334 6790
rect 63404 6700 63652 6790
rect 63722 6700 63970 6790
rect 64040 6700 64288 6790
rect 64358 6700 64606 6790
rect 64676 6700 64924 6790
rect 64994 6700 65242 6790
rect 65312 6700 65560 6790
rect 65630 6700 65878 6790
rect 65948 6700 66196 6790
rect 66266 6700 66514 6790
rect 66584 6700 66832 6790
rect 66902 6700 67150 6790
rect 67220 6700 67468 6790
rect 67538 6700 67786 6790
rect 67856 6700 68104 6790
rect 68174 6700 68422 6790
rect 68492 6700 68740 6790
rect 68810 6700 69058 6790
rect 69128 6700 69376 6790
rect 69446 6700 69694 6790
rect 69764 6700 70012 6790
rect 70082 6700 70330 6790
rect 70400 6700 70648 6790
rect 70718 6700 70966 6790
rect 71036 6700 71284 6790
rect 71354 6700 71602 6790
rect 71672 6700 71920 6790
rect 71990 6700 72238 6790
rect 72308 6700 72556 6790
rect 72626 6700 72874 6790
rect 72944 6700 73192 6790
rect 73262 6700 73510 6790
rect 73580 6700 73828 6790
rect 73898 6700 74146 6790
rect 74216 6700 74464 6790
rect 74534 6700 74782 6790
rect 74852 6700 75100 6790
rect 75170 6700 75418 6790
rect 75488 6700 75736 6790
rect 75806 6700 76054 6790
rect 76124 6700 76372 6790
rect 76442 6700 76690 6790
rect 76760 6700 77008 6790
rect 77078 6700 77326 6790
rect 77396 6700 77644 6790
rect 77714 6700 77962 6790
rect 78032 6700 78280 6790
rect 78350 6700 78598 6790
rect 78668 6700 78916 6790
rect 78986 6700 79234 6790
rect 79304 6700 79552 6790
rect 79622 6700 79870 6790
rect 79940 6700 80188 6790
rect 80258 6700 80320 6790
rect 48680 -1074 48706 -880
rect 48776 -1074 49024 -880
rect 49094 -1074 49342 -880
rect 49412 -1074 49660 -880
rect 49730 -1074 49978 -880
rect 50048 -1074 50296 -880
rect 50366 -1074 50614 -880
rect 50684 -1074 50932 -880
rect 51002 -1074 51250 -880
rect 51320 -1074 51568 -880
rect 51638 -1074 51886 -880
rect 51956 -1074 52204 -880
rect 52274 -1074 52522 -880
rect 52592 -1074 52840 -880
rect 52910 -1074 53158 -880
rect 53228 -1074 53476 -880
rect 53546 -1074 53794 -880
rect 53864 -1074 54112 -880
rect 54182 -1074 54430 -880
rect 54500 -1074 54748 -880
rect 54818 -1074 55066 -880
rect 55136 -1074 55384 -880
rect 55454 -1074 55702 -880
rect 55772 -1074 56020 -880
rect 56090 -1074 56338 -880
rect 56408 -1074 56656 -880
rect 56726 -1074 56974 -880
rect 57044 -1074 57292 -880
rect 57362 -1074 57610 -880
rect 57680 -1074 57928 -880
rect 57998 -1074 58246 -880
rect 58316 -1074 58564 -880
rect 58634 -1074 58882 -880
rect 58952 -1074 59200 -880
rect 59270 -1074 59518 -880
rect 59588 -1074 59836 -880
rect 59906 -1074 60154 -880
rect 60224 -1074 60472 -880
rect 60542 -1074 60790 -880
rect 60860 -1074 61108 -880
rect 61178 -1074 61426 -880
rect 61496 -1074 61744 -880
rect 61814 -1074 62062 -880
rect 62132 -1074 62380 -880
rect 62450 -1074 62698 -880
rect 62768 -1074 63016 -880
rect 63086 -1074 63334 -880
rect 63404 -1074 63652 -880
rect 63722 -1074 63970 -880
rect 64040 -1074 64288 -880
rect 64358 -1074 64606 -880
rect 64676 -1074 64924 -880
rect 64994 -1074 65242 -880
rect 65312 -1074 65560 -880
rect 65630 -1074 65878 -880
rect 65948 -1074 66196 -880
rect 66266 -1074 66514 -880
rect 66584 -1074 66832 -880
rect 66902 -1074 67150 -880
rect 67220 -1074 67468 -880
rect 67538 -1074 67786 -880
rect 67856 -1074 68104 -880
rect 68174 -1074 68422 -880
rect 68492 -1074 68740 -880
rect 68810 -1074 69058 -880
rect 69128 -1074 69376 -880
rect 69446 -1074 69694 -880
rect 69764 -1074 70012 -880
rect 70082 -1074 70330 -880
rect 70400 -1074 70648 -880
rect 70718 -1074 70966 -880
rect 71036 -1074 71284 -880
rect 71354 -1074 71602 -880
rect 71672 -1074 71920 -880
rect 71990 -1074 72238 -880
rect 72308 -1074 72556 -880
rect 72626 -1074 72874 -880
rect 72944 -1074 73192 -880
rect 73262 -1074 73510 -880
rect 73580 -1074 73828 -880
rect 73898 -1074 74146 -880
rect 74216 -1074 74464 -880
rect 74534 -1074 74782 -880
rect 74852 -1074 75100 -880
rect 75170 -1074 75418 -880
rect 75488 -1074 75736 -880
rect 75806 -1074 76054 -880
rect 76124 -1074 76372 -880
rect 76442 -1074 76690 -880
rect 76760 -1074 77008 -880
rect 77078 -1074 77326 -880
rect 77396 -1074 77644 -880
rect 77714 -1074 77962 -880
rect 78032 -1074 78280 -880
rect 78350 -1074 78598 -880
rect 78668 -1074 78916 -880
rect 78986 -1074 79234 -880
rect 79304 -1074 79552 -880
rect 79622 -1074 79870 -880
rect 79940 -1074 80188 -880
rect 80258 -1074 80300 -880
rect 48680 -1080 80300 -1074
rect 48576 -1170 48610 -1108
rect 80354 -1170 80388 -1108
rect 48576 -1204 48672 -1170
rect 80292 -1204 80388 -1170
rect 48580 -1240 48640 -1204
<< viali >>
rect 48722 14503 48760 14900
rect 49040 14503 49078 14900
rect 49358 14503 49396 14900
rect 49676 14503 49714 14900
rect 49994 14503 50032 14900
rect 50312 14503 50350 14900
rect 50630 14503 50668 14900
rect 50948 14503 50986 14900
rect 51266 14503 51304 14900
rect 51584 14503 51622 14900
rect 51902 14503 51940 14900
rect 52220 14503 52258 14900
rect 52538 14503 52576 14900
rect 52856 14503 52894 14900
rect 53174 14503 53212 14900
rect 53492 14503 53530 14900
rect 53810 14503 53848 14900
rect 54128 14503 54166 14900
rect 54446 14503 54484 14900
rect 54764 14503 54802 14900
rect 55082 14503 55120 14900
rect 55400 14503 55438 14900
rect 55718 14503 55756 14900
rect 56036 14503 56074 14900
rect 56354 14503 56392 14900
rect 56672 14503 56710 14900
rect 56990 14503 57028 14900
rect 57308 14503 57346 14900
rect 57626 14503 57664 14900
rect 57944 14503 57982 14900
rect 58262 14503 58300 14900
rect 58580 14503 58618 14900
rect 58898 14503 58936 14900
rect 59216 14503 59254 14900
rect 59534 14503 59572 14900
rect 59852 14503 59890 14900
rect 60170 14503 60208 14900
rect 60488 14503 60526 14900
rect 60806 14503 60844 14900
rect 61124 14503 61162 14900
rect 61442 14503 61480 14900
rect 61760 14503 61798 14900
rect 62078 14503 62116 14900
rect 62396 14503 62434 14900
rect 62714 14503 62752 14900
rect 63032 14503 63070 14900
rect 63350 14503 63388 14900
rect 63668 14503 63706 14900
rect 63986 14503 64024 14900
rect 64304 14503 64342 14900
rect 64622 14503 64660 14900
rect 64940 14503 64978 14900
rect 65258 14503 65296 14900
rect 65576 14503 65614 14900
rect 65894 14503 65932 14900
rect 66212 14503 66250 14900
rect 66530 14503 66568 14900
rect 66848 14503 66886 14900
rect 67166 14503 67204 14900
rect 67484 14503 67522 14900
rect 67802 14503 67840 14900
rect 68120 14503 68158 14900
rect 68438 14503 68476 14900
rect 68756 14503 68794 14900
rect 69074 14503 69112 14900
rect 69392 14503 69430 14900
rect 69710 14503 69748 14900
rect 70028 14503 70066 14900
rect 70346 14503 70384 14900
rect 70664 14503 70702 14900
rect 70982 14503 71020 14900
rect 71300 14503 71338 14900
rect 71618 14503 71656 14900
rect 71936 14503 71974 14900
rect 72254 14503 72292 14900
rect 72572 14503 72610 14900
rect 72890 14503 72928 14900
rect 73208 14503 73246 14900
rect 73526 14503 73564 14900
rect 73844 14503 73882 14900
rect 74162 14503 74200 14900
rect 74480 14503 74518 14900
rect 74798 14503 74836 14900
rect 75116 14503 75154 14900
rect 75434 14503 75472 14900
rect 75752 14503 75790 14900
rect 76070 14503 76108 14900
rect 76388 14503 76426 14900
rect 76706 14503 76744 14900
rect 77024 14503 77062 14900
rect 77342 14503 77380 14900
rect 77660 14503 77698 14900
rect 77978 14503 78016 14900
rect 78296 14503 78334 14900
rect 78614 14503 78652 14900
rect 78932 14503 78970 14900
rect 79250 14503 79288 14900
rect 79568 14503 79606 14900
rect 79886 14503 79924 14900
rect 80204 14503 80242 14900
rect 48722 7072 48760 7469
rect 49040 7072 49078 7469
rect 49358 7072 49396 7469
rect 49676 7072 49714 7469
rect 49994 7072 50032 7469
rect 50312 7072 50350 7469
rect 50630 7072 50668 7469
rect 50948 7072 50986 7469
rect 51266 7072 51304 7469
rect 51584 7072 51622 7469
rect 51902 7072 51940 7469
rect 52220 7072 52258 7469
rect 52538 7072 52576 7469
rect 52856 7072 52894 7469
rect 53174 7072 53212 7469
rect 53492 7072 53530 7469
rect 53810 7072 53848 7469
rect 54128 7072 54166 7469
rect 54446 7072 54484 7469
rect 54764 7072 54802 7469
rect 55082 7072 55120 7469
rect 55400 7072 55438 7469
rect 55718 7072 55756 7469
rect 56036 7072 56074 7469
rect 56354 7072 56392 7469
rect 56672 7072 56710 7469
rect 56990 7072 57028 7469
rect 57308 7072 57346 7469
rect 57626 7072 57664 7469
rect 57944 7072 57982 7469
rect 58262 7072 58300 7469
rect 58580 7072 58618 7469
rect 58898 7072 58936 7469
rect 59216 7072 59254 7469
rect 59534 7072 59572 7469
rect 59852 7072 59890 7469
rect 60170 7072 60208 7469
rect 60488 7072 60526 7469
rect 60806 7072 60844 7469
rect 61124 7072 61162 7469
rect 61442 7072 61480 7469
rect 61760 7072 61798 7469
rect 62078 7072 62116 7469
rect 62396 7072 62434 7469
rect 62714 7072 62752 7469
rect 63032 7072 63070 7469
rect 63350 7072 63388 7469
rect 63668 7072 63706 7469
rect 63986 7072 64024 7469
rect 64304 7072 64342 7469
rect 64622 7072 64660 7469
rect 64940 7072 64978 7469
rect 65258 7072 65296 7469
rect 65576 7072 65614 7469
rect 65894 7072 65932 7469
rect 66212 7072 66250 7469
rect 66530 7072 66568 7469
rect 66848 7072 66886 7469
rect 67166 7072 67204 7469
rect 67484 7072 67522 7469
rect 67802 7072 67840 7469
rect 68120 7072 68158 7469
rect 68438 7072 68476 7469
rect 68756 7072 68794 7469
rect 69074 7072 69112 7469
rect 69392 7072 69430 7469
rect 69710 7072 69748 7469
rect 70028 7072 70066 7469
rect 70346 7072 70384 7469
rect 70664 7072 70702 7469
rect 70982 7072 71020 7469
rect 71300 7072 71338 7469
rect 71618 7072 71656 7469
rect 71936 7072 71974 7469
rect 72254 7072 72292 7469
rect 72572 7072 72610 7469
rect 72890 7072 72928 7469
rect 73208 7072 73246 7469
rect 73526 7072 73564 7469
rect 73844 7072 73882 7469
rect 74162 7072 74200 7469
rect 74480 7072 74518 7469
rect 74798 7072 74836 7469
rect 75116 7072 75154 7469
rect 75434 7072 75472 7469
rect 75752 7072 75790 7469
rect 76070 7072 76108 7469
rect 76388 7072 76426 7469
rect 76706 7072 76744 7469
rect 77024 7072 77062 7469
rect 77342 7072 77380 7469
rect 77660 7072 77698 7469
rect 77978 7072 78016 7469
rect 78296 7072 78334 7469
rect 78614 7072 78652 7469
rect 78932 7072 78970 7469
rect 79250 7072 79288 7469
rect 79568 7072 79606 7469
rect 79886 7072 79924 7469
rect 80204 7072 80242 7469
rect 48722 6375 48760 6772
rect 49040 6375 49078 6772
rect 49358 6375 49396 6772
rect 49676 6375 49714 6772
rect 49994 6375 50032 6772
rect 50312 6375 50350 6772
rect 50630 6375 50668 6772
rect 50948 6375 50986 6772
rect 51266 6375 51304 6772
rect 51584 6375 51622 6772
rect 51902 6375 51940 6772
rect 52220 6375 52258 6772
rect 52538 6375 52576 6772
rect 52856 6375 52894 6772
rect 53174 6375 53212 6772
rect 53492 6375 53530 6772
rect 53810 6375 53848 6772
rect 54128 6375 54166 6772
rect 54446 6375 54484 6772
rect 54764 6375 54802 6772
rect 55082 6375 55120 6772
rect 55400 6375 55438 6772
rect 55718 6375 55756 6772
rect 56036 6375 56074 6772
rect 56354 6375 56392 6772
rect 56672 6375 56710 6772
rect 56990 6375 57028 6772
rect 57308 6375 57346 6772
rect 57626 6375 57664 6772
rect 57944 6375 57982 6772
rect 58262 6375 58300 6772
rect 58580 6375 58618 6772
rect 58898 6375 58936 6772
rect 59216 6375 59254 6772
rect 59534 6375 59572 6772
rect 59852 6375 59890 6772
rect 60170 6375 60208 6772
rect 60488 6375 60526 6772
rect 60806 6375 60844 6772
rect 61124 6375 61162 6772
rect 61442 6375 61480 6772
rect 61760 6375 61798 6772
rect 62078 6375 62116 6772
rect 62396 6375 62434 6772
rect 62714 6375 62752 6772
rect 63032 6375 63070 6772
rect 63350 6375 63388 6772
rect 63668 6375 63706 6772
rect 63986 6375 64024 6772
rect 64304 6375 64342 6772
rect 64622 6375 64660 6772
rect 64940 6375 64978 6772
rect 65258 6375 65296 6772
rect 65576 6375 65614 6772
rect 65894 6375 65932 6772
rect 66212 6375 66250 6772
rect 66530 6375 66568 6772
rect 66848 6375 66886 6772
rect 67166 6375 67204 6772
rect 67484 6375 67522 6772
rect 67802 6375 67840 6772
rect 68120 6375 68158 6772
rect 68438 6375 68476 6772
rect 68756 6375 68794 6772
rect 69074 6375 69112 6772
rect 69392 6375 69430 6772
rect 69710 6375 69748 6772
rect 70028 6375 70066 6772
rect 70346 6375 70384 6772
rect 70664 6375 70702 6772
rect 70982 6375 71020 6772
rect 71300 6375 71338 6772
rect 71618 6375 71656 6772
rect 71936 6375 71974 6772
rect 72254 6375 72292 6772
rect 72572 6375 72610 6772
rect 72890 6375 72928 6772
rect 73208 6375 73246 6772
rect 73526 6375 73564 6772
rect 73844 6375 73882 6772
rect 74162 6375 74200 6772
rect 74480 6375 74518 6772
rect 74798 6375 74836 6772
rect 75116 6375 75154 6772
rect 75434 6375 75472 6772
rect 75752 6375 75790 6772
rect 76070 6375 76108 6772
rect 76388 6375 76426 6772
rect 76706 6375 76744 6772
rect 77024 6375 77062 6772
rect 77342 6375 77380 6772
rect 77660 6375 77698 6772
rect 77978 6375 78016 6772
rect 78296 6375 78334 6772
rect 78614 6375 78652 6772
rect 78932 6375 78970 6772
rect 79250 6375 79288 6772
rect 79568 6375 79606 6772
rect 79886 6375 79924 6772
rect 80204 6375 80242 6772
rect 48722 -1056 48760 -659
rect 49040 -1056 49078 -659
rect 49358 -1056 49396 -659
rect 49676 -1056 49714 -659
rect 49994 -1056 50032 -659
rect 50312 -1056 50350 -659
rect 50630 -1056 50668 -659
rect 50948 -1056 50986 -659
rect 51266 -1056 51304 -659
rect 51584 -1056 51622 -659
rect 51902 -1056 51940 -659
rect 52220 -1056 52258 -659
rect 52538 -1056 52576 -659
rect 52856 -1056 52894 -659
rect 53174 -1056 53212 -659
rect 53492 -1056 53530 -659
rect 53810 -1056 53848 -659
rect 54128 -1056 54166 -659
rect 54446 -1056 54484 -659
rect 54764 -1056 54802 -659
rect 55082 -1056 55120 -659
rect 55400 -1056 55438 -659
rect 55718 -1056 55756 -659
rect 56036 -1056 56074 -659
rect 56354 -1056 56392 -659
rect 56672 -1056 56710 -659
rect 56990 -1056 57028 -659
rect 57308 -1056 57346 -659
rect 57626 -1056 57664 -659
rect 57944 -1056 57982 -659
rect 58262 -1056 58300 -659
rect 58580 -1056 58618 -659
rect 58898 -1056 58936 -659
rect 59216 -1056 59254 -659
rect 59534 -1056 59572 -659
rect 59852 -1056 59890 -659
rect 60170 -1056 60208 -659
rect 60488 -1056 60526 -659
rect 60806 -1056 60844 -659
rect 61124 -1056 61162 -659
rect 61442 -1056 61480 -659
rect 61760 -1056 61798 -659
rect 62078 -1056 62116 -659
rect 62396 -1056 62434 -659
rect 62714 -1056 62752 -659
rect 63032 -1056 63070 -659
rect 63350 -1056 63388 -659
rect 63668 -1056 63706 -659
rect 63986 -1056 64024 -659
rect 64304 -1056 64342 -659
rect 64622 -1056 64660 -659
rect 64940 -1056 64978 -659
rect 65258 -1056 65296 -659
rect 65576 -1056 65614 -659
rect 65894 -1056 65932 -659
rect 66212 -1056 66250 -659
rect 66530 -1056 66568 -659
rect 66848 -1056 66886 -659
rect 67166 -1056 67204 -659
rect 67484 -1056 67522 -659
rect 67802 -1056 67840 -659
rect 68120 -1056 68158 -659
rect 68438 -1056 68476 -659
rect 68756 -1056 68794 -659
rect 69074 -1056 69112 -659
rect 69392 -1056 69430 -659
rect 69710 -1056 69748 -659
rect 70028 -1056 70066 -659
rect 70346 -1056 70384 -659
rect 70664 -1056 70702 -659
rect 70982 -1056 71020 -659
rect 71300 -1056 71338 -659
rect 71618 -1056 71656 -659
rect 71936 -1056 71974 -659
rect 72254 -1056 72292 -659
rect 72572 -1056 72610 -659
rect 72890 -1056 72928 -659
rect 73208 -1056 73246 -659
rect 73526 -1056 73564 -659
rect 73844 -1056 73882 -659
rect 74162 -1056 74200 -659
rect 74480 -1056 74518 -659
rect 74798 -1056 74836 -659
rect 75116 -1056 75154 -659
rect 75434 -1056 75472 -659
rect 75752 -1056 75790 -659
rect 76070 -1056 76108 -659
rect 76388 -1056 76426 -659
rect 76706 -1056 76744 -659
rect 77024 -1056 77062 -659
rect 77342 -1056 77380 -659
rect 77660 -1056 77698 -659
rect 77978 -1056 78016 -659
rect 78296 -1056 78334 -659
rect 78614 -1056 78652 -659
rect 78932 -1056 78970 -659
rect 79250 -1056 79288 -659
rect 79568 -1056 79606 -659
rect 79886 -1056 79924 -659
rect 80204 -1056 80242 -659
<< metal1 >>
rect 48716 14900 48766 14912
rect 48716 14503 48722 14900
rect 48760 14503 48766 14900
rect 48716 14491 48766 14503
rect 49034 14900 49084 14912
rect 49034 14503 49040 14900
rect 49078 14503 49084 14900
rect 49034 14491 49084 14503
rect 49352 14900 49402 14912
rect 49352 14503 49358 14900
rect 49396 14503 49402 14900
rect 49352 14491 49402 14503
rect 49670 14900 49720 14912
rect 49670 14503 49676 14900
rect 49714 14503 49720 14900
rect 49670 14491 49720 14503
rect 49988 14900 50038 14912
rect 49988 14503 49994 14900
rect 50032 14503 50038 14900
rect 49988 14491 50038 14503
rect 50306 14900 50356 14912
rect 50306 14503 50312 14900
rect 50350 14503 50356 14900
rect 50306 14491 50356 14503
rect 50624 14900 50674 14912
rect 50624 14503 50630 14900
rect 50668 14503 50674 14900
rect 50624 14491 50674 14503
rect 50942 14900 50992 14912
rect 50942 14503 50948 14900
rect 50986 14503 50992 14900
rect 50942 14491 50992 14503
rect 51260 14900 51310 14912
rect 51260 14503 51266 14900
rect 51304 14503 51310 14900
rect 51260 14491 51310 14503
rect 51578 14900 51628 14912
rect 51578 14503 51584 14900
rect 51622 14503 51628 14900
rect 51578 14491 51628 14503
rect 51896 14900 51946 14912
rect 51896 14503 51902 14900
rect 51940 14503 51946 14900
rect 51896 14491 51946 14503
rect 52214 14900 52264 14912
rect 52214 14503 52220 14900
rect 52258 14503 52264 14900
rect 52214 14491 52264 14503
rect 52532 14900 52582 14912
rect 52532 14503 52538 14900
rect 52576 14503 52582 14900
rect 52532 14491 52582 14503
rect 52850 14900 52900 14912
rect 52850 14503 52856 14900
rect 52894 14503 52900 14900
rect 52850 14491 52900 14503
rect 53168 14900 53218 14912
rect 53168 14503 53174 14900
rect 53212 14503 53218 14900
rect 53168 14491 53218 14503
rect 53486 14900 53536 14912
rect 53486 14503 53492 14900
rect 53530 14503 53536 14900
rect 53486 14491 53536 14503
rect 53804 14900 53854 14912
rect 53804 14503 53810 14900
rect 53848 14503 53854 14900
rect 53804 14491 53854 14503
rect 54122 14900 54172 14912
rect 54122 14503 54128 14900
rect 54166 14503 54172 14900
rect 54122 14491 54172 14503
rect 54440 14900 54490 14912
rect 54440 14503 54446 14900
rect 54484 14503 54490 14900
rect 54440 14491 54490 14503
rect 54758 14900 54808 14912
rect 54758 14503 54764 14900
rect 54802 14503 54808 14900
rect 54758 14491 54808 14503
rect 55076 14900 55126 14912
rect 55076 14503 55082 14900
rect 55120 14503 55126 14900
rect 55076 14491 55126 14503
rect 55394 14900 55444 14912
rect 55394 14503 55400 14900
rect 55438 14503 55444 14900
rect 55394 14491 55444 14503
rect 55712 14900 55762 14912
rect 55712 14503 55718 14900
rect 55756 14503 55762 14900
rect 55712 14491 55762 14503
rect 56030 14900 56080 14912
rect 56030 14503 56036 14900
rect 56074 14503 56080 14900
rect 56030 14491 56080 14503
rect 56348 14900 56398 14912
rect 56348 14503 56354 14900
rect 56392 14503 56398 14900
rect 56348 14491 56398 14503
rect 56666 14900 56716 14912
rect 56666 14503 56672 14900
rect 56710 14503 56716 14900
rect 56666 14491 56716 14503
rect 56984 14900 57034 14912
rect 56984 14503 56990 14900
rect 57028 14503 57034 14900
rect 56984 14491 57034 14503
rect 57302 14900 57352 14912
rect 57302 14503 57308 14900
rect 57346 14503 57352 14900
rect 57302 14491 57352 14503
rect 57620 14900 57670 14912
rect 57620 14503 57626 14900
rect 57664 14503 57670 14900
rect 57620 14491 57670 14503
rect 57938 14900 57988 14912
rect 57938 14503 57944 14900
rect 57982 14503 57988 14900
rect 57938 14491 57988 14503
rect 58256 14900 58306 14912
rect 58256 14503 58262 14900
rect 58300 14503 58306 14900
rect 58256 14491 58306 14503
rect 58574 14900 58624 14912
rect 58574 14503 58580 14900
rect 58618 14503 58624 14900
rect 58574 14491 58624 14503
rect 58892 14900 58942 14912
rect 58892 14503 58898 14900
rect 58936 14503 58942 14900
rect 58892 14491 58942 14503
rect 59210 14900 59260 14912
rect 59210 14503 59216 14900
rect 59254 14503 59260 14900
rect 59210 14491 59260 14503
rect 59528 14900 59578 14912
rect 59528 14503 59534 14900
rect 59572 14503 59578 14900
rect 59528 14491 59578 14503
rect 59846 14900 59896 14912
rect 59846 14503 59852 14900
rect 59890 14503 59896 14900
rect 59846 14491 59896 14503
rect 60164 14900 60214 14912
rect 60164 14503 60170 14900
rect 60208 14503 60214 14900
rect 60164 14491 60214 14503
rect 60482 14900 60532 14912
rect 60482 14503 60488 14900
rect 60526 14503 60532 14900
rect 60482 14491 60532 14503
rect 60800 14900 60850 14912
rect 60800 14503 60806 14900
rect 60844 14503 60850 14900
rect 60800 14491 60850 14503
rect 61118 14900 61168 14912
rect 61118 14503 61124 14900
rect 61162 14503 61168 14900
rect 61118 14491 61168 14503
rect 61436 14900 61486 14912
rect 61436 14503 61442 14900
rect 61480 14503 61486 14900
rect 61436 14491 61486 14503
rect 61754 14900 61804 14912
rect 61754 14503 61760 14900
rect 61798 14503 61804 14900
rect 61754 14491 61804 14503
rect 62072 14900 62122 14912
rect 62072 14503 62078 14900
rect 62116 14503 62122 14900
rect 62072 14491 62122 14503
rect 62390 14900 62440 14912
rect 62390 14503 62396 14900
rect 62434 14503 62440 14900
rect 62390 14491 62440 14503
rect 62708 14900 62758 14912
rect 62708 14503 62714 14900
rect 62752 14503 62758 14900
rect 62708 14491 62758 14503
rect 63026 14900 63076 14912
rect 63026 14503 63032 14900
rect 63070 14503 63076 14900
rect 63026 14491 63076 14503
rect 63344 14900 63394 14912
rect 63344 14503 63350 14900
rect 63388 14503 63394 14900
rect 63344 14491 63394 14503
rect 63662 14900 63712 14912
rect 63662 14503 63668 14900
rect 63706 14503 63712 14900
rect 63662 14491 63712 14503
rect 63980 14900 64030 14912
rect 63980 14503 63986 14900
rect 64024 14503 64030 14900
rect 63980 14491 64030 14503
rect 64298 14900 64348 14912
rect 64298 14503 64304 14900
rect 64342 14503 64348 14900
rect 64298 14491 64348 14503
rect 64616 14900 64666 14912
rect 64616 14503 64622 14900
rect 64660 14503 64666 14900
rect 64616 14491 64666 14503
rect 64934 14900 64984 14912
rect 64934 14503 64940 14900
rect 64978 14503 64984 14900
rect 64934 14491 64984 14503
rect 65252 14900 65302 14912
rect 65252 14503 65258 14900
rect 65296 14503 65302 14900
rect 65252 14491 65302 14503
rect 65570 14900 65620 14912
rect 65570 14503 65576 14900
rect 65614 14503 65620 14900
rect 65570 14491 65620 14503
rect 65888 14900 65938 14912
rect 65888 14503 65894 14900
rect 65932 14503 65938 14900
rect 65888 14491 65938 14503
rect 66206 14900 66256 14912
rect 66206 14503 66212 14900
rect 66250 14503 66256 14900
rect 66206 14491 66256 14503
rect 66524 14900 66574 14912
rect 66524 14503 66530 14900
rect 66568 14503 66574 14900
rect 66524 14491 66574 14503
rect 66842 14900 66892 14912
rect 66842 14503 66848 14900
rect 66886 14503 66892 14900
rect 66842 14491 66892 14503
rect 67160 14900 67210 14912
rect 67160 14503 67166 14900
rect 67204 14503 67210 14900
rect 67160 14491 67210 14503
rect 67478 14900 67528 14912
rect 67478 14503 67484 14900
rect 67522 14503 67528 14900
rect 67478 14491 67528 14503
rect 67796 14900 67846 14912
rect 67796 14503 67802 14900
rect 67840 14503 67846 14900
rect 67796 14491 67846 14503
rect 68114 14900 68164 14912
rect 68114 14503 68120 14900
rect 68158 14503 68164 14900
rect 68114 14491 68164 14503
rect 68432 14900 68482 14912
rect 68432 14503 68438 14900
rect 68476 14503 68482 14900
rect 68432 14491 68482 14503
rect 68750 14900 68800 14912
rect 68750 14503 68756 14900
rect 68794 14503 68800 14900
rect 68750 14491 68800 14503
rect 69068 14900 69118 14912
rect 69068 14503 69074 14900
rect 69112 14503 69118 14900
rect 69068 14491 69118 14503
rect 69386 14900 69436 14912
rect 69386 14503 69392 14900
rect 69430 14503 69436 14900
rect 69386 14491 69436 14503
rect 69704 14900 69754 14912
rect 69704 14503 69710 14900
rect 69748 14503 69754 14900
rect 69704 14491 69754 14503
rect 70022 14900 70072 14912
rect 70022 14503 70028 14900
rect 70066 14503 70072 14900
rect 70022 14491 70072 14503
rect 70340 14900 70390 14912
rect 70340 14503 70346 14900
rect 70384 14503 70390 14900
rect 70340 14491 70390 14503
rect 70658 14900 70708 14912
rect 70658 14503 70664 14900
rect 70702 14503 70708 14900
rect 70658 14491 70708 14503
rect 70976 14900 71026 14912
rect 70976 14503 70982 14900
rect 71020 14503 71026 14900
rect 70976 14491 71026 14503
rect 71294 14900 71344 14912
rect 71294 14503 71300 14900
rect 71338 14503 71344 14900
rect 71294 14491 71344 14503
rect 71612 14900 71662 14912
rect 71612 14503 71618 14900
rect 71656 14503 71662 14900
rect 71612 14491 71662 14503
rect 71930 14900 71980 14912
rect 71930 14503 71936 14900
rect 71974 14503 71980 14900
rect 71930 14491 71980 14503
rect 72248 14900 72298 14912
rect 72248 14503 72254 14900
rect 72292 14503 72298 14900
rect 72248 14491 72298 14503
rect 72566 14900 72616 14912
rect 72566 14503 72572 14900
rect 72610 14503 72616 14900
rect 72566 14491 72616 14503
rect 72884 14900 72934 14912
rect 72884 14503 72890 14900
rect 72928 14503 72934 14900
rect 72884 14491 72934 14503
rect 73202 14900 73252 14912
rect 73202 14503 73208 14900
rect 73246 14503 73252 14900
rect 73202 14491 73252 14503
rect 73520 14900 73570 14912
rect 73520 14503 73526 14900
rect 73564 14503 73570 14900
rect 73520 14491 73570 14503
rect 73838 14900 73888 14912
rect 73838 14503 73844 14900
rect 73882 14503 73888 14900
rect 73838 14491 73888 14503
rect 74156 14900 74206 14912
rect 74156 14503 74162 14900
rect 74200 14503 74206 14900
rect 74156 14491 74206 14503
rect 74474 14900 74524 14912
rect 74474 14503 74480 14900
rect 74518 14503 74524 14900
rect 74474 14491 74524 14503
rect 74792 14900 74842 14912
rect 74792 14503 74798 14900
rect 74836 14503 74842 14900
rect 74792 14491 74842 14503
rect 75110 14900 75160 14912
rect 75110 14503 75116 14900
rect 75154 14503 75160 14900
rect 75110 14491 75160 14503
rect 75428 14900 75478 14912
rect 75428 14503 75434 14900
rect 75472 14503 75478 14900
rect 75428 14491 75478 14503
rect 75746 14900 75796 14912
rect 75746 14503 75752 14900
rect 75790 14503 75796 14900
rect 75746 14491 75796 14503
rect 76064 14900 76114 14912
rect 76064 14503 76070 14900
rect 76108 14503 76114 14900
rect 76064 14491 76114 14503
rect 76382 14900 76432 14912
rect 76382 14503 76388 14900
rect 76426 14503 76432 14900
rect 76382 14491 76432 14503
rect 76700 14900 76750 14912
rect 76700 14503 76706 14900
rect 76744 14503 76750 14900
rect 76700 14491 76750 14503
rect 77018 14900 77068 14912
rect 77018 14503 77024 14900
rect 77062 14503 77068 14900
rect 77018 14491 77068 14503
rect 77336 14900 77386 14912
rect 77336 14503 77342 14900
rect 77380 14503 77386 14900
rect 77336 14491 77386 14503
rect 77654 14900 77704 14912
rect 77654 14503 77660 14900
rect 77698 14503 77704 14900
rect 77654 14491 77704 14503
rect 77972 14900 78022 14912
rect 77972 14503 77978 14900
rect 78016 14503 78022 14900
rect 77972 14491 78022 14503
rect 78290 14900 78340 14912
rect 78290 14503 78296 14900
rect 78334 14503 78340 14900
rect 78290 14491 78340 14503
rect 78608 14900 78658 14912
rect 78608 14503 78614 14900
rect 78652 14503 78658 14900
rect 78608 14491 78658 14503
rect 78926 14900 78976 14912
rect 78926 14503 78932 14900
rect 78970 14503 78976 14900
rect 78926 14491 78976 14503
rect 79244 14900 79294 14912
rect 79244 14503 79250 14900
rect 79288 14503 79294 14900
rect 79244 14491 79294 14503
rect 79562 14900 79612 14912
rect 79562 14503 79568 14900
rect 79606 14503 79612 14900
rect 79562 14491 79612 14503
rect 79880 14900 79930 14912
rect 79880 14503 79886 14900
rect 79924 14503 79930 14900
rect 79880 14491 79930 14503
rect 80198 14900 80248 14912
rect 80198 14503 80204 14900
rect 80242 14503 80248 14900
rect 80198 14491 80248 14503
rect 48716 7469 48766 7481
rect 48716 7072 48722 7469
rect 48760 7072 48766 7469
rect 48716 7060 48766 7072
rect 49034 7469 49084 7481
rect 49034 7072 49040 7469
rect 49078 7072 49084 7469
rect 49034 7060 49084 7072
rect 49352 7469 49402 7481
rect 49352 7072 49358 7469
rect 49396 7072 49402 7469
rect 49352 7060 49402 7072
rect 49670 7469 49720 7481
rect 49670 7072 49676 7469
rect 49714 7072 49720 7469
rect 49670 7060 49720 7072
rect 49988 7469 50038 7481
rect 49988 7072 49994 7469
rect 50032 7072 50038 7469
rect 49988 7060 50038 7072
rect 50306 7469 50356 7481
rect 50306 7072 50312 7469
rect 50350 7072 50356 7469
rect 50306 7060 50356 7072
rect 50624 7469 50674 7481
rect 50624 7072 50630 7469
rect 50668 7072 50674 7469
rect 50624 7060 50674 7072
rect 50942 7469 50992 7481
rect 50942 7072 50948 7469
rect 50986 7072 50992 7469
rect 50942 7060 50992 7072
rect 51260 7469 51310 7481
rect 51260 7072 51266 7469
rect 51304 7072 51310 7469
rect 51260 7060 51310 7072
rect 51578 7469 51628 7481
rect 51578 7072 51584 7469
rect 51622 7072 51628 7469
rect 51578 7060 51628 7072
rect 51896 7469 51946 7481
rect 51896 7072 51902 7469
rect 51940 7072 51946 7469
rect 51896 7060 51946 7072
rect 52214 7469 52264 7481
rect 52214 7072 52220 7469
rect 52258 7072 52264 7469
rect 52214 7060 52264 7072
rect 52532 7469 52582 7481
rect 52532 7072 52538 7469
rect 52576 7072 52582 7469
rect 52532 7060 52582 7072
rect 52850 7469 52900 7481
rect 52850 7072 52856 7469
rect 52894 7072 52900 7469
rect 52850 7060 52900 7072
rect 53168 7469 53218 7481
rect 53168 7072 53174 7469
rect 53212 7072 53218 7469
rect 53168 7060 53218 7072
rect 53486 7469 53536 7481
rect 53486 7072 53492 7469
rect 53530 7072 53536 7469
rect 53486 7060 53536 7072
rect 53804 7469 53854 7481
rect 53804 7072 53810 7469
rect 53848 7072 53854 7469
rect 53804 7060 53854 7072
rect 54122 7469 54172 7481
rect 54122 7072 54128 7469
rect 54166 7072 54172 7469
rect 54122 7060 54172 7072
rect 54440 7469 54490 7481
rect 54440 7072 54446 7469
rect 54484 7072 54490 7469
rect 54440 7060 54490 7072
rect 54758 7469 54808 7481
rect 54758 7072 54764 7469
rect 54802 7072 54808 7469
rect 54758 7060 54808 7072
rect 55076 7469 55126 7481
rect 55076 7072 55082 7469
rect 55120 7072 55126 7469
rect 55076 7060 55126 7072
rect 55394 7469 55444 7481
rect 55394 7072 55400 7469
rect 55438 7072 55444 7469
rect 55394 7060 55444 7072
rect 55712 7469 55762 7481
rect 55712 7072 55718 7469
rect 55756 7072 55762 7469
rect 55712 7060 55762 7072
rect 56030 7469 56080 7481
rect 56030 7072 56036 7469
rect 56074 7072 56080 7469
rect 56030 7060 56080 7072
rect 56348 7469 56398 7481
rect 56348 7072 56354 7469
rect 56392 7072 56398 7469
rect 56348 7060 56398 7072
rect 56666 7469 56716 7481
rect 56666 7072 56672 7469
rect 56710 7072 56716 7469
rect 56666 7060 56716 7072
rect 56984 7469 57034 7481
rect 56984 7072 56990 7469
rect 57028 7072 57034 7469
rect 56984 7060 57034 7072
rect 57302 7469 57352 7481
rect 57302 7072 57308 7469
rect 57346 7072 57352 7469
rect 57302 7060 57352 7072
rect 57620 7469 57670 7481
rect 57620 7072 57626 7469
rect 57664 7072 57670 7469
rect 57620 7060 57670 7072
rect 57938 7469 57988 7481
rect 57938 7072 57944 7469
rect 57982 7072 57988 7469
rect 57938 7060 57988 7072
rect 58256 7469 58306 7481
rect 58256 7072 58262 7469
rect 58300 7072 58306 7469
rect 58256 7060 58306 7072
rect 58574 7469 58624 7481
rect 58574 7072 58580 7469
rect 58618 7072 58624 7469
rect 58574 7060 58624 7072
rect 58892 7469 58942 7481
rect 58892 7072 58898 7469
rect 58936 7072 58942 7469
rect 58892 7060 58942 7072
rect 59210 7469 59260 7481
rect 59210 7072 59216 7469
rect 59254 7072 59260 7469
rect 59210 7060 59260 7072
rect 59528 7469 59578 7481
rect 59528 7072 59534 7469
rect 59572 7072 59578 7469
rect 59528 7060 59578 7072
rect 59846 7469 59896 7481
rect 59846 7072 59852 7469
rect 59890 7072 59896 7469
rect 59846 7060 59896 7072
rect 60164 7469 60214 7481
rect 60164 7072 60170 7469
rect 60208 7072 60214 7469
rect 60164 7060 60214 7072
rect 60482 7469 60532 7481
rect 60482 7072 60488 7469
rect 60526 7072 60532 7469
rect 60482 7060 60532 7072
rect 60800 7469 60850 7481
rect 60800 7072 60806 7469
rect 60844 7072 60850 7469
rect 60800 7060 60850 7072
rect 61118 7469 61168 7481
rect 61118 7072 61124 7469
rect 61162 7072 61168 7469
rect 61118 7060 61168 7072
rect 61436 7469 61486 7481
rect 61436 7072 61442 7469
rect 61480 7072 61486 7469
rect 61436 7060 61486 7072
rect 61754 7469 61804 7481
rect 61754 7072 61760 7469
rect 61798 7072 61804 7469
rect 61754 7060 61804 7072
rect 62072 7469 62122 7481
rect 62072 7072 62078 7469
rect 62116 7072 62122 7469
rect 62072 7060 62122 7072
rect 62390 7469 62440 7481
rect 62390 7072 62396 7469
rect 62434 7072 62440 7469
rect 62390 7060 62440 7072
rect 62708 7469 62758 7481
rect 62708 7072 62714 7469
rect 62752 7072 62758 7469
rect 62708 7060 62758 7072
rect 63026 7469 63076 7481
rect 63026 7072 63032 7469
rect 63070 7072 63076 7469
rect 63026 7060 63076 7072
rect 63344 7469 63394 7481
rect 63344 7072 63350 7469
rect 63388 7072 63394 7469
rect 63344 7060 63394 7072
rect 63662 7469 63712 7481
rect 63662 7072 63668 7469
rect 63706 7072 63712 7469
rect 63662 7060 63712 7072
rect 63980 7469 64030 7481
rect 63980 7072 63986 7469
rect 64024 7072 64030 7469
rect 63980 7060 64030 7072
rect 64298 7469 64348 7481
rect 64298 7072 64304 7469
rect 64342 7072 64348 7469
rect 64298 7060 64348 7072
rect 64616 7469 64666 7481
rect 64616 7072 64622 7469
rect 64660 7072 64666 7469
rect 64616 7060 64666 7072
rect 64934 7469 64984 7481
rect 64934 7072 64940 7469
rect 64978 7072 64984 7469
rect 64934 7060 64984 7072
rect 65252 7469 65302 7481
rect 65252 7072 65258 7469
rect 65296 7072 65302 7469
rect 65252 7060 65302 7072
rect 65570 7469 65620 7481
rect 65570 7072 65576 7469
rect 65614 7072 65620 7469
rect 65570 7060 65620 7072
rect 65888 7469 65938 7481
rect 65888 7072 65894 7469
rect 65932 7072 65938 7469
rect 65888 7060 65938 7072
rect 66206 7469 66256 7481
rect 66206 7072 66212 7469
rect 66250 7072 66256 7469
rect 66206 7060 66256 7072
rect 66524 7469 66574 7481
rect 66524 7072 66530 7469
rect 66568 7072 66574 7469
rect 66524 7060 66574 7072
rect 66842 7469 66892 7481
rect 66842 7072 66848 7469
rect 66886 7072 66892 7469
rect 66842 7060 66892 7072
rect 67160 7469 67210 7481
rect 67160 7072 67166 7469
rect 67204 7072 67210 7469
rect 67160 7060 67210 7072
rect 67478 7469 67528 7481
rect 67478 7072 67484 7469
rect 67522 7072 67528 7469
rect 67478 7060 67528 7072
rect 67796 7469 67846 7481
rect 67796 7072 67802 7469
rect 67840 7072 67846 7469
rect 67796 7060 67846 7072
rect 68114 7469 68164 7481
rect 68114 7072 68120 7469
rect 68158 7072 68164 7469
rect 68114 7060 68164 7072
rect 68432 7469 68482 7481
rect 68432 7072 68438 7469
rect 68476 7072 68482 7469
rect 68432 7060 68482 7072
rect 68750 7469 68800 7481
rect 68750 7072 68756 7469
rect 68794 7072 68800 7469
rect 68750 7060 68800 7072
rect 69068 7469 69118 7481
rect 69068 7072 69074 7469
rect 69112 7072 69118 7469
rect 69068 7060 69118 7072
rect 69386 7469 69436 7481
rect 69386 7072 69392 7469
rect 69430 7072 69436 7469
rect 69386 7060 69436 7072
rect 69704 7469 69754 7481
rect 69704 7072 69710 7469
rect 69748 7072 69754 7469
rect 69704 7060 69754 7072
rect 70022 7469 70072 7481
rect 70022 7072 70028 7469
rect 70066 7072 70072 7469
rect 70022 7060 70072 7072
rect 70340 7469 70390 7481
rect 70340 7072 70346 7469
rect 70384 7072 70390 7469
rect 70340 7060 70390 7072
rect 70658 7469 70708 7481
rect 70658 7072 70664 7469
rect 70702 7072 70708 7469
rect 70658 7060 70708 7072
rect 70976 7469 71026 7481
rect 70976 7072 70982 7469
rect 71020 7072 71026 7469
rect 70976 7060 71026 7072
rect 71294 7469 71344 7481
rect 71294 7072 71300 7469
rect 71338 7072 71344 7469
rect 71294 7060 71344 7072
rect 71612 7469 71662 7481
rect 71612 7072 71618 7469
rect 71656 7072 71662 7469
rect 71612 7060 71662 7072
rect 71930 7469 71980 7481
rect 71930 7072 71936 7469
rect 71974 7072 71980 7469
rect 71930 7060 71980 7072
rect 72248 7469 72298 7481
rect 72248 7072 72254 7469
rect 72292 7072 72298 7469
rect 72248 7060 72298 7072
rect 72566 7469 72616 7481
rect 72566 7072 72572 7469
rect 72610 7072 72616 7469
rect 72566 7060 72616 7072
rect 72884 7469 72934 7481
rect 72884 7072 72890 7469
rect 72928 7072 72934 7469
rect 72884 7060 72934 7072
rect 73202 7469 73252 7481
rect 73202 7072 73208 7469
rect 73246 7072 73252 7469
rect 73202 7060 73252 7072
rect 73520 7469 73570 7481
rect 73520 7072 73526 7469
rect 73564 7072 73570 7469
rect 73520 7060 73570 7072
rect 73838 7469 73888 7481
rect 73838 7072 73844 7469
rect 73882 7072 73888 7469
rect 73838 7060 73888 7072
rect 74156 7469 74206 7481
rect 74156 7072 74162 7469
rect 74200 7072 74206 7469
rect 74156 7060 74206 7072
rect 74474 7469 74524 7481
rect 74474 7072 74480 7469
rect 74518 7072 74524 7469
rect 74474 7060 74524 7072
rect 74792 7469 74842 7481
rect 74792 7072 74798 7469
rect 74836 7072 74842 7469
rect 74792 7060 74842 7072
rect 75110 7469 75160 7481
rect 75110 7072 75116 7469
rect 75154 7072 75160 7469
rect 75110 7060 75160 7072
rect 75428 7469 75478 7481
rect 75428 7072 75434 7469
rect 75472 7072 75478 7469
rect 75428 7060 75478 7072
rect 75746 7469 75796 7481
rect 75746 7072 75752 7469
rect 75790 7072 75796 7469
rect 75746 7060 75796 7072
rect 76064 7469 76114 7481
rect 76064 7072 76070 7469
rect 76108 7072 76114 7469
rect 76064 7060 76114 7072
rect 76382 7469 76432 7481
rect 76382 7072 76388 7469
rect 76426 7072 76432 7469
rect 76382 7060 76432 7072
rect 76700 7469 76750 7481
rect 76700 7072 76706 7469
rect 76744 7072 76750 7469
rect 76700 7060 76750 7072
rect 77018 7469 77068 7481
rect 77018 7072 77024 7469
rect 77062 7072 77068 7469
rect 77018 7060 77068 7072
rect 77336 7469 77386 7481
rect 77336 7072 77342 7469
rect 77380 7072 77386 7469
rect 77336 7060 77386 7072
rect 77654 7469 77704 7481
rect 77654 7072 77660 7469
rect 77698 7072 77704 7469
rect 77654 7060 77704 7072
rect 77972 7469 78022 7481
rect 77972 7072 77978 7469
rect 78016 7072 78022 7469
rect 77972 7060 78022 7072
rect 78290 7469 78340 7481
rect 78290 7072 78296 7469
rect 78334 7072 78340 7469
rect 78290 7060 78340 7072
rect 78608 7469 78658 7481
rect 78608 7072 78614 7469
rect 78652 7072 78658 7469
rect 78608 7060 78658 7072
rect 78926 7469 78976 7481
rect 78926 7072 78932 7469
rect 78970 7072 78976 7469
rect 78926 7060 78976 7072
rect 79244 7469 79294 7481
rect 79244 7072 79250 7469
rect 79288 7072 79294 7469
rect 79244 7060 79294 7072
rect 79562 7469 79612 7481
rect 79562 7072 79568 7469
rect 79606 7072 79612 7469
rect 79562 7060 79612 7072
rect 79880 7469 79930 7481
rect 79880 7072 79886 7469
rect 79924 7072 79930 7469
rect 79880 7060 79930 7072
rect 80198 7469 80248 7481
rect 80198 7072 80204 7469
rect 80242 7072 80248 7469
rect 80198 7060 80248 7072
rect 48716 6772 48766 6784
rect 48716 6375 48722 6772
rect 48760 6375 48766 6772
rect 48716 6363 48766 6375
rect 49034 6772 49084 6784
rect 49034 6375 49040 6772
rect 49078 6375 49084 6772
rect 49034 6363 49084 6375
rect 49352 6772 49402 6784
rect 49352 6375 49358 6772
rect 49396 6375 49402 6772
rect 49352 6363 49402 6375
rect 49670 6772 49720 6784
rect 49670 6375 49676 6772
rect 49714 6375 49720 6772
rect 49670 6363 49720 6375
rect 49988 6772 50038 6784
rect 49988 6375 49994 6772
rect 50032 6375 50038 6772
rect 49988 6363 50038 6375
rect 50306 6772 50356 6784
rect 50306 6375 50312 6772
rect 50350 6375 50356 6772
rect 50306 6363 50356 6375
rect 50624 6772 50674 6784
rect 50624 6375 50630 6772
rect 50668 6375 50674 6772
rect 50624 6363 50674 6375
rect 50942 6772 50992 6784
rect 50942 6375 50948 6772
rect 50986 6375 50992 6772
rect 50942 6363 50992 6375
rect 51260 6772 51310 6784
rect 51260 6375 51266 6772
rect 51304 6375 51310 6772
rect 51260 6363 51310 6375
rect 51578 6772 51628 6784
rect 51578 6375 51584 6772
rect 51622 6375 51628 6772
rect 51578 6363 51628 6375
rect 51896 6772 51946 6784
rect 51896 6375 51902 6772
rect 51940 6375 51946 6772
rect 51896 6363 51946 6375
rect 52214 6772 52264 6784
rect 52214 6375 52220 6772
rect 52258 6375 52264 6772
rect 52214 6363 52264 6375
rect 52532 6772 52582 6784
rect 52532 6375 52538 6772
rect 52576 6375 52582 6772
rect 52532 6363 52582 6375
rect 52850 6772 52900 6784
rect 52850 6375 52856 6772
rect 52894 6375 52900 6772
rect 52850 6363 52900 6375
rect 53168 6772 53218 6784
rect 53168 6375 53174 6772
rect 53212 6375 53218 6772
rect 53168 6363 53218 6375
rect 53486 6772 53536 6784
rect 53486 6375 53492 6772
rect 53530 6375 53536 6772
rect 53486 6363 53536 6375
rect 53804 6772 53854 6784
rect 53804 6375 53810 6772
rect 53848 6375 53854 6772
rect 53804 6363 53854 6375
rect 54122 6772 54172 6784
rect 54122 6375 54128 6772
rect 54166 6375 54172 6772
rect 54122 6363 54172 6375
rect 54440 6772 54490 6784
rect 54440 6375 54446 6772
rect 54484 6375 54490 6772
rect 54440 6363 54490 6375
rect 54758 6772 54808 6784
rect 54758 6375 54764 6772
rect 54802 6375 54808 6772
rect 54758 6363 54808 6375
rect 55076 6772 55126 6784
rect 55076 6375 55082 6772
rect 55120 6375 55126 6772
rect 55076 6363 55126 6375
rect 55394 6772 55444 6784
rect 55394 6375 55400 6772
rect 55438 6375 55444 6772
rect 55394 6363 55444 6375
rect 55712 6772 55762 6784
rect 55712 6375 55718 6772
rect 55756 6375 55762 6772
rect 55712 6363 55762 6375
rect 56030 6772 56080 6784
rect 56030 6375 56036 6772
rect 56074 6375 56080 6772
rect 56030 6363 56080 6375
rect 56348 6772 56398 6784
rect 56348 6375 56354 6772
rect 56392 6375 56398 6772
rect 56348 6363 56398 6375
rect 56666 6772 56716 6784
rect 56666 6375 56672 6772
rect 56710 6375 56716 6772
rect 56666 6363 56716 6375
rect 56984 6772 57034 6784
rect 56984 6375 56990 6772
rect 57028 6375 57034 6772
rect 56984 6363 57034 6375
rect 57302 6772 57352 6784
rect 57302 6375 57308 6772
rect 57346 6375 57352 6772
rect 57302 6363 57352 6375
rect 57620 6772 57670 6784
rect 57620 6375 57626 6772
rect 57664 6375 57670 6772
rect 57620 6363 57670 6375
rect 57938 6772 57988 6784
rect 57938 6375 57944 6772
rect 57982 6375 57988 6772
rect 57938 6363 57988 6375
rect 58256 6772 58306 6784
rect 58256 6375 58262 6772
rect 58300 6375 58306 6772
rect 58256 6363 58306 6375
rect 58574 6772 58624 6784
rect 58574 6375 58580 6772
rect 58618 6375 58624 6772
rect 58574 6363 58624 6375
rect 58892 6772 58942 6784
rect 58892 6375 58898 6772
rect 58936 6375 58942 6772
rect 58892 6363 58942 6375
rect 59210 6772 59260 6784
rect 59210 6375 59216 6772
rect 59254 6375 59260 6772
rect 59210 6363 59260 6375
rect 59528 6772 59578 6784
rect 59528 6375 59534 6772
rect 59572 6375 59578 6772
rect 59528 6363 59578 6375
rect 59846 6772 59896 6784
rect 59846 6375 59852 6772
rect 59890 6375 59896 6772
rect 59846 6363 59896 6375
rect 60164 6772 60214 6784
rect 60164 6375 60170 6772
rect 60208 6375 60214 6772
rect 60164 6363 60214 6375
rect 60482 6772 60532 6784
rect 60482 6375 60488 6772
rect 60526 6375 60532 6772
rect 60482 6363 60532 6375
rect 60800 6772 60850 6784
rect 60800 6375 60806 6772
rect 60844 6375 60850 6772
rect 60800 6363 60850 6375
rect 61118 6772 61168 6784
rect 61118 6375 61124 6772
rect 61162 6375 61168 6772
rect 61118 6363 61168 6375
rect 61436 6772 61486 6784
rect 61436 6375 61442 6772
rect 61480 6375 61486 6772
rect 61436 6363 61486 6375
rect 61754 6772 61804 6784
rect 61754 6375 61760 6772
rect 61798 6375 61804 6772
rect 61754 6363 61804 6375
rect 62072 6772 62122 6784
rect 62072 6375 62078 6772
rect 62116 6375 62122 6772
rect 62072 6363 62122 6375
rect 62390 6772 62440 6784
rect 62390 6375 62396 6772
rect 62434 6375 62440 6772
rect 62390 6363 62440 6375
rect 62708 6772 62758 6784
rect 62708 6375 62714 6772
rect 62752 6375 62758 6772
rect 62708 6363 62758 6375
rect 63026 6772 63076 6784
rect 63026 6375 63032 6772
rect 63070 6375 63076 6772
rect 63026 6363 63076 6375
rect 63344 6772 63394 6784
rect 63344 6375 63350 6772
rect 63388 6375 63394 6772
rect 63344 6363 63394 6375
rect 63662 6772 63712 6784
rect 63662 6375 63668 6772
rect 63706 6375 63712 6772
rect 63662 6363 63712 6375
rect 63980 6772 64030 6784
rect 63980 6375 63986 6772
rect 64024 6375 64030 6772
rect 63980 6363 64030 6375
rect 64298 6772 64348 6784
rect 64298 6375 64304 6772
rect 64342 6375 64348 6772
rect 64298 6363 64348 6375
rect 64616 6772 64666 6784
rect 64616 6375 64622 6772
rect 64660 6375 64666 6772
rect 64616 6363 64666 6375
rect 64934 6772 64984 6784
rect 64934 6375 64940 6772
rect 64978 6375 64984 6772
rect 64934 6363 64984 6375
rect 65252 6772 65302 6784
rect 65252 6375 65258 6772
rect 65296 6375 65302 6772
rect 65252 6363 65302 6375
rect 65570 6772 65620 6784
rect 65570 6375 65576 6772
rect 65614 6375 65620 6772
rect 65570 6363 65620 6375
rect 65888 6772 65938 6784
rect 65888 6375 65894 6772
rect 65932 6375 65938 6772
rect 65888 6363 65938 6375
rect 66206 6772 66256 6784
rect 66206 6375 66212 6772
rect 66250 6375 66256 6772
rect 66206 6363 66256 6375
rect 66524 6772 66574 6784
rect 66524 6375 66530 6772
rect 66568 6375 66574 6772
rect 66524 6363 66574 6375
rect 66842 6772 66892 6784
rect 66842 6375 66848 6772
rect 66886 6375 66892 6772
rect 66842 6363 66892 6375
rect 67160 6772 67210 6784
rect 67160 6375 67166 6772
rect 67204 6375 67210 6772
rect 67160 6363 67210 6375
rect 67478 6772 67528 6784
rect 67478 6375 67484 6772
rect 67522 6375 67528 6772
rect 67478 6363 67528 6375
rect 67796 6772 67846 6784
rect 67796 6375 67802 6772
rect 67840 6375 67846 6772
rect 67796 6363 67846 6375
rect 68114 6772 68164 6784
rect 68114 6375 68120 6772
rect 68158 6375 68164 6772
rect 68114 6363 68164 6375
rect 68432 6772 68482 6784
rect 68432 6375 68438 6772
rect 68476 6375 68482 6772
rect 68432 6363 68482 6375
rect 68750 6772 68800 6784
rect 68750 6375 68756 6772
rect 68794 6375 68800 6772
rect 68750 6363 68800 6375
rect 69068 6772 69118 6784
rect 69068 6375 69074 6772
rect 69112 6375 69118 6772
rect 69068 6363 69118 6375
rect 69386 6772 69436 6784
rect 69386 6375 69392 6772
rect 69430 6375 69436 6772
rect 69386 6363 69436 6375
rect 69704 6772 69754 6784
rect 69704 6375 69710 6772
rect 69748 6375 69754 6772
rect 69704 6363 69754 6375
rect 70022 6772 70072 6784
rect 70022 6375 70028 6772
rect 70066 6375 70072 6772
rect 70022 6363 70072 6375
rect 70340 6772 70390 6784
rect 70340 6375 70346 6772
rect 70384 6375 70390 6772
rect 70340 6363 70390 6375
rect 70658 6772 70708 6784
rect 70658 6375 70664 6772
rect 70702 6375 70708 6772
rect 70658 6363 70708 6375
rect 70976 6772 71026 6784
rect 70976 6375 70982 6772
rect 71020 6375 71026 6772
rect 70976 6363 71026 6375
rect 71294 6772 71344 6784
rect 71294 6375 71300 6772
rect 71338 6375 71344 6772
rect 71294 6363 71344 6375
rect 71612 6772 71662 6784
rect 71612 6375 71618 6772
rect 71656 6375 71662 6772
rect 71612 6363 71662 6375
rect 71930 6772 71980 6784
rect 71930 6375 71936 6772
rect 71974 6375 71980 6772
rect 71930 6363 71980 6375
rect 72248 6772 72298 6784
rect 72248 6375 72254 6772
rect 72292 6375 72298 6772
rect 72248 6363 72298 6375
rect 72566 6772 72616 6784
rect 72566 6375 72572 6772
rect 72610 6375 72616 6772
rect 72566 6363 72616 6375
rect 72884 6772 72934 6784
rect 72884 6375 72890 6772
rect 72928 6375 72934 6772
rect 72884 6363 72934 6375
rect 73202 6772 73252 6784
rect 73202 6375 73208 6772
rect 73246 6375 73252 6772
rect 73202 6363 73252 6375
rect 73520 6772 73570 6784
rect 73520 6375 73526 6772
rect 73564 6375 73570 6772
rect 73520 6363 73570 6375
rect 73838 6772 73888 6784
rect 73838 6375 73844 6772
rect 73882 6375 73888 6772
rect 73838 6363 73888 6375
rect 74156 6772 74206 6784
rect 74156 6375 74162 6772
rect 74200 6375 74206 6772
rect 74156 6363 74206 6375
rect 74474 6772 74524 6784
rect 74474 6375 74480 6772
rect 74518 6375 74524 6772
rect 74474 6363 74524 6375
rect 74792 6772 74842 6784
rect 74792 6375 74798 6772
rect 74836 6375 74842 6772
rect 74792 6363 74842 6375
rect 75110 6772 75160 6784
rect 75110 6375 75116 6772
rect 75154 6375 75160 6772
rect 75110 6363 75160 6375
rect 75428 6772 75478 6784
rect 75428 6375 75434 6772
rect 75472 6375 75478 6772
rect 75428 6363 75478 6375
rect 75746 6772 75796 6784
rect 75746 6375 75752 6772
rect 75790 6375 75796 6772
rect 75746 6363 75796 6375
rect 76064 6772 76114 6784
rect 76064 6375 76070 6772
rect 76108 6375 76114 6772
rect 76064 6363 76114 6375
rect 76382 6772 76432 6784
rect 76382 6375 76388 6772
rect 76426 6375 76432 6772
rect 76382 6363 76432 6375
rect 76700 6772 76750 6784
rect 76700 6375 76706 6772
rect 76744 6375 76750 6772
rect 76700 6363 76750 6375
rect 77018 6772 77068 6784
rect 77018 6375 77024 6772
rect 77062 6375 77068 6772
rect 77018 6363 77068 6375
rect 77336 6772 77386 6784
rect 77336 6375 77342 6772
rect 77380 6375 77386 6772
rect 77336 6363 77386 6375
rect 77654 6772 77704 6784
rect 77654 6375 77660 6772
rect 77698 6375 77704 6772
rect 77654 6363 77704 6375
rect 77972 6772 78022 6784
rect 77972 6375 77978 6772
rect 78016 6375 78022 6772
rect 77972 6363 78022 6375
rect 78290 6772 78340 6784
rect 78290 6375 78296 6772
rect 78334 6375 78340 6772
rect 78290 6363 78340 6375
rect 78608 6772 78658 6784
rect 78608 6375 78614 6772
rect 78652 6375 78658 6772
rect 78608 6363 78658 6375
rect 78926 6772 78976 6784
rect 78926 6375 78932 6772
rect 78970 6375 78976 6772
rect 78926 6363 78976 6375
rect 79244 6772 79294 6784
rect 79244 6375 79250 6772
rect 79288 6375 79294 6772
rect 79244 6363 79294 6375
rect 79562 6772 79612 6784
rect 79562 6375 79568 6772
rect 79606 6375 79612 6772
rect 79562 6363 79612 6375
rect 79880 6772 79930 6784
rect 79880 6375 79886 6772
rect 79924 6375 79930 6772
rect 79880 6363 79930 6375
rect 80198 6772 80248 6784
rect 80198 6375 80204 6772
rect 80242 6375 80248 6772
rect 80198 6363 80248 6375
rect 48716 -659 48766 -647
rect 48716 -1056 48722 -659
rect 48760 -1056 48766 -659
rect 48716 -1068 48766 -1056
rect 49034 -659 49084 -647
rect 49034 -1056 49040 -659
rect 49078 -1056 49084 -659
rect 49034 -1068 49084 -1056
rect 49352 -659 49402 -647
rect 49352 -1056 49358 -659
rect 49396 -1056 49402 -659
rect 49352 -1068 49402 -1056
rect 49670 -659 49720 -647
rect 49670 -1056 49676 -659
rect 49714 -1056 49720 -659
rect 49670 -1068 49720 -1056
rect 49988 -659 50038 -647
rect 49988 -1056 49994 -659
rect 50032 -1056 50038 -659
rect 49988 -1068 50038 -1056
rect 50306 -659 50356 -647
rect 50306 -1056 50312 -659
rect 50350 -1056 50356 -659
rect 50306 -1068 50356 -1056
rect 50624 -659 50674 -647
rect 50624 -1056 50630 -659
rect 50668 -1056 50674 -659
rect 50624 -1068 50674 -1056
rect 50942 -659 50992 -647
rect 50942 -1056 50948 -659
rect 50986 -1056 50992 -659
rect 50942 -1068 50992 -1056
rect 51260 -659 51310 -647
rect 51260 -1056 51266 -659
rect 51304 -1056 51310 -659
rect 51260 -1068 51310 -1056
rect 51578 -659 51628 -647
rect 51578 -1056 51584 -659
rect 51622 -1056 51628 -659
rect 51578 -1068 51628 -1056
rect 51896 -659 51946 -647
rect 51896 -1056 51902 -659
rect 51940 -1056 51946 -659
rect 51896 -1068 51946 -1056
rect 52214 -659 52264 -647
rect 52214 -1056 52220 -659
rect 52258 -1056 52264 -659
rect 52214 -1068 52264 -1056
rect 52532 -659 52582 -647
rect 52532 -1056 52538 -659
rect 52576 -1056 52582 -659
rect 52532 -1068 52582 -1056
rect 52850 -659 52900 -647
rect 52850 -1056 52856 -659
rect 52894 -1056 52900 -659
rect 52850 -1068 52900 -1056
rect 53168 -659 53218 -647
rect 53168 -1056 53174 -659
rect 53212 -1056 53218 -659
rect 53168 -1068 53218 -1056
rect 53486 -659 53536 -647
rect 53486 -1056 53492 -659
rect 53530 -1056 53536 -659
rect 53486 -1068 53536 -1056
rect 53804 -659 53854 -647
rect 53804 -1056 53810 -659
rect 53848 -1056 53854 -659
rect 53804 -1068 53854 -1056
rect 54122 -659 54172 -647
rect 54122 -1056 54128 -659
rect 54166 -1056 54172 -659
rect 54122 -1068 54172 -1056
rect 54440 -659 54490 -647
rect 54440 -1056 54446 -659
rect 54484 -1056 54490 -659
rect 54440 -1068 54490 -1056
rect 54758 -659 54808 -647
rect 54758 -1056 54764 -659
rect 54802 -1056 54808 -659
rect 54758 -1068 54808 -1056
rect 55076 -659 55126 -647
rect 55076 -1056 55082 -659
rect 55120 -1056 55126 -659
rect 55076 -1068 55126 -1056
rect 55394 -659 55444 -647
rect 55394 -1056 55400 -659
rect 55438 -1056 55444 -659
rect 55394 -1068 55444 -1056
rect 55712 -659 55762 -647
rect 55712 -1056 55718 -659
rect 55756 -1056 55762 -659
rect 55712 -1068 55762 -1056
rect 56030 -659 56080 -647
rect 56030 -1056 56036 -659
rect 56074 -1056 56080 -659
rect 56030 -1068 56080 -1056
rect 56348 -659 56398 -647
rect 56348 -1056 56354 -659
rect 56392 -1056 56398 -659
rect 56348 -1068 56398 -1056
rect 56666 -659 56716 -647
rect 56666 -1056 56672 -659
rect 56710 -1056 56716 -659
rect 56666 -1068 56716 -1056
rect 56984 -659 57034 -647
rect 56984 -1056 56990 -659
rect 57028 -1056 57034 -659
rect 56984 -1068 57034 -1056
rect 57302 -659 57352 -647
rect 57302 -1056 57308 -659
rect 57346 -1056 57352 -659
rect 57302 -1068 57352 -1056
rect 57620 -659 57670 -647
rect 57620 -1056 57626 -659
rect 57664 -1056 57670 -659
rect 57620 -1068 57670 -1056
rect 57938 -659 57988 -647
rect 57938 -1056 57944 -659
rect 57982 -1056 57988 -659
rect 57938 -1068 57988 -1056
rect 58256 -659 58306 -647
rect 58256 -1056 58262 -659
rect 58300 -1056 58306 -659
rect 58256 -1068 58306 -1056
rect 58574 -659 58624 -647
rect 58574 -1056 58580 -659
rect 58618 -1056 58624 -659
rect 58574 -1068 58624 -1056
rect 58892 -659 58942 -647
rect 58892 -1056 58898 -659
rect 58936 -1056 58942 -659
rect 58892 -1068 58942 -1056
rect 59210 -659 59260 -647
rect 59210 -1056 59216 -659
rect 59254 -1056 59260 -659
rect 59210 -1068 59260 -1056
rect 59528 -659 59578 -647
rect 59528 -1056 59534 -659
rect 59572 -1056 59578 -659
rect 59528 -1068 59578 -1056
rect 59846 -659 59896 -647
rect 59846 -1056 59852 -659
rect 59890 -1056 59896 -659
rect 59846 -1068 59896 -1056
rect 60164 -659 60214 -647
rect 60164 -1056 60170 -659
rect 60208 -1056 60214 -659
rect 60164 -1068 60214 -1056
rect 60482 -659 60532 -647
rect 60482 -1056 60488 -659
rect 60526 -1056 60532 -659
rect 60482 -1068 60532 -1056
rect 60800 -659 60850 -647
rect 60800 -1056 60806 -659
rect 60844 -1056 60850 -659
rect 60800 -1068 60850 -1056
rect 61118 -659 61168 -647
rect 61118 -1056 61124 -659
rect 61162 -1056 61168 -659
rect 61118 -1068 61168 -1056
rect 61436 -659 61486 -647
rect 61436 -1056 61442 -659
rect 61480 -1056 61486 -659
rect 61436 -1068 61486 -1056
rect 61754 -659 61804 -647
rect 61754 -1056 61760 -659
rect 61798 -1056 61804 -659
rect 61754 -1068 61804 -1056
rect 62072 -659 62122 -647
rect 62072 -1056 62078 -659
rect 62116 -1056 62122 -659
rect 62072 -1068 62122 -1056
rect 62390 -659 62440 -647
rect 62390 -1056 62396 -659
rect 62434 -1056 62440 -659
rect 62390 -1068 62440 -1056
rect 62708 -659 62758 -647
rect 62708 -1056 62714 -659
rect 62752 -1056 62758 -659
rect 62708 -1068 62758 -1056
rect 63026 -659 63076 -647
rect 63026 -1056 63032 -659
rect 63070 -1056 63076 -659
rect 63026 -1068 63076 -1056
rect 63344 -659 63394 -647
rect 63344 -1056 63350 -659
rect 63388 -1056 63394 -659
rect 63344 -1068 63394 -1056
rect 63662 -659 63712 -647
rect 63662 -1056 63668 -659
rect 63706 -1056 63712 -659
rect 63662 -1068 63712 -1056
rect 63980 -659 64030 -647
rect 63980 -1056 63986 -659
rect 64024 -1056 64030 -659
rect 63980 -1068 64030 -1056
rect 64298 -659 64348 -647
rect 64298 -1056 64304 -659
rect 64342 -1056 64348 -659
rect 64298 -1068 64348 -1056
rect 64616 -659 64666 -647
rect 64616 -1056 64622 -659
rect 64660 -1056 64666 -659
rect 64616 -1068 64666 -1056
rect 64934 -659 64984 -647
rect 64934 -1056 64940 -659
rect 64978 -1056 64984 -659
rect 64934 -1068 64984 -1056
rect 65252 -659 65302 -647
rect 65252 -1056 65258 -659
rect 65296 -1056 65302 -659
rect 65252 -1068 65302 -1056
rect 65570 -659 65620 -647
rect 65570 -1056 65576 -659
rect 65614 -1056 65620 -659
rect 65570 -1068 65620 -1056
rect 65888 -659 65938 -647
rect 65888 -1056 65894 -659
rect 65932 -1056 65938 -659
rect 65888 -1068 65938 -1056
rect 66206 -659 66256 -647
rect 66206 -1056 66212 -659
rect 66250 -1056 66256 -659
rect 66206 -1068 66256 -1056
rect 66524 -659 66574 -647
rect 66524 -1056 66530 -659
rect 66568 -1056 66574 -659
rect 66524 -1068 66574 -1056
rect 66842 -659 66892 -647
rect 66842 -1056 66848 -659
rect 66886 -1056 66892 -659
rect 66842 -1068 66892 -1056
rect 67160 -659 67210 -647
rect 67160 -1056 67166 -659
rect 67204 -1056 67210 -659
rect 67160 -1068 67210 -1056
rect 67478 -659 67528 -647
rect 67478 -1056 67484 -659
rect 67522 -1056 67528 -659
rect 67478 -1068 67528 -1056
rect 67796 -659 67846 -647
rect 67796 -1056 67802 -659
rect 67840 -1056 67846 -659
rect 67796 -1068 67846 -1056
rect 68114 -659 68164 -647
rect 68114 -1056 68120 -659
rect 68158 -1056 68164 -659
rect 68114 -1068 68164 -1056
rect 68432 -659 68482 -647
rect 68432 -1056 68438 -659
rect 68476 -1056 68482 -659
rect 68432 -1068 68482 -1056
rect 68750 -659 68800 -647
rect 68750 -1056 68756 -659
rect 68794 -1056 68800 -659
rect 68750 -1068 68800 -1056
rect 69068 -659 69118 -647
rect 69068 -1056 69074 -659
rect 69112 -1056 69118 -659
rect 69068 -1068 69118 -1056
rect 69386 -659 69436 -647
rect 69386 -1056 69392 -659
rect 69430 -1056 69436 -659
rect 69386 -1068 69436 -1056
rect 69704 -659 69754 -647
rect 69704 -1056 69710 -659
rect 69748 -1056 69754 -659
rect 69704 -1068 69754 -1056
rect 70022 -659 70072 -647
rect 70022 -1056 70028 -659
rect 70066 -1056 70072 -659
rect 70022 -1068 70072 -1056
rect 70340 -659 70390 -647
rect 70340 -1056 70346 -659
rect 70384 -1056 70390 -659
rect 70340 -1068 70390 -1056
rect 70658 -659 70708 -647
rect 70658 -1056 70664 -659
rect 70702 -1056 70708 -659
rect 70658 -1068 70708 -1056
rect 70976 -659 71026 -647
rect 70976 -1056 70982 -659
rect 71020 -1056 71026 -659
rect 70976 -1068 71026 -1056
rect 71294 -659 71344 -647
rect 71294 -1056 71300 -659
rect 71338 -1056 71344 -659
rect 71294 -1068 71344 -1056
rect 71612 -659 71662 -647
rect 71612 -1056 71618 -659
rect 71656 -1056 71662 -659
rect 71612 -1068 71662 -1056
rect 71930 -659 71980 -647
rect 71930 -1056 71936 -659
rect 71974 -1056 71980 -659
rect 71930 -1068 71980 -1056
rect 72248 -659 72298 -647
rect 72248 -1056 72254 -659
rect 72292 -1056 72298 -659
rect 72248 -1068 72298 -1056
rect 72566 -659 72616 -647
rect 72566 -1056 72572 -659
rect 72610 -1056 72616 -659
rect 72566 -1068 72616 -1056
rect 72884 -659 72934 -647
rect 72884 -1056 72890 -659
rect 72928 -1056 72934 -659
rect 72884 -1068 72934 -1056
rect 73202 -659 73252 -647
rect 73202 -1056 73208 -659
rect 73246 -1056 73252 -659
rect 73202 -1068 73252 -1056
rect 73520 -659 73570 -647
rect 73520 -1056 73526 -659
rect 73564 -1056 73570 -659
rect 73520 -1068 73570 -1056
rect 73838 -659 73888 -647
rect 73838 -1056 73844 -659
rect 73882 -1056 73888 -659
rect 73838 -1068 73888 -1056
rect 74156 -659 74206 -647
rect 74156 -1056 74162 -659
rect 74200 -1056 74206 -659
rect 74156 -1068 74206 -1056
rect 74474 -659 74524 -647
rect 74474 -1056 74480 -659
rect 74518 -1056 74524 -659
rect 74474 -1068 74524 -1056
rect 74792 -659 74842 -647
rect 74792 -1056 74798 -659
rect 74836 -1056 74842 -659
rect 74792 -1068 74842 -1056
rect 75110 -659 75160 -647
rect 75110 -1056 75116 -659
rect 75154 -1056 75160 -659
rect 75110 -1068 75160 -1056
rect 75428 -659 75478 -647
rect 75428 -1056 75434 -659
rect 75472 -1056 75478 -659
rect 75428 -1068 75478 -1056
rect 75746 -659 75796 -647
rect 75746 -1056 75752 -659
rect 75790 -1056 75796 -659
rect 75746 -1068 75796 -1056
rect 76064 -659 76114 -647
rect 76064 -1056 76070 -659
rect 76108 -1056 76114 -659
rect 76064 -1068 76114 -1056
rect 76382 -659 76432 -647
rect 76382 -1056 76388 -659
rect 76426 -1056 76432 -659
rect 76382 -1068 76432 -1056
rect 76700 -659 76750 -647
rect 76700 -1056 76706 -659
rect 76744 -1056 76750 -659
rect 76700 -1068 76750 -1056
rect 77018 -659 77068 -647
rect 77018 -1056 77024 -659
rect 77062 -1056 77068 -659
rect 77018 -1068 77068 -1056
rect 77336 -659 77386 -647
rect 77336 -1056 77342 -659
rect 77380 -1056 77386 -659
rect 77336 -1068 77386 -1056
rect 77654 -659 77704 -647
rect 77654 -1056 77660 -659
rect 77698 -1056 77704 -659
rect 77654 -1068 77704 -1056
rect 77972 -659 78022 -647
rect 77972 -1056 77978 -659
rect 78016 -1056 78022 -659
rect 77972 -1068 78022 -1056
rect 78290 -659 78340 -647
rect 78290 -1056 78296 -659
rect 78334 -1056 78340 -659
rect 78290 -1068 78340 -1056
rect 78608 -659 78658 -647
rect 78608 -1056 78614 -659
rect 78652 -1056 78658 -659
rect 78608 -1068 78658 -1056
rect 78926 -659 78976 -647
rect 78926 -1056 78932 -659
rect 78970 -1056 78976 -659
rect 78926 -1068 78976 -1056
rect 79244 -659 79294 -647
rect 79244 -1056 79250 -659
rect 79288 -1056 79294 -659
rect 79244 -1068 79294 -1056
rect 79562 -659 79612 -647
rect 79562 -1056 79568 -659
rect 79606 -1056 79612 -659
rect 79562 -1068 79612 -1056
rect 79880 -659 79930 -647
rect 79880 -1056 79886 -659
rect 79924 -1056 79930 -659
rect 79880 -1068 79930 -1056
rect 80198 -659 80248 -647
rect 80198 -1056 80204 -659
rect 80242 -1056 80248 -659
rect 80198 -1068 80248 -1056
<< labels >>
rlabel locali 48580 -1200 48600 -1180 1 gnd
port 4 n
rlabel locali 48840 14660 48900 14720 1 A
port 1 n
rlabel locali 48880 6820 48940 6880 1 B
port 2 n
rlabel locali 48900 -1040 48960 -980 1 C
port 3 n
<< end >>
