* SPICE3 file created from p1_8.ext - technology: sky130A

.option scale=10000u

.subckt p1_8 D G S B SUB
X0 S G a1 B sky130_fd_pr__pfet_01v8_lvt ad=15000 pd=700 as=30000 ps=1400 w=300 l=800
X1 D G a7 B sky130_fd_pr__pfet_01v8_lvt ad=15000 pd=700 as=30000 ps=1400 w=300 l=800
X2 a4 G a5 B sky130_fd_pr__pfet_01v8_lvt ad=30000 pd=1400 as=30000 ps=1400 w=300 l=800
X3 a6 G a5 B sky130_fd_pr__pfet_01v8_lvt ad=30000 pd=1400 as=0 ps=0 w=300 l=800
X4 a2 G a3 B sky130_fd_pr__pfet_01v8_lvt ad=30000 pd=1400 as=30000 ps=1400 w=300 l=800
X5 a6 G a7 B sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=300 l=800
X6 a4 G a3 B sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=300 l=800
X7 a2 G a1 B sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=300 l=800
.ends
