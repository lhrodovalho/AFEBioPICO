* FD-OTA netlist


