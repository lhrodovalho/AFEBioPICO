magic
tech sky130A
timestamp 1634337365
<< pwell >>
rect 0 1150 940 1230
rect 0 1120 850 1150
rect 860 1120 940 1150
rect 0 0 940 1120
<< nmoslvt >>
rect 70 990 870 1090
rect 70 860 870 960
rect 70 730 870 830
rect 70 600 870 700
rect 70 470 870 570
rect 70 340 870 440
rect 70 210 870 310
rect 70 80 870 180
<< ndiff >>
rect 20 1080 70 1090
rect 20 1000 30 1080
rect 60 1000 70 1080
rect 20 990 70 1000
rect 870 1080 920 1090
rect 870 1000 880 1080
rect 910 1000 920 1080
rect 870 990 920 1000
rect 20 950 70 960
rect 20 870 30 950
rect 60 870 70 950
rect 20 860 70 870
rect 870 950 920 960
rect 870 870 880 950
rect 910 870 920 950
rect 870 860 920 870
rect 20 820 70 830
rect 20 740 30 820
rect 60 740 70 820
rect 20 730 70 740
rect 870 820 920 830
rect 870 740 880 820
rect 910 740 920 820
rect 870 730 920 740
rect 20 690 70 700
rect 20 610 30 690
rect 60 610 70 690
rect 20 600 70 610
rect 870 690 920 700
rect 870 610 880 690
rect 910 610 920 690
rect 870 600 920 610
rect 20 560 70 570
rect 20 480 30 560
rect 60 480 70 560
rect 20 470 70 480
rect 870 560 920 570
rect 870 480 880 560
rect 910 480 920 560
rect 870 470 920 480
rect 20 430 70 440
rect 20 350 30 430
rect 60 350 70 430
rect 20 340 70 350
rect 870 430 920 440
rect 870 350 880 430
rect 910 350 920 430
rect 870 340 920 350
rect 20 300 70 310
rect 20 220 30 300
rect 60 220 70 300
rect 20 210 70 220
rect 870 300 920 310
rect 870 220 880 300
rect 910 220 920 300
rect 870 210 920 220
rect 20 170 70 180
rect 20 90 30 170
rect 60 90 70 170
rect 20 80 70 90
rect 870 170 920 180
rect 870 90 880 170
rect 910 90 920 170
rect 870 80 920 90
<< ndiffc >>
rect 30 1000 60 1080
rect 880 1000 910 1080
rect 30 870 60 950
rect 880 870 910 950
rect 30 740 60 820
rect 880 740 910 820
rect 30 610 60 690
rect 880 610 910 690
rect 30 480 60 560
rect 880 480 910 560
rect 30 350 60 430
rect 880 350 910 430
rect 30 220 60 300
rect 880 220 910 300
rect 30 90 60 170
rect 880 90 910 170
<< psubdiff >>
rect 0 1180 70 1210
rect 870 1180 940 1210
rect 0 20 70 50
rect 870 20 940 50
<< psubdiffcont >>
rect 70 1180 870 1210
rect 70 20 870 50
<< poly >>
rect 70 1150 870 1160
rect 70 1120 90 1150
rect 850 1120 870 1150
rect 70 1090 870 1120
rect 70 960 870 990
rect 70 830 870 860
rect 70 700 870 730
rect 70 570 870 600
rect 70 440 870 470
rect 70 310 870 340
rect 70 180 870 210
rect 70 60 870 80
<< polycont >>
rect 90 1120 850 1150
<< locali >>
rect 0 1180 70 1210
rect 870 1180 940 1210
rect 80 1120 90 1150
rect 850 1120 860 1150
rect 30 1080 60 1090
rect 30 990 60 1000
rect 880 1080 910 1090
rect 30 950 60 960
rect 30 820 60 870
rect 880 950 910 1000
rect 880 860 910 870
rect 30 730 60 740
rect 880 820 910 830
rect 30 690 60 700
rect 30 560 60 610
rect 880 690 910 740
rect 880 600 910 610
rect 30 470 60 480
rect 880 560 910 570
rect 30 430 60 440
rect 30 300 60 350
rect 880 430 910 480
rect 880 340 910 350
rect 30 210 60 220
rect 880 300 910 310
rect 30 170 60 180
rect 30 80 60 90
rect 880 170 910 220
rect 880 80 910 90
rect 0 20 70 50
rect 870 20 940 50
<< viali >>
rect 760 1120 790 1150
rect 30 1000 60 1080
rect 30 90 60 170
<< metal1 >>
rect 30 1090 60 1230
rect 760 1160 790 1230
rect 750 1150 800 1160
rect 750 1120 760 1150
rect 790 1120 800 1150
rect 750 1110 800 1120
rect 20 1080 70 1090
rect 20 1000 30 1080
rect 60 1000 70 1080
rect 20 990 70 1000
rect 20 170 70 180
rect 20 90 30 170
rect 60 90 70 170
rect 20 80 70 90
rect 30 0 60 80
<< labels >>
rlabel metal1 30 1220 60 1230 5 D
port 1 s
rlabel metal1 30 0 60 10 1 S
port 3 n
rlabel metal1 760 1220 790 1230 5 G
port 2 s
rlabel locali 890 190 900 200 1 a1
rlabel locali 40 320 50 330 1 a2
rlabel locali 890 450 900 460 1 a3
rlabel locali 40 580 50 590 1 a4
rlabel locali 890 710 900 720 1 a5
rlabel locali 40 840 50 850 1 a6
rlabel locali 890 970 900 980 1 a7
rlabel locali 0 20 10 50 3 B
port 4 e
<< end >>
