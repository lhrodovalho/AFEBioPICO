magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< pwell >>
rect -12906 3574 14906 3706
rect -12906 1466 -12774 3574
rect 14774 1466 14906 3574
rect -12906 1334 14906 1466
<< psubdiff >>
rect -12880 3657 14880 3680
rect -12880 3623 -12719 3657
rect -12685 3623 -12651 3657
rect -12617 3623 -12583 3657
rect -12549 3623 -12515 3657
rect -12481 3623 -12447 3657
rect -12413 3623 -12379 3657
rect -12345 3623 -12311 3657
rect -12277 3623 -12243 3657
rect -12209 3623 -12175 3657
rect -12141 3623 -12107 3657
rect -12073 3623 -12039 3657
rect -12005 3623 -11971 3657
rect -11937 3623 -11903 3657
rect -11869 3623 -11835 3657
rect -11801 3623 -11767 3657
rect -11733 3623 -11699 3657
rect -11665 3623 -11631 3657
rect -11597 3623 -11563 3657
rect -11529 3623 -11495 3657
rect -11461 3623 -11427 3657
rect -11393 3623 -11359 3657
rect -11325 3623 -11291 3657
rect -11257 3623 -11223 3657
rect -11189 3623 -11155 3657
rect -11121 3623 -11087 3657
rect -11053 3623 -11019 3657
rect -10985 3623 -10951 3657
rect -10917 3623 -10883 3657
rect -10849 3623 -10815 3657
rect -10781 3623 -10747 3657
rect -10713 3623 -10679 3657
rect -10645 3623 -10611 3657
rect -10577 3623 -10543 3657
rect -10509 3623 -10475 3657
rect -10441 3623 -10407 3657
rect -10373 3623 -10339 3657
rect -10305 3623 -10271 3657
rect -10237 3623 -10203 3657
rect -10169 3623 -10135 3657
rect -10101 3623 -10067 3657
rect -10033 3623 -9999 3657
rect -9965 3623 -9931 3657
rect -9897 3623 -9863 3657
rect -9829 3623 -9795 3657
rect -9761 3623 -9727 3657
rect -9693 3623 -9659 3657
rect -9625 3623 -9591 3657
rect -9557 3623 -9523 3657
rect -9489 3623 -9455 3657
rect -9421 3623 -9387 3657
rect -9353 3623 -9319 3657
rect -9285 3623 -9251 3657
rect -9217 3623 -9183 3657
rect -9149 3623 -9115 3657
rect -9081 3623 -9047 3657
rect -9013 3623 -8979 3657
rect -8945 3623 -8911 3657
rect -8877 3623 -8843 3657
rect -8809 3623 -8775 3657
rect -8741 3623 -8707 3657
rect -8673 3623 -8639 3657
rect -8605 3623 -8571 3657
rect -8537 3623 -8503 3657
rect -8469 3623 -8435 3657
rect -8401 3623 -8367 3657
rect -8333 3623 -8299 3657
rect -8265 3623 -8231 3657
rect -8197 3623 -8163 3657
rect -8129 3623 -8095 3657
rect -8061 3623 -8027 3657
rect -7993 3623 -7959 3657
rect -7925 3623 -7891 3657
rect -7857 3623 -7823 3657
rect -7789 3623 -7755 3657
rect -7721 3623 -7687 3657
rect -7653 3623 -7619 3657
rect -7585 3623 -7551 3657
rect -7517 3623 -7483 3657
rect -7449 3623 -7415 3657
rect -7381 3623 -7347 3657
rect -7313 3623 -7279 3657
rect -7245 3623 -7211 3657
rect -7177 3623 -7143 3657
rect -7109 3623 -7075 3657
rect -7041 3623 -7007 3657
rect -6973 3623 -6939 3657
rect -6905 3623 -6871 3657
rect -6837 3623 -6803 3657
rect -6769 3623 -6735 3657
rect -6701 3623 -6667 3657
rect -6633 3623 -6599 3657
rect -6565 3623 -6531 3657
rect -6497 3623 -6463 3657
rect -6429 3623 -6395 3657
rect -6361 3623 -6327 3657
rect -6293 3623 -6259 3657
rect -6225 3623 -6191 3657
rect -6157 3623 -6123 3657
rect -6089 3623 -6055 3657
rect -6021 3623 -5987 3657
rect -5953 3623 -5919 3657
rect -5885 3623 -5851 3657
rect -5817 3623 -5783 3657
rect -5749 3623 -5715 3657
rect -5681 3623 -5647 3657
rect -5613 3623 -5579 3657
rect -5545 3623 -5511 3657
rect -5477 3623 -5443 3657
rect -5409 3623 -5375 3657
rect -5341 3623 -5307 3657
rect -5273 3623 -5239 3657
rect -5205 3623 -5171 3657
rect -5137 3623 -5103 3657
rect -5069 3623 -5035 3657
rect -5001 3623 -4967 3657
rect -4933 3623 -4899 3657
rect -4865 3623 -4831 3657
rect -4797 3623 -4763 3657
rect -4729 3623 -4695 3657
rect -4661 3623 -4627 3657
rect -4593 3623 -4559 3657
rect -4525 3623 -4491 3657
rect -4457 3623 -4423 3657
rect -4389 3623 -4355 3657
rect -4321 3623 -4287 3657
rect -4253 3623 -4219 3657
rect -4185 3623 -4151 3657
rect -4117 3623 -4083 3657
rect -4049 3623 -4015 3657
rect -3981 3623 -3947 3657
rect -3913 3623 -3879 3657
rect -3845 3623 -3811 3657
rect -3777 3623 -3743 3657
rect -3709 3623 -3675 3657
rect -3641 3623 -3607 3657
rect -3573 3623 -3539 3657
rect -3505 3623 -3471 3657
rect -3437 3623 -3403 3657
rect -3369 3623 -3335 3657
rect -3301 3623 -3267 3657
rect -3233 3623 -3199 3657
rect -3165 3623 -3131 3657
rect -3097 3623 -3063 3657
rect -3029 3623 -2995 3657
rect -2961 3623 -2927 3657
rect -2893 3623 -2859 3657
rect -2825 3623 -2791 3657
rect -2757 3623 -2723 3657
rect -2689 3623 -2655 3657
rect -2621 3623 -2587 3657
rect -2553 3623 -2519 3657
rect -2485 3623 -2451 3657
rect -2417 3623 -2383 3657
rect -2349 3623 -2315 3657
rect -2281 3623 -2247 3657
rect -2213 3623 -2179 3657
rect -2145 3623 -2111 3657
rect -2077 3623 -2043 3657
rect -2009 3623 -1975 3657
rect -1941 3623 -1907 3657
rect -1873 3623 -1839 3657
rect -1805 3623 -1771 3657
rect -1737 3623 -1703 3657
rect -1669 3623 -1635 3657
rect -1601 3623 -1567 3657
rect -1533 3623 -1499 3657
rect -1465 3623 -1431 3657
rect -1397 3623 -1363 3657
rect -1329 3623 -1295 3657
rect -1261 3623 -1227 3657
rect -1193 3623 -1159 3657
rect -1125 3623 -1091 3657
rect -1057 3623 -1023 3657
rect -989 3623 -955 3657
rect -921 3623 -887 3657
rect -853 3623 -819 3657
rect -785 3623 -751 3657
rect -717 3623 -683 3657
rect -649 3623 -615 3657
rect -581 3623 -547 3657
rect -513 3623 -479 3657
rect -445 3623 -411 3657
rect -377 3623 -343 3657
rect -309 3623 -275 3657
rect -241 3623 -207 3657
rect -173 3623 -139 3657
rect -105 3623 -71 3657
rect -37 3623 -3 3657
rect 31 3623 65 3657
rect 99 3623 133 3657
rect 167 3623 201 3657
rect 235 3623 269 3657
rect 303 3623 337 3657
rect 371 3623 405 3657
rect 439 3623 473 3657
rect 507 3623 541 3657
rect 575 3623 609 3657
rect 643 3623 677 3657
rect 711 3623 745 3657
rect 779 3623 813 3657
rect 847 3623 881 3657
rect 915 3623 949 3657
rect 983 3623 1017 3657
rect 1051 3623 1085 3657
rect 1119 3623 1153 3657
rect 1187 3623 1221 3657
rect 1255 3623 1289 3657
rect 1323 3623 1357 3657
rect 1391 3623 1425 3657
rect 1459 3623 1493 3657
rect 1527 3623 1561 3657
rect 1595 3623 1629 3657
rect 1663 3623 1697 3657
rect 1731 3623 1765 3657
rect 1799 3623 1833 3657
rect 1867 3623 1901 3657
rect 1935 3623 1969 3657
rect 2003 3623 2037 3657
rect 2071 3623 2105 3657
rect 2139 3623 2173 3657
rect 2207 3623 2241 3657
rect 2275 3623 2309 3657
rect 2343 3623 2377 3657
rect 2411 3623 2445 3657
rect 2479 3623 2513 3657
rect 2547 3623 2581 3657
rect 2615 3623 2649 3657
rect 2683 3623 2717 3657
rect 2751 3623 2785 3657
rect 2819 3623 2853 3657
rect 2887 3623 2921 3657
rect 2955 3623 2989 3657
rect 3023 3623 3057 3657
rect 3091 3623 3125 3657
rect 3159 3623 3193 3657
rect 3227 3623 3261 3657
rect 3295 3623 3329 3657
rect 3363 3623 3397 3657
rect 3431 3623 3465 3657
rect 3499 3623 3533 3657
rect 3567 3623 3601 3657
rect 3635 3623 3669 3657
rect 3703 3623 3737 3657
rect 3771 3623 3805 3657
rect 3839 3623 3873 3657
rect 3907 3623 3941 3657
rect 3975 3623 4009 3657
rect 4043 3623 4077 3657
rect 4111 3623 4145 3657
rect 4179 3623 4213 3657
rect 4247 3623 4281 3657
rect 4315 3623 4349 3657
rect 4383 3623 4417 3657
rect 4451 3623 4485 3657
rect 4519 3623 4553 3657
rect 4587 3623 4621 3657
rect 4655 3623 4689 3657
rect 4723 3623 4757 3657
rect 4791 3623 4825 3657
rect 4859 3623 4893 3657
rect 4927 3623 4961 3657
rect 4995 3623 5029 3657
rect 5063 3623 5097 3657
rect 5131 3623 5165 3657
rect 5199 3623 5233 3657
rect 5267 3623 5301 3657
rect 5335 3623 5369 3657
rect 5403 3623 5437 3657
rect 5471 3623 5505 3657
rect 5539 3623 5573 3657
rect 5607 3623 5641 3657
rect 5675 3623 5709 3657
rect 5743 3623 5777 3657
rect 5811 3623 5845 3657
rect 5879 3623 5913 3657
rect 5947 3623 5981 3657
rect 6015 3623 6049 3657
rect 6083 3623 6117 3657
rect 6151 3623 6185 3657
rect 6219 3623 6253 3657
rect 6287 3623 6321 3657
rect 6355 3623 6389 3657
rect 6423 3623 6457 3657
rect 6491 3623 6525 3657
rect 6559 3623 6593 3657
rect 6627 3623 6661 3657
rect 6695 3623 6729 3657
rect 6763 3623 6797 3657
rect 6831 3623 6865 3657
rect 6899 3623 6933 3657
rect 6967 3623 7001 3657
rect 7035 3623 7069 3657
rect 7103 3623 7137 3657
rect 7171 3623 7205 3657
rect 7239 3623 7273 3657
rect 7307 3623 7341 3657
rect 7375 3623 7409 3657
rect 7443 3623 7477 3657
rect 7511 3623 7545 3657
rect 7579 3623 7613 3657
rect 7647 3623 7681 3657
rect 7715 3623 7749 3657
rect 7783 3623 7817 3657
rect 7851 3623 7885 3657
rect 7919 3623 7953 3657
rect 7987 3623 8021 3657
rect 8055 3623 8089 3657
rect 8123 3623 8157 3657
rect 8191 3623 8225 3657
rect 8259 3623 8293 3657
rect 8327 3623 8361 3657
rect 8395 3623 8429 3657
rect 8463 3623 8497 3657
rect 8531 3623 8565 3657
rect 8599 3623 8633 3657
rect 8667 3623 8701 3657
rect 8735 3623 8769 3657
rect 8803 3623 8837 3657
rect 8871 3623 8905 3657
rect 8939 3623 8973 3657
rect 9007 3623 9041 3657
rect 9075 3623 9109 3657
rect 9143 3623 9177 3657
rect 9211 3623 9245 3657
rect 9279 3623 9313 3657
rect 9347 3623 9381 3657
rect 9415 3623 9449 3657
rect 9483 3623 9517 3657
rect 9551 3623 9585 3657
rect 9619 3623 9653 3657
rect 9687 3623 9721 3657
rect 9755 3623 9789 3657
rect 9823 3623 9857 3657
rect 9891 3623 9925 3657
rect 9959 3623 9993 3657
rect 10027 3623 10061 3657
rect 10095 3623 10129 3657
rect 10163 3623 10197 3657
rect 10231 3623 10265 3657
rect 10299 3623 10333 3657
rect 10367 3623 10401 3657
rect 10435 3623 10469 3657
rect 10503 3623 10537 3657
rect 10571 3623 10605 3657
rect 10639 3623 10673 3657
rect 10707 3623 10741 3657
rect 10775 3623 10809 3657
rect 10843 3623 10877 3657
rect 10911 3623 10945 3657
rect 10979 3623 11013 3657
rect 11047 3623 11081 3657
rect 11115 3623 11149 3657
rect 11183 3623 11217 3657
rect 11251 3623 11285 3657
rect 11319 3623 11353 3657
rect 11387 3623 11421 3657
rect 11455 3623 11489 3657
rect 11523 3623 11557 3657
rect 11591 3623 11625 3657
rect 11659 3623 11693 3657
rect 11727 3623 11761 3657
rect 11795 3623 11829 3657
rect 11863 3623 11897 3657
rect 11931 3623 11965 3657
rect 11999 3623 12033 3657
rect 12067 3623 12101 3657
rect 12135 3623 12169 3657
rect 12203 3623 12237 3657
rect 12271 3623 12305 3657
rect 12339 3623 12373 3657
rect 12407 3623 12441 3657
rect 12475 3623 12509 3657
rect 12543 3623 12577 3657
rect 12611 3623 12645 3657
rect 12679 3623 12713 3657
rect 12747 3623 12781 3657
rect 12815 3623 12849 3657
rect 12883 3623 12917 3657
rect 12951 3623 12985 3657
rect 13019 3623 13053 3657
rect 13087 3623 13121 3657
rect 13155 3623 13189 3657
rect 13223 3623 13257 3657
rect 13291 3623 13325 3657
rect 13359 3623 13393 3657
rect 13427 3623 13461 3657
rect 13495 3623 13529 3657
rect 13563 3623 13597 3657
rect 13631 3623 13665 3657
rect 13699 3623 13733 3657
rect 13767 3623 13801 3657
rect 13835 3623 13869 3657
rect 13903 3623 13937 3657
rect 13971 3623 14005 3657
rect 14039 3623 14073 3657
rect 14107 3623 14141 3657
rect 14175 3623 14209 3657
rect 14243 3623 14277 3657
rect 14311 3623 14345 3657
rect 14379 3623 14413 3657
rect 14447 3623 14481 3657
rect 14515 3623 14549 3657
rect 14583 3623 14617 3657
rect 14651 3623 14685 3657
rect 14719 3623 14880 3657
rect -12880 3600 14880 3623
rect -12880 3489 -12800 3600
rect -12880 3455 -12857 3489
rect -12823 3455 -12800 3489
rect -12880 3421 -12800 3455
rect -12880 3387 -12857 3421
rect -12823 3387 -12800 3421
rect -12880 3353 -12800 3387
rect -12880 3319 -12857 3353
rect -12823 3319 -12800 3353
rect -12880 3285 -12800 3319
rect -12880 3251 -12857 3285
rect -12823 3251 -12800 3285
rect -12880 3217 -12800 3251
rect -12880 3183 -12857 3217
rect -12823 3183 -12800 3217
rect -12880 3149 -12800 3183
rect -12880 3115 -12857 3149
rect -12823 3115 -12800 3149
rect -12880 3081 -12800 3115
rect -12880 3047 -12857 3081
rect -12823 3047 -12800 3081
rect -12880 3013 -12800 3047
rect -12880 2979 -12857 3013
rect -12823 2979 -12800 3013
rect -12880 2945 -12800 2979
rect -12880 2911 -12857 2945
rect -12823 2911 -12800 2945
rect -12880 2877 -12800 2911
rect -12880 2843 -12857 2877
rect -12823 2843 -12800 2877
rect -12880 2809 -12800 2843
rect -12880 2775 -12857 2809
rect -12823 2775 -12800 2809
rect -12880 2741 -12800 2775
rect -12880 2707 -12857 2741
rect -12823 2707 -12800 2741
rect -12880 2673 -12800 2707
rect -12880 2639 -12857 2673
rect -12823 2639 -12800 2673
rect -12880 2605 -12800 2639
rect -12880 2571 -12857 2605
rect -12823 2571 -12800 2605
rect -12880 2537 -12800 2571
rect -12880 2503 -12857 2537
rect -12823 2503 -12800 2537
rect -12880 2469 -12800 2503
rect -12880 2435 -12857 2469
rect -12823 2435 -12800 2469
rect -12880 2401 -12800 2435
rect -12880 2367 -12857 2401
rect -12823 2367 -12800 2401
rect -12880 2333 -12800 2367
rect -12880 2299 -12857 2333
rect -12823 2299 -12800 2333
rect -12880 2265 -12800 2299
rect -12880 2231 -12857 2265
rect -12823 2231 -12800 2265
rect -12880 2197 -12800 2231
rect -12880 2163 -12857 2197
rect -12823 2163 -12800 2197
rect -12880 2129 -12800 2163
rect -12880 2095 -12857 2129
rect -12823 2095 -12800 2129
rect -12880 2061 -12800 2095
rect -12880 2027 -12857 2061
rect -12823 2027 -12800 2061
rect -12880 1993 -12800 2027
rect -12880 1959 -12857 1993
rect -12823 1959 -12800 1993
rect -12880 1925 -12800 1959
rect -12880 1891 -12857 1925
rect -12823 1891 -12800 1925
rect -12880 1857 -12800 1891
rect -12880 1823 -12857 1857
rect -12823 1823 -12800 1857
rect -12880 1789 -12800 1823
rect -12880 1755 -12857 1789
rect -12823 1755 -12800 1789
rect -12880 1721 -12800 1755
rect -12880 1687 -12857 1721
rect -12823 1687 -12800 1721
rect -12880 1653 -12800 1687
rect -12880 1619 -12857 1653
rect -12823 1619 -12800 1653
rect -12880 1585 -12800 1619
rect -12880 1551 -12857 1585
rect -12823 1551 -12800 1585
rect -12880 1440 -12800 1551
rect 14800 3489 14880 3600
rect 14800 3455 14823 3489
rect 14857 3455 14880 3489
rect 14800 3421 14880 3455
rect 14800 3387 14823 3421
rect 14857 3387 14880 3421
rect 14800 3353 14880 3387
rect 14800 3319 14823 3353
rect 14857 3319 14880 3353
rect 14800 3285 14880 3319
rect 14800 3251 14823 3285
rect 14857 3251 14880 3285
rect 14800 3217 14880 3251
rect 14800 3183 14823 3217
rect 14857 3183 14880 3217
rect 14800 3149 14880 3183
rect 14800 3115 14823 3149
rect 14857 3115 14880 3149
rect 14800 3081 14880 3115
rect 14800 3047 14823 3081
rect 14857 3047 14880 3081
rect 14800 3013 14880 3047
rect 14800 2979 14823 3013
rect 14857 2979 14880 3013
rect 14800 2945 14880 2979
rect 14800 2911 14823 2945
rect 14857 2911 14880 2945
rect 14800 2877 14880 2911
rect 14800 2843 14823 2877
rect 14857 2843 14880 2877
rect 14800 2809 14880 2843
rect 14800 2775 14823 2809
rect 14857 2775 14880 2809
rect 14800 2741 14880 2775
rect 14800 2707 14823 2741
rect 14857 2707 14880 2741
rect 14800 2673 14880 2707
rect 14800 2639 14823 2673
rect 14857 2639 14880 2673
rect 14800 2605 14880 2639
rect 14800 2571 14823 2605
rect 14857 2571 14880 2605
rect 14800 2537 14880 2571
rect 14800 2503 14823 2537
rect 14857 2503 14880 2537
rect 14800 2469 14880 2503
rect 14800 2435 14823 2469
rect 14857 2435 14880 2469
rect 14800 2401 14880 2435
rect 14800 2367 14823 2401
rect 14857 2367 14880 2401
rect 14800 2333 14880 2367
rect 14800 2299 14823 2333
rect 14857 2299 14880 2333
rect 14800 2265 14880 2299
rect 14800 2231 14823 2265
rect 14857 2231 14880 2265
rect 14800 2197 14880 2231
rect 14800 2163 14823 2197
rect 14857 2163 14880 2197
rect 14800 2129 14880 2163
rect 14800 2095 14823 2129
rect 14857 2095 14880 2129
rect 14800 2061 14880 2095
rect 14800 2027 14823 2061
rect 14857 2027 14880 2061
rect 14800 1993 14880 2027
rect 14800 1959 14823 1993
rect 14857 1959 14880 1993
rect 14800 1925 14880 1959
rect 14800 1891 14823 1925
rect 14857 1891 14880 1925
rect 14800 1857 14880 1891
rect 14800 1823 14823 1857
rect 14857 1823 14880 1857
rect 14800 1789 14880 1823
rect 14800 1755 14823 1789
rect 14857 1755 14880 1789
rect 14800 1721 14880 1755
rect 14800 1687 14823 1721
rect 14857 1687 14880 1721
rect 14800 1653 14880 1687
rect 14800 1619 14823 1653
rect 14857 1619 14880 1653
rect 14800 1585 14880 1619
rect 14800 1551 14823 1585
rect 14857 1551 14880 1585
rect 14800 1440 14880 1551
rect -12880 1417 14880 1440
rect -12880 1383 -12719 1417
rect -12685 1383 -12651 1417
rect -12617 1383 -12583 1417
rect -12549 1383 -12515 1417
rect -12481 1383 -12447 1417
rect -12413 1383 -12379 1417
rect -12345 1383 -12311 1417
rect -12277 1383 -12243 1417
rect -12209 1383 -12175 1417
rect -12141 1383 -12107 1417
rect -12073 1383 -12039 1417
rect -12005 1383 -11971 1417
rect -11937 1383 -11903 1417
rect -11869 1383 -11835 1417
rect -11801 1383 -11767 1417
rect -11733 1383 -11699 1417
rect -11665 1383 -11631 1417
rect -11597 1383 -11563 1417
rect -11529 1383 -11495 1417
rect -11461 1383 -11427 1417
rect -11393 1383 -11359 1417
rect -11325 1383 -11291 1417
rect -11257 1383 -11223 1417
rect -11189 1383 -11155 1417
rect -11121 1383 -11087 1417
rect -11053 1383 -11019 1417
rect -10985 1383 -10951 1417
rect -10917 1383 -10883 1417
rect -10849 1383 -10815 1417
rect -10781 1383 -10747 1417
rect -10713 1383 -10679 1417
rect -10645 1383 -10611 1417
rect -10577 1383 -10543 1417
rect -10509 1383 -10475 1417
rect -10441 1383 -10407 1417
rect -10373 1383 -10339 1417
rect -10305 1383 -10271 1417
rect -10237 1383 -10203 1417
rect -10169 1383 -10135 1417
rect -10101 1383 -10067 1417
rect -10033 1383 -9999 1417
rect -9965 1383 -9931 1417
rect -9897 1383 -9863 1417
rect -9829 1383 -9795 1417
rect -9761 1383 -9727 1417
rect -9693 1383 -9659 1417
rect -9625 1383 -9591 1417
rect -9557 1383 -9523 1417
rect -9489 1383 -9455 1417
rect -9421 1383 -9387 1417
rect -9353 1383 -9319 1417
rect -9285 1383 -9251 1417
rect -9217 1383 -9183 1417
rect -9149 1383 -9115 1417
rect -9081 1383 -9047 1417
rect -9013 1383 -8979 1417
rect -8945 1383 -8911 1417
rect -8877 1383 -8843 1417
rect -8809 1383 -8775 1417
rect -8741 1383 -8707 1417
rect -8673 1383 -8639 1417
rect -8605 1383 -8571 1417
rect -8537 1383 -8503 1417
rect -8469 1383 -8435 1417
rect -8401 1383 -8367 1417
rect -8333 1383 -8299 1417
rect -8265 1383 -8231 1417
rect -8197 1383 -8163 1417
rect -8129 1383 -8095 1417
rect -8061 1383 -8027 1417
rect -7993 1383 -7959 1417
rect -7925 1383 -7891 1417
rect -7857 1383 -7823 1417
rect -7789 1383 -7755 1417
rect -7721 1383 -7687 1417
rect -7653 1383 -7619 1417
rect -7585 1383 -7551 1417
rect -7517 1383 -7483 1417
rect -7449 1383 -7415 1417
rect -7381 1383 -7347 1417
rect -7313 1383 -7279 1417
rect -7245 1383 -7211 1417
rect -7177 1383 -7143 1417
rect -7109 1383 -7075 1417
rect -7041 1383 -7007 1417
rect -6973 1383 -6939 1417
rect -6905 1383 -6871 1417
rect -6837 1383 -6803 1417
rect -6769 1383 -6735 1417
rect -6701 1383 -6667 1417
rect -6633 1383 -6599 1417
rect -6565 1383 -6531 1417
rect -6497 1383 -6463 1417
rect -6429 1383 -6395 1417
rect -6361 1383 -6327 1417
rect -6293 1383 -6259 1417
rect -6225 1383 -6191 1417
rect -6157 1383 -6123 1417
rect -6089 1383 -6055 1417
rect -6021 1383 -5987 1417
rect -5953 1383 -5919 1417
rect -5885 1383 -5851 1417
rect -5817 1383 -5783 1417
rect -5749 1383 -5715 1417
rect -5681 1383 -5647 1417
rect -5613 1383 -5579 1417
rect -5545 1383 -5511 1417
rect -5477 1383 -5443 1417
rect -5409 1383 -5375 1417
rect -5341 1383 -5307 1417
rect -5273 1383 -5239 1417
rect -5205 1383 -5171 1417
rect -5137 1383 -5103 1417
rect -5069 1383 -5035 1417
rect -5001 1383 -4967 1417
rect -4933 1383 -4899 1417
rect -4865 1383 -4831 1417
rect -4797 1383 -4763 1417
rect -4729 1383 -4695 1417
rect -4661 1383 -4627 1417
rect -4593 1383 -4559 1417
rect -4525 1383 -4491 1417
rect -4457 1383 -4423 1417
rect -4389 1383 -4355 1417
rect -4321 1383 -4287 1417
rect -4253 1383 -4219 1417
rect -4185 1383 -4151 1417
rect -4117 1383 -4083 1417
rect -4049 1383 -4015 1417
rect -3981 1383 -3947 1417
rect -3913 1383 -3879 1417
rect -3845 1383 -3811 1417
rect -3777 1383 -3743 1417
rect -3709 1383 -3675 1417
rect -3641 1383 -3607 1417
rect -3573 1383 -3539 1417
rect -3505 1383 -3471 1417
rect -3437 1383 -3403 1417
rect -3369 1383 -3335 1417
rect -3301 1383 -3267 1417
rect -3233 1383 -3199 1417
rect -3165 1383 -3131 1417
rect -3097 1383 -3063 1417
rect -3029 1383 -2995 1417
rect -2961 1383 -2927 1417
rect -2893 1383 -2859 1417
rect -2825 1383 -2791 1417
rect -2757 1383 -2723 1417
rect -2689 1383 -2655 1417
rect -2621 1383 -2587 1417
rect -2553 1383 -2519 1417
rect -2485 1383 -2451 1417
rect -2417 1383 -2383 1417
rect -2349 1383 -2315 1417
rect -2281 1383 -2247 1417
rect -2213 1383 -2179 1417
rect -2145 1383 -2111 1417
rect -2077 1383 -2043 1417
rect -2009 1383 -1975 1417
rect -1941 1383 -1907 1417
rect -1873 1383 -1839 1417
rect -1805 1383 -1771 1417
rect -1737 1383 -1703 1417
rect -1669 1383 -1635 1417
rect -1601 1383 -1567 1417
rect -1533 1383 -1499 1417
rect -1465 1383 -1431 1417
rect -1397 1383 -1363 1417
rect -1329 1383 -1295 1417
rect -1261 1383 -1227 1417
rect -1193 1383 -1159 1417
rect -1125 1383 -1091 1417
rect -1057 1383 -1023 1417
rect -989 1383 -955 1417
rect -921 1383 -887 1417
rect -853 1383 -819 1417
rect -785 1383 -751 1417
rect -717 1383 -683 1417
rect -649 1383 -615 1417
rect -581 1383 -547 1417
rect -513 1383 -479 1417
rect -445 1383 -411 1417
rect -377 1383 -343 1417
rect -309 1383 -275 1417
rect -241 1383 -207 1417
rect -173 1383 -139 1417
rect -105 1383 -71 1417
rect -37 1383 -3 1417
rect 31 1383 65 1417
rect 99 1383 133 1417
rect 167 1383 201 1417
rect 235 1383 269 1417
rect 303 1383 337 1417
rect 371 1383 405 1417
rect 439 1383 473 1417
rect 507 1383 541 1417
rect 575 1383 609 1417
rect 643 1383 677 1417
rect 711 1383 745 1417
rect 779 1383 813 1417
rect 847 1383 881 1417
rect 915 1383 949 1417
rect 983 1383 1017 1417
rect 1051 1383 1085 1417
rect 1119 1383 1153 1417
rect 1187 1383 1221 1417
rect 1255 1383 1289 1417
rect 1323 1383 1357 1417
rect 1391 1383 1425 1417
rect 1459 1383 1493 1417
rect 1527 1383 1561 1417
rect 1595 1383 1629 1417
rect 1663 1383 1697 1417
rect 1731 1383 1765 1417
rect 1799 1383 1833 1417
rect 1867 1383 1901 1417
rect 1935 1383 1969 1417
rect 2003 1383 2037 1417
rect 2071 1383 2105 1417
rect 2139 1383 2173 1417
rect 2207 1383 2241 1417
rect 2275 1383 2309 1417
rect 2343 1383 2377 1417
rect 2411 1383 2445 1417
rect 2479 1383 2513 1417
rect 2547 1383 2581 1417
rect 2615 1383 2649 1417
rect 2683 1383 2717 1417
rect 2751 1383 2785 1417
rect 2819 1383 2853 1417
rect 2887 1383 2921 1417
rect 2955 1383 2989 1417
rect 3023 1383 3057 1417
rect 3091 1383 3125 1417
rect 3159 1383 3193 1417
rect 3227 1383 3261 1417
rect 3295 1383 3329 1417
rect 3363 1383 3397 1417
rect 3431 1383 3465 1417
rect 3499 1383 3533 1417
rect 3567 1383 3601 1417
rect 3635 1383 3669 1417
rect 3703 1383 3737 1417
rect 3771 1383 3805 1417
rect 3839 1383 3873 1417
rect 3907 1383 3941 1417
rect 3975 1383 4009 1417
rect 4043 1383 4077 1417
rect 4111 1383 4145 1417
rect 4179 1383 4213 1417
rect 4247 1383 4281 1417
rect 4315 1383 4349 1417
rect 4383 1383 4417 1417
rect 4451 1383 4485 1417
rect 4519 1383 4553 1417
rect 4587 1383 4621 1417
rect 4655 1383 4689 1417
rect 4723 1383 4757 1417
rect 4791 1383 4825 1417
rect 4859 1383 4893 1417
rect 4927 1383 4961 1417
rect 4995 1383 5029 1417
rect 5063 1383 5097 1417
rect 5131 1383 5165 1417
rect 5199 1383 5233 1417
rect 5267 1383 5301 1417
rect 5335 1383 5369 1417
rect 5403 1383 5437 1417
rect 5471 1383 5505 1417
rect 5539 1383 5573 1417
rect 5607 1383 5641 1417
rect 5675 1383 5709 1417
rect 5743 1383 5777 1417
rect 5811 1383 5845 1417
rect 5879 1383 5913 1417
rect 5947 1383 5981 1417
rect 6015 1383 6049 1417
rect 6083 1383 6117 1417
rect 6151 1383 6185 1417
rect 6219 1383 6253 1417
rect 6287 1383 6321 1417
rect 6355 1383 6389 1417
rect 6423 1383 6457 1417
rect 6491 1383 6525 1417
rect 6559 1383 6593 1417
rect 6627 1383 6661 1417
rect 6695 1383 6729 1417
rect 6763 1383 6797 1417
rect 6831 1383 6865 1417
rect 6899 1383 6933 1417
rect 6967 1383 7001 1417
rect 7035 1383 7069 1417
rect 7103 1383 7137 1417
rect 7171 1383 7205 1417
rect 7239 1383 7273 1417
rect 7307 1383 7341 1417
rect 7375 1383 7409 1417
rect 7443 1383 7477 1417
rect 7511 1383 7545 1417
rect 7579 1383 7613 1417
rect 7647 1383 7681 1417
rect 7715 1383 7749 1417
rect 7783 1383 7817 1417
rect 7851 1383 7885 1417
rect 7919 1383 7953 1417
rect 7987 1383 8021 1417
rect 8055 1383 8089 1417
rect 8123 1383 8157 1417
rect 8191 1383 8225 1417
rect 8259 1383 8293 1417
rect 8327 1383 8361 1417
rect 8395 1383 8429 1417
rect 8463 1383 8497 1417
rect 8531 1383 8565 1417
rect 8599 1383 8633 1417
rect 8667 1383 8701 1417
rect 8735 1383 8769 1417
rect 8803 1383 8837 1417
rect 8871 1383 8905 1417
rect 8939 1383 8973 1417
rect 9007 1383 9041 1417
rect 9075 1383 9109 1417
rect 9143 1383 9177 1417
rect 9211 1383 9245 1417
rect 9279 1383 9313 1417
rect 9347 1383 9381 1417
rect 9415 1383 9449 1417
rect 9483 1383 9517 1417
rect 9551 1383 9585 1417
rect 9619 1383 9653 1417
rect 9687 1383 9721 1417
rect 9755 1383 9789 1417
rect 9823 1383 9857 1417
rect 9891 1383 9925 1417
rect 9959 1383 9993 1417
rect 10027 1383 10061 1417
rect 10095 1383 10129 1417
rect 10163 1383 10197 1417
rect 10231 1383 10265 1417
rect 10299 1383 10333 1417
rect 10367 1383 10401 1417
rect 10435 1383 10469 1417
rect 10503 1383 10537 1417
rect 10571 1383 10605 1417
rect 10639 1383 10673 1417
rect 10707 1383 10741 1417
rect 10775 1383 10809 1417
rect 10843 1383 10877 1417
rect 10911 1383 10945 1417
rect 10979 1383 11013 1417
rect 11047 1383 11081 1417
rect 11115 1383 11149 1417
rect 11183 1383 11217 1417
rect 11251 1383 11285 1417
rect 11319 1383 11353 1417
rect 11387 1383 11421 1417
rect 11455 1383 11489 1417
rect 11523 1383 11557 1417
rect 11591 1383 11625 1417
rect 11659 1383 11693 1417
rect 11727 1383 11761 1417
rect 11795 1383 11829 1417
rect 11863 1383 11897 1417
rect 11931 1383 11965 1417
rect 11999 1383 12033 1417
rect 12067 1383 12101 1417
rect 12135 1383 12169 1417
rect 12203 1383 12237 1417
rect 12271 1383 12305 1417
rect 12339 1383 12373 1417
rect 12407 1383 12441 1417
rect 12475 1383 12509 1417
rect 12543 1383 12577 1417
rect 12611 1383 12645 1417
rect 12679 1383 12713 1417
rect 12747 1383 12781 1417
rect 12815 1383 12849 1417
rect 12883 1383 12917 1417
rect 12951 1383 12985 1417
rect 13019 1383 13053 1417
rect 13087 1383 13121 1417
rect 13155 1383 13189 1417
rect 13223 1383 13257 1417
rect 13291 1383 13325 1417
rect 13359 1383 13393 1417
rect 13427 1383 13461 1417
rect 13495 1383 13529 1417
rect 13563 1383 13597 1417
rect 13631 1383 13665 1417
rect 13699 1383 13733 1417
rect 13767 1383 13801 1417
rect 13835 1383 13869 1417
rect 13903 1383 13937 1417
rect 13971 1383 14005 1417
rect 14039 1383 14073 1417
rect 14107 1383 14141 1417
rect 14175 1383 14209 1417
rect 14243 1383 14277 1417
rect 14311 1383 14345 1417
rect 14379 1383 14413 1417
rect 14447 1383 14481 1417
rect 14515 1383 14549 1417
rect 14583 1383 14617 1417
rect 14651 1383 14685 1417
rect 14719 1383 14880 1417
rect -12880 1360 14880 1383
<< psubdiffcont >>
rect -12719 3623 -12685 3657
rect -12651 3623 -12617 3657
rect -12583 3623 -12549 3657
rect -12515 3623 -12481 3657
rect -12447 3623 -12413 3657
rect -12379 3623 -12345 3657
rect -12311 3623 -12277 3657
rect -12243 3623 -12209 3657
rect -12175 3623 -12141 3657
rect -12107 3623 -12073 3657
rect -12039 3623 -12005 3657
rect -11971 3623 -11937 3657
rect -11903 3623 -11869 3657
rect -11835 3623 -11801 3657
rect -11767 3623 -11733 3657
rect -11699 3623 -11665 3657
rect -11631 3623 -11597 3657
rect -11563 3623 -11529 3657
rect -11495 3623 -11461 3657
rect -11427 3623 -11393 3657
rect -11359 3623 -11325 3657
rect -11291 3623 -11257 3657
rect -11223 3623 -11189 3657
rect -11155 3623 -11121 3657
rect -11087 3623 -11053 3657
rect -11019 3623 -10985 3657
rect -10951 3623 -10917 3657
rect -10883 3623 -10849 3657
rect -10815 3623 -10781 3657
rect -10747 3623 -10713 3657
rect -10679 3623 -10645 3657
rect -10611 3623 -10577 3657
rect -10543 3623 -10509 3657
rect -10475 3623 -10441 3657
rect -10407 3623 -10373 3657
rect -10339 3623 -10305 3657
rect -10271 3623 -10237 3657
rect -10203 3623 -10169 3657
rect -10135 3623 -10101 3657
rect -10067 3623 -10033 3657
rect -9999 3623 -9965 3657
rect -9931 3623 -9897 3657
rect -9863 3623 -9829 3657
rect -9795 3623 -9761 3657
rect -9727 3623 -9693 3657
rect -9659 3623 -9625 3657
rect -9591 3623 -9557 3657
rect -9523 3623 -9489 3657
rect -9455 3623 -9421 3657
rect -9387 3623 -9353 3657
rect -9319 3623 -9285 3657
rect -9251 3623 -9217 3657
rect -9183 3623 -9149 3657
rect -9115 3623 -9081 3657
rect -9047 3623 -9013 3657
rect -8979 3623 -8945 3657
rect -8911 3623 -8877 3657
rect -8843 3623 -8809 3657
rect -8775 3623 -8741 3657
rect -8707 3623 -8673 3657
rect -8639 3623 -8605 3657
rect -8571 3623 -8537 3657
rect -8503 3623 -8469 3657
rect -8435 3623 -8401 3657
rect -8367 3623 -8333 3657
rect -8299 3623 -8265 3657
rect -8231 3623 -8197 3657
rect -8163 3623 -8129 3657
rect -8095 3623 -8061 3657
rect -8027 3623 -7993 3657
rect -7959 3623 -7925 3657
rect -7891 3623 -7857 3657
rect -7823 3623 -7789 3657
rect -7755 3623 -7721 3657
rect -7687 3623 -7653 3657
rect -7619 3623 -7585 3657
rect -7551 3623 -7517 3657
rect -7483 3623 -7449 3657
rect -7415 3623 -7381 3657
rect -7347 3623 -7313 3657
rect -7279 3623 -7245 3657
rect -7211 3623 -7177 3657
rect -7143 3623 -7109 3657
rect -7075 3623 -7041 3657
rect -7007 3623 -6973 3657
rect -6939 3623 -6905 3657
rect -6871 3623 -6837 3657
rect -6803 3623 -6769 3657
rect -6735 3623 -6701 3657
rect -6667 3623 -6633 3657
rect -6599 3623 -6565 3657
rect -6531 3623 -6497 3657
rect -6463 3623 -6429 3657
rect -6395 3623 -6361 3657
rect -6327 3623 -6293 3657
rect -6259 3623 -6225 3657
rect -6191 3623 -6157 3657
rect -6123 3623 -6089 3657
rect -6055 3623 -6021 3657
rect -5987 3623 -5953 3657
rect -5919 3623 -5885 3657
rect -5851 3623 -5817 3657
rect -5783 3623 -5749 3657
rect -5715 3623 -5681 3657
rect -5647 3623 -5613 3657
rect -5579 3623 -5545 3657
rect -5511 3623 -5477 3657
rect -5443 3623 -5409 3657
rect -5375 3623 -5341 3657
rect -5307 3623 -5273 3657
rect -5239 3623 -5205 3657
rect -5171 3623 -5137 3657
rect -5103 3623 -5069 3657
rect -5035 3623 -5001 3657
rect -4967 3623 -4933 3657
rect -4899 3623 -4865 3657
rect -4831 3623 -4797 3657
rect -4763 3623 -4729 3657
rect -4695 3623 -4661 3657
rect -4627 3623 -4593 3657
rect -4559 3623 -4525 3657
rect -4491 3623 -4457 3657
rect -4423 3623 -4389 3657
rect -4355 3623 -4321 3657
rect -4287 3623 -4253 3657
rect -4219 3623 -4185 3657
rect -4151 3623 -4117 3657
rect -4083 3623 -4049 3657
rect -4015 3623 -3981 3657
rect -3947 3623 -3913 3657
rect -3879 3623 -3845 3657
rect -3811 3623 -3777 3657
rect -3743 3623 -3709 3657
rect -3675 3623 -3641 3657
rect -3607 3623 -3573 3657
rect -3539 3623 -3505 3657
rect -3471 3623 -3437 3657
rect -3403 3623 -3369 3657
rect -3335 3623 -3301 3657
rect -3267 3623 -3233 3657
rect -3199 3623 -3165 3657
rect -3131 3623 -3097 3657
rect -3063 3623 -3029 3657
rect -2995 3623 -2961 3657
rect -2927 3623 -2893 3657
rect -2859 3623 -2825 3657
rect -2791 3623 -2757 3657
rect -2723 3623 -2689 3657
rect -2655 3623 -2621 3657
rect -2587 3623 -2553 3657
rect -2519 3623 -2485 3657
rect -2451 3623 -2417 3657
rect -2383 3623 -2349 3657
rect -2315 3623 -2281 3657
rect -2247 3623 -2213 3657
rect -2179 3623 -2145 3657
rect -2111 3623 -2077 3657
rect -2043 3623 -2009 3657
rect -1975 3623 -1941 3657
rect -1907 3623 -1873 3657
rect -1839 3623 -1805 3657
rect -1771 3623 -1737 3657
rect -1703 3623 -1669 3657
rect -1635 3623 -1601 3657
rect -1567 3623 -1533 3657
rect -1499 3623 -1465 3657
rect -1431 3623 -1397 3657
rect -1363 3623 -1329 3657
rect -1295 3623 -1261 3657
rect -1227 3623 -1193 3657
rect -1159 3623 -1125 3657
rect -1091 3623 -1057 3657
rect -1023 3623 -989 3657
rect -955 3623 -921 3657
rect -887 3623 -853 3657
rect -819 3623 -785 3657
rect -751 3623 -717 3657
rect -683 3623 -649 3657
rect -615 3623 -581 3657
rect -547 3623 -513 3657
rect -479 3623 -445 3657
rect -411 3623 -377 3657
rect -343 3623 -309 3657
rect -275 3623 -241 3657
rect -207 3623 -173 3657
rect -139 3623 -105 3657
rect -71 3623 -37 3657
rect -3 3623 31 3657
rect 65 3623 99 3657
rect 133 3623 167 3657
rect 201 3623 235 3657
rect 269 3623 303 3657
rect 337 3623 371 3657
rect 405 3623 439 3657
rect 473 3623 507 3657
rect 541 3623 575 3657
rect 609 3623 643 3657
rect 677 3623 711 3657
rect 745 3623 779 3657
rect 813 3623 847 3657
rect 881 3623 915 3657
rect 949 3623 983 3657
rect 1017 3623 1051 3657
rect 1085 3623 1119 3657
rect 1153 3623 1187 3657
rect 1221 3623 1255 3657
rect 1289 3623 1323 3657
rect 1357 3623 1391 3657
rect 1425 3623 1459 3657
rect 1493 3623 1527 3657
rect 1561 3623 1595 3657
rect 1629 3623 1663 3657
rect 1697 3623 1731 3657
rect 1765 3623 1799 3657
rect 1833 3623 1867 3657
rect 1901 3623 1935 3657
rect 1969 3623 2003 3657
rect 2037 3623 2071 3657
rect 2105 3623 2139 3657
rect 2173 3623 2207 3657
rect 2241 3623 2275 3657
rect 2309 3623 2343 3657
rect 2377 3623 2411 3657
rect 2445 3623 2479 3657
rect 2513 3623 2547 3657
rect 2581 3623 2615 3657
rect 2649 3623 2683 3657
rect 2717 3623 2751 3657
rect 2785 3623 2819 3657
rect 2853 3623 2887 3657
rect 2921 3623 2955 3657
rect 2989 3623 3023 3657
rect 3057 3623 3091 3657
rect 3125 3623 3159 3657
rect 3193 3623 3227 3657
rect 3261 3623 3295 3657
rect 3329 3623 3363 3657
rect 3397 3623 3431 3657
rect 3465 3623 3499 3657
rect 3533 3623 3567 3657
rect 3601 3623 3635 3657
rect 3669 3623 3703 3657
rect 3737 3623 3771 3657
rect 3805 3623 3839 3657
rect 3873 3623 3907 3657
rect 3941 3623 3975 3657
rect 4009 3623 4043 3657
rect 4077 3623 4111 3657
rect 4145 3623 4179 3657
rect 4213 3623 4247 3657
rect 4281 3623 4315 3657
rect 4349 3623 4383 3657
rect 4417 3623 4451 3657
rect 4485 3623 4519 3657
rect 4553 3623 4587 3657
rect 4621 3623 4655 3657
rect 4689 3623 4723 3657
rect 4757 3623 4791 3657
rect 4825 3623 4859 3657
rect 4893 3623 4927 3657
rect 4961 3623 4995 3657
rect 5029 3623 5063 3657
rect 5097 3623 5131 3657
rect 5165 3623 5199 3657
rect 5233 3623 5267 3657
rect 5301 3623 5335 3657
rect 5369 3623 5403 3657
rect 5437 3623 5471 3657
rect 5505 3623 5539 3657
rect 5573 3623 5607 3657
rect 5641 3623 5675 3657
rect 5709 3623 5743 3657
rect 5777 3623 5811 3657
rect 5845 3623 5879 3657
rect 5913 3623 5947 3657
rect 5981 3623 6015 3657
rect 6049 3623 6083 3657
rect 6117 3623 6151 3657
rect 6185 3623 6219 3657
rect 6253 3623 6287 3657
rect 6321 3623 6355 3657
rect 6389 3623 6423 3657
rect 6457 3623 6491 3657
rect 6525 3623 6559 3657
rect 6593 3623 6627 3657
rect 6661 3623 6695 3657
rect 6729 3623 6763 3657
rect 6797 3623 6831 3657
rect 6865 3623 6899 3657
rect 6933 3623 6967 3657
rect 7001 3623 7035 3657
rect 7069 3623 7103 3657
rect 7137 3623 7171 3657
rect 7205 3623 7239 3657
rect 7273 3623 7307 3657
rect 7341 3623 7375 3657
rect 7409 3623 7443 3657
rect 7477 3623 7511 3657
rect 7545 3623 7579 3657
rect 7613 3623 7647 3657
rect 7681 3623 7715 3657
rect 7749 3623 7783 3657
rect 7817 3623 7851 3657
rect 7885 3623 7919 3657
rect 7953 3623 7987 3657
rect 8021 3623 8055 3657
rect 8089 3623 8123 3657
rect 8157 3623 8191 3657
rect 8225 3623 8259 3657
rect 8293 3623 8327 3657
rect 8361 3623 8395 3657
rect 8429 3623 8463 3657
rect 8497 3623 8531 3657
rect 8565 3623 8599 3657
rect 8633 3623 8667 3657
rect 8701 3623 8735 3657
rect 8769 3623 8803 3657
rect 8837 3623 8871 3657
rect 8905 3623 8939 3657
rect 8973 3623 9007 3657
rect 9041 3623 9075 3657
rect 9109 3623 9143 3657
rect 9177 3623 9211 3657
rect 9245 3623 9279 3657
rect 9313 3623 9347 3657
rect 9381 3623 9415 3657
rect 9449 3623 9483 3657
rect 9517 3623 9551 3657
rect 9585 3623 9619 3657
rect 9653 3623 9687 3657
rect 9721 3623 9755 3657
rect 9789 3623 9823 3657
rect 9857 3623 9891 3657
rect 9925 3623 9959 3657
rect 9993 3623 10027 3657
rect 10061 3623 10095 3657
rect 10129 3623 10163 3657
rect 10197 3623 10231 3657
rect 10265 3623 10299 3657
rect 10333 3623 10367 3657
rect 10401 3623 10435 3657
rect 10469 3623 10503 3657
rect 10537 3623 10571 3657
rect 10605 3623 10639 3657
rect 10673 3623 10707 3657
rect 10741 3623 10775 3657
rect 10809 3623 10843 3657
rect 10877 3623 10911 3657
rect 10945 3623 10979 3657
rect 11013 3623 11047 3657
rect 11081 3623 11115 3657
rect 11149 3623 11183 3657
rect 11217 3623 11251 3657
rect 11285 3623 11319 3657
rect 11353 3623 11387 3657
rect 11421 3623 11455 3657
rect 11489 3623 11523 3657
rect 11557 3623 11591 3657
rect 11625 3623 11659 3657
rect 11693 3623 11727 3657
rect 11761 3623 11795 3657
rect 11829 3623 11863 3657
rect 11897 3623 11931 3657
rect 11965 3623 11999 3657
rect 12033 3623 12067 3657
rect 12101 3623 12135 3657
rect 12169 3623 12203 3657
rect 12237 3623 12271 3657
rect 12305 3623 12339 3657
rect 12373 3623 12407 3657
rect 12441 3623 12475 3657
rect 12509 3623 12543 3657
rect 12577 3623 12611 3657
rect 12645 3623 12679 3657
rect 12713 3623 12747 3657
rect 12781 3623 12815 3657
rect 12849 3623 12883 3657
rect 12917 3623 12951 3657
rect 12985 3623 13019 3657
rect 13053 3623 13087 3657
rect 13121 3623 13155 3657
rect 13189 3623 13223 3657
rect 13257 3623 13291 3657
rect 13325 3623 13359 3657
rect 13393 3623 13427 3657
rect 13461 3623 13495 3657
rect 13529 3623 13563 3657
rect 13597 3623 13631 3657
rect 13665 3623 13699 3657
rect 13733 3623 13767 3657
rect 13801 3623 13835 3657
rect 13869 3623 13903 3657
rect 13937 3623 13971 3657
rect 14005 3623 14039 3657
rect 14073 3623 14107 3657
rect 14141 3623 14175 3657
rect 14209 3623 14243 3657
rect 14277 3623 14311 3657
rect 14345 3623 14379 3657
rect 14413 3623 14447 3657
rect 14481 3623 14515 3657
rect 14549 3623 14583 3657
rect 14617 3623 14651 3657
rect 14685 3623 14719 3657
rect -12857 3455 -12823 3489
rect -12857 3387 -12823 3421
rect -12857 3319 -12823 3353
rect -12857 3251 -12823 3285
rect -12857 3183 -12823 3217
rect -12857 3115 -12823 3149
rect -12857 3047 -12823 3081
rect -12857 2979 -12823 3013
rect -12857 2911 -12823 2945
rect -12857 2843 -12823 2877
rect -12857 2775 -12823 2809
rect -12857 2707 -12823 2741
rect -12857 2639 -12823 2673
rect -12857 2571 -12823 2605
rect -12857 2503 -12823 2537
rect -12857 2435 -12823 2469
rect -12857 2367 -12823 2401
rect -12857 2299 -12823 2333
rect -12857 2231 -12823 2265
rect -12857 2163 -12823 2197
rect -12857 2095 -12823 2129
rect -12857 2027 -12823 2061
rect -12857 1959 -12823 1993
rect -12857 1891 -12823 1925
rect -12857 1823 -12823 1857
rect -12857 1755 -12823 1789
rect -12857 1687 -12823 1721
rect -12857 1619 -12823 1653
rect -12857 1551 -12823 1585
rect 14823 3455 14857 3489
rect 14823 3387 14857 3421
rect 14823 3319 14857 3353
rect 14823 3251 14857 3285
rect 14823 3183 14857 3217
rect 14823 3115 14857 3149
rect 14823 3047 14857 3081
rect 14823 2979 14857 3013
rect 14823 2911 14857 2945
rect 14823 2843 14857 2877
rect 14823 2775 14857 2809
rect 14823 2707 14857 2741
rect 14823 2639 14857 2673
rect 14823 2571 14857 2605
rect 14823 2503 14857 2537
rect 14823 2435 14857 2469
rect 14823 2367 14857 2401
rect 14823 2299 14857 2333
rect 14823 2231 14857 2265
rect 14823 2163 14857 2197
rect 14823 2095 14857 2129
rect 14823 2027 14857 2061
rect 14823 1959 14857 1993
rect 14823 1891 14857 1925
rect 14823 1823 14857 1857
rect 14823 1755 14857 1789
rect 14823 1687 14857 1721
rect 14823 1619 14857 1653
rect 14823 1551 14857 1585
rect -12719 1383 -12685 1417
rect -12651 1383 -12617 1417
rect -12583 1383 -12549 1417
rect -12515 1383 -12481 1417
rect -12447 1383 -12413 1417
rect -12379 1383 -12345 1417
rect -12311 1383 -12277 1417
rect -12243 1383 -12209 1417
rect -12175 1383 -12141 1417
rect -12107 1383 -12073 1417
rect -12039 1383 -12005 1417
rect -11971 1383 -11937 1417
rect -11903 1383 -11869 1417
rect -11835 1383 -11801 1417
rect -11767 1383 -11733 1417
rect -11699 1383 -11665 1417
rect -11631 1383 -11597 1417
rect -11563 1383 -11529 1417
rect -11495 1383 -11461 1417
rect -11427 1383 -11393 1417
rect -11359 1383 -11325 1417
rect -11291 1383 -11257 1417
rect -11223 1383 -11189 1417
rect -11155 1383 -11121 1417
rect -11087 1383 -11053 1417
rect -11019 1383 -10985 1417
rect -10951 1383 -10917 1417
rect -10883 1383 -10849 1417
rect -10815 1383 -10781 1417
rect -10747 1383 -10713 1417
rect -10679 1383 -10645 1417
rect -10611 1383 -10577 1417
rect -10543 1383 -10509 1417
rect -10475 1383 -10441 1417
rect -10407 1383 -10373 1417
rect -10339 1383 -10305 1417
rect -10271 1383 -10237 1417
rect -10203 1383 -10169 1417
rect -10135 1383 -10101 1417
rect -10067 1383 -10033 1417
rect -9999 1383 -9965 1417
rect -9931 1383 -9897 1417
rect -9863 1383 -9829 1417
rect -9795 1383 -9761 1417
rect -9727 1383 -9693 1417
rect -9659 1383 -9625 1417
rect -9591 1383 -9557 1417
rect -9523 1383 -9489 1417
rect -9455 1383 -9421 1417
rect -9387 1383 -9353 1417
rect -9319 1383 -9285 1417
rect -9251 1383 -9217 1417
rect -9183 1383 -9149 1417
rect -9115 1383 -9081 1417
rect -9047 1383 -9013 1417
rect -8979 1383 -8945 1417
rect -8911 1383 -8877 1417
rect -8843 1383 -8809 1417
rect -8775 1383 -8741 1417
rect -8707 1383 -8673 1417
rect -8639 1383 -8605 1417
rect -8571 1383 -8537 1417
rect -8503 1383 -8469 1417
rect -8435 1383 -8401 1417
rect -8367 1383 -8333 1417
rect -8299 1383 -8265 1417
rect -8231 1383 -8197 1417
rect -8163 1383 -8129 1417
rect -8095 1383 -8061 1417
rect -8027 1383 -7993 1417
rect -7959 1383 -7925 1417
rect -7891 1383 -7857 1417
rect -7823 1383 -7789 1417
rect -7755 1383 -7721 1417
rect -7687 1383 -7653 1417
rect -7619 1383 -7585 1417
rect -7551 1383 -7517 1417
rect -7483 1383 -7449 1417
rect -7415 1383 -7381 1417
rect -7347 1383 -7313 1417
rect -7279 1383 -7245 1417
rect -7211 1383 -7177 1417
rect -7143 1383 -7109 1417
rect -7075 1383 -7041 1417
rect -7007 1383 -6973 1417
rect -6939 1383 -6905 1417
rect -6871 1383 -6837 1417
rect -6803 1383 -6769 1417
rect -6735 1383 -6701 1417
rect -6667 1383 -6633 1417
rect -6599 1383 -6565 1417
rect -6531 1383 -6497 1417
rect -6463 1383 -6429 1417
rect -6395 1383 -6361 1417
rect -6327 1383 -6293 1417
rect -6259 1383 -6225 1417
rect -6191 1383 -6157 1417
rect -6123 1383 -6089 1417
rect -6055 1383 -6021 1417
rect -5987 1383 -5953 1417
rect -5919 1383 -5885 1417
rect -5851 1383 -5817 1417
rect -5783 1383 -5749 1417
rect -5715 1383 -5681 1417
rect -5647 1383 -5613 1417
rect -5579 1383 -5545 1417
rect -5511 1383 -5477 1417
rect -5443 1383 -5409 1417
rect -5375 1383 -5341 1417
rect -5307 1383 -5273 1417
rect -5239 1383 -5205 1417
rect -5171 1383 -5137 1417
rect -5103 1383 -5069 1417
rect -5035 1383 -5001 1417
rect -4967 1383 -4933 1417
rect -4899 1383 -4865 1417
rect -4831 1383 -4797 1417
rect -4763 1383 -4729 1417
rect -4695 1383 -4661 1417
rect -4627 1383 -4593 1417
rect -4559 1383 -4525 1417
rect -4491 1383 -4457 1417
rect -4423 1383 -4389 1417
rect -4355 1383 -4321 1417
rect -4287 1383 -4253 1417
rect -4219 1383 -4185 1417
rect -4151 1383 -4117 1417
rect -4083 1383 -4049 1417
rect -4015 1383 -3981 1417
rect -3947 1383 -3913 1417
rect -3879 1383 -3845 1417
rect -3811 1383 -3777 1417
rect -3743 1383 -3709 1417
rect -3675 1383 -3641 1417
rect -3607 1383 -3573 1417
rect -3539 1383 -3505 1417
rect -3471 1383 -3437 1417
rect -3403 1383 -3369 1417
rect -3335 1383 -3301 1417
rect -3267 1383 -3233 1417
rect -3199 1383 -3165 1417
rect -3131 1383 -3097 1417
rect -3063 1383 -3029 1417
rect -2995 1383 -2961 1417
rect -2927 1383 -2893 1417
rect -2859 1383 -2825 1417
rect -2791 1383 -2757 1417
rect -2723 1383 -2689 1417
rect -2655 1383 -2621 1417
rect -2587 1383 -2553 1417
rect -2519 1383 -2485 1417
rect -2451 1383 -2417 1417
rect -2383 1383 -2349 1417
rect -2315 1383 -2281 1417
rect -2247 1383 -2213 1417
rect -2179 1383 -2145 1417
rect -2111 1383 -2077 1417
rect -2043 1383 -2009 1417
rect -1975 1383 -1941 1417
rect -1907 1383 -1873 1417
rect -1839 1383 -1805 1417
rect -1771 1383 -1737 1417
rect -1703 1383 -1669 1417
rect -1635 1383 -1601 1417
rect -1567 1383 -1533 1417
rect -1499 1383 -1465 1417
rect -1431 1383 -1397 1417
rect -1363 1383 -1329 1417
rect -1295 1383 -1261 1417
rect -1227 1383 -1193 1417
rect -1159 1383 -1125 1417
rect -1091 1383 -1057 1417
rect -1023 1383 -989 1417
rect -955 1383 -921 1417
rect -887 1383 -853 1417
rect -819 1383 -785 1417
rect -751 1383 -717 1417
rect -683 1383 -649 1417
rect -615 1383 -581 1417
rect -547 1383 -513 1417
rect -479 1383 -445 1417
rect -411 1383 -377 1417
rect -343 1383 -309 1417
rect -275 1383 -241 1417
rect -207 1383 -173 1417
rect -139 1383 -105 1417
rect -71 1383 -37 1417
rect -3 1383 31 1417
rect 65 1383 99 1417
rect 133 1383 167 1417
rect 201 1383 235 1417
rect 269 1383 303 1417
rect 337 1383 371 1417
rect 405 1383 439 1417
rect 473 1383 507 1417
rect 541 1383 575 1417
rect 609 1383 643 1417
rect 677 1383 711 1417
rect 745 1383 779 1417
rect 813 1383 847 1417
rect 881 1383 915 1417
rect 949 1383 983 1417
rect 1017 1383 1051 1417
rect 1085 1383 1119 1417
rect 1153 1383 1187 1417
rect 1221 1383 1255 1417
rect 1289 1383 1323 1417
rect 1357 1383 1391 1417
rect 1425 1383 1459 1417
rect 1493 1383 1527 1417
rect 1561 1383 1595 1417
rect 1629 1383 1663 1417
rect 1697 1383 1731 1417
rect 1765 1383 1799 1417
rect 1833 1383 1867 1417
rect 1901 1383 1935 1417
rect 1969 1383 2003 1417
rect 2037 1383 2071 1417
rect 2105 1383 2139 1417
rect 2173 1383 2207 1417
rect 2241 1383 2275 1417
rect 2309 1383 2343 1417
rect 2377 1383 2411 1417
rect 2445 1383 2479 1417
rect 2513 1383 2547 1417
rect 2581 1383 2615 1417
rect 2649 1383 2683 1417
rect 2717 1383 2751 1417
rect 2785 1383 2819 1417
rect 2853 1383 2887 1417
rect 2921 1383 2955 1417
rect 2989 1383 3023 1417
rect 3057 1383 3091 1417
rect 3125 1383 3159 1417
rect 3193 1383 3227 1417
rect 3261 1383 3295 1417
rect 3329 1383 3363 1417
rect 3397 1383 3431 1417
rect 3465 1383 3499 1417
rect 3533 1383 3567 1417
rect 3601 1383 3635 1417
rect 3669 1383 3703 1417
rect 3737 1383 3771 1417
rect 3805 1383 3839 1417
rect 3873 1383 3907 1417
rect 3941 1383 3975 1417
rect 4009 1383 4043 1417
rect 4077 1383 4111 1417
rect 4145 1383 4179 1417
rect 4213 1383 4247 1417
rect 4281 1383 4315 1417
rect 4349 1383 4383 1417
rect 4417 1383 4451 1417
rect 4485 1383 4519 1417
rect 4553 1383 4587 1417
rect 4621 1383 4655 1417
rect 4689 1383 4723 1417
rect 4757 1383 4791 1417
rect 4825 1383 4859 1417
rect 4893 1383 4927 1417
rect 4961 1383 4995 1417
rect 5029 1383 5063 1417
rect 5097 1383 5131 1417
rect 5165 1383 5199 1417
rect 5233 1383 5267 1417
rect 5301 1383 5335 1417
rect 5369 1383 5403 1417
rect 5437 1383 5471 1417
rect 5505 1383 5539 1417
rect 5573 1383 5607 1417
rect 5641 1383 5675 1417
rect 5709 1383 5743 1417
rect 5777 1383 5811 1417
rect 5845 1383 5879 1417
rect 5913 1383 5947 1417
rect 5981 1383 6015 1417
rect 6049 1383 6083 1417
rect 6117 1383 6151 1417
rect 6185 1383 6219 1417
rect 6253 1383 6287 1417
rect 6321 1383 6355 1417
rect 6389 1383 6423 1417
rect 6457 1383 6491 1417
rect 6525 1383 6559 1417
rect 6593 1383 6627 1417
rect 6661 1383 6695 1417
rect 6729 1383 6763 1417
rect 6797 1383 6831 1417
rect 6865 1383 6899 1417
rect 6933 1383 6967 1417
rect 7001 1383 7035 1417
rect 7069 1383 7103 1417
rect 7137 1383 7171 1417
rect 7205 1383 7239 1417
rect 7273 1383 7307 1417
rect 7341 1383 7375 1417
rect 7409 1383 7443 1417
rect 7477 1383 7511 1417
rect 7545 1383 7579 1417
rect 7613 1383 7647 1417
rect 7681 1383 7715 1417
rect 7749 1383 7783 1417
rect 7817 1383 7851 1417
rect 7885 1383 7919 1417
rect 7953 1383 7987 1417
rect 8021 1383 8055 1417
rect 8089 1383 8123 1417
rect 8157 1383 8191 1417
rect 8225 1383 8259 1417
rect 8293 1383 8327 1417
rect 8361 1383 8395 1417
rect 8429 1383 8463 1417
rect 8497 1383 8531 1417
rect 8565 1383 8599 1417
rect 8633 1383 8667 1417
rect 8701 1383 8735 1417
rect 8769 1383 8803 1417
rect 8837 1383 8871 1417
rect 8905 1383 8939 1417
rect 8973 1383 9007 1417
rect 9041 1383 9075 1417
rect 9109 1383 9143 1417
rect 9177 1383 9211 1417
rect 9245 1383 9279 1417
rect 9313 1383 9347 1417
rect 9381 1383 9415 1417
rect 9449 1383 9483 1417
rect 9517 1383 9551 1417
rect 9585 1383 9619 1417
rect 9653 1383 9687 1417
rect 9721 1383 9755 1417
rect 9789 1383 9823 1417
rect 9857 1383 9891 1417
rect 9925 1383 9959 1417
rect 9993 1383 10027 1417
rect 10061 1383 10095 1417
rect 10129 1383 10163 1417
rect 10197 1383 10231 1417
rect 10265 1383 10299 1417
rect 10333 1383 10367 1417
rect 10401 1383 10435 1417
rect 10469 1383 10503 1417
rect 10537 1383 10571 1417
rect 10605 1383 10639 1417
rect 10673 1383 10707 1417
rect 10741 1383 10775 1417
rect 10809 1383 10843 1417
rect 10877 1383 10911 1417
rect 10945 1383 10979 1417
rect 11013 1383 11047 1417
rect 11081 1383 11115 1417
rect 11149 1383 11183 1417
rect 11217 1383 11251 1417
rect 11285 1383 11319 1417
rect 11353 1383 11387 1417
rect 11421 1383 11455 1417
rect 11489 1383 11523 1417
rect 11557 1383 11591 1417
rect 11625 1383 11659 1417
rect 11693 1383 11727 1417
rect 11761 1383 11795 1417
rect 11829 1383 11863 1417
rect 11897 1383 11931 1417
rect 11965 1383 11999 1417
rect 12033 1383 12067 1417
rect 12101 1383 12135 1417
rect 12169 1383 12203 1417
rect 12237 1383 12271 1417
rect 12305 1383 12339 1417
rect 12373 1383 12407 1417
rect 12441 1383 12475 1417
rect 12509 1383 12543 1417
rect 12577 1383 12611 1417
rect 12645 1383 12679 1417
rect 12713 1383 12747 1417
rect 12781 1383 12815 1417
rect 12849 1383 12883 1417
rect 12917 1383 12951 1417
rect 12985 1383 13019 1417
rect 13053 1383 13087 1417
rect 13121 1383 13155 1417
rect 13189 1383 13223 1417
rect 13257 1383 13291 1417
rect 13325 1383 13359 1417
rect 13393 1383 13427 1417
rect 13461 1383 13495 1417
rect 13529 1383 13563 1417
rect 13597 1383 13631 1417
rect 13665 1383 13699 1417
rect 13733 1383 13767 1417
rect 13801 1383 13835 1417
rect 13869 1383 13903 1417
rect 13937 1383 13971 1417
rect 14005 1383 14039 1417
rect 14073 1383 14107 1417
rect 14141 1383 14175 1417
rect 14209 1383 14243 1417
rect 14277 1383 14311 1417
rect 14345 1383 14379 1417
rect 14413 1383 14447 1417
rect 14481 1383 14515 1417
rect 14549 1383 14583 1417
rect 14617 1383 14651 1417
rect 14685 1383 14719 1417
<< locali >>
rect -12880 3657 14880 3680
rect -12880 3623 -12719 3657
rect -12685 3623 -12651 3657
rect -12617 3623 -12583 3657
rect -12549 3623 -12515 3657
rect -12481 3623 -12447 3657
rect -12413 3623 -12379 3657
rect -12345 3623 -12311 3657
rect -12277 3623 -12243 3657
rect -12209 3623 -12175 3657
rect -12141 3623 -12107 3657
rect -12073 3623 -12039 3657
rect -12005 3623 -11971 3657
rect -11937 3623 -11903 3657
rect -11869 3623 -11835 3657
rect -11801 3623 -11767 3657
rect -11733 3623 -11699 3657
rect -11665 3623 -11631 3657
rect -11597 3623 -11563 3657
rect -11529 3623 -11495 3657
rect -11461 3623 -11427 3657
rect -11393 3623 -11359 3657
rect -11325 3623 -11291 3657
rect -11257 3623 -11223 3657
rect -11189 3623 -11155 3657
rect -11121 3623 -11087 3657
rect -11053 3623 -11019 3657
rect -10985 3623 -10951 3657
rect -10917 3623 -10883 3657
rect -10849 3623 -10815 3657
rect -10781 3623 -10747 3657
rect -10713 3623 -10679 3657
rect -10645 3623 -10611 3657
rect -10577 3623 -10543 3657
rect -10509 3623 -10475 3657
rect -10441 3623 -10407 3657
rect -10373 3623 -10339 3657
rect -10305 3623 -10271 3657
rect -10237 3623 -10203 3657
rect -10169 3623 -10135 3657
rect -10101 3623 -10067 3657
rect -10033 3623 -9999 3657
rect -9965 3623 -9931 3657
rect -9897 3623 -9863 3657
rect -9829 3623 -9795 3657
rect -9761 3623 -9727 3657
rect -9693 3623 -9659 3657
rect -9625 3623 -9591 3657
rect -9557 3623 -9523 3657
rect -9489 3623 -9455 3657
rect -9421 3623 -9387 3657
rect -9353 3623 -9319 3657
rect -9285 3623 -9251 3657
rect -9217 3623 -9183 3657
rect -9149 3623 -9115 3657
rect -9081 3623 -9047 3657
rect -9013 3623 -8979 3657
rect -8945 3623 -8911 3657
rect -8877 3623 -8843 3657
rect -8809 3623 -8775 3657
rect -8741 3623 -8707 3657
rect -8673 3623 -8639 3657
rect -8605 3623 -8571 3657
rect -8537 3623 -8503 3657
rect -8469 3623 -8435 3657
rect -8401 3623 -8367 3657
rect -8333 3623 -8299 3657
rect -8265 3623 -8231 3657
rect -8197 3623 -8163 3657
rect -8129 3623 -8095 3657
rect -8061 3623 -8027 3657
rect -7993 3623 -7959 3657
rect -7925 3623 -7891 3657
rect -7857 3623 -7823 3657
rect -7789 3623 -7755 3657
rect -7721 3623 -7687 3657
rect -7653 3623 -7619 3657
rect -7585 3623 -7551 3657
rect -7517 3623 -7483 3657
rect -7449 3623 -7415 3657
rect -7381 3623 -7347 3657
rect -7313 3623 -7279 3657
rect -7245 3623 -7211 3657
rect -7177 3623 -7143 3657
rect -7109 3623 -7075 3657
rect -7041 3623 -7007 3657
rect -6973 3623 -6939 3657
rect -6905 3623 -6871 3657
rect -6837 3623 -6803 3657
rect -6769 3623 -6735 3657
rect -6701 3623 -6667 3657
rect -6633 3623 -6599 3657
rect -6565 3623 -6531 3657
rect -6497 3623 -6463 3657
rect -6429 3623 -6395 3657
rect -6361 3623 -6327 3657
rect -6293 3623 -6259 3657
rect -6225 3623 -6191 3657
rect -6157 3623 -6123 3657
rect -6089 3623 -6055 3657
rect -6021 3623 -5987 3657
rect -5953 3623 -5919 3657
rect -5885 3623 -5851 3657
rect -5817 3623 -5783 3657
rect -5749 3623 -5715 3657
rect -5681 3623 -5647 3657
rect -5613 3623 -5579 3657
rect -5545 3623 -5511 3657
rect -5477 3623 -5443 3657
rect -5409 3623 -5375 3657
rect -5341 3623 -5307 3657
rect -5273 3623 -5239 3657
rect -5205 3623 -5171 3657
rect -5137 3623 -5103 3657
rect -5069 3623 -5035 3657
rect -5001 3623 -4967 3657
rect -4933 3623 -4899 3657
rect -4865 3623 -4831 3657
rect -4797 3623 -4763 3657
rect -4729 3623 -4695 3657
rect -4661 3623 -4627 3657
rect -4593 3623 -4559 3657
rect -4525 3623 -4491 3657
rect -4457 3623 -4423 3657
rect -4389 3623 -4355 3657
rect -4321 3623 -4287 3657
rect -4253 3623 -4219 3657
rect -4185 3623 -4151 3657
rect -4117 3623 -4083 3657
rect -4049 3623 -4015 3657
rect -3981 3623 -3947 3657
rect -3913 3623 -3879 3657
rect -3845 3623 -3811 3657
rect -3777 3623 -3743 3657
rect -3709 3623 -3675 3657
rect -3641 3623 -3607 3657
rect -3573 3623 -3539 3657
rect -3505 3623 -3471 3657
rect -3437 3623 -3403 3657
rect -3369 3623 -3335 3657
rect -3301 3623 -3267 3657
rect -3233 3623 -3199 3657
rect -3165 3623 -3131 3657
rect -3097 3623 -3063 3657
rect -3029 3623 -2995 3657
rect -2961 3623 -2927 3657
rect -2893 3623 -2859 3657
rect -2825 3623 -2791 3657
rect -2757 3623 -2723 3657
rect -2689 3623 -2655 3657
rect -2621 3623 -2587 3657
rect -2553 3623 -2519 3657
rect -2485 3623 -2451 3657
rect -2417 3623 -2383 3657
rect -2349 3623 -2315 3657
rect -2281 3623 -2247 3657
rect -2213 3623 -2179 3657
rect -2145 3623 -2111 3657
rect -2077 3623 -2043 3657
rect -2009 3623 -1975 3657
rect -1941 3623 -1907 3657
rect -1873 3623 -1839 3657
rect -1805 3623 -1771 3657
rect -1737 3623 -1703 3657
rect -1669 3623 -1635 3657
rect -1601 3623 -1567 3657
rect -1533 3623 -1499 3657
rect -1465 3623 -1431 3657
rect -1397 3623 -1363 3657
rect -1329 3623 -1295 3657
rect -1261 3623 -1227 3657
rect -1193 3623 -1159 3657
rect -1125 3623 -1091 3657
rect -1057 3623 -1023 3657
rect -989 3623 -955 3657
rect -921 3623 -887 3657
rect -853 3623 -819 3657
rect -785 3623 -751 3657
rect -717 3623 -683 3657
rect -649 3623 -615 3657
rect -581 3623 -547 3657
rect -513 3623 -479 3657
rect -445 3623 -411 3657
rect -377 3623 -343 3657
rect -309 3623 -275 3657
rect -241 3623 -207 3657
rect -173 3623 -139 3657
rect -105 3623 -71 3657
rect -37 3623 -3 3657
rect 31 3623 65 3657
rect 99 3623 133 3657
rect 167 3623 201 3657
rect 235 3623 269 3657
rect 303 3623 337 3657
rect 371 3623 405 3657
rect 439 3623 473 3657
rect 507 3623 541 3657
rect 575 3623 609 3657
rect 643 3623 677 3657
rect 711 3623 745 3657
rect 779 3623 813 3657
rect 847 3623 881 3657
rect 915 3623 949 3657
rect 983 3623 1017 3657
rect 1051 3623 1085 3657
rect 1119 3623 1153 3657
rect 1187 3623 1221 3657
rect 1255 3623 1289 3657
rect 1323 3623 1357 3657
rect 1391 3623 1425 3657
rect 1459 3623 1493 3657
rect 1527 3623 1561 3657
rect 1595 3623 1629 3657
rect 1663 3623 1697 3657
rect 1731 3623 1765 3657
rect 1799 3623 1833 3657
rect 1867 3623 1901 3657
rect 1935 3623 1969 3657
rect 2003 3623 2037 3657
rect 2071 3623 2105 3657
rect 2139 3623 2173 3657
rect 2207 3623 2241 3657
rect 2275 3623 2309 3657
rect 2343 3623 2377 3657
rect 2411 3623 2445 3657
rect 2479 3623 2513 3657
rect 2547 3623 2581 3657
rect 2615 3623 2649 3657
rect 2683 3623 2717 3657
rect 2751 3623 2785 3657
rect 2819 3623 2853 3657
rect 2887 3623 2921 3657
rect 2955 3623 2989 3657
rect 3023 3623 3057 3657
rect 3091 3623 3125 3657
rect 3159 3623 3193 3657
rect 3227 3623 3261 3657
rect 3295 3623 3329 3657
rect 3363 3623 3397 3657
rect 3431 3623 3465 3657
rect 3499 3623 3533 3657
rect 3567 3623 3601 3657
rect 3635 3623 3669 3657
rect 3703 3623 3737 3657
rect 3771 3623 3805 3657
rect 3839 3623 3873 3657
rect 3907 3623 3941 3657
rect 3975 3623 4009 3657
rect 4043 3623 4077 3657
rect 4111 3623 4145 3657
rect 4179 3623 4213 3657
rect 4247 3623 4281 3657
rect 4315 3623 4349 3657
rect 4383 3623 4417 3657
rect 4451 3623 4485 3657
rect 4519 3623 4553 3657
rect 4587 3623 4621 3657
rect 4655 3623 4689 3657
rect 4723 3623 4757 3657
rect 4791 3623 4825 3657
rect 4859 3623 4893 3657
rect 4927 3623 4961 3657
rect 4995 3623 5029 3657
rect 5063 3623 5097 3657
rect 5131 3623 5165 3657
rect 5199 3623 5233 3657
rect 5267 3623 5301 3657
rect 5335 3623 5369 3657
rect 5403 3623 5437 3657
rect 5471 3623 5505 3657
rect 5539 3623 5573 3657
rect 5607 3623 5641 3657
rect 5675 3623 5709 3657
rect 5743 3623 5777 3657
rect 5811 3623 5845 3657
rect 5879 3623 5913 3657
rect 5947 3623 5981 3657
rect 6015 3623 6049 3657
rect 6083 3623 6117 3657
rect 6151 3623 6185 3657
rect 6219 3623 6253 3657
rect 6287 3623 6321 3657
rect 6355 3623 6389 3657
rect 6423 3623 6457 3657
rect 6491 3623 6525 3657
rect 6559 3623 6593 3657
rect 6627 3623 6661 3657
rect 6695 3623 6729 3657
rect 6763 3623 6797 3657
rect 6831 3623 6865 3657
rect 6899 3623 6933 3657
rect 6967 3623 7001 3657
rect 7035 3623 7069 3657
rect 7103 3623 7137 3657
rect 7171 3623 7205 3657
rect 7239 3623 7273 3657
rect 7307 3623 7341 3657
rect 7375 3623 7409 3657
rect 7443 3623 7477 3657
rect 7511 3623 7545 3657
rect 7579 3623 7613 3657
rect 7647 3623 7681 3657
rect 7715 3623 7749 3657
rect 7783 3623 7817 3657
rect 7851 3623 7885 3657
rect 7919 3623 7953 3657
rect 7987 3623 8021 3657
rect 8055 3623 8089 3657
rect 8123 3623 8157 3657
rect 8191 3623 8225 3657
rect 8259 3623 8293 3657
rect 8327 3623 8361 3657
rect 8395 3623 8429 3657
rect 8463 3623 8497 3657
rect 8531 3623 8565 3657
rect 8599 3623 8633 3657
rect 8667 3623 8701 3657
rect 8735 3623 8769 3657
rect 8803 3623 8837 3657
rect 8871 3623 8905 3657
rect 8939 3623 8973 3657
rect 9007 3623 9041 3657
rect 9075 3623 9109 3657
rect 9143 3623 9177 3657
rect 9211 3623 9245 3657
rect 9279 3623 9313 3657
rect 9347 3623 9381 3657
rect 9415 3623 9449 3657
rect 9483 3623 9517 3657
rect 9551 3623 9585 3657
rect 9619 3623 9653 3657
rect 9687 3623 9721 3657
rect 9755 3623 9789 3657
rect 9823 3623 9857 3657
rect 9891 3623 9925 3657
rect 9959 3623 9993 3657
rect 10027 3623 10061 3657
rect 10095 3623 10129 3657
rect 10163 3623 10197 3657
rect 10231 3623 10265 3657
rect 10299 3623 10333 3657
rect 10367 3623 10401 3657
rect 10435 3623 10469 3657
rect 10503 3623 10537 3657
rect 10571 3623 10605 3657
rect 10639 3623 10673 3657
rect 10707 3623 10741 3657
rect 10775 3623 10809 3657
rect 10843 3623 10877 3657
rect 10911 3623 10945 3657
rect 10979 3623 11013 3657
rect 11047 3623 11081 3657
rect 11115 3623 11149 3657
rect 11183 3623 11217 3657
rect 11251 3623 11285 3657
rect 11319 3623 11353 3657
rect 11387 3623 11421 3657
rect 11455 3623 11489 3657
rect 11523 3623 11557 3657
rect 11591 3623 11625 3657
rect 11659 3623 11693 3657
rect 11727 3623 11761 3657
rect 11795 3623 11829 3657
rect 11863 3623 11897 3657
rect 11931 3623 11965 3657
rect 11999 3623 12033 3657
rect 12067 3623 12101 3657
rect 12135 3623 12169 3657
rect 12203 3623 12237 3657
rect 12271 3623 12305 3657
rect 12339 3623 12373 3657
rect 12407 3623 12441 3657
rect 12475 3623 12509 3657
rect 12543 3623 12577 3657
rect 12611 3623 12645 3657
rect 12679 3623 12713 3657
rect 12747 3623 12781 3657
rect 12815 3623 12849 3657
rect 12883 3623 12917 3657
rect 12951 3623 12985 3657
rect 13019 3623 13053 3657
rect 13087 3623 13121 3657
rect 13155 3623 13189 3657
rect 13223 3623 13257 3657
rect 13291 3623 13325 3657
rect 13359 3623 13393 3657
rect 13427 3623 13461 3657
rect 13495 3623 13529 3657
rect 13563 3623 13597 3657
rect 13631 3623 13665 3657
rect 13699 3623 13733 3657
rect 13767 3623 13801 3657
rect 13835 3623 13869 3657
rect 13903 3623 13937 3657
rect 13971 3623 14005 3657
rect 14039 3623 14073 3657
rect 14107 3623 14141 3657
rect 14175 3623 14209 3657
rect 14243 3623 14277 3657
rect 14311 3623 14345 3657
rect 14379 3623 14413 3657
rect 14447 3623 14481 3657
rect 14515 3623 14549 3657
rect 14583 3623 14617 3657
rect 14651 3623 14685 3657
rect 14719 3623 14880 3657
rect -12880 3600 14880 3623
rect -12880 3489 -12800 3600
rect -12880 3455 -12857 3489
rect -12823 3455 -12800 3489
rect -12880 3421 -12800 3455
rect -12880 3387 -12857 3421
rect -12823 3387 -12800 3421
rect -12880 3353 -12800 3387
rect -12880 3319 -12857 3353
rect -12823 3319 -12800 3353
rect -12880 3285 -12800 3319
rect -12880 3251 -12857 3285
rect -12823 3251 -12800 3285
rect -12880 3217 -12800 3251
rect -12880 3183 -12857 3217
rect -12823 3183 -12800 3217
rect -12880 3149 -12800 3183
rect -12880 3115 -12857 3149
rect -12823 3115 -12800 3149
rect -12880 3081 -12800 3115
rect -12880 3047 -12857 3081
rect -12823 3047 -12800 3081
rect -12880 3013 -12800 3047
rect -12880 2979 -12857 3013
rect -12823 2979 -12800 3013
rect -12880 2945 -12800 2979
rect -12880 2911 -12857 2945
rect -12823 2911 -12800 2945
rect -12880 2877 -12800 2911
rect -12880 2843 -12857 2877
rect -12823 2843 -12800 2877
rect -12880 2809 -12800 2843
rect -12880 2775 -12857 2809
rect -12823 2775 -12800 2809
rect -12880 2741 -12800 2775
rect -12880 2707 -12857 2741
rect -12823 2707 -12800 2741
rect -12880 2673 -12800 2707
rect -12880 2639 -12857 2673
rect -12823 2639 -12800 2673
rect -12880 2605 -12800 2639
rect -12880 2571 -12857 2605
rect -12823 2571 -12800 2605
rect -12880 2537 -12800 2571
rect -12880 2503 -12857 2537
rect -12823 2503 -12800 2537
rect -12880 2469 -12800 2503
rect -12880 2435 -12857 2469
rect -12823 2435 -12800 2469
rect -12880 2401 -12800 2435
rect -12880 2367 -12857 2401
rect -12823 2367 -12800 2401
rect -12880 2333 -12800 2367
rect -12880 2299 -12857 2333
rect -12823 2299 -12800 2333
rect -12880 2265 -12800 2299
rect -12880 2231 -12857 2265
rect -12823 2231 -12800 2265
rect -12880 2197 -12800 2231
rect -12880 2163 -12857 2197
rect -12823 2163 -12800 2197
rect -12880 2129 -12800 2163
rect -12880 2095 -12857 2129
rect -12823 2095 -12800 2129
rect -12880 2061 -12800 2095
rect -12880 2027 -12857 2061
rect -12823 2027 -12800 2061
rect -12880 1993 -12800 2027
rect -12880 1959 -12857 1993
rect -12823 1959 -12800 1993
rect -12880 1925 -12800 1959
rect -12880 1891 -12857 1925
rect -12823 1891 -12800 1925
rect -12880 1857 -12800 1891
rect -12880 1823 -12857 1857
rect -12823 1823 -12800 1857
rect -12880 1789 -12800 1823
rect -12880 1755 -12857 1789
rect -12823 1755 -12800 1789
rect -12880 1721 -12800 1755
rect -12880 1687 -12857 1721
rect -12823 1687 -12800 1721
rect -12880 1653 -12800 1687
rect -12880 1619 -12857 1653
rect -12823 1619 -12800 1653
rect -12880 1585 -12800 1619
rect -12880 1551 -12857 1585
rect -12823 1551 -12800 1585
rect -12880 1440 -12800 1551
rect 14800 3489 14880 3600
rect 14800 3455 14823 3489
rect 14857 3455 14880 3489
rect 14800 3421 14880 3455
rect 14800 3387 14823 3421
rect 14857 3387 14880 3421
rect 14800 3353 14880 3387
rect 14800 3319 14823 3353
rect 14857 3319 14880 3353
rect 14800 3285 14880 3319
rect 14800 3251 14823 3285
rect 14857 3251 14880 3285
rect 14800 3217 14880 3251
rect 14800 3183 14823 3217
rect 14857 3183 14880 3217
rect 14800 3149 14880 3183
rect 14800 3115 14823 3149
rect 14857 3115 14880 3149
rect 14800 3081 14880 3115
rect 14800 3047 14823 3081
rect 14857 3047 14880 3081
rect 14800 3013 14880 3047
rect 14800 2979 14823 3013
rect 14857 2979 14880 3013
rect 14800 2945 14880 2979
rect 14800 2911 14823 2945
rect 14857 2911 14880 2945
rect 14800 2877 14880 2911
rect 14800 2843 14823 2877
rect 14857 2843 14880 2877
rect 14800 2809 14880 2843
rect 14800 2775 14823 2809
rect 14857 2775 14880 2809
rect 14800 2741 14880 2775
rect 14800 2707 14823 2741
rect 14857 2707 14880 2741
rect 14800 2673 14880 2707
rect 14800 2639 14823 2673
rect 14857 2639 14880 2673
rect 14800 2605 14880 2639
rect 14800 2571 14823 2605
rect 14857 2571 14880 2605
rect 14800 2537 14880 2571
rect 14800 2503 14823 2537
rect 14857 2503 14880 2537
rect 14800 2469 14880 2503
rect 14800 2435 14823 2469
rect 14857 2435 14880 2469
rect 14800 2401 14880 2435
rect 14800 2367 14823 2401
rect 14857 2367 14880 2401
rect 14800 2333 14880 2367
rect 14800 2299 14823 2333
rect 14857 2299 14880 2333
rect 14800 2265 14880 2299
rect 14800 2231 14823 2265
rect 14857 2231 14880 2265
rect 14800 2197 14880 2231
rect 14800 2163 14823 2197
rect 14857 2163 14880 2197
rect 14800 2129 14880 2163
rect 14800 2095 14823 2129
rect 14857 2095 14880 2129
rect 14800 2061 14880 2095
rect 14800 2027 14823 2061
rect 14857 2027 14880 2061
rect 14800 1993 14880 2027
rect 14800 1959 14823 1993
rect 14857 1959 14880 1993
rect 14800 1925 14880 1959
rect 14800 1891 14823 1925
rect 14857 1891 14880 1925
rect 14800 1857 14880 1891
rect 14800 1823 14823 1857
rect 14857 1823 14880 1857
rect 14800 1789 14880 1823
rect 14800 1755 14823 1789
rect 14857 1755 14880 1789
rect 14800 1721 14880 1755
rect 14800 1687 14823 1721
rect 14857 1687 14880 1721
rect 14800 1653 14880 1687
rect 14800 1619 14823 1653
rect 14857 1619 14880 1653
rect 14800 1585 14880 1619
rect 14800 1551 14823 1585
rect 14857 1551 14880 1585
rect 14800 1440 14880 1551
rect -12880 1417 14880 1440
rect -12880 1383 -12719 1417
rect -12685 1383 -12651 1417
rect -12617 1383 -12583 1417
rect -12549 1383 -12515 1417
rect -12481 1383 -12447 1417
rect -12413 1383 -12379 1417
rect -12345 1383 -12311 1417
rect -12277 1383 -12243 1417
rect -12209 1383 -12175 1417
rect -12141 1383 -12107 1417
rect -12073 1383 -12039 1417
rect -12005 1383 -11971 1417
rect -11937 1383 -11903 1417
rect -11869 1383 -11835 1417
rect -11801 1383 -11767 1417
rect -11733 1383 -11699 1417
rect -11665 1383 -11631 1417
rect -11597 1383 -11563 1417
rect -11529 1383 -11495 1417
rect -11461 1383 -11427 1417
rect -11393 1383 -11359 1417
rect -11325 1383 -11291 1417
rect -11257 1383 -11223 1417
rect -11189 1383 -11155 1417
rect -11121 1383 -11087 1417
rect -11053 1383 -11019 1417
rect -10985 1383 -10951 1417
rect -10917 1383 -10883 1417
rect -10849 1383 -10815 1417
rect -10781 1383 -10747 1417
rect -10713 1383 -10679 1417
rect -10645 1383 -10611 1417
rect -10577 1383 -10543 1417
rect -10509 1383 -10475 1417
rect -10441 1383 -10407 1417
rect -10373 1383 -10339 1417
rect -10305 1383 -10271 1417
rect -10237 1383 -10203 1417
rect -10169 1383 -10135 1417
rect -10101 1383 -10067 1417
rect -10033 1383 -9999 1417
rect -9965 1383 -9931 1417
rect -9897 1383 -9863 1417
rect -9829 1383 -9795 1417
rect -9761 1383 -9727 1417
rect -9693 1383 -9659 1417
rect -9625 1383 -9591 1417
rect -9557 1383 -9523 1417
rect -9489 1383 -9455 1417
rect -9421 1383 -9387 1417
rect -9353 1383 -9319 1417
rect -9285 1383 -9251 1417
rect -9217 1383 -9183 1417
rect -9149 1383 -9115 1417
rect -9081 1383 -9047 1417
rect -9013 1383 -8979 1417
rect -8945 1383 -8911 1417
rect -8877 1383 -8843 1417
rect -8809 1383 -8775 1417
rect -8741 1383 -8707 1417
rect -8673 1383 -8639 1417
rect -8605 1383 -8571 1417
rect -8537 1383 -8503 1417
rect -8469 1383 -8435 1417
rect -8401 1383 -8367 1417
rect -8333 1383 -8299 1417
rect -8265 1383 -8231 1417
rect -8197 1383 -8163 1417
rect -8129 1383 -8095 1417
rect -8061 1383 -8027 1417
rect -7993 1383 -7959 1417
rect -7925 1383 -7891 1417
rect -7857 1383 -7823 1417
rect -7789 1383 -7755 1417
rect -7721 1383 -7687 1417
rect -7653 1383 -7619 1417
rect -7585 1383 -7551 1417
rect -7517 1383 -7483 1417
rect -7449 1383 -7415 1417
rect -7381 1383 -7347 1417
rect -7313 1383 -7279 1417
rect -7245 1383 -7211 1417
rect -7177 1383 -7143 1417
rect -7109 1383 -7075 1417
rect -7041 1383 -7007 1417
rect -6973 1383 -6939 1417
rect -6905 1383 -6871 1417
rect -6837 1383 -6803 1417
rect -6769 1383 -6735 1417
rect -6701 1383 -6667 1417
rect -6633 1383 -6599 1417
rect -6565 1383 -6531 1417
rect -6497 1383 -6463 1417
rect -6429 1383 -6395 1417
rect -6361 1383 -6327 1417
rect -6293 1383 -6259 1417
rect -6225 1383 -6191 1417
rect -6157 1383 -6123 1417
rect -6089 1383 -6055 1417
rect -6021 1383 -5987 1417
rect -5953 1383 -5919 1417
rect -5885 1383 -5851 1417
rect -5817 1383 -5783 1417
rect -5749 1383 -5715 1417
rect -5681 1383 -5647 1417
rect -5613 1383 -5579 1417
rect -5545 1383 -5511 1417
rect -5477 1383 -5443 1417
rect -5409 1383 -5375 1417
rect -5341 1383 -5307 1417
rect -5273 1383 -5239 1417
rect -5205 1383 -5171 1417
rect -5137 1383 -5103 1417
rect -5069 1383 -5035 1417
rect -5001 1383 -4967 1417
rect -4933 1383 -4899 1417
rect -4865 1383 -4831 1417
rect -4797 1383 -4763 1417
rect -4729 1383 -4695 1417
rect -4661 1383 -4627 1417
rect -4593 1383 -4559 1417
rect -4525 1383 -4491 1417
rect -4457 1383 -4423 1417
rect -4389 1383 -4355 1417
rect -4321 1383 -4287 1417
rect -4253 1383 -4219 1417
rect -4185 1383 -4151 1417
rect -4117 1383 -4083 1417
rect -4049 1383 -4015 1417
rect -3981 1383 -3947 1417
rect -3913 1383 -3879 1417
rect -3845 1383 -3811 1417
rect -3777 1383 -3743 1417
rect -3709 1383 -3675 1417
rect -3641 1383 -3607 1417
rect -3573 1383 -3539 1417
rect -3505 1383 -3471 1417
rect -3437 1383 -3403 1417
rect -3369 1383 -3335 1417
rect -3301 1383 -3267 1417
rect -3233 1383 -3199 1417
rect -3165 1383 -3131 1417
rect -3097 1383 -3063 1417
rect -3029 1383 -2995 1417
rect -2961 1383 -2927 1417
rect -2893 1383 -2859 1417
rect -2825 1383 -2791 1417
rect -2757 1383 -2723 1417
rect -2689 1383 -2655 1417
rect -2621 1383 -2587 1417
rect -2553 1383 -2519 1417
rect -2485 1383 -2451 1417
rect -2417 1383 -2383 1417
rect -2349 1383 -2315 1417
rect -2281 1383 -2247 1417
rect -2213 1383 -2179 1417
rect -2145 1383 -2111 1417
rect -2077 1383 -2043 1417
rect -2009 1383 -1975 1417
rect -1941 1383 -1907 1417
rect -1873 1383 -1839 1417
rect -1805 1383 -1771 1417
rect -1737 1383 -1703 1417
rect -1669 1383 -1635 1417
rect -1601 1383 -1567 1417
rect -1533 1383 -1499 1417
rect -1465 1383 -1431 1417
rect -1397 1383 -1363 1417
rect -1329 1383 -1295 1417
rect -1261 1383 -1227 1417
rect -1193 1383 -1159 1417
rect -1125 1383 -1091 1417
rect -1057 1383 -1023 1417
rect -989 1383 -955 1417
rect -921 1383 -887 1417
rect -853 1383 -819 1417
rect -785 1383 -751 1417
rect -717 1383 -683 1417
rect -649 1383 -615 1417
rect -581 1383 -547 1417
rect -513 1383 -479 1417
rect -445 1383 -411 1417
rect -377 1383 -343 1417
rect -309 1383 -275 1417
rect -241 1383 -207 1417
rect -173 1383 -139 1417
rect -105 1383 -71 1417
rect -37 1383 -3 1417
rect 31 1383 65 1417
rect 99 1383 133 1417
rect 167 1383 201 1417
rect 235 1383 269 1417
rect 303 1383 337 1417
rect 371 1383 405 1417
rect 439 1383 473 1417
rect 507 1383 541 1417
rect 575 1383 609 1417
rect 643 1383 677 1417
rect 711 1383 745 1417
rect 779 1383 813 1417
rect 847 1383 881 1417
rect 915 1383 949 1417
rect 983 1383 1017 1417
rect 1051 1383 1085 1417
rect 1119 1383 1153 1417
rect 1187 1383 1221 1417
rect 1255 1383 1289 1417
rect 1323 1383 1357 1417
rect 1391 1383 1425 1417
rect 1459 1383 1493 1417
rect 1527 1383 1561 1417
rect 1595 1383 1629 1417
rect 1663 1383 1697 1417
rect 1731 1383 1765 1417
rect 1799 1383 1833 1417
rect 1867 1383 1901 1417
rect 1935 1383 1969 1417
rect 2003 1383 2037 1417
rect 2071 1383 2105 1417
rect 2139 1383 2173 1417
rect 2207 1383 2241 1417
rect 2275 1383 2309 1417
rect 2343 1383 2377 1417
rect 2411 1383 2445 1417
rect 2479 1383 2513 1417
rect 2547 1383 2581 1417
rect 2615 1383 2649 1417
rect 2683 1383 2717 1417
rect 2751 1383 2785 1417
rect 2819 1383 2853 1417
rect 2887 1383 2921 1417
rect 2955 1383 2989 1417
rect 3023 1383 3057 1417
rect 3091 1383 3125 1417
rect 3159 1383 3193 1417
rect 3227 1383 3261 1417
rect 3295 1383 3329 1417
rect 3363 1383 3397 1417
rect 3431 1383 3465 1417
rect 3499 1383 3533 1417
rect 3567 1383 3601 1417
rect 3635 1383 3669 1417
rect 3703 1383 3737 1417
rect 3771 1383 3805 1417
rect 3839 1383 3873 1417
rect 3907 1383 3941 1417
rect 3975 1383 4009 1417
rect 4043 1383 4077 1417
rect 4111 1383 4145 1417
rect 4179 1383 4213 1417
rect 4247 1383 4281 1417
rect 4315 1383 4349 1417
rect 4383 1383 4417 1417
rect 4451 1383 4485 1417
rect 4519 1383 4553 1417
rect 4587 1383 4621 1417
rect 4655 1383 4689 1417
rect 4723 1383 4757 1417
rect 4791 1383 4825 1417
rect 4859 1383 4893 1417
rect 4927 1383 4961 1417
rect 4995 1383 5029 1417
rect 5063 1383 5097 1417
rect 5131 1383 5165 1417
rect 5199 1383 5233 1417
rect 5267 1383 5301 1417
rect 5335 1383 5369 1417
rect 5403 1383 5437 1417
rect 5471 1383 5505 1417
rect 5539 1383 5573 1417
rect 5607 1383 5641 1417
rect 5675 1383 5709 1417
rect 5743 1383 5777 1417
rect 5811 1383 5845 1417
rect 5879 1383 5913 1417
rect 5947 1383 5981 1417
rect 6015 1383 6049 1417
rect 6083 1383 6117 1417
rect 6151 1383 6185 1417
rect 6219 1383 6253 1417
rect 6287 1383 6321 1417
rect 6355 1383 6389 1417
rect 6423 1383 6457 1417
rect 6491 1383 6525 1417
rect 6559 1383 6593 1417
rect 6627 1383 6661 1417
rect 6695 1383 6729 1417
rect 6763 1383 6797 1417
rect 6831 1383 6865 1417
rect 6899 1383 6933 1417
rect 6967 1383 7001 1417
rect 7035 1383 7069 1417
rect 7103 1383 7137 1417
rect 7171 1383 7205 1417
rect 7239 1383 7273 1417
rect 7307 1383 7341 1417
rect 7375 1383 7409 1417
rect 7443 1383 7477 1417
rect 7511 1383 7545 1417
rect 7579 1383 7613 1417
rect 7647 1383 7681 1417
rect 7715 1383 7749 1417
rect 7783 1383 7817 1417
rect 7851 1383 7885 1417
rect 7919 1383 7953 1417
rect 7987 1383 8021 1417
rect 8055 1383 8089 1417
rect 8123 1383 8157 1417
rect 8191 1383 8225 1417
rect 8259 1383 8293 1417
rect 8327 1383 8361 1417
rect 8395 1383 8429 1417
rect 8463 1383 8497 1417
rect 8531 1383 8565 1417
rect 8599 1383 8633 1417
rect 8667 1383 8701 1417
rect 8735 1383 8769 1417
rect 8803 1383 8837 1417
rect 8871 1383 8905 1417
rect 8939 1383 8973 1417
rect 9007 1383 9041 1417
rect 9075 1383 9109 1417
rect 9143 1383 9177 1417
rect 9211 1383 9245 1417
rect 9279 1383 9313 1417
rect 9347 1383 9381 1417
rect 9415 1383 9449 1417
rect 9483 1383 9517 1417
rect 9551 1383 9585 1417
rect 9619 1383 9653 1417
rect 9687 1383 9721 1417
rect 9755 1383 9789 1417
rect 9823 1383 9857 1417
rect 9891 1383 9925 1417
rect 9959 1383 9993 1417
rect 10027 1383 10061 1417
rect 10095 1383 10129 1417
rect 10163 1383 10197 1417
rect 10231 1383 10265 1417
rect 10299 1383 10333 1417
rect 10367 1383 10401 1417
rect 10435 1383 10469 1417
rect 10503 1383 10537 1417
rect 10571 1383 10605 1417
rect 10639 1383 10673 1417
rect 10707 1383 10741 1417
rect 10775 1383 10809 1417
rect 10843 1383 10877 1417
rect 10911 1383 10945 1417
rect 10979 1383 11013 1417
rect 11047 1383 11081 1417
rect 11115 1383 11149 1417
rect 11183 1383 11217 1417
rect 11251 1383 11285 1417
rect 11319 1383 11353 1417
rect 11387 1383 11421 1417
rect 11455 1383 11489 1417
rect 11523 1383 11557 1417
rect 11591 1383 11625 1417
rect 11659 1383 11693 1417
rect 11727 1383 11761 1417
rect 11795 1383 11829 1417
rect 11863 1383 11897 1417
rect 11931 1383 11965 1417
rect 11999 1383 12033 1417
rect 12067 1383 12101 1417
rect 12135 1383 12169 1417
rect 12203 1383 12237 1417
rect 12271 1383 12305 1417
rect 12339 1383 12373 1417
rect 12407 1383 12441 1417
rect 12475 1383 12509 1417
rect 12543 1383 12577 1417
rect 12611 1383 12645 1417
rect 12679 1383 12713 1417
rect 12747 1383 12781 1417
rect 12815 1383 12849 1417
rect 12883 1383 12917 1417
rect 12951 1383 12985 1417
rect 13019 1383 13053 1417
rect 13087 1383 13121 1417
rect 13155 1383 13189 1417
rect 13223 1383 13257 1417
rect 13291 1383 13325 1417
rect 13359 1383 13393 1417
rect 13427 1383 13461 1417
rect 13495 1383 13529 1417
rect 13563 1383 13597 1417
rect 13631 1383 13665 1417
rect 13699 1383 13733 1417
rect 13767 1383 13801 1417
rect 13835 1383 13869 1417
rect 13903 1383 13937 1417
rect 13971 1383 14005 1417
rect 14039 1383 14073 1417
rect 14107 1383 14141 1417
rect 14175 1383 14209 1417
rect 14243 1383 14277 1417
rect 14311 1383 14345 1417
rect 14379 1383 14413 1417
rect 14447 1383 14481 1417
rect 14515 1383 14549 1417
rect 14583 1383 14617 1417
rect 14651 1383 14685 1417
rect 14719 1383 14880 1417
rect -12880 1360 14880 1383
<< metal3 >>
rect -12720 3512 -12640 3520
rect -12720 3448 -12712 3512
rect -12648 3448 -12640 3512
rect -12720 3192 -12640 3448
rect -12720 3128 -12712 3192
rect -12648 3128 -12640 3192
rect -12720 2872 -12640 3128
rect -12720 2808 -12712 2872
rect -12648 2808 -12640 2872
rect -12720 2720 -12640 2808
rect -12560 3512 -12480 3520
rect -12560 3448 -12552 3512
rect -12488 3448 -12480 3512
rect -12560 3192 -12480 3448
rect -12560 3128 -12552 3192
rect -12488 3128 -12480 3192
rect -12560 2872 -12480 3128
rect -12560 2808 -12552 2872
rect -12488 2808 -12480 2872
rect -12560 2720 -12480 2808
rect -12400 3512 -12320 3520
rect -12400 3448 -12392 3512
rect -12328 3448 -12320 3512
rect -12400 3192 -12320 3448
rect 14320 3512 14400 3520
rect 14320 3448 14328 3512
rect 14392 3448 14400 3512
rect -12400 3128 -12392 3192
rect -12328 3128 -12320 3192
rect -12400 2872 -12320 3128
rect -11040 3352 -10960 3360
rect -11040 3288 -11032 3352
rect -10968 3288 -10960 3352
rect -12400 2808 -12392 2872
rect -12328 2808 -12320 2872
rect -12400 2720 -12320 2808
rect -12720 2320 -12320 2720
rect -12720 2232 -12640 2320
rect -12720 2168 -12712 2232
rect -12648 2168 -12640 2232
rect -12720 1912 -12640 2168
rect -12720 1848 -12712 1912
rect -12648 1848 -12640 1912
rect -12720 1592 -12640 1848
rect -12720 1528 -12712 1592
rect -12648 1528 -12640 1592
rect -12720 1520 -12640 1528
rect -12560 2232 -12480 2320
rect -12560 2168 -12552 2232
rect -12488 2168 -12480 2232
rect -12560 1912 -12480 2168
rect -12560 1848 -12552 1912
rect -12488 1848 -12480 1912
rect -12560 1592 -12480 1848
rect -12560 1528 -12552 1592
rect -12488 1528 -12480 1592
rect -12560 1520 -12480 1528
rect -12400 2232 -12320 2320
rect -12400 2168 -12392 2232
rect -12328 2168 -12320 2232
rect -12400 1912 -12320 2168
rect -12240 2872 -12160 2880
rect -12240 2808 -12232 2872
rect -12168 2808 -12160 2872
rect -12240 2232 -12160 2808
rect -11040 2720 -10960 3288
rect -8640 3352 -8560 3360
rect -8640 3288 -8632 3352
rect -8568 3288 -8560 3352
rect -9840 2872 -9760 2880
rect -9840 2808 -9832 2872
rect -9768 2808 -9760 2872
rect -12080 2320 -9920 2720
rect -12240 2168 -12232 2232
rect -12168 2168 -12160 2232
rect -12240 2160 -12160 2168
rect -12400 1848 -12392 1912
rect -12328 1848 -12320 1912
rect -12400 1592 -12320 1848
rect -11040 1752 -10960 2320
rect -9840 2232 -9760 2808
rect -8640 2720 -8560 3288
rect -6240 3352 -6160 3360
rect -6240 3288 -6232 3352
rect -6168 3288 -6160 3352
rect -7440 2872 -7360 2880
rect -7440 2808 -7432 2872
rect -7368 2808 -7360 2872
rect -9680 2320 -7520 2720
rect -9840 2168 -9832 2232
rect -9768 2168 -9760 2232
rect -9840 2160 -9760 2168
rect -11040 1688 -11032 1752
rect -10968 1688 -10960 1752
rect -11040 1680 -10960 1688
rect -8640 1752 -8560 2320
rect -7440 2232 -7360 2808
rect -6240 2720 -6160 3288
rect -3840 3352 -3760 3360
rect -3840 3288 -3832 3352
rect -3768 3288 -3760 3352
rect -5040 2872 -4960 2880
rect -5040 2808 -5032 2872
rect -4968 2808 -4960 2872
rect -7280 2320 -5120 2720
rect -7440 2168 -7432 2232
rect -7368 2168 -7360 2232
rect -7440 2160 -7360 2168
rect -8640 1688 -8632 1752
rect -8568 1688 -8560 1752
rect -8640 1680 -8560 1688
rect -6240 1752 -6160 2320
rect -5040 2232 -4960 2808
rect -3840 2720 -3760 3288
rect -1440 3352 -1360 3360
rect -1440 3288 -1432 3352
rect -1368 3288 -1360 3352
rect -2640 2872 -2560 2880
rect -2640 2808 -2632 2872
rect -2568 2808 -2560 2872
rect -4880 2320 -2720 2720
rect -5040 2168 -5032 2232
rect -4968 2168 -4960 2232
rect -5040 2160 -4960 2168
rect -6240 1688 -6232 1752
rect -6168 1688 -6160 1752
rect -6240 1680 -6160 1688
rect -3840 1752 -3760 2320
rect -2640 2232 -2560 2808
rect -1440 2720 -1360 3288
rect 3360 3352 3440 3360
rect 3360 3288 3368 3352
rect 3432 3288 3440 3352
rect 960 3032 1040 3040
rect 960 2968 968 3032
rect 1032 2968 1040 3032
rect -240 2872 -160 2880
rect -240 2808 -232 2872
rect -168 2808 -160 2872
rect -2480 2320 -320 2720
rect -2640 2168 -2632 2232
rect -2568 2168 -2560 2232
rect -2640 2160 -2560 2168
rect -3840 1688 -3832 1752
rect -3768 1688 -3760 1752
rect -3840 1680 -3760 1688
rect -1440 1752 -1360 2320
rect -240 2232 -160 2808
rect 960 2720 1040 2968
rect 2160 2872 2240 2880
rect 2160 2808 2168 2872
rect 2232 2808 2240 2872
rect -80 2320 2080 2720
rect -240 2168 -232 2232
rect -168 2168 -160 2232
rect -240 2160 -160 2168
rect 960 2072 1040 2320
rect 2160 2232 2240 2808
rect 3360 2720 3440 3288
rect 5760 3352 5840 3360
rect 5760 3288 5768 3352
rect 5832 3288 5840 3352
rect 4560 2872 4640 2880
rect 4560 2808 4568 2872
rect 4632 2808 4640 2872
rect 2320 2320 4480 2720
rect 2160 2168 2168 2232
rect 2232 2168 2240 2232
rect 2160 2160 2240 2168
rect 960 2008 968 2072
rect 1032 2008 1040 2072
rect 960 2000 1040 2008
rect -1440 1688 -1432 1752
rect -1368 1688 -1360 1752
rect -1440 1680 -1360 1688
rect 3360 1752 3440 2320
rect 4560 2232 4640 2808
rect 5760 2720 5840 3288
rect 8160 3352 8240 3360
rect 8160 3288 8168 3352
rect 8232 3288 8240 3352
rect 6960 2872 7040 2880
rect 6960 2808 6968 2872
rect 7032 2808 7040 2872
rect 4720 2320 6880 2720
rect 4560 2168 4568 2232
rect 4632 2168 4640 2232
rect 4560 2160 4640 2168
rect 3360 1688 3368 1752
rect 3432 1688 3440 1752
rect 3360 1680 3440 1688
rect 5760 1752 5840 2320
rect 6960 2232 7040 2808
rect 8160 2720 8240 3288
rect 10560 3352 10640 3360
rect 10560 3288 10568 3352
rect 10632 3288 10640 3352
rect 9360 2872 9440 2880
rect 9360 2808 9368 2872
rect 9432 2808 9440 2872
rect 7120 2320 9280 2720
rect 6960 2168 6968 2232
rect 7032 2168 7040 2232
rect 6960 2160 7040 2168
rect 5760 1688 5768 1752
rect 5832 1688 5840 1752
rect 5760 1680 5840 1688
rect 8160 1752 8240 2320
rect 9360 2232 9440 2808
rect 10560 2720 10640 3288
rect 12960 3352 13040 3360
rect 12960 3288 12968 3352
rect 13032 3288 13040 3352
rect 11760 2872 11840 2880
rect 11760 2808 11768 2872
rect 11832 2808 11840 2872
rect 9520 2320 11680 2720
rect 9360 2168 9368 2232
rect 9432 2168 9440 2232
rect 9360 2160 9440 2168
rect 8160 1688 8168 1752
rect 8232 1688 8240 1752
rect 8160 1680 8240 1688
rect 10560 1752 10640 2320
rect 11760 2232 11840 2808
rect 12960 2720 13040 3288
rect 14320 3352 14400 3448
rect 14320 3288 14328 3352
rect 14392 3288 14400 3352
rect 14320 3192 14400 3288
rect 14320 3128 14328 3192
rect 14392 3128 14400 3192
rect 14320 3032 14400 3128
rect 14320 2968 14328 3032
rect 14392 2968 14400 3032
rect 14160 2872 14240 2880
rect 14160 2808 14168 2872
rect 14232 2808 14240 2872
rect 11920 2320 14080 2720
rect 11760 2168 11768 2232
rect 11832 2168 11840 2232
rect 11760 2160 11840 2168
rect 10560 1688 10568 1752
rect 10632 1688 10640 1752
rect 10560 1680 10640 1688
rect 12960 1752 13040 2320
rect 14160 2232 14240 2808
rect 14160 2168 14168 2232
rect 14232 2168 14240 2232
rect 14160 2160 14240 2168
rect 14320 2872 14400 2968
rect 14320 2808 14328 2872
rect 14392 2808 14400 2872
rect 14320 2720 14400 2808
rect 14480 3512 14560 3520
rect 14480 3448 14488 3512
rect 14552 3448 14560 3512
rect 14480 3352 14560 3448
rect 14480 3288 14488 3352
rect 14552 3288 14560 3352
rect 14480 3192 14560 3288
rect 14480 3128 14488 3192
rect 14552 3128 14560 3192
rect 14480 3032 14560 3128
rect 14480 2968 14488 3032
rect 14552 2968 14560 3032
rect 14480 2872 14560 2968
rect 14480 2808 14488 2872
rect 14552 2808 14560 2872
rect 14480 2720 14560 2808
rect 14640 3512 14720 3520
rect 14640 3448 14648 3512
rect 14712 3448 14720 3512
rect 14640 3352 14720 3448
rect 14640 3288 14648 3352
rect 14712 3288 14720 3352
rect 14640 3192 14720 3288
rect 14640 3128 14648 3192
rect 14712 3128 14720 3192
rect 14640 3032 14720 3128
rect 14640 2968 14648 3032
rect 14712 2968 14720 3032
rect 14640 2872 14720 2968
rect 14640 2808 14648 2872
rect 14712 2808 14720 2872
rect 14640 2720 14720 2808
rect 14320 2320 14720 2720
rect 14320 2232 14400 2320
rect 14320 2168 14328 2232
rect 14392 2168 14400 2232
rect 12960 1688 12968 1752
rect 13032 1688 13040 1752
rect 12960 1680 13040 1688
rect 14320 2072 14400 2168
rect 14320 2008 14328 2072
rect 14392 2008 14400 2072
rect 14320 1912 14400 2008
rect 14320 1848 14328 1912
rect 14392 1848 14400 1912
rect 14320 1752 14400 1848
rect 14320 1688 14328 1752
rect 14392 1688 14400 1752
rect -12400 1528 -12392 1592
rect -12328 1528 -12320 1592
rect -12400 1520 -12320 1528
rect 14320 1592 14400 1688
rect 14320 1528 14328 1592
rect 14392 1528 14400 1592
rect 14320 1520 14400 1528
rect 14480 2232 14560 2320
rect 14480 2168 14488 2232
rect 14552 2168 14560 2232
rect 14480 2072 14560 2168
rect 14480 2008 14488 2072
rect 14552 2008 14560 2072
rect 14480 1912 14560 2008
rect 14480 1848 14488 1912
rect 14552 1848 14560 1912
rect 14480 1752 14560 1848
rect 14480 1688 14488 1752
rect 14552 1688 14560 1752
rect 14480 1592 14560 1688
rect 14480 1528 14488 1592
rect 14552 1528 14560 1592
rect 14480 1520 14560 1528
rect 14640 2232 14720 2320
rect 14640 2168 14648 2232
rect 14712 2168 14720 2232
rect 14640 2072 14720 2168
rect 14640 2008 14648 2072
rect 14712 2008 14720 2072
rect 14640 1912 14720 2008
rect 14640 1848 14648 1912
rect 14712 1848 14720 1912
rect 14640 1752 14720 1848
rect 14640 1688 14648 1752
rect 14712 1688 14720 1752
rect 14640 1592 14720 1688
rect 14640 1528 14648 1592
rect 14712 1528 14720 1592
rect 14640 1520 14720 1528
<< via3 >>
rect -12712 3448 -12648 3512
rect -12712 3128 -12648 3192
rect -12712 2808 -12648 2872
rect -12552 3448 -12488 3512
rect -12552 3128 -12488 3192
rect -12552 2808 -12488 2872
rect -12392 3448 -12328 3512
rect 14328 3448 14392 3512
rect -12392 3128 -12328 3192
rect -11032 3288 -10968 3352
rect -12392 2808 -12328 2872
rect -12712 2168 -12648 2232
rect -12712 1848 -12648 1912
rect -12712 1528 -12648 1592
rect -12552 2168 -12488 2232
rect -12552 1848 -12488 1912
rect -12552 1528 -12488 1592
rect -12392 2168 -12328 2232
rect -12232 2808 -12168 2872
rect -8632 3288 -8568 3352
rect -9832 2808 -9768 2872
rect -12232 2168 -12168 2232
rect -12392 1848 -12328 1912
rect -6232 3288 -6168 3352
rect -7432 2808 -7368 2872
rect -9832 2168 -9768 2232
rect -11032 1688 -10968 1752
rect -3832 3288 -3768 3352
rect -5032 2808 -4968 2872
rect -7432 2168 -7368 2232
rect -8632 1688 -8568 1752
rect -1432 3288 -1368 3352
rect -2632 2808 -2568 2872
rect -5032 2168 -4968 2232
rect -6232 1688 -6168 1752
rect 3368 3288 3432 3352
rect 968 2968 1032 3032
rect -232 2808 -168 2872
rect -2632 2168 -2568 2232
rect -3832 1688 -3768 1752
rect 2168 2808 2232 2872
rect -232 2168 -168 2232
rect 5768 3288 5832 3352
rect 4568 2808 4632 2872
rect 2168 2168 2232 2232
rect 968 2008 1032 2072
rect -1432 1688 -1368 1752
rect 8168 3288 8232 3352
rect 6968 2808 7032 2872
rect 4568 2168 4632 2232
rect 3368 1688 3432 1752
rect 10568 3288 10632 3352
rect 9368 2808 9432 2872
rect 6968 2168 7032 2232
rect 5768 1688 5832 1752
rect 12968 3288 13032 3352
rect 11768 2808 11832 2872
rect 9368 2168 9432 2232
rect 8168 1688 8232 1752
rect 14328 3288 14392 3352
rect 14328 3128 14392 3192
rect 14328 2968 14392 3032
rect 14168 2808 14232 2872
rect 11768 2168 11832 2232
rect 10568 1688 10632 1752
rect 14168 2168 14232 2232
rect 14328 2808 14392 2872
rect 14488 3448 14552 3512
rect 14488 3288 14552 3352
rect 14488 3128 14552 3192
rect 14488 2968 14552 3032
rect 14488 2808 14552 2872
rect 14648 3448 14712 3512
rect 14648 3288 14712 3352
rect 14648 3128 14712 3192
rect 14648 2968 14712 3032
rect 14648 2808 14712 2872
rect 14328 2168 14392 2232
rect 12968 1688 13032 1752
rect 14328 2008 14392 2072
rect 14328 1848 14392 1912
rect 14328 1688 14392 1752
rect -12392 1528 -12328 1592
rect 14328 1528 14392 1592
rect 14488 2168 14552 2232
rect 14488 2008 14552 2072
rect 14488 1848 14552 1912
rect 14488 1688 14552 1752
rect 14488 1528 14552 1592
rect 14648 2168 14712 2232
rect 14648 2008 14712 2072
rect 14648 1848 14712 1912
rect 14648 1688 14712 1752
rect 14648 1528 14712 1592
<< mimcap >>
rect -12640 2552 -12400 2640
rect -12640 2488 -12552 2552
rect -12488 2488 -12400 2552
rect -12640 2400 -12400 2488
rect -12000 2552 -10000 2640
rect -12000 2488 -11912 2552
rect -10088 2488 -10000 2552
rect -12000 2400 -10000 2488
rect -9600 2552 -7600 2640
rect -9600 2488 -9512 2552
rect -7688 2488 -7600 2552
rect -9600 2400 -7600 2488
rect -7200 2552 -5200 2640
rect -7200 2488 -7112 2552
rect -5288 2488 -5200 2552
rect -7200 2400 -5200 2488
rect -4800 2552 -2800 2640
rect -4800 2488 -4712 2552
rect -2888 2488 -2800 2552
rect -4800 2400 -2800 2488
rect -2400 2552 -400 2640
rect -2400 2488 -2312 2552
rect -488 2488 -400 2552
rect -2400 2400 -400 2488
rect 0 2552 2000 2640
rect 0 2488 88 2552
rect 1912 2488 2000 2552
rect 0 2400 2000 2488
rect 2400 2552 4400 2640
rect 2400 2488 2488 2552
rect 4312 2488 4400 2552
rect 2400 2400 4400 2488
rect 4800 2552 6800 2640
rect 4800 2488 4888 2552
rect 6712 2488 6800 2552
rect 4800 2400 6800 2488
rect 7200 2552 9200 2640
rect 7200 2488 7288 2552
rect 9112 2488 9200 2552
rect 7200 2400 9200 2488
rect 9600 2552 11600 2640
rect 9600 2488 9688 2552
rect 11512 2488 11600 2552
rect 9600 2400 11600 2488
rect 12000 2552 14000 2640
rect 12000 2488 12088 2552
rect 13912 2488 14000 2552
rect 12000 2400 14000 2488
rect 14400 2552 14640 2640
rect 14400 2488 14488 2552
rect 14552 2488 14640 2552
rect 14400 2400 14640 2488
<< mimcapcontact >>
rect -12552 2488 -12488 2552
rect -11912 2488 -10088 2552
rect -9512 2488 -7688 2552
rect -7112 2488 -5288 2552
rect -4712 2488 -2888 2552
rect -2312 2488 -488 2552
rect 88 2488 1912 2552
rect 2488 2488 4312 2552
rect 4888 2488 6712 2552
rect 7288 2488 9112 2552
rect 9688 2488 11512 2552
rect 12088 2488 13912 2552
rect 14488 2488 14552 2552
<< metal4 >>
rect -12720 3512 14880 3520
rect -12720 3448 -12712 3512
rect -12648 3448 -12552 3512
rect -12488 3448 -12392 3512
rect -12328 3448 14328 3512
rect 14392 3448 14488 3512
rect 14552 3448 14648 3512
rect 14712 3448 14880 3512
rect -12720 3440 14880 3448
rect -12720 3352 14880 3360
rect -12720 3288 -11032 3352
rect -10968 3288 -8632 3352
rect -8568 3288 -6232 3352
rect -6168 3288 -3832 3352
rect -3768 3288 -1432 3352
rect -1368 3288 3368 3352
rect 3432 3288 5768 3352
rect 5832 3288 8168 3352
rect 8232 3288 10568 3352
rect 10632 3288 12968 3352
rect 13032 3288 14328 3352
rect 14392 3288 14488 3352
rect 14552 3288 14648 3352
rect 14712 3288 14880 3352
rect -12720 3280 14880 3288
rect -11040 3200 -10960 3280
rect -8640 3200 -8560 3280
rect -6240 3200 -6160 3280
rect -3840 3200 -3760 3280
rect -1440 3200 -1360 3280
rect 3360 3200 3440 3280
rect 5760 3200 5840 3280
rect 8160 3200 8240 3280
rect 10560 3200 10640 3280
rect 12960 3200 13040 3280
rect -12720 3192 14880 3200
rect -12720 3128 -12712 3192
rect -12648 3128 -12552 3192
rect -12488 3128 -12392 3192
rect -12328 3128 14328 3192
rect 14392 3128 14488 3192
rect 14552 3128 14648 3192
rect 14712 3128 14880 3192
rect -12720 3120 14880 3128
rect -11040 3040 -10960 3120
rect -8640 3040 -8560 3120
rect -6240 3040 -6160 3120
rect -3840 3040 -3760 3120
rect -1440 3040 -1360 3120
rect 3360 3040 3440 3120
rect 5760 3040 5840 3120
rect 8160 3040 8240 3120
rect 10560 3040 10640 3120
rect 12960 3040 13040 3120
rect -12720 3032 14880 3040
rect -12720 2968 968 3032
rect 1032 2968 14328 3032
rect 14392 2968 14488 3032
rect 14552 2968 14648 3032
rect 14712 2968 14880 3032
rect -12720 2960 14880 2968
rect -11040 2880 -10960 2960
rect -8640 2880 -8560 2960
rect -6240 2880 -6160 2960
rect -3840 2880 -3760 2960
rect -1440 2880 -1360 2960
rect 960 2880 1040 2960
rect 3360 2880 3440 2960
rect 5760 2880 5840 2960
rect 8160 2880 8240 2960
rect 10560 2880 10640 2960
rect 12960 2880 13040 2960
rect -12720 2872 14880 2880
rect -12720 2808 -12712 2872
rect -12648 2808 -12552 2872
rect -12488 2808 -12392 2872
rect -12328 2808 -12232 2872
rect -12168 2808 -9832 2872
rect -9768 2808 -7432 2872
rect -7368 2808 -5032 2872
rect -4968 2808 -2632 2872
rect -2568 2808 -232 2872
rect -168 2808 2168 2872
rect 2232 2808 4568 2872
rect 4632 2808 6968 2872
rect 7032 2808 9368 2872
rect 9432 2808 11768 2872
rect 11832 2808 14168 2872
rect 14232 2808 14328 2872
rect 14392 2808 14488 2872
rect 14552 2808 14648 2872
rect 14712 2808 14880 2872
rect -12720 2800 14880 2808
rect -12720 2720 -12640 2800
rect -12560 2720 -12480 2800
rect -12400 2720 -12320 2800
rect -12720 2552 -12320 2720
rect -12720 2488 -12552 2552
rect -12488 2488 -12320 2552
rect -12720 2320 -12320 2488
rect -12720 2240 -12640 2320
rect -12560 2240 -12480 2320
rect -12400 2240 -12320 2320
rect -12240 2240 -12160 2800
rect -11040 2720 -10960 2800
rect -12080 2552 -9920 2720
rect -12080 2488 -11912 2552
rect -10088 2488 -9920 2552
rect -12080 2320 -9920 2488
rect -11040 2240 -10960 2320
rect -9840 2240 -9760 2800
rect -8640 2720 -8560 2800
rect -9680 2552 -7520 2720
rect -9680 2488 -9512 2552
rect -7688 2488 -7520 2552
rect -9680 2320 -7520 2488
rect -8640 2240 -8560 2320
rect -7440 2240 -7360 2800
rect -6240 2720 -6160 2800
rect -7280 2552 -5120 2720
rect -7280 2488 -7112 2552
rect -5288 2488 -5120 2552
rect -7280 2320 -5120 2488
rect -6240 2240 -6160 2320
rect -5040 2240 -4960 2800
rect -3840 2720 -3760 2800
rect -4880 2552 -2720 2720
rect -4880 2488 -4712 2552
rect -2888 2488 -2720 2552
rect -4880 2320 -2720 2488
rect -3840 2240 -3760 2320
rect -2640 2240 -2560 2800
rect -1440 2720 -1360 2800
rect -2480 2552 -320 2720
rect -2480 2488 -2312 2552
rect -488 2488 -320 2552
rect -2480 2320 -320 2488
rect -1440 2240 -1360 2320
rect -240 2240 -160 2800
rect 960 2720 1040 2800
rect -80 2552 2080 2720
rect -80 2488 88 2552
rect 1912 2488 2080 2552
rect -80 2320 2080 2488
rect 960 2240 1040 2320
rect 2160 2240 2240 2800
rect 3360 2720 3440 2800
rect 2320 2552 4480 2720
rect 2320 2488 2488 2552
rect 4312 2488 4480 2552
rect 2320 2320 4480 2488
rect 3360 2240 3440 2320
rect 4560 2240 4640 2800
rect 5760 2720 5840 2800
rect 4720 2552 6880 2720
rect 4720 2488 4888 2552
rect 6712 2488 6880 2552
rect 4720 2320 6880 2488
rect 5760 2240 5840 2320
rect 6960 2240 7040 2800
rect 8160 2720 8240 2800
rect 7120 2552 9280 2720
rect 7120 2488 7288 2552
rect 9112 2488 9280 2552
rect 7120 2320 9280 2488
rect 8160 2240 8240 2320
rect 9360 2240 9440 2800
rect 10560 2720 10640 2800
rect 9520 2552 11680 2720
rect 9520 2488 9688 2552
rect 11512 2488 11680 2552
rect 9520 2320 11680 2488
rect 10560 2240 10640 2320
rect 11760 2240 11840 2800
rect 12960 2720 13040 2800
rect 11920 2552 14080 2720
rect 11920 2488 12088 2552
rect 13912 2488 14080 2552
rect 11920 2320 14080 2488
rect 12960 2240 13040 2320
rect 14160 2240 14240 2800
rect 14320 2720 14400 2800
rect 14480 2720 14560 2800
rect 14640 2720 14720 2800
rect 14320 2552 14720 2720
rect 14320 2488 14488 2552
rect 14552 2488 14720 2552
rect 14320 2320 14720 2488
rect 14320 2240 14400 2320
rect 14480 2240 14560 2320
rect 14640 2240 14720 2320
rect -12800 2232 14880 2240
rect -12800 2168 -12712 2232
rect -12648 2168 -12552 2232
rect -12488 2168 -12392 2232
rect -12328 2168 -12232 2232
rect -12168 2168 -9832 2232
rect -9768 2168 -7432 2232
rect -7368 2168 -5032 2232
rect -4968 2168 -2632 2232
rect -2568 2168 -232 2232
rect -168 2168 2168 2232
rect 2232 2168 4568 2232
rect 4632 2168 6968 2232
rect 7032 2168 9368 2232
rect 9432 2168 11768 2232
rect 11832 2168 14168 2232
rect 14232 2168 14328 2232
rect 14392 2168 14488 2232
rect 14552 2168 14648 2232
rect 14712 2168 14880 2232
rect -12800 2160 14880 2168
rect -11040 2080 -10960 2160
rect -8640 2080 -8560 2160
rect -6240 2080 -6160 2160
rect -3840 2080 -3760 2160
rect -1440 2080 -1360 2160
rect 960 2080 1040 2160
rect 3360 2080 3440 2160
rect 5760 2080 5840 2160
rect 8160 2080 8240 2160
rect 10560 2080 10640 2160
rect 12960 2080 13040 2160
rect -12800 2072 14880 2080
rect -12800 2008 968 2072
rect 1032 2008 14328 2072
rect 14392 2008 14488 2072
rect 14552 2008 14648 2072
rect 14712 2008 14880 2072
rect -12800 2000 14880 2008
rect -11040 1920 -10960 2000
rect -8640 1920 -8560 2000
rect -6240 1920 -6160 2000
rect -3840 1920 -3760 2000
rect -1440 1920 -1360 2000
rect 3360 1920 3440 2000
rect 5760 1920 5840 2000
rect 8160 1920 8240 2000
rect 10560 1920 10640 2000
rect 12960 1920 13040 2000
rect -12800 1912 14880 1920
rect -12800 1848 -12712 1912
rect -12648 1848 -12552 1912
rect -12488 1848 -12392 1912
rect -12328 1848 14328 1912
rect 14392 1848 14488 1912
rect 14552 1848 14648 1912
rect 14712 1848 14880 1912
rect -12800 1840 14880 1848
rect -11040 1760 -10960 1840
rect -8640 1760 -8560 1840
rect -6240 1760 -6160 1840
rect -3840 1760 -3760 1840
rect -1440 1760 -1360 1840
rect 3360 1760 3440 1840
rect 5760 1760 5840 1840
rect 8160 1760 8240 1840
rect 10560 1760 10640 1840
rect 12960 1760 13040 1840
rect -12800 1752 14880 1760
rect -12800 1688 -11032 1752
rect -10968 1688 -8632 1752
rect -8568 1688 -6232 1752
rect -6168 1688 -3832 1752
rect -3768 1688 -1432 1752
rect -1368 1688 3368 1752
rect 3432 1688 5768 1752
rect 5832 1688 8168 1752
rect 8232 1688 10568 1752
rect 10632 1688 12968 1752
rect 13032 1688 14328 1752
rect 14392 1688 14488 1752
rect 14552 1688 14648 1752
rect 14712 1688 14880 1752
rect -12800 1680 14880 1688
rect -12800 1592 14880 1600
rect -12800 1528 -12712 1592
rect -12648 1528 -12552 1592
rect -12488 1528 -12392 1592
rect -12328 1528 14328 1592
rect 14392 1528 14488 1592
rect 14552 1528 14648 1592
rect 14712 1528 14880 1592
rect -12800 1520 14880 1528
<< labels >>
rlabel metal4 s 14800 3440 14880 3520 4 gnda
port 1 nsew
rlabel locali s 14800 3600 14880 3680 4 vssa
port 2 nsew
<< end >>
