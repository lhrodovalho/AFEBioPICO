* fully-differential single stage OTA open-loop testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
*.include "../mag/ota_core.spice"
.include "../mag/ota.spice"

* supply voltages
vdda  vdda 0 1.8
vssa  vssa 0 0.0

* DUT
x0 im ip op om ib q vdda gnda vssa ota
IB vdda ib 10n

egnda gnda vssa q vssa 1
vin in gnda dc 0 ac 1 
eip ip gnda in gnda  0.5
eim im gnda in gnda -0.5

clp op gnda 10p
clm om gnda 10p

*.save v(in) v(out) v(ib) i(vdda)
.option gmin=1e-12
.control

	op
	print i(vdda) v(op) v(om) v(q) v(vddx)
	
	dc vin -100m 100m 1m
	plot ip im op om x0.vddx vdda
	
	ac dec 10 1 1Meg
	plot vdb(op,ip)

	noise v(op,om) vin dec 10 1 100
	print inoise_total onoise_total	

.endc

.end
