* NGSPICE file created from p1_8.ext - technology: sky130A

.subckt p1_8 D G S B
X0 x4 G x3 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X1 S G x1 B sky130_fd_pr__pfet_01v8_lvt ad=1.5e+12p pd=7e+06u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X2 x6 G x5 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X3 x2 G x1 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=0p ps=0u w=3e+06u l=8e+06u
X4 x6 G x7 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X5 x2 G x3 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X6 x4 G x5 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X7 D G x7 B sky130_fd_pr__pfet_01v8_lvt ad=1.5e+12p pd=7e+06u as=0p ps=0u w=3e+06u l=8e+06u
.ends

