magic
tech sky130A
timestamp 1637806411
<< mvnmos >>
rect 0 -960 200 -860
rect 320 -960 520 -860
rect 640 -960 840 -860
rect 960 -960 1160 -860
rect 1280 -960 1480 -860
rect 1600 -960 1800 -860
rect 1920 -960 2120 -860
rect 2240 -960 2440 -860
rect 2560 -960 2760 -860
rect 2880 -960 3080 -860
rect 3200 -960 3400 -860
rect 3520 -960 3720 -860
rect 3840 -960 4040 -860
rect 4160 -960 4360 -860
rect 4480 -960 4680 -860
rect 4800 -960 5000 -860
rect 0 -1240 200 -1140
rect 320 -1240 520 -1140
rect 640 -1240 840 -1140
rect 960 -1240 1160 -1140
rect 1280 -1240 1480 -1140
rect 1600 -1240 1800 -1140
rect 1920 -1240 2120 -1140
rect 2240 -1240 2440 -1140
rect 2560 -1240 2760 -1140
rect 2880 -1240 3080 -1140
rect 3200 -1240 3400 -1140
rect 3520 -1240 3720 -1140
rect 3840 -1240 4040 -1140
rect 4160 -1240 4360 -1140
rect 4480 -1240 4680 -1140
rect 4800 -1240 5000 -1140
rect 0 -1440 200 -1340
rect 320 -1440 520 -1340
rect 640 -1440 840 -1340
rect 960 -1440 1160 -1340
rect 1280 -1440 1480 -1340
rect 1600 -1440 1800 -1340
rect 1920 -1440 2120 -1340
rect 2240 -1440 2440 -1340
rect 2560 -1440 2760 -1340
rect 2880 -1440 3080 -1340
rect 3200 -1440 3400 -1340
rect 3520 -1440 3720 -1340
rect 3840 -1440 4040 -1340
rect 4160 -1440 4360 -1340
rect 4480 -1440 4680 -1340
rect 4800 -1440 5000 -1340
<< mvndiff >>
rect -80 -870 0 -860
rect -80 -950 -75 -870
rect -45 -950 0 -870
rect -80 -960 0 -950
rect 200 -870 320 -860
rect 200 -950 245 -870
rect 275 -950 320 -870
rect 200 -960 320 -950
rect 520 -870 640 -860
rect 520 -950 565 -870
rect 595 -950 640 -870
rect 520 -960 640 -950
rect 840 -870 960 -860
rect 840 -950 885 -870
rect 915 -950 960 -870
rect 840 -960 960 -950
rect 1160 -870 1280 -860
rect 1160 -950 1205 -870
rect 1235 -950 1280 -870
rect 1160 -960 1280 -950
rect 1480 -870 1600 -860
rect 1480 -950 1525 -870
rect 1555 -950 1600 -870
rect 1480 -960 1600 -950
rect 1800 -870 1920 -860
rect 1800 -950 1845 -870
rect 1875 -950 1920 -870
rect 1800 -960 1920 -950
rect 2120 -870 2240 -860
rect 2120 -950 2165 -870
rect 2195 -950 2240 -870
rect 2120 -960 2240 -950
rect 2440 -870 2560 -860
rect 2440 -950 2485 -870
rect 2515 -950 2560 -870
rect 2440 -960 2560 -950
rect 2760 -870 2880 -860
rect 2760 -950 2805 -870
rect 2835 -950 2880 -870
rect 2760 -960 2880 -950
rect 3080 -870 3200 -860
rect 3080 -950 3125 -870
rect 3155 -950 3200 -870
rect 3080 -960 3200 -950
rect 3400 -870 3520 -860
rect 3400 -950 3445 -870
rect 3475 -950 3520 -870
rect 3400 -960 3520 -950
rect 3720 -870 3840 -860
rect 3720 -950 3765 -870
rect 3795 -950 3840 -870
rect 3720 -960 3840 -950
rect 4040 -870 4160 -860
rect 4040 -950 4085 -870
rect 4115 -950 4160 -870
rect 4040 -960 4160 -950
rect 4360 -870 4480 -860
rect 4360 -950 4405 -870
rect 4435 -950 4480 -870
rect 4360 -960 4480 -950
rect 4680 -870 4800 -860
rect 4680 -950 4725 -870
rect 4755 -950 4800 -870
rect 4680 -960 4800 -950
rect 5000 -870 5080 -860
rect 5000 -950 5045 -870
rect 5075 -950 5080 -870
rect 5000 -960 5080 -950
rect -80 -1150 0 -1140
rect -80 -1230 -75 -1150
rect -45 -1230 0 -1150
rect -80 -1240 0 -1230
rect 200 -1150 320 -1140
rect 200 -1230 245 -1150
rect 275 -1230 320 -1150
rect 200 -1240 320 -1230
rect 520 -1150 640 -1140
rect 520 -1230 565 -1150
rect 595 -1230 640 -1150
rect 520 -1240 640 -1230
rect 840 -1150 960 -1140
rect 840 -1230 885 -1150
rect 915 -1230 960 -1150
rect 840 -1240 960 -1230
rect 1160 -1150 1280 -1140
rect 1160 -1230 1205 -1150
rect 1235 -1230 1280 -1150
rect 1160 -1240 1280 -1230
rect 1480 -1150 1600 -1140
rect 1480 -1230 1525 -1150
rect 1555 -1230 1600 -1150
rect 1480 -1240 1600 -1230
rect 1800 -1150 1920 -1140
rect 1800 -1230 1845 -1150
rect 1875 -1230 1920 -1150
rect 1800 -1240 1920 -1230
rect 2120 -1150 2240 -1140
rect 2120 -1230 2165 -1150
rect 2195 -1230 2240 -1150
rect 2120 -1240 2240 -1230
rect 2440 -1150 2560 -1140
rect 2440 -1230 2485 -1150
rect 2515 -1230 2560 -1150
rect 2440 -1240 2560 -1230
rect 2760 -1150 2880 -1140
rect 2760 -1230 2805 -1150
rect 2835 -1230 2880 -1150
rect 2760 -1240 2880 -1230
rect 3080 -1150 3200 -1140
rect 3080 -1230 3125 -1150
rect 3155 -1230 3200 -1150
rect 3080 -1240 3200 -1230
rect 3400 -1150 3520 -1140
rect 3400 -1230 3445 -1150
rect 3475 -1230 3520 -1150
rect 3400 -1240 3520 -1230
rect 3720 -1150 3840 -1140
rect 3720 -1230 3765 -1150
rect 3795 -1230 3840 -1150
rect 3720 -1240 3840 -1230
rect 4040 -1150 4160 -1140
rect 4040 -1230 4085 -1150
rect 4115 -1230 4160 -1150
rect 4040 -1240 4160 -1230
rect 4360 -1150 4480 -1140
rect 4360 -1230 4405 -1150
rect 4435 -1230 4480 -1150
rect 4360 -1240 4480 -1230
rect 4680 -1150 4800 -1140
rect 4680 -1230 4725 -1150
rect 4755 -1230 4800 -1150
rect 4680 -1240 4800 -1230
rect 5000 -1150 5080 -1140
rect 5000 -1230 5045 -1150
rect 5075 -1230 5080 -1150
rect 5000 -1240 5080 -1230
rect -80 -1350 0 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 0 -1350
rect -80 -1440 0 -1430
rect 200 -1350 320 -1340
rect 200 -1430 245 -1350
rect 275 -1430 320 -1350
rect 200 -1440 320 -1430
rect 520 -1350 640 -1340
rect 520 -1430 565 -1350
rect 595 -1430 640 -1350
rect 520 -1440 640 -1430
rect 840 -1350 960 -1340
rect 840 -1430 885 -1350
rect 915 -1430 960 -1350
rect 840 -1440 960 -1430
rect 1160 -1350 1280 -1340
rect 1160 -1430 1205 -1350
rect 1235 -1430 1280 -1350
rect 1160 -1440 1280 -1430
rect 1480 -1350 1600 -1340
rect 1480 -1430 1525 -1350
rect 1555 -1430 1600 -1350
rect 1480 -1440 1600 -1430
rect 1800 -1350 1920 -1340
rect 1800 -1430 1845 -1350
rect 1875 -1430 1920 -1350
rect 1800 -1440 1920 -1430
rect 2120 -1350 2240 -1340
rect 2120 -1430 2165 -1350
rect 2195 -1430 2240 -1350
rect 2120 -1440 2240 -1430
rect 2440 -1350 2560 -1340
rect 2440 -1430 2485 -1350
rect 2515 -1430 2560 -1350
rect 2440 -1440 2560 -1430
rect 2760 -1350 2880 -1340
rect 2760 -1430 2805 -1350
rect 2835 -1430 2880 -1350
rect 2760 -1440 2880 -1430
rect 3080 -1350 3200 -1340
rect 3080 -1430 3125 -1350
rect 3155 -1430 3200 -1350
rect 3080 -1440 3200 -1430
rect 3400 -1350 3520 -1340
rect 3400 -1430 3445 -1350
rect 3475 -1430 3520 -1350
rect 3400 -1440 3520 -1430
rect 3720 -1350 3840 -1340
rect 3720 -1430 3765 -1350
rect 3795 -1430 3840 -1350
rect 3720 -1440 3840 -1430
rect 4040 -1350 4160 -1340
rect 4040 -1430 4085 -1350
rect 4115 -1430 4160 -1350
rect 4040 -1440 4160 -1430
rect 4360 -1350 4480 -1340
rect 4360 -1430 4405 -1350
rect 4435 -1430 4480 -1350
rect 4360 -1440 4480 -1430
rect 4680 -1350 4800 -1340
rect 4680 -1430 4725 -1350
rect 4755 -1430 4800 -1350
rect 4680 -1440 4800 -1430
rect 5000 -1350 5080 -1340
rect 5000 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5000 -1440 5080 -1430
<< mvndiffc >>
rect -75 -950 -45 -870
rect 245 -950 275 -870
rect 565 -950 595 -870
rect 885 -950 915 -870
rect 1205 -950 1235 -870
rect 1525 -950 1555 -870
rect 1845 -950 1875 -870
rect 2165 -950 2195 -870
rect 2485 -950 2515 -870
rect 2805 -950 2835 -870
rect 3125 -950 3155 -870
rect 3445 -950 3475 -870
rect 3765 -950 3795 -870
rect 4085 -950 4115 -870
rect 4405 -950 4435 -870
rect 4725 -950 4755 -870
rect 5045 -950 5075 -870
rect -75 -1230 -45 -1150
rect 245 -1230 275 -1150
rect 565 -1230 595 -1150
rect 885 -1230 915 -1150
rect 1205 -1230 1235 -1150
rect 1525 -1230 1555 -1150
rect 1845 -1230 1875 -1150
rect 2165 -1230 2195 -1150
rect 2485 -1230 2515 -1150
rect 2805 -1230 2835 -1150
rect 3125 -1230 3155 -1150
rect 3445 -1230 3475 -1150
rect 3765 -1230 3795 -1150
rect 4085 -1230 4115 -1150
rect 4405 -1230 4435 -1150
rect 4725 -1230 4755 -1150
rect 5045 -1230 5075 -1150
rect -75 -1430 -45 -1350
rect 245 -1430 275 -1350
rect 565 -1430 595 -1350
rect 885 -1430 915 -1350
rect 1205 -1430 1235 -1350
rect 1525 -1430 1555 -1350
rect 1845 -1430 1875 -1350
rect 2165 -1430 2195 -1350
rect 2485 -1430 2515 -1350
rect 2805 -1430 2835 -1350
rect 3125 -1430 3155 -1350
rect 3445 -1430 3475 -1350
rect 3765 -1430 3795 -1350
rect 4085 -1430 4115 -1350
rect 4405 -1430 4435 -1350
rect 4725 -1430 4755 -1350
rect 5045 -1430 5075 -1350
<< psubdiff >>
rect -240 -760 -180 -720
rect 5180 -760 5240 -720
rect -240 -780 -200 -760
rect 5200 -780 5240 -760
rect -200 -1040 -180 -1000
rect 5180 -1040 5200 -1000
rect -240 -1480 -200 -1460
rect 5200 -1480 5240 -1460
rect -240 -1520 -180 -1480
rect 5180 -1520 5240 -1480
<< psubdiffcont >>
rect -180 -760 5180 -720
rect -240 -1460 -200 -780
rect -180 -1040 5180 -1000
rect 5200 -1460 5240 -780
rect -180 -1520 5180 -1480
<< poly >>
rect 0 -805 200 -800
rect 0 -835 10 -805
rect 190 -835 200 -805
rect 0 -860 200 -835
rect 320 -805 520 -800
rect 320 -835 330 -805
rect 510 -835 520 -805
rect 320 -860 520 -835
rect 640 -805 840 -800
rect 640 -835 650 -805
rect 830 -835 840 -805
rect 640 -860 840 -835
rect 960 -805 1160 -800
rect 960 -835 970 -805
rect 1150 -835 1160 -805
rect 960 -860 1160 -835
rect 1280 -805 1480 -800
rect 1280 -835 1290 -805
rect 1470 -835 1480 -805
rect 1280 -860 1480 -835
rect 1600 -805 1800 -800
rect 1600 -835 1610 -805
rect 1790 -835 1800 -805
rect 1600 -860 1800 -835
rect 1920 -805 2120 -800
rect 1920 -835 1930 -805
rect 2110 -835 2120 -805
rect 1920 -860 2120 -835
rect 2240 -805 2440 -800
rect 2240 -835 2250 -805
rect 2430 -835 2440 -805
rect 2240 -860 2440 -835
rect 2560 -805 2760 -800
rect 2560 -835 2570 -805
rect 2750 -835 2760 -805
rect 2560 -860 2760 -835
rect 2880 -805 3080 -800
rect 2880 -835 2890 -805
rect 3070 -835 3080 -805
rect 2880 -860 3080 -835
rect 3200 -805 3400 -800
rect 3200 -835 3210 -805
rect 3390 -835 3400 -805
rect 3200 -860 3400 -835
rect 3520 -805 3720 -800
rect 3520 -835 3530 -805
rect 3710 -835 3720 -805
rect 3520 -860 3720 -835
rect 3840 -805 4040 -800
rect 3840 -835 3850 -805
rect 4030 -835 4040 -805
rect 3840 -860 4040 -835
rect 4160 -805 4360 -800
rect 4160 -835 4170 -805
rect 4350 -835 4360 -805
rect 4160 -860 4360 -835
rect 4480 -805 4680 -800
rect 4480 -835 4490 -805
rect 4670 -835 4680 -805
rect 4480 -860 4680 -835
rect 4800 -805 5000 -800
rect 4800 -835 4810 -805
rect 4990 -835 5000 -805
rect 4800 -860 5000 -835
rect 0 -980 200 -960
rect 320 -980 520 -960
rect 640 -980 840 -960
rect 960 -980 1160 -960
rect 1280 -980 1480 -960
rect 1600 -980 1800 -960
rect 1920 -980 2120 -960
rect 2240 -980 2440 -960
rect 2560 -980 2760 -960
rect 2880 -980 3080 -960
rect 3200 -980 3400 -960
rect 3520 -980 3720 -960
rect 3840 -980 4040 -960
rect 4160 -980 4360 -960
rect 4480 -980 4680 -960
rect 4800 -980 5000 -960
rect 0 -1085 200 -1080
rect 0 -1115 10 -1085
rect 190 -1115 200 -1085
rect 0 -1140 200 -1115
rect 320 -1085 520 -1080
rect 320 -1115 330 -1085
rect 510 -1115 520 -1085
rect 320 -1140 520 -1115
rect 640 -1085 840 -1080
rect 640 -1115 650 -1085
rect 830 -1115 840 -1085
rect 640 -1140 840 -1115
rect 960 -1085 1160 -1080
rect 960 -1115 970 -1085
rect 1150 -1115 1160 -1085
rect 960 -1140 1160 -1115
rect 1280 -1085 1480 -1080
rect 1280 -1115 1290 -1085
rect 1470 -1115 1480 -1085
rect 1280 -1140 1480 -1115
rect 1600 -1085 1800 -1080
rect 1600 -1115 1610 -1085
rect 1790 -1115 1800 -1085
rect 1600 -1140 1800 -1115
rect 1920 -1085 2120 -1080
rect 1920 -1115 1930 -1085
rect 2110 -1115 2120 -1085
rect 1920 -1140 2120 -1115
rect 2240 -1085 2440 -1080
rect 2240 -1115 2250 -1085
rect 2430 -1115 2440 -1085
rect 2240 -1140 2440 -1115
rect 2560 -1085 2760 -1080
rect 2560 -1115 2570 -1085
rect 2750 -1115 2760 -1085
rect 2560 -1140 2760 -1115
rect 2880 -1085 3080 -1080
rect 2880 -1115 2890 -1085
rect 3070 -1115 3080 -1085
rect 2880 -1140 3080 -1115
rect 3200 -1085 3400 -1080
rect 3200 -1115 3210 -1085
rect 3390 -1115 3400 -1085
rect 3200 -1140 3400 -1115
rect 3520 -1085 3720 -1080
rect 3520 -1115 3530 -1085
rect 3710 -1115 3720 -1085
rect 3520 -1140 3720 -1115
rect 3840 -1085 4040 -1080
rect 3840 -1115 3850 -1085
rect 4030 -1115 4040 -1085
rect 3840 -1140 4040 -1115
rect 4160 -1085 4360 -1080
rect 4160 -1115 4170 -1085
rect 4350 -1115 4360 -1085
rect 4160 -1140 4360 -1115
rect 4480 -1085 4680 -1080
rect 4480 -1115 4490 -1085
rect 4670 -1115 4680 -1085
rect 4480 -1140 4680 -1115
rect 4800 -1085 5000 -1080
rect 4800 -1115 4810 -1085
rect 4990 -1115 5000 -1085
rect 4800 -1140 5000 -1115
rect 0 -1340 200 -1240
rect 320 -1340 520 -1240
rect 640 -1340 840 -1240
rect 960 -1340 1160 -1240
rect 1280 -1340 1480 -1240
rect 1600 -1340 1800 -1240
rect 1920 -1340 2120 -1240
rect 2240 -1340 2440 -1240
rect 2560 -1340 2760 -1240
rect 2880 -1340 3080 -1240
rect 3200 -1340 3400 -1240
rect 3520 -1340 3720 -1240
rect 3840 -1340 4040 -1240
rect 4160 -1340 4360 -1240
rect 4480 -1340 4680 -1240
rect 4800 -1340 5000 -1240
rect 0 -1460 200 -1440
rect 320 -1460 520 -1440
rect 640 -1460 840 -1440
rect 960 -1460 1160 -1440
rect 1280 -1460 1480 -1440
rect 1600 -1460 1800 -1440
rect 1920 -1460 2120 -1440
rect 2240 -1460 2440 -1440
rect 2560 -1460 2760 -1440
rect 2880 -1460 3080 -1440
rect 3200 -1460 3400 -1440
rect 3520 -1460 3720 -1440
rect 3840 -1460 4040 -1440
rect 4160 -1460 4360 -1440
rect 4480 -1460 4680 -1440
rect 4800 -1460 5000 -1440
<< polycont >>
rect 10 -835 190 -805
rect 330 -835 510 -805
rect 650 -835 830 -805
rect 970 -835 1150 -805
rect 1290 -835 1470 -805
rect 1610 -835 1790 -805
rect 1930 -835 2110 -805
rect 2250 -835 2430 -805
rect 2570 -835 2750 -805
rect 2890 -835 3070 -805
rect 3210 -835 3390 -805
rect 3530 -835 3710 -805
rect 3850 -835 4030 -805
rect 4170 -835 4350 -805
rect 4490 -835 4670 -805
rect 4810 -835 4990 -805
rect 10 -1115 190 -1085
rect 330 -1115 510 -1085
rect 650 -1115 830 -1085
rect 970 -1115 1150 -1085
rect 1290 -1115 1470 -1085
rect 1610 -1115 1790 -1085
rect 1930 -1115 2110 -1085
rect 2250 -1115 2430 -1085
rect 2570 -1115 2750 -1085
rect 2890 -1115 3070 -1085
rect 3210 -1115 3390 -1085
rect 3530 -1115 3710 -1085
rect 3850 -1115 4030 -1085
rect 4170 -1115 4350 -1085
rect 4490 -1115 4670 -1085
rect 4810 -1115 4990 -1085
<< locali >>
rect -240 -760 -180 -720
rect 5180 -760 5240 -720
rect -240 -780 -200 -760
rect 5200 -780 5240 -760
rect 0 -805 200 -800
rect 0 -835 10 -805
rect 190 -835 200 -805
rect 0 -840 200 -835
rect 320 -805 520 -800
rect 320 -835 330 -805
rect 510 -835 520 -805
rect 320 -840 520 -835
rect 640 -805 840 -800
rect 640 -835 650 -805
rect 830 -835 840 -805
rect 640 -840 840 -835
rect 960 -805 1160 -800
rect 960 -835 970 -805
rect 1150 -835 1160 -805
rect 960 -840 1160 -835
rect 1280 -805 1480 -800
rect 1280 -835 1290 -805
rect 1470 -835 1480 -805
rect 1280 -840 1480 -835
rect 1600 -805 1800 -800
rect 1600 -835 1610 -805
rect 1790 -835 1800 -805
rect 1600 -840 1800 -835
rect 1920 -805 2120 -800
rect 1920 -835 1930 -805
rect 2110 -835 2120 -805
rect 1920 -840 2120 -835
rect 2240 -805 2440 -800
rect 2240 -835 2250 -805
rect 2430 -835 2440 -805
rect 2240 -840 2440 -835
rect 2560 -805 2760 -800
rect 2560 -835 2570 -805
rect 2750 -835 2760 -805
rect 2560 -840 2760 -835
rect 2880 -805 3080 -800
rect 2880 -835 2890 -805
rect 3070 -835 3080 -805
rect 2880 -840 3080 -835
rect 3200 -805 3400 -800
rect 3200 -835 3210 -805
rect 3390 -835 3400 -805
rect 3200 -840 3400 -835
rect 3520 -805 3720 -800
rect 3520 -835 3530 -805
rect 3710 -835 3720 -805
rect 3520 -840 3720 -835
rect 3840 -805 4040 -800
rect 3840 -835 3850 -805
rect 4030 -835 4040 -805
rect 3840 -840 4040 -835
rect 4160 -805 4360 -800
rect 4160 -835 4170 -805
rect 4350 -835 4360 -805
rect 4160 -840 4360 -835
rect 4480 -805 4680 -800
rect 4480 -835 4490 -805
rect 4670 -835 4680 -805
rect 4480 -840 4680 -835
rect 4800 -805 5000 -800
rect 4800 -835 4810 -805
rect 4990 -835 5000 -805
rect 4800 -840 5000 -835
rect -80 -870 -40 -860
rect -80 -950 -75 -870
rect -45 -950 -40 -870
rect -80 -960 -40 -950
rect 240 -870 280 -860
rect 240 -950 245 -870
rect 275 -950 280 -870
rect 240 -960 280 -950
rect 560 -870 600 -860
rect 560 -950 565 -870
rect 595 -950 600 -870
rect 560 -960 600 -950
rect 880 -870 920 -860
rect 880 -950 885 -870
rect 915 -950 920 -870
rect 880 -960 920 -950
rect 1200 -870 1240 -860
rect 1200 -950 1205 -870
rect 1235 -950 1240 -870
rect 1200 -960 1240 -950
rect 1520 -870 1560 -860
rect 1520 -950 1525 -870
rect 1555 -950 1560 -870
rect 1520 -960 1560 -950
rect 1840 -870 1880 -860
rect 1840 -950 1845 -870
rect 1875 -950 1880 -870
rect 1840 -960 1880 -950
rect 2160 -870 2200 -860
rect 2160 -950 2165 -870
rect 2195 -950 2200 -870
rect 2160 -960 2200 -950
rect 2480 -870 2520 -860
rect 2480 -950 2485 -870
rect 2515 -950 2520 -870
rect 2480 -960 2520 -950
rect 2800 -870 2840 -860
rect 2800 -950 2805 -870
rect 2835 -950 2840 -870
rect 2800 -960 2840 -950
rect 3120 -870 3160 -860
rect 3120 -950 3125 -870
rect 3155 -950 3160 -870
rect 3120 -960 3160 -950
rect 3440 -870 3480 -860
rect 3440 -950 3445 -870
rect 3475 -950 3480 -870
rect 3440 -960 3480 -950
rect 3760 -870 3800 -860
rect 3760 -950 3765 -870
rect 3795 -950 3800 -870
rect 3760 -960 3800 -950
rect 4080 -870 4120 -860
rect 4080 -950 4085 -870
rect 4115 -950 4120 -870
rect 4080 -960 4120 -950
rect 4400 -870 4440 -860
rect 4400 -950 4405 -870
rect 4435 -950 4440 -870
rect 4400 -960 4440 -950
rect 4720 -870 4760 -860
rect 4720 -950 4725 -870
rect 4755 -950 4760 -870
rect 4720 -960 4760 -950
rect 5040 -870 5080 -860
rect 5040 -950 5045 -870
rect 5075 -950 5080 -870
rect 5040 -960 5080 -950
rect -200 -1040 -180 -1000
rect 5180 -1040 5200 -1000
rect 0 -1085 200 -1080
rect 0 -1115 10 -1085
rect 190 -1115 200 -1085
rect 0 -1120 200 -1115
rect 320 -1085 520 -1080
rect 320 -1115 330 -1085
rect 510 -1115 520 -1085
rect 320 -1120 520 -1115
rect 640 -1085 840 -1080
rect 640 -1115 650 -1085
rect 830 -1115 840 -1085
rect 640 -1120 840 -1115
rect 960 -1085 1160 -1080
rect 960 -1115 970 -1085
rect 1150 -1115 1160 -1085
rect 960 -1120 1160 -1115
rect 1280 -1085 1480 -1080
rect 1280 -1115 1290 -1085
rect 1470 -1115 1480 -1085
rect 1280 -1120 1480 -1115
rect 1600 -1085 1800 -1080
rect 1600 -1115 1610 -1085
rect 1790 -1115 1800 -1085
rect 1600 -1120 1800 -1115
rect 1920 -1085 2120 -1080
rect 1920 -1115 1930 -1085
rect 2110 -1115 2120 -1085
rect 1920 -1120 2120 -1115
rect 2240 -1085 2440 -1080
rect 2240 -1115 2250 -1085
rect 2430 -1115 2440 -1085
rect 2240 -1120 2440 -1115
rect 2560 -1085 2760 -1080
rect 2560 -1115 2570 -1085
rect 2750 -1115 2760 -1085
rect 2560 -1120 2760 -1115
rect 2880 -1085 3080 -1080
rect 2880 -1115 2890 -1085
rect 3070 -1115 3080 -1085
rect 2880 -1120 3080 -1115
rect 3200 -1085 3400 -1080
rect 3200 -1115 3210 -1085
rect 3390 -1115 3400 -1085
rect 3200 -1120 3400 -1115
rect 3520 -1085 3720 -1080
rect 3520 -1115 3530 -1085
rect 3710 -1115 3720 -1085
rect 3520 -1120 3720 -1115
rect 3840 -1085 4040 -1080
rect 3840 -1115 3850 -1085
rect 4030 -1115 4040 -1085
rect 3840 -1120 4040 -1115
rect 4160 -1085 4360 -1080
rect 4160 -1115 4170 -1085
rect 4350 -1115 4360 -1085
rect 4160 -1120 4360 -1115
rect 4480 -1085 4680 -1080
rect 4480 -1115 4490 -1085
rect 4670 -1115 4680 -1085
rect 4480 -1120 4680 -1115
rect 4800 -1085 5000 -1080
rect 4800 -1115 4810 -1085
rect 4990 -1115 5000 -1085
rect 4800 -1120 5000 -1115
rect -80 -1150 -40 -1140
rect -80 -1230 -75 -1150
rect -45 -1230 -40 -1150
rect -80 -1240 -40 -1230
rect 240 -1150 280 -1140
rect 240 -1230 245 -1150
rect 275 -1230 280 -1150
rect 240 -1280 280 -1230
rect 560 -1150 600 -1140
rect 560 -1230 565 -1150
rect 595 -1230 600 -1150
rect 560 -1240 600 -1230
rect 880 -1150 920 -1140
rect 880 -1230 885 -1150
rect 915 -1230 920 -1150
rect 880 -1280 920 -1230
rect 1200 -1150 1240 -1140
rect 1200 -1230 1205 -1150
rect 1235 -1230 1240 -1150
rect 1200 -1240 1240 -1230
rect 1520 -1150 1560 -1140
rect 1520 -1230 1525 -1150
rect 1555 -1230 1560 -1150
rect 1520 -1280 1560 -1230
rect 1840 -1150 1880 -1140
rect 1840 -1230 1845 -1150
rect 1875 -1230 1880 -1150
rect 1840 -1240 1880 -1230
rect 2160 -1150 2200 -1140
rect 2160 -1230 2165 -1150
rect 2195 -1230 2200 -1150
rect 2160 -1280 2200 -1230
rect 2480 -1150 2520 -1140
rect 2480 -1230 2485 -1150
rect 2515 -1230 2520 -1150
rect 2480 -1240 2520 -1230
rect 2800 -1150 2840 -1140
rect 2800 -1230 2805 -1150
rect 2835 -1230 2840 -1150
rect 2800 -1280 2840 -1230
rect 3120 -1150 3160 -1140
rect 3120 -1230 3125 -1150
rect 3155 -1230 3160 -1150
rect 3120 -1240 3160 -1230
rect 3440 -1150 3480 -1140
rect 3440 -1230 3445 -1150
rect 3475 -1230 3480 -1150
rect 3440 -1280 3480 -1230
rect 3760 -1150 3800 -1140
rect 3760 -1230 3765 -1150
rect 3795 -1230 3800 -1150
rect 3760 -1240 3800 -1230
rect 4080 -1150 4120 -1140
rect 4080 -1230 4085 -1150
rect 4115 -1230 4120 -1150
rect 4080 -1280 4120 -1230
rect 4400 -1150 4440 -1140
rect 4400 -1230 4405 -1150
rect 4435 -1230 4440 -1150
rect 4400 -1240 4440 -1230
rect 4720 -1150 4760 -1140
rect 4720 -1230 4725 -1150
rect 4755 -1230 4760 -1150
rect 4720 -1280 4760 -1230
rect 5040 -1150 5080 -1140
rect 5040 -1230 5045 -1150
rect 5075 -1230 5080 -1150
rect 5040 -1240 5080 -1230
rect -80 -1320 5080 -1280
rect -240 -1480 -200 -1460
rect -80 -1350 -40 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 -40 -1350
rect -80 -1480 -40 -1430
rect 240 -1350 280 -1340
rect 240 -1430 245 -1350
rect 275 -1430 280 -1350
rect 240 -1440 280 -1430
rect 560 -1350 600 -1320
rect 560 -1430 565 -1350
rect 595 -1430 600 -1350
rect 560 -1440 600 -1430
rect 880 -1350 920 -1340
rect 880 -1430 885 -1350
rect 915 -1430 920 -1350
rect 880 -1440 920 -1430
rect 1200 -1350 1240 -1340
rect 1200 -1430 1205 -1350
rect 1235 -1430 1240 -1350
rect 1200 -1480 1240 -1430
rect 1520 -1350 1560 -1340
rect 1520 -1430 1525 -1350
rect 1555 -1430 1560 -1350
rect 1520 -1440 1560 -1430
rect 1840 -1350 1880 -1320
rect 1840 -1430 1845 -1350
rect 1875 -1430 1880 -1350
rect 1840 -1440 1880 -1430
rect 2160 -1350 2200 -1340
rect 2160 -1430 2165 -1350
rect 2195 -1430 2200 -1350
rect 2160 -1440 2200 -1430
rect 2480 -1350 2520 -1340
rect 2480 -1430 2485 -1350
rect 2515 -1430 2520 -1350
rect 2480 -1480 2520 -1430
rect 2800 -1350 2840 -1340
rect 2800 -1430 2805 -1350
rect 2835 -1430 2840 -1350
rect 2800 -1440 2840 -1430
rect 3120 -1350 3160 -1320
rect 3120 -1430 3125 -1350
rect 3155 -1430 3160 -1350
rect 3120 -1440 3160 -1430
rect 3440 -1350 3480 -1340
rect 3440 -1430 3445 -1350
rect 3475 -1430 3480 -1350
rect 3440 -1440 3480 -1430
rect 3760 -1350 3800 -1340
rect 3760 -1430 3765 -1350
rect 3795 -1430 3800 -1350
rect 3760 -1480 3800 -1430
rect 4080 -1350 4120 -1340
rect 4080 -1430 4085 -1350
rect 4115 -1430 4120 -1350
rect 4080 -1440 4120 -1430
rect 4400 -1350 4440 -1320
rect 4400 -1430 4405 -1350
rect 4435 -1430 4440 -1350
rect 4400 -1440 4440 -1430
rect 4720 -1350 4760 -1340
rect 4720 -1430 4725 -1350
rect 4755 -1430 4760 -1350
rect 4720 -1440 4760 -1430
rect 5040 -1350 5080 -1340
rect 5040 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5040 -1480 5080 -1430
rect 5200 -1480 5240 -1460
rect -240 -1520 -180 -1480
rect 5180 -1520 5240 -1480
<< viali >>
rect 10 -835 190 -805
rect 330 -835 510 -805
rect 650 -835 830 -805
rect 970 -835 1150 -805
rect 1290 -835 1470 -805
rect 1610 -835 1790 -805
rect 1930 -835 2110 -805
rect 2250 -835 2430 -805
rect 2570 -835 2750 -805
rect 2890 -835 3070 -805
rect 3210 -835 3390 -805
rect 3530 -835 3710 -805
rect 3850 -835 4030 -805
rect 4170 -835 4350 -805
rect 4490 -835 4670 -805
rect 4810 -835 4990 -805
rect -75 -950 -45 -870
rect 245 -950 275 -870
rect 565 -950 595 -870
rect 885 -950 915 -870
rect 1205 -950 1235 -870
rect 1525 -950 1555 -870
rect 1845 -950 1875 -870
rect 2165 -950 2195 -870
rect 2485 -950 2515 -870
rect 2805 -950 2835 -870
rect 3125 -950 3155 -870
rect 3445 -950 3475 -870
rect 3765 -950 3795 -870
rect 4085 -950 4115 -870
rect 4405 -950 4435 -870
rect 4725 -950 4755 -870
rect 5045 -950 5075 -870
rect 10 -1115 190 -1085
rect 330 -1115 510 -1085
rect 650 -1115 830 -1085
rect 970 -1115 1150 -1085
rect 1290 -1115 1470 -1085
rect 1610 -1115 1790 -1085
rect 1930 -1115 2110 -1085
rect 2250 -1115 2430 -1085
rect 2570 -1115 2750 -1085
rect 2890 -1115 3070 -1085
rect 3210 -1115 3390 -1085
rect 3530 -1115 3710 -1085
rect 3850 -1115 4030 -1085
rect 4170 -1115 4350 -1085
rect 4490 -1115 4670 -1085
rect 4810 -1115 4990 -1085
rect -75 -1230 -45 -1150
rect 245 -1230 275 -1150
rect 565 -1230 595 -1150
rect 885 -1230 915 -1150
rect 1205 -1230 1235 -1150
rect 1525 -1230 1555 -1150
rect 1845 -1230 1875 -1150
rect 2165 -1230 2195 -1150
rect 2485 -1230 2515 -1150
rect 2805 -1230 2835 -1150
rect 3125 -1230 3155 -1150
rect 3445 -1230 3475 -1150
rect 3765 -1230 3795 -1150
rect 4085 -1230 4115 -1150
rect 4405 -1230 4435 -1150
rect 4725 -1230 4755 -1150
rect 5045 -1230 5075 -1150
rect -75 -1430 -45 -1350
rect 245 -1430 275 -1350
rect 565 -1430 595 -1350
rect 885 -1430 915 -1350
rect 1205 -1430 1235 -1350
rect 1525 -1430 1555 -1350
rect 1845 -1430 1875 -1350
rect 2165 -1430 2195 -1350
rect 2485 -1430 2515 -1350
rect 2805 -1430 2835 -1350
rect 3125 -1430 3155 -1350
rect 3445 -1430 3475 -1350
rect 3765 -1430 3795 -1350
rect 4085 -1430 4115 -1350
rect 4405 -1430 4435 -1350
rect 4725 -1430 4755 -1350
rect 5045 -1430 5075 -1350
<< metal1 >>
rect 0 -805 200 -800
rect 0 -835 10 -805
rect 190 -835 200 -805
rect 0 -840 200 -835
rect 240 -805 280 -800
rect 240 -835 245 -805
rect 275 -835 280 -805
rect -80 -870 -40 -860
rect -80 -950 -75 -870
rect -45 -950 -40 -870
rect -80 -1085 -40 -950
rect 240 -870 280 -835
rect 320 -805 520 -800
rect 320 -835 330 -805
rect 510 -835 520 -805
rect 320 -840 520 -835
rect 640 -805 840 -800
rect 640 -835 650 -805
rect 830 -835 840 -805
rect 640 -840 840 -835
rect 880 -805 920 -800
rect 880 -835 885 -805
rect 915 -835 920 -805
rect 240 -950 245 -870
rect 275 -950 280 -870
rect 240 -960 280 -950
rect 560 -870 600 -860
rect 560 -950 565 -870
rect 595 -950 600 -870
rect -80 -1115 -75 -1085
rect -45 -1115 -40 -1085
rect -80 -1150 -40 -1115
rect 0 -1085 200 -1080
rect 0 -1115 10 -1085
rect 190 -1115 200 -1085
rect 0 -1120 200 -1115
rect 320 -1085 520 -1080
rect 320 -1115 330 -1085
rect 510 -1115 520 -1085
rect 320 -1120 520 -1115
rect 560 -1085 600 -950
rect 880 -870 920 -835
rect 960 -805 1160 -800
rect 960 -835 970 -805
rect 1150 -835 1160 -805
rect 960 -840 1160 -835
rect 1280 -805 1480 -800
rect 1280 -835 1290 -805
rect 1470 -835 1480 -805
rect 1280 -840 1480 -835
rect 1520 -805 1560 -800
rect 1520 -835 1525 -805
rect 1555 -835 1560 -805
rect 880 -950 885 -870
rect 915 -950 920 -870
rect 880 -960 920 -950
rect 1200 -870 1240 -860
rect 1200 -950 1205 -870
rect 1235 -950 1240 -870
rect 560 -1115 565 -1085
rect 595 -1115 600 -1085
rect -80 -1230 -75 -1150
rect -45 -1230 -40 -1150
rect -80 -1240 -40 -1230
rect 240 -1150 280 -1140
rect 240 -1230 245 -1150
rect 275 -1230 280 -1150
rect 240 -1240 280 -1230
rect 560 -1150 600 -1115
rect 640 -1085 840 -1080
rect 640 -1115 650 -1085
rect 830 -1115 840 -1085
rect 640 -1120 840 -1115
rect 960 -1085 1160 -1080
rect 960 -1115 970 -1085
rect 1150 -1115 1160 -1085
rect 960 -1120 1160 -1115
rect 1200 -1085 1240 -950
rect 1520 -870 1560 -835
rect 1600 -805 1800 -800
rect 1600 -835 1610 -805
rect 1790 -835 1800 -805
rect 1600 -840 1800 -835
rect 1920 -805 2120 -800
rect 1920 -835 1930 -805
rect 2110 -835 2120 -805
rect 1920 -840 2120 -835
rect 2160 -805 2200 -800
rect 2160 -835 2165 -805
rect 2195 -835 2200 -805
rect 1520 -950 1525 -870
rect 1555 -950 1560 -870
rect 1520 -960 1560 -950
rect 1840 -870 1880 -860
rect 1840 -950 1845 -870
rect 1875 -950 1880 -870
rect 1200 -1115 1205 -1085
rect 1235 -1115 1240 -1085
rect 560 -1230 565 -1150
rect 595 -1230 600 -1150
rect 560 -1240 600 -1230
rect 880 -1150 920 -1140
rect 880 -1230 885 -1150
rect 915 -1230 920 -1150
rect 880 -1240 920 -1230
rect 1200 -1150 1240 -1115
rect 1280 -1085 1480 -1080
rect 1280 -1115 1290 -1085
rect 1470 -1115 1480 -1085
rect 1280 -1120 1480 -1115
rect 1600 -1085 1800 -1080
rect 1600 -1115 1610 -1085
rect 1790 -1115 1800 -1085
rect 1600 -1120 1800 -1115
rect 1840 -1085 1880 -950
rect 2160 -870 2200 -835
rect 2240 -805 2440 -800
rect 2240 -835 2250 -805
rect 2430 -835 2440 -805
rect 2240 -840 2440 -835
rect 2560 -805 2760 -800
rect 2560 -835 2570 -805
rect 2750 -835 2760 -805
rect 2560 -840 2760 -835
rect 2800 -805 2840 -800
rect 2800 -835 2805 -805
rect 2835 -835 2840 -805
rect 2160 -950 2165 -870
rect 2195 -950 2200 -870
rect 2160 -960 2200 -950
rect 2480 -870 2520 -860
rect 2480 -950 2485 -870
rect 2515 -950 2520 -870
rect 1840 -1115 1845 -1085
rect 1875 -1115 1880 -1085
rect 1200 -1230 1205 -1150
rect 1235 -1230 1240 -1150
rect 1200 -1240 1240 -1230
rect 1520 -1150 1560 -1140
rect 1520 -1230 1525 -1150
rect 1555 -1230 1560 -1150
rect 1520 -1240 1560 -1230
rect 1840 -1150 1880 -1115
rect 1920 -1085 2120 -1080
rect 1920 -1115 1930 -1085
rect 2110 -1115 2120 -1085
rect 1920 -1120 2120 -1115
rect 2240 -1085 2440 -1080
rect 2240 -1115 2250 -1085
rect 2430 -1115 2440 -1085
rect 2240 -1120 2440 -1115
rect 2480 -1085 2520 -950
rect 2800 -870 2840 -835
rect 2880 -805 3080 -800
rect 2880 -835 2890 -805
rect 3070 -835 3080 -805
rect 2880 -840 3080 -835
rect 3200 -805 3400 -800
rect 3200 -835 3210 -805
rect 3390 -835 3400 -805
rect 3200 -840 3400 -835
rect 3440 -805 3480 -800
rect 3440 -835 3445 -805
rect 3475 -835 3480 -805
rect 2800 -950 2805 -870
rect 2835 -950 2840 -870
rect 2800 -960 2840 -950
rect 3120 -870 3160 -860
rect 3120 -950 3125 -870
rect 3155 -950 3160 -870
rect 2480 -1115 2485 -1085
rect 2515 -1115 2520 -1085
rect 1840 -1230 1845 -1150
rect 1875 -1230 1880 -1150
rect 1840 -1240 1880 -1230
rect 2160 -1150 2200 -1140
rect 2160 -1230 2165 -1150
rect 2195 -1230 2200 -1150
rect 2160 -1240 2200 -1230
rect 2480 -1150 2520 -1115
rect 2560 -1085 2760 -1080
rect 2560 -1115 2570 -1085
rect 2750 -1115 2760 -1085
rect 2560 -1120 2760 -1115
rect 2880 -1085 3080 -1080
rect 2880 -1115 2890 -1085
rect 3070 -1115 3080 -1085
rect 2880 -1120 3080 -1115
rect 3120 -1085 3160 -950
rect 3440 -870 3480 -835
rect 3520 -805 3720 -800
rect 3520 -835 3530 -805
rect 3710 -835 3720 -805
rect 3520 -840 3720 -835
rect 3840 -805 4040 -800
rect 3840 -835 3850 -805
rect 4030 -835 4040 -805
rect 3840 -840 4040 -835
rect 4080 -805 4120 -800
rect 4080 -835 4085 -805
rect 4115 -835 4120 -805
rect 3440 -950 3445 -870
rect 3475 -950 3480 -870
rect 3440 -960 3480 -950
rect 3760 -870 3800 -860
rect 3760 -950 3765 -870
rect 3795 -950 3800 -870
rect 3120 -1115 3125 -1085
rect 3155 -1115 3160 -1085
rect 2480 -1230 2485 -1150
rect 2515 -1230 2520 -1150
rect 2480 -1240 2520 -1230
rect 2800 -1150 2840 -1140
rect 2800 -1230 2805 -1150
rect 2835 -1230 2840 -1150
rect 2800 -1240 2840 -1230
rect 3120 -1150 3160 -1115
rect 3200 -1085 3400 -1080
rect 3200 -1115 3210 -1085
rect 3390 -1115 3400 -1085
rect 3200 -1120 3400 -1115
rect 3520 -1085 3720 -1080
rect 3520 -1115 3530 -1085
rect 3710 -1115 3720 -1085
rect 3520 -1120 3720 -1115
rect 3760 -1085 3800 -950
rect 4080 -870 4120 -835
rect 4160 -805 4360 -800
rect 4160 -835 4170 -805
rect 4350 -835 4360 -805
rect 4160 -840 4360 -835
rect 4480 -805 4680 -800
rect 4480 -835 4490 -805
rect 4670 -835 4680 -805
rect 4480 -840 4680 -835
rect 4720 -805 4760 -800
rect 4720 -835 4725 -805
rect 4755 -835 4760 -805
rect 4080 -950 4085 -870
rect 4115 -950 4120 -870
rect 4080 -960 4120 -950
rect 4400 -870 4440 -860
rect 4400 -950 4405 -870
rect 4435 -950 4440 -870
rect 3760 -1115 3765 -1085
rect 3795 -1115 3800 -1085
rect 3120 -1230 3125 -1150
rect 3155 -1230 3160 -1150
rect 3120 -1240 3160 -1230
rect 3440 -1150 3480 -1140
rect 3440 -1230 3445 -1150
rect 3475 -1230 3480 -1150
rect 3440 -1240 3480 -1230
rect 3760 -1150 3800 -1115
rect 3840 -1085 4040 -1080
rect 3840 -1115 3850 -1085
rect 4030 -1115 4040 -1085
rect 3840 -1120 4040 -1115
rect 4160 -1085 4360 -1080
rect 4160 -1115 4170 -1085
rect 4350 -1115 4360 -1085
rect 4160 -1120 4360 -1115
rect 4400 -1085 4440 -950
rect 4720 -870 4760 -835
rect 4800 -805 5000 -800
rect 4800 -835 4810 -805
rect 4990 -835 5000 -805
rect 4800 -840 5000 -835
rect 4720 -950 4725 -870
rect 4755 -950 4760 -870
rect 4720 -960 4760 -950
rect 5040 -870 5080 -860
rect 5040 -950 5045 -870
rect 5075 -950 5080 -870
rect 4400 -1115 4405 -1085
rect 4435 -1115 4440 -1085
rect 3760 -1230 3765 -1150
rect 3795 -1230 3800 -1150
rect 3760 -1240 3800 -1230
rect 4080 -1150 4120 -1140
rect 4080 -1230 4085 -1150
rect 4115 -1230 4120 -1150
rect 4080 -1240 4120 -1230
rect 4400 -1150 4440 -1115
rect 4480 -1085 4680 -1080
rect 4480 -1115 4490 -1085
rect 4670 -1115 4680 -1085
rect 4480 -1120 4680 -1115
rect 4800 -1085 5000 -1080
rect 4800 -1115 4810 -1085
rect 4990 -1115 5000 -1085
rect 4800 -1120 5000 -1115
rect 5040 -1085 5080 -950
rect 5040 -1115 5045 -1085
rect 5075 -1115 5080 -1085
rect 4400 -1230 4405 -1150
rect 4435 -1230 4440 -1150
rect 4400 -1240 4440 -1230
rect 4720 -1150 4760 -1140
rect 4720 -1230 4725 -1150
rect 4755 -1230 4760 -1150
rect 4720 -1240 4760 -1230
rect 5040 -1150 5080 -1115
rect 5040 -1230 5045 -1150
rect 5075 -1230 5080 -1150
rect 5040 -1240 5080 -1230
rect -80 -1350 -40 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 -40 -1350
rect -80 -1440 -40 -1430
rect 240 -1350 280 -1340
rect 240 -1430 245 -1350
rect 275 -1430 280 -1350
rect 240 -1440 280 -1430
rect 560 -1350 600 -1340
rect 560 -1430 565 -1350
rect 595 -1430 600 -1350
rect 560 -1440 600 -1430
rect 880 -1350 920 -1340
rect 880 -1430 885 -1350
rect 915 -1430 920 -1350
rect 880 -1440 920 -1430
rect 1200 -1350 1240 -1340
rect 1200 -1430 1205 -1350
rect 1235 -1430 1240 -1350
rect 1200 -1440 1240 -1430
rect 1520 -1350 1560 -1340
rect 1520 -1430 1525 -1350
rect 1555 -1430 1560 -1350
rect 1520 -1440 1560 -1430
rect 1840 -1350 1880 -1340
rect 1840 -1430 1845 -1350
rect 1875 -1430 1880 -1350
rect 1840 -1440 1880 -1430
rect 2160 -1350 2200 -1340
rect 2160 -1430 2165 -1350
rect 2195 -1430 2200 -1350
rect 2160 -1440 2200 -1430
rect 2480 -1350 2520 -1340
rect 2480 -1430 2485 -1350
rect 2515 -1430 2520 -1350
rect 2480 -1440 2520 -1430
rect 2800 -1350 2840 -1340
rect 2800 -1430 2805 -1350
rect 2835 -1430 2840 -1350
rect 2800 -1440 2840 -1430
rect 3120 -1350 3160 -1340
rect 3120 -1430 3125 -1350
rect 3155 -1430 3160 -1350
rect 3120 -1440 3160 -1430
rect 3440 -1350 3480 -1340
rect 3440 -1430 3445 -1350
rect 3475 -1430 3480 -1350
rect 3440 -1440 3480 -1430
rect 3760 -1350 3800 -1340
rect 3760 -1430 3765 -1350
rect 3795 -1430 3800 -1350
rect 3760 -1440 3800 -1430
rect 4080 -1350 4120 -1340
rect 4080 -1430 4085 -1350
rect 4115 -1430 4120 -1350
rect 4080 -1440 4120 -1430
rect 4400 -1350 4440 -1340
rect 4400 -1430 4405 -1350
rect 4435 -1430 4440 -1350
rect 4400 -1440 4440 -1430
rect 4720 -1350 4760 -1340
rect 4720 -1430 4725 -1350
rect 4755 -1430 4760 -1350
rect 4720 -1440 4760 -1430
rect 5040 -1350 5080 -1340
rect 5040 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5040 -1440 5080 -1430
<< via1 >>
rect 10 -835 190 -805
rect 245 -835 275 -805
rect 330 -835 510 -805
rect 650 -835 830 -805
rect 885 -835 915 -805
rect -75 -1115 -45 -1085
rect 10 -1115 190 -1085
rect 330 -1115 510 -1085
rect 970 -835 1150 -805
rect 1290 -835 1470 -805
rect 1525 -835 1555 -805
rect 565 -1115 595 -1085
rect 650 -1115 830 -1085
rect 970 -1115 1150 -1085
rect 1610 -835 1790 -805
rect 1930 -835 2110 -805
rect 2165 -835 2195 -805
rect 1205 -1115 1235 -1085
rect 1290 -1115 1470 -1085
rect 1610 -1115 1790 -1085
rect 2250 -835 2430 -805
rect 2570 -835 2750 -805
rect 2805 -835 2835 -805
rect 1845 -1115 1875 -1085
rect 1930 -1115 2110 -1085
rect 2250 -1115 2430 -1085
rect 2890 -835 3070 -805
rect 3210 -835 3390 -805
rect 3445 -835 3475 -805
rect 2485 -1115 2515 -1085
rect 2570 -1115 2750 -1085
rect 2890 -1115 3070 -1085
rect 3530 -835 3710 -805
rect 3850 -835 4030 -805
rect 4085 -835 4115 -805
rect 3125 -1115 3155 -1085
rect 3210 -1115 3390 -1085
rect 3530 -1115 3710 -1085
rect 4170 -835 4350 -805
rect 4490 -835 4670 -805
rect 4725 -835 4755 -805
rect 3765 -1115 3795 -1085
rect 3850 -1115 4030 -1085
rect 4170 -1115 4350 -1085
rect 4810 -835 4990 -805
rect 4405 -1115 4435 -1085
rect 4490 -1115 4670 -1085
rect 4810 -1115 4990 -1085
rect 5045 -1115 5075 -1085
rect -75 -1430 -45 -1360
rect 1205 -1430 1235 -1360
rect 2485 -1430 2515 -1360
rect 3765 -1430 3795 -1360
rect 5045 -1430 5075 -1360
<< metal2 >>
rect -240 -725 5240 -720
rect -240 -755 -235 -725
rect -205 -755 -155 -725
rect -125 -755 -75 -725
rect -45 -755 5 -725
rect 35 -755 85 -725
rect 115 -755 165 -725
rect 195 -755 245 -725
rect 275 -755 325 -725
rect 355 -755 405 -725
rect 435 -755 485 -725
rect 515 -755 565 -725
rect 595 -755 645 -725
rect 675 -755 725 -725
rect 755 -755 805 -725
rect 835 -755 885 -725
rect 915 -755 965 -725
rect 995 -755 1045 -725
rect 1075 -755 1125 -725
rect 1155 -755 1205 -725
rect 1235 -755 1285 -725
rect 1315 -755 1365 -725
rect 1395 -755 1445 -725
rect 1475 -755 1525 -725
rect 1555 -755 1605 -725
rect 1635 -755 1685 -725
rect 1715 -755 1765 -725
rect 1795 -755 1845 -725
rect 1875 -755 1925 -725
rect 1955 -755 2005 -725
rect 2035 -755 2085 -725
rect 2115 -755 2165 -725
rect 2195 -755 2245 -725
rect 2275 -755 2325 -725
rect 2355 -755 2405 -725
rect 2435 -755 2485 -725
rect 2515 -755 2565 -725
rect 2595 -755 2645 -725
rect 2675 -755 2725 -725
rect 2755 -755 2805 -725
rect 2835 -755 2885 -725
rect 2915 -755 2965 -725
rect 2995 -755 3045 -725
rect 3075 -755 3125 -725
rect 3155 -755 3205 -725
rect 3235 -755 3285 -725
rect 3315 -755 3365 -725
rect 3395 -755 3445 -725
rect 3475 -755 3525 -725
rect 3555 -755 3605 -725
rect 3635 -755 3685 -725
rect 3715 -755 3765 -725
rect 3795 -755 3845 -725
rect 3875 -755 3925 -725
rect 3955 -755 4005 -725
rect 4035 -755 4085 -725
rect 4115 -755 4165 -725
rect 4195 -755 4245 -725
rect 4275 -755 4325 -725
rect 4355 -755 4405 -725
rect 4435 -755 4485 -725
rect 4515 -755 4565 -725
rect 4595 -755 4645 -725
rect 4675 -755 4725 -725
rect 4755 -755 4805 -725
rect 4835 -755 4885 -725
rect 4915 -755 4965 -725
rect 4995 -755 5045 -725
rect 5075 -755 5125 -725
rect 5155 -755 5205 -725
rect 5235 -755 5240 -725
rect -240 -760 5240 -755
rect -240 -805 5240 -800
rect -240 -835 10 -805
rect 190 -835 245 -805
rect 275 -835 330 -805
rect 510 -835 650 -805
rect 830 -835 885 -805
rect 915 -835 970 -805
rect 1150 -835 1290 -805
rect 1470 -835 1525 -805
rect 1555 -835 1610 -805
rect 1790 -835 1930 -805
rect 2110 -835 2165 -805
rect 2195 -835 2250 -805
rect 2430 -835 2570 -805
rect 2750 -835 2805 -805
rect 2835 -835 2890 -805
rect 3070 -835 3210 -805
rect 3390 -835 3445 -805
rect 3475 -835 3530 -805
rect 3710 -835 3850 -805
rect 4030 -835 4085 -805
rect 4115 -835 4170 -805
rect 4350 -835 4490 -805
rect 4670 -835 4725 -805
rect 4755 -835 4810 -805
rect 4990 -835 5240 -805
rect -240 -840 5240 -835
rect -240 -885 5240 -880
rect -240 -915 -235 -885
rect -205 -915 -155 -885
rect -125 -915 -75 -885
rect -45 -915 5 -885
rect 35 -915 85 -885
rect 115 -915 165 -885
rect 195 -915 245 -885
rect 275 -915 325 -885
rect 355 -915 405 -885
rect 435 -915 485 -885
rect 515 -915 565 -885
rect 595 -915 645 -885
rect 675 -915 725 -885
rect 755 -915 805 -885
rect 835 -915 885 -885
rect 915 -915 965 -885
rect 995 -915 1045 -885
rect 1075 -915 1125 -885
rect 1155 -915 1205 -885
rect 1235 -915 1285 -885
rect 1315 -915 1365 -885
rect 1395 -915 1445 -885
rect 1475 -915 1525 -885
rect 1555 -915 1605 -885
rect 1635 -915 1685 -885
rect 1715 -915 1765 -885
rect 1795 -915 1845 -885
rect 1875 -915 1925 -885
rect 1955 -915 2005 -885
rect 2035 -915 2085 -885
rect 2115 -915 2165 -885
rect 2195 -915 2245 -885
rect 2275 -915 2325 -885
rect 2355 -915 2405 -885
rect 2435 -915 2485 -885
rect 2515 -915 2565 -885
rect 2595 -915 2645 -885
rect 2675 -915 2725 -885
rect 2755 -915 2805 -885
rect 2835 -915 2885 -885
rect 2915 -915 2965 -885
rect 2995 -915 3045 -885
rect 3075 -915 3125 -885
rect 3155 -915 3205 -885
rect 3235 -915 3285 -885
rect 3315 -915 3365 -885
rect 3395 -915 3445 -885
rect 3475 -915 3525 -885
rect 3555 -915 3605 -885
rect 3635 -915 3685 -885
rect 3715 -915 3765 -885
rect 3795 -915 3845 -885
rect 3875 -915 3925 -885
rect 3955 -915 4005 -885
rect 4035 -915 4085 -885
rect 4115 -915 4165 -885
rect 4195 -915 4245 -885
rect 4275 -915 4325 -885
rect 4355 -915 4405 -885
rect 4435 -915 4485 -885
rect 4515 -915 4565 -885
rect 4595 -915 4645 -885
rect 4675 -915 4725 -885
rect 4755 -915 4805 -885
rect 4835 -915 4885 -885
rect 4915 -915 4965 -885
rect 4995 -915 5045 -885
rect 5075 -915 5125 -885
rect 5155 -915 5205 -885
rect 5235 -915 5240 -885
rect -240 -920 5240 -915
rect -240 -1005 5240 -1000
rect -240 -1035 -235 -1005
rect -205 -1035 -155 -1005
rect -125 -1035 -75 -1005
rect -45 -1035 5 -1005
rect 35 -1035 85 -1005
rect 115 -1035 165 -1005
rect 195 -1035 245 -1005
rect 275 -1035 325 -1005
rect 355 -1035 405 -1005
rect 435 -1035 485 -1005
rect 515 -1035 565 -1005
rect 595 -1035 645 -1005
rect 675 -1035 725 -1005
rect 755 -1035 805 -1005
rect 835 -1035 885 -1005
rect 915 -1035 965 -1005
rect 995 -1035 1045 -1005
rect 1075 -1035 1125 -1005
rect 1155 -1035 1205 -1005
rect 1235 -1035 1285 -1005
rect 1315 -1035 1365 -1005
rect 1395 -1035 1445 -1005
rect 1475 -1035 1525 -1005
rect 1555 -1035 1605 -1005
rect 1635 -1035 1685 -1005
rect 1715 -1035 1765 -1005
rect 1795 -1035 1845 -1005
rect 1875 -1035 1925 -1005
rect 1955 -1035 2005 -1005
rect 2035 -1035 2085 -1005
rect 2115 -1035 2165 -1005
rect 2195 -1035 2245 -1005
rect 2275 -1035 2325 -1005
rect 2355 -1035 2405 -1005
rect 2435 -1035 2485 -1005
rect 2515 -1035 2565 -1005
rect 2595 -1035 2645 -1005
rect 2675 -1035 2725 -1005
rect 2755 -1035 2805 -1005
rect 2835 -1035 2885 -1005
rect 2915 -1035 2965 -1005
rect 2995 -1035 3045 -1005
rect 3075 -1035 3125 -1005
rect 3155 -1035 3205 -1005
rect 3235 -1035 3285 -1005
rect 3315 -1035 3365 -1005
rect 3395 -1035 3445 -1005
rect 3475 -1035 3525 -1005
rect 3555 -1035 3605 -1005
rect 3635 -1035 3685 -1005
rect 3715 -1035 3765 -1005
rect 3795 -1035 3845 -1005
rect 3875 -1035 3925 -1005
rect 3955 -1035 4005 -1005
rect 4035 -1035 4085 -1005
rect 4115 -1035 4165 -1005
rect 4195 -1035 4245 -1005
rect 4275 -1035 4325 -1005
rect 4355 -1035 4405 -1005
rect 4435 -1035 4485 -1005
rect 4515 -1035 4565 -1005
rect 4595 -1035 4645 -1005
rect 4675 -1035 4725 -1005
rect 4755 -1035 4805 -1005
rect 4835 -1035 4885 -1005
rect 4915 -1035 4965 -1005
rect 4995 -1035 5045 -1005
rect 5075 -1035 5125 -1005
rect 5155 -1035 5240 -1005
rect -240 -1040 5240 -1035
rect -240 -1085 5240 -1080
rect -240 -1115 -75 -1085
rect -45 -1115 10 -1085
rect 190 -1115 330 -1085
rect 510 -1115 565 -1085
rect 595 -1115 650 -1085
rect 830 -1115 970 -1085
rect 1150 -1115 1205 -1085
rect 1235 -1115 1290 -1085
rect 1470 -1115 1610 -1085
rect 1790 -1115 1845 -1085
rect 1875 -1115 1930 -1085
rect 2110 -1115 2250 -1085
rect 2430 -1115 2485 -1085
rect 2515 -1115 2570 -1085
rect 2750 -1115 2890 -1085
rect 3070 -1115 3125 -1085
rect 3155 -1115 3210 -1085
rect 3390 -1115 3530 -1085
rect 3710 -1115 3765 -1085
rect 3795 -1115 3850 -1085
rect 4030 -1115 4170 -1085
rect 4350 -1115 4405 -1085
rect 4435 -1115 4490 -1085
rect 4670 -1115 4810 -1085
rect 4990 -1115 5045 -1085
rect 5075 -1115 5240 -1085
rect -240 -1120 5240 -1115
rect -240 -1165 5240 -1160
rect -240 -1195 -235 -1165
rect -205 -1195 -155 -1165
rect -125 -1195 -75 -1165
rect -45 -1195 5 -1165
rect 35 -1195 85 -1165
rect 115 -1195 165 -1165
rect 195 -1195 245 -1165
rect 275 -1195 325 -1165
rect 355 -1195 405 -1165
rect 435 -1195 485 -1165
rect 515 -1195 565 -1165
rect 595 -1195 645 -1165
rect 675 -1195 725 -1165
rect 755 -1195 805 -1165
rect 835 -1195 885 -1165
rect 915 -1195 965 -1165
rect 995 -1195 1045 -1165
rect 1075 -1195 1125 -1165
rect 1155 -1195 1205 -1165
rect 1235 -1195 1285 -1165
rect 1315 -1195 1365 -1165
rect 1395 -1195 1445 -1165
rect 1475 -1195 1525 -1165
rect 1555 -1195 1605 -1165
rect 1635 -1195 1685 -1165
rect 1715 -1195 1765 -1165
rect 1795 -1195 1845 -1165
rect 1875 -1195 1925 -1165
rect 1955 -1195 2005 -1165
rect 2035 -1195 2085 -1165
rect 2115 -1195 2165 -1165
rect 2195 -1195 2245 -1165
rect 2275 -1195 2325 -1165
rect 2355 -1195 2405 -1165
rect 2435 -1195 2485 -1165
rect 2515 -1195 2565 -1165
rect 2595 -1195 2645 -1165
rect 2675 -1195 2725 -1165
rect 2755 -1195 2805 -1165
rect 2835 -1195 2885 -1165
rect 2915 -1195 2965 -1165
rect 2995 -1195 3045 -1165
rect 3075 -1195 3125 -1165
rect 3155 -1195 3205 -1165
rect 3235 -1195 3285 -1165
rect 3315 -1195 3365 -1165
rect 3395 -1195 3445 -1165
rect 3475 -1195 3525 -1165
rect 3555 -1195 3605 -1165
rect 3635 -1195 3685 -1165
rect 3715 -1195 3765 -1165
rect 3795 -1195 3845 -1165
rect 3875 -1195 3925 -1165
rect 3955 -1195 4005 -1165
rect 4035 -1195 4085 -1165
rect 4115 -1195 4165 -1165
rect 4195 -1195 4245 -1165
rect 4275 -1195 4325 -1165
rect 4355 -1195 4405 -1165
rect 4435 -1195 4485 -1165
rect 4515 -1195 4565 -1165
rect 4595 -1195 4645 -1165
rect 4675 -1195 4725 -1165
rect 4755 -1195 4805 -1165
rect 4835 -1195 4885 -1165
rect 4915 -1195 4965 -1165
rect 4995 -1195 5045 -1165
rect 5075 -1195 5125 -1165
rect 5155 -1195 5205 -1165
rect 5235 -1195 5240 -1165
rect -240 -1200 5240 -1195
rect -80 -1430 -75 -1360
rect -45 -1430 -40 -1360
rect -80 -1440 -40 -1430
rect 1200 -1430 1205 -1360
rect 1235 -1430 1240 -1360
rect 1200 -1440 1240 -1430
rect 2480 -1430 2485 -1360
rect 2515 -1430 2520 -1360
rect 2480 -1440 2520 -1430
rect 3760 -1430 3765 -1360
rect 3795 -1430 3800 -1360
rect 3760 -1440 3800 -1430
rect 5040 -1430 5045 -1360
rect 5075 -1430 5080 -1360
rect 5040 -1440 5080 -1430
<< via2 >>
rect -235 -755 -205 -725
rect -155 -755 -125 -725
rect -75 -755 -45 -725
rect 5 -755 35 -725
rect 85 -755 115 -725
rect 165 -755 195 -725
rect 245 -755 275 -725
rect 325 -755 355 -725
rect 405 -755 435 -725
rect 485 -755 515 -725
rect 565 -755 595 -725
rect 645 -755 675 -725
rect 725 -755 755 -725
rect 805 -755 835 -725
rect 885 -755 915 -725
rect 965 -755 995 -725
rect 1045 -755 1075 -725
rect 1125 -755 1155 -725
rect 1205 -755 1235 -725
rect 1285 -755 1315 -725
rect 1365 -755 1395 -725
rect 1445 -755 1475 -725
rect 1525 -755 1555 -725
rect 1605 -755 1635 -725
rect 1685 -755 1715 -725
rect 1765 -755 1795 -725
rect 1845 -755 1875 -725
rect 1925 -755 1955 -725
rect 2005 -755 2035 -725
rect 2085 -755 2115 -725
rect 2165 -755 2195 -725
rect 2245 -755 2275 -725
rect 2325 -755 2355 -725
rect 2405 -755 2435 -725
rect 2485 -755 2515 -725
rect 2565 -755 2595 -725
rect 2645 -755 2675 -725
rect 2725 -755 2755 -725
rect 2805 -755 2835 -725
rect 2885 -755 2915 -725
rect 2965 -755 2995 -725
rect 3045 -755 3075 -725
rect 3125 -755 3155 -725
rect 3205 -755 3235 -725
rect 3285 -755 3315 -725
rect 3365 -755 3395 -725
rect 3445 -755 3475 -725
rect 3525 -755 3555 -725
rect 3605 -755 3635 -725
rect 3685 -755 3715 -725
rect 3765 -755 3795 -725
rect 3845 -755 3875 -725
rect 3925 -755 3955 -725
rect 4005 -755 4035 -725
rect 4085 -755 4115 -725
rect 4165 -755 4195 -725
rect 4245 -755 4275 -725
rect 4325 -755 4355 -725
rect 4405 -755 4435 -725
rect 4485 -755 4515 -725
rect 4565 -755 4595 -725
rect 4645 -755 4675 -725
rect 4725 -755 4755 -725
rect 4805 -755 4835 -725
rect 4885 -755 4915 -725
rect 4965 -755 4995 -725
rect 5045 -755 5075 -725
rect 5125 -755 5155 -725
rect 5205 -755 5235 -725
rect -235 -915 -205 -885
rect -155 -915 -125 -885
rect -75 -915 -45 -885
rect 5 -915 35 -885
rect 85 -915 115 -885
rect 165 -915 195 -885
rect 245 -915 275 -885
rect 325 -915 355 -885
rect 405 -915 435 -885
rect 485 -915 515 -885
rect 565 -915 595 -885
rect 645 -915 675 -885
rect 725 -915 755 -885
rect 805 -915 835 -885
rect 885 -915 915 -885
rect 965 -915 995 -885
rect 1045 -915 1075 -885
rect 1125 -915 1155 -885
rect 1205 -915 1235 -885
rect 1285 -915 1315 -885
rect 1365 -915 1395 -885
rect 1445 -915 1475 -885
rect 1525 -915 1555 -885
rect 1605 -915 1635 -885
rect 1685 -915 1715 -885
rect 1765 -915 1795 -885
rect 1845 -915 1875 -885
rect 1925 -915 1955 -885
rect 2005 -915 2035 -885
rect 2085 -915 2115 -885
rect 2165 -915 2195 -885
rect 2245 -915 2275 -885
rect 2325 -915 2355 -885
rect 2405 -915 2435 -885
rect 2485 -915 2515 -885
rect 2565 -915 2595 -885
rect 2645 -915 2675 -885
rect 2725 -915 2755 -885
rect 2805 -915 2835 -885
rect 2885 -915 2915 -885
rect 2965 -915 2995 -885
rect 3045 -915 3075 -885
rect 3125 -915 3155 -885
rect 3205 -915 3235 -885
rect 3285 -915 3315 -885
rect 3365 -915 3395 -885
rect 3445 -915 3475 -885
rect 3525 -915 3555 -885
rect 3605 -915 3635 -885
rect 3685 -915 3715 -885
rect 3765 -915 3795 -885
rect 3845 -915 3875 -885
rect 3925 -915 3955 -885
rect 4005 -915 4035 -885
rect 4085 -915 4115 -885
rect 4165 -915 4195 -885
rect 4245 -915 4275 -885
rect 4325 -915 4355 -885
rect 4405 -915 4435 -885
rect 4485 -915 4515 -885
rect 4565 -915 4595 -885
rect 4645 -915 4675 -885
rect 4725 -915 4755 -885
rect 4805 -915 4835 -885
rect 4885 -915 4915 -885
rect 4965 -915 4995 -885
rect 5045 -915 5075 -885
rect 5125 -915 5155 -885
rect 5205 -915 5235 -885
rect -235 -1035 -205 -1005
rect -155 -1035 -125 -1005
rect -75 -1035 -45 -1005
rect 5 -1035 35 -1005
rect 85 -1035 115 -1005
rect 165 -1035 195 -1005
rect 245 -1035 275 -1005
rect 325 -1035 355 -1005
rect 405 -1035 435 -1005
rect 485 -1035 515 -1005
rect 565 -1035 595 -1005
rect 645 -1035 675 -1005
rect 725 -1035 755 -1005
rect 805 -1035 835 -1005
rect 885 -1035 915 -1005
rect 965 -1035 995 -1005
rect 1045 -1035 1075 -1005
rect 1125 -1035 1155 -1005
rect 1205 -1035 1235 -1005
rect 1285 -1035 1315 -1005
rect 1365 -1035 1395 -1005
rect 1445 -1035 1475 -1005
rect 1525 -1035 1555 -1005
rect 1605 -1035 1635 -1005
rect 1685 -1035 1715 -1005
rect 1765 -1035 1795 -1005
rect 1845 -1035 1875 -1005
rect 1925 -1035 1955 -1005
rect 2005 -1035 2035 -1005
rect 2085 -1035 2115 -1005
rect 2165 -1035 2195 -1005
rect 2245 -1035 2275 -1005
rect 2325 -1035 2355 -1005
rect 2405 -1035 2435 -1005
rect 2485 -1035 2515 -1005
rect 2565 -1035 2595 -1005
rect 2645 -1035 2675 -1005
rect 2725 -1035 2755 -1005
rect 2805 -1035 2835 -1005
rect 2885 -1035 2915 -1005
rect 2965 -1035 2995 -1005
rect 3045 -1035 3075 -1005
rect 3125 -1035 3155 -1005
rect 3205 -1035 3235 -1005
rect 3285 -1035 3315 -1005
rect 3365 -1035 3395 -1005
rect 3445 -1035 3475 -1005
rect 3525 -1035 3555 -1005
rect 3605 -1035 3635 -1005
rect 3685 -1035 3715 -1005
rect 3765 -1035 3795 -1005
rect 3845 -1035 3875 -1005
rect 3925 -1035 3955 -1005
rect 4005 -1035 4035 -1005
rect 4085 -1035 4115 -1005
rect 4165 -1035 4195 -1005
rect 4245 -1035 4275 -1005
rect 4325 -1035 4355 -1005
rect 4405 -1035 4435 -1005
rect 4485 -1035 4515 -1005
rect 4565 -1035 4595 -1005
rect 4645 -1035 4675 -1005
rect 4725 -1035 4755 -1005
rect 4805 -1035 4835 -1005
rect 4885 -1035 4915 -1005
rect 4965 -1035 4995 -1005
rect 5045 -1035 5075 -1005
rect 5125 -1035 5155 -1005
rect -235 -1195 -205 -1165
rect -155 -1195 -125 -1165
rect -75 -1195 -45 -1165
rect 5 -1195 35 -1165
rect 85 -1195 115 -1165
rect 165 -1195 195 -1165
rect 245 -1195 275 -1165
rect 325 -1195 355 -1165
rect 405 -1195 435 -1165
rect 485 -1195 515 -1165
rect 565 -1195 595 -1165
rect 645 -1195 675 -1165
rect 725 -1195 755 -1165
rect 805 -1195 835 -1165
rect 885 -1195 915 -1165
rect 965 -1195 995 -1165
rect 1045 -1195 1075 -1165
rect 1125 -1195 1155 -1165
rect 1205 -1195 1235 -1165
rect 1285 -1195 1315 -1165
rect 1365 -1195 1395 -1165
rect 1445 -1195 1475 -1165
rect 1525 -1195 1555 -1165
rect 1605 -1195 1635 -1165
rect 1685 -1195 1715 -1165
rect 1765 -1195 1795 -1165
rect 1845 -1195 1875 -1165
rect 1925 -1195 1955 -1165
rect 2005 -1195 2035 -1165
rect 2085 -1195 2115 -1165
rect 2165 -1195 2195 -1165
rect 2245 -1195 2275 -1165
rect 2325 -1195 2355 -1165
rect 2405 -1195 2435 -1165
rect 2485 -1195 2515 -1165
rect 2565 -1195 2595 -1165
rect 2645 -1195 2675 -1165
rect 2725 -1195 2755 -1165
rect 2805 -1195 2835 -1165
rect 2885 -1195 2915 -1165
rect 2965 -1195 2995 -1165
rect 3045 -1195 3075 -1165
rect 3125 -1195 3155 -1165
rect 3205 -1195 3235 -1165
rect 3285 -1195 3315 -1165
rect 3365 -1195 3395 -1165
rect 3445 -1195 3475 -1165
rect 3525 -1195 3555 -1165
rect 3605 -1195 3635 -1165
rect 3685 -1195 3715 -1165
rect 3765 -1195 3795 -1165
rect 3845 -1195 3875 -1165
rect 3925 -1195 3955 -1165
rect 4005 -1195 4035 -1165
rect 4085 -1195 4115 -1165
rect 4165 -1195 4195 -1165
rect 4245 -1195 4275 -1165
rect 4325 -1195 4355 -1165
rect 4405 -1195 4435 -1165
rect 4485 -1195 4515 -1165
rect 4565 -1195 4595 -1165
rect 4645 -1195 4675 -1165
rect 4725 -1195 4755 -1165
rect 4805 -1195 4835 -1165
rect 4885 -1195 4915 -1165
rect 4965 -1195 4995 -1165
rect 5045 -1195 5075 -1165
rect 5125 -1195 5155 -1165
rect 5205 -1195 5235 -1165
rect -75 -1430 -45 -1360
rect 1205 -1430 1235 -1360
rect 2485 -1430 2515 -1360
rect 3765 -1430 3795 -1360
rect 5045 -1430 5075 -1360
<< metal3 >>
rect -240 -725 -200 -720
rect -240 -755 -235 -725
rect -205 -755 -200 -725
rect -240 -885 -200 -755
rect -240 -915 -235 -885
rect -205 -915 -200 -885
rect -240 -1005 -200 -915
rect -240 -1035 -235 -1005
rect -205 -1035 -200 -1005
rect -240 -1165 -200 -1035
rect -240 -1195 -235 -1165
rect -205 -1195 -200 -1165
rect -240 -1360 -200 -1195
rect -160 -725 -120 -720
rect -160 -755 -155 -725
rect -125 -755 -120 -725
rect -160 -885 -120 -755
rect -160 -915 -155 -885
rect -125 -915 -120 -885
rect -160 -1005 -120 -915
rect -160 -1035 -155 -1005
rect -125 -1035 -120 -1005
rect -160 -1165 -120 -1035
rect -160 -1195 -155 -1165
rect -125 -1195 -120 -1165
rect -160 -1360 -120 -1195
rect -80 -725 -40 -720
rect -80 -755 -75 -725
rect -45 -755 -40 -725
rect -80 -885 -40 -755
rect -80 -915 -75 -885
rect -45 -915 -40 -885
rect -80 -1005 -40 -915
rect -80 -1035 -75 -1005
rect -45 -1035 -40 -1005
rect -80 -1165 -40 -1035
rect -80 -1195 -75 -1165
rect -45 -1195 -40 -1165
rect -80 -1349 -40 -1195
rect -80 -1431 -76 -1349
rect -44 -1431 -40 -1349
rect 0 -725 40 -720
rect 0 -755 5 -725
rect 35 -755 40 -725
rect 0 -885 40 -755
rect 0 -915 5 -885
rect 35 -915 40 -885
rect 0 -1005 40 -915
rect 0 -1035 5 -1005
rect 35 -1035 40 -1005
rect 0 -1165 40 -1035
rect 0 -1195 5 -1165
rect 35 -1195 40 -1165
rect 0 -1360 40 -1195
rect 80 -725 120 -720
rect 80 -755 85 -725
rect 115 -755 120 -725
rect 80 -885 120 -755
rect 80 -915 85 -885
rect 115 -915 120 -885
rect 80 -1005 120 -915
rect 80 -1035 85 -1005
rect 115 -1035 120 -1005
rect 80 -1165 120 -1035
rect 80 -1195 85 -1165
rect 115 -1195 120 -1165
rect 80 -1360 120 -1195
rect 160 -725 200 -720
rect 160 -755 165 -725
rect 195 -755 200 -725
rect 160 -885 200 -755
rect 160 -915 165 -885
rect 195 -915 200 -885
rect 160 -1005 200 -915
rect 160 -1035 165 -1005
rect 195 -1035 200 -1005
rect 160 -1165 200 -1035
rect 160 -1195 165 -1165
rect 195 -1195 200 -1165
rect 160 -1360 200 -1195
rect 240 -725 280 -720
rect 240 -755 245 -725
rect 275 -755 280 -725
rect 240 -885 280 -755
rect 240 -915 245 -885
rect 275 -915 280 -885
rect 240 -1005 280 -915
rect 240 -1035 245 -1005
rect 275 -1035 280 -1005
rect 240 -1165 280 -1035
rect 240 -1195 245 -1165
rect 275 -1195 280 -1165
rect 240 -1360 280 -1195
rect 320 -725 360 -720
rect 320 -755 325 -725
rect 355 -755 360 -725
rect 320 -885 360 -755
rect 320 -915 325 -885
rect 355 -915 360 -885
rect 320 -1005 360 -915
rect 320 -1035 325 -1005
rect 355 -1035 360 -1005
rect 320 -1165 360 -1035
rect 320 -1195 325 -1165
rect 355 -1195 360 -1165
rect 320 -1360 360 -1195
rect 400 -725 440 -720
rect 400 -755 405 -725
rect 435 -755 440 -725
rect 400 -885 440 -755
rect 400 -915 405 -885
rect 435 -915 440 -885
rect 400 -1005 440 -915
rect 400 -1035 405 -1005
rect 435 -1035 440 -1005
rect 400 -1165 440 -1035
rect 400 -1195 405 -1165
rect 435 -1195 440 -1165
rect 400 -1360 440 -1195
rect 480 -725 520 -720
rect 480 -755 485 -725
rect 515 -755 520 -725
rect 480 -885 520 -755
rect 480 -915 485 -885
rect 515 -915 520 -885
rect 480 -1005 520 -915
rect 560 -725 600 -720
rect 560 -755 565 -725
rect 595 -755 600 -725
rect 560 -885 600 -755
rect 560 -915 565 -885
rect 595 -915 600 -885
rect 560 -920 600 -915
rect 640 -725 680 -720
rect 640 -755 645 -725
rect 675 -755 680 -725
rect 640 -885 680 -755
rect 640 -915 645 -885
rect 675 -915 680 -885
rect 480 -1035 485 -1005
rect 515 -1035 520 -1005
rect 480 -1165 520 -1035
rect 480 -1195 485 -1165
rect 515 -1195 520 -1165
rect 480 -1360 520 -1195
rect 560 -1005 600 -960
rect 560 -1035 565 -1005
rect 595 -1035 600 -1005
rect 560 -1165 600 -1035
rect 560 -1195 565 -1165
rect 595 -1195 600 -1165
rect 560 -1200 600 -1195
rect 640 -1005 680 -915
rect 640 -1035 645 -1005
rect 675 -1035 680 -1005
rect 640 -1165 680 -1035
rect 640 -1195 645 -1165
rect 675 -1195 680 -1165
rect 640 -1360 680 -1195
rect 720 -725 760 -720
rect 720 -755 725 -725
rect 755 -755 760 -725
rect 720 -885 760 -755
rect 720 -915 725 -885
rect 755 -915 760 -885
rect 720 -1005 760 -915
rect 720 -1035 725 -1005
rect 755 -1035 760 -1005
rect 720 -1165 760 -1035
rect 720 -1195 725 -1165
rect 755 -1195 760 -1165
rect 720 -1360 760 -1195
rect 800 -725 840 -720
rect 800 -755 805 -725
rect 835 -755 840 -725
rect 800 -885 840 -755
rect 800 -915 805 -885
rect 835 -915 840 -885
rect 800 -1005 840 -915
rect 800 -1035 805 -1005
rect 835 -1035 840 -1005
rect 800 -1165 840 -1035
rect 800 -1195 805 -1165
rect 835 -1195 840 -1165
rect 800 -1360 840 -1195
rect 880 -725 920 -720
rect 880 -755 885 -725
rect 915 -755 920 -725
rect 880 -885 920 -755
rect 880 -915 885 -885
rect 915 -915 920 -885
rect 880 -1005 920 -915
rect 880 -1035 885 -1005
rect 915 -1035 920 -1005
rect 880 -1165 920 -1035
rect 880 -1195 885 -1165
rect 915 -1195 920 -1165
rect 880 -1360 920 -1195
rect 960 -725 1000 -720
rect 960 -755 965 -725
rect 995 -755 1000 -725
rect 960 -885 1000 -755
rect 960 -915 965 -885
rect 995 -915 1000 -885
rect 960 -1005 1000 -915
rect 960 -1035 965 -1005
rect 995 -1035 1000 -1005
rect 960 -1165 1000 -1035
rect 960 -1195 965 -1165
rect 995 -1195 1000 -1165
rect 960 -1360 1000 -1195
rect 1040 -725 1080 -720
rect 1040 -755 1045 -725
rect 1075 -755 1080 -725
rect 1040 -885 1080 -755
rect 1040 -915 1045 -885
rect 1075 -915 1080 -885
rect 1040 -1005 1080 -915
rect 1040 -1035 1045 -1005
rect 1075 -1035 1080 -1005
rect 1040 -1165 1080 -1035
rect 1040 -1195 1045 -1165
rect 1075 -1195 1080 -1165
rect 1040 -1360 1080 -1195
rect 1120 -725 1160 -720
rect 1120 -755 1125 -725
rect 1155 -755 1160 -725
rect 1120 -885 1160 -755
rect 1120 -915 1125 -885
rect 1155 -915 1160 -885
rect 1120 -1005 1160 -915
rect 1200 -725 1240 -720
rect 1200 -755 1205 -725
rect 1235 -755 1240 -725
rect 1200 -885 1240 -755
rect 1200 -915 1205 -885
rect 1235 -915 1240 -885
rect 1200 -920 1240 -915
rect 1280 -725 1320 -720
rect 1280 -755 1285 -725
rect 1315 -755 1320 -725
rect 1280 -885 1320 -755
rect 1280 -915 1285 -885
rect 1315 -915 1320 -885
rect 1120 -1035 1125 -1005
rect 1155 -1035 1160 -1005
rect 1120 -1165 1160 -1035
rect 1120 -1195 1125 -1165
rect 1155 -1195 1160 -1165
rect 1120 -1360 1160 -1195
rect 1200 -1005 1240 -960
rect 1200 -1035 1205 -1005
rect 1235 -1035 1240 -1005
rect 1200 -1165 1240 -1035
rect 1200 -1195 1205 -1165
rect 1235 -1195 1240 -1165
rect 1200 -1200 1240 -1195
rect 1280 -1005 1320 -915
rect 1280 -1035 1285 -1005
rect 1315 -1035 1320 -1005
rect 1280 -1165 1320 -1035
rect 1280 -1195 1285 -1165
rect 1315 -1195 1320 -1165
rect 1200 -1349 1240 -1320
rect -80 -1440 -40 -1431
rect 1200 -1431 1204 -1349
rect 1236 -1431 1240 -1349
rect 1280 -1360 1320 -1195
rect 1360 -725 1400 -720
rect 1360 -755 1365 -725
rect 1395 -755 1400 -725
rect 1360 -885 1400 -755
rect 1360 -915 1365 -885
rect 1395 -915 1400 -885
rect 1360 -1005 1400 -915
rect 1360 -1035 1365 -1005
rect 1395 -1035 1400 -1005
rect 1360 -1165 1400 -1035
rect 1360 -1195 1365 -1165
rect 1395 -1195 1400 -1165
rect 1360 -1360 1400 -1195
rect 1440 -725 1480 -720
rect 1440 -755 1445 -725
rect 1475 -755 1480 -725
rect 1440 -885 1480 -755
rect 1440 -915 1445 -885
rect 1475 -915 1480 -885
rect 1440 -1005 1480 -915
rect 1440 -1035 1445 -1005
rect 1475 -1035 1480 -1005
rect 1440 -1165 1480 -1035
rect 1440 -1195 1445 -1165
rect 1475 -1195 1480 -1165
rect 1440 -1360 1480 -1195
rect 1520 -725 1560 -720
rect 1520 -755 1525 -725
rect 1555 -755 1560 -725
rect 1520 -885 1560 -755
rect 1520 -915 1525 -885
rect 1555 -915 1560 -885
rect 1520 -1005 1560 -915
rect 1520 -1035 1525 -1005
rect 1555 -1035 1560 -1005
rect 1520 -1165 1560 -1035
rect 1520 -1195 1525 -1165
rect 1555 -1195 1560 -1165
rect 1520 -1360 1560 -1195
rect 1600 -725 1640 -720
rect 1600 -755 1605 -725
rect 1635 -755 1640 -725
rect 1600 -885 1640 -755
rect 1600 -915 1605 -885
rect 1635 -915 1640 -885
rect 1600 -1005 1640 -915
rect 1600 -1035 1605 -1005
rect 1635 -1035 1640 -1005
rect 1600 -1165 1640 -1035
rect 1600 -1195 1605 -1165
rect 1635 -1195 1640 -1165
rect 1600 -1360 1640 -1195
rect 1680 -725 1720 -720
rect 1680 -755 1685 -725
rect 1715 -755 1720 -725
rect 1680 -885 1720 -755
rect 1680 -915 1685 -885
rect 1715 -915 1720 -885
rect 1680 -1005 1720 -915
rect 1680 -1035 1685 -1005
rect 1715 -1035 1720 -1005
rect 1680 -1165 1720 -1035
rect 1680 -1195 1685 -1165
rect 1715 -1195 1720 -1165
rect 1680 -1360 1720 -1195
rect 1760 -725 1800 -720
rect 1760 -755 1765 -725
rect 1795 -755 1800 -725
rect 1760 -885 1800 -755
rect 1760 -915 1765 -885
rect 1795 -915 1800 -885
rect 1760 -1005 1800 -915
rect 1840 -725 1880 -720
rect 1840 -755 1845 -725
rect 1875 -755 1880 -725
rect 1840 -885 1880 -755
rect 1840 -915 1845 -885
rect 1875 -915 1880 -885
rect 1840 -920 1880 -915
rect 1920 -725 1960 -720
rect 1920 -755 1925 -725
rect 1955 -755 1960 -725
rect 1920 -885 1960 -755
rect 1920 -915 1925 -885
rect 1955 -915 1960 -885
rect 1760 -1035 1765 -1005
rect 1795 -1035 1800 -1005
rect 1760 -1165 1800 -1035
rect 1760 -1195 1765 -1165
rect 1795 -1195 1800 -1165
rect 1760 -1360 1800 -1195
rect 1840 -1005 1880 -960
rect 1840 -1035 1845 -1005
rect 1875 -1035 1880 -1005
rect 1840 -1165 1880 -1035
rect 1840 -1195 1845 -1165
rect 1875 -1195 1880 -1165
rect 1840 -1200 1880 -1195
rect 1920 -1005 1960 -915
rect 1920 -1035 1925 -1005
rect 1955 -1035 1960 -1005
rect 1920 -1165 1960 -1035
rect 1920 -1195 1925 -1165
rect 1955 -1195 1960 -1165
rect 1920 -1360 1960 -1195
rect 2000 -725 2040 -720
rect 2000 -755 2005 -725
rect 2035 -755 2040 -725
rect 2000 -885 2040 -755
rect 2000 -915 2005 -885
rect 2035 -915 2040 -885
rect 2000 -1005 2040 -915
rect 2000 -1035 2005 -1005
rect 2035 -1035 2040 -1005
rect 2000 -1165 2040 -1035
rect 2000 -1195 2005 -1165
rect 2035 -1195 2040 -1165
rect 2000 -1360 2040 -1195
rect 2080 -725 2120 -720
rect 2080 -755 2085 -725
rect 2115 -755 2120 -725
rect 2080 -885 2120 -755
rect 2080 -915 2085 -885
rect 2115 -915 2120 -885
rect 2080 -1005 2120 -915
rect 2080 -1035 2085 -1005
rect 2115 -1035 2120 -1005
rect 2080 -1165 2120 -1035
rect 2080 -1195 2085 -1165
rect 2115 -1195 2120 -1165
rect 2080 -1360 2120 -1195
rect 2160 -725 2200 -720
rect 2160 -755 2165 -725
rect 2195 -755 2200 -725
rect 2160 -885 2200 -755
rect 2160 -915 2165 -885
rect 2195 -915 2200 -885
rect 2160 -1005 2200 -915
rect 2160 -1035 2165 -1005
rect 2195 -1035 2200 -1005
rect 2160 -1165 2200 -1035
rect 2160 -1195 2165 -1165
rect 2195 -1195 2200 -1165
rect 2160 -1360 2200 -1195
rect 2240 -725 2280 -720
rect 2240 -755 2245 -725
rect 2275 -755 2280 -725
rect 2240 -885 2280 -755
rect 2240 -915 2245 -885
rect 2275 -915 2280 -885
rect 2240 -1005 2280 -915
rect 2240 -1035 2245 -1005
rect 2275 -1035 2280 -1005
rect 2240 -1165 2280 -1035
rect 2240 -1195 2245 -1165
rect 2275 -1195 2280 -1165
rect 2240 -1360 2280 -1195
rect 2320 -725 2360 -720
rect 2320 -755 2325 -725
rect 2355 -755 2360 -725
rect 2320 -885 2360 -755
rect 2320 -915 2325 -885
rect 2355 -915 2360 -885
rect 2320 -1005 2360 -915
rect 2320 -1035 2325 -1005
rect 2355 -1035 2360 -1005
rect 2320 -1165 2360 -1035
rect 2320 -1195 2325 -1165
rect 2355 -1195 2360 -1165
rect 2320 -1360 2360 -1195
rect 2400 -725 2440 -720
rect 2400 -755 2405 -725
rect 2435 -755 2440 -725
rect 2400 -885 2440 -755
rect 2400 -915 2405 -885
rect 2435 -915 2440 -885
rect 2400 -1005 2440 -915
rect 2480 -725 2520 -720
rect 2480 -755 2485 -725
rect 2515 -755 2520 -725
rect 2480 -885 2520 -755
rect 2480 -915 2485 -885
rect 2515 -915 2520 -885
rect 2480 -920 2520 -915
rect 2560 -725 2600 -720
rect 2560 -755 2565 -725
rect 2595 -755 2600 -725
rect 2560 -885 2600 -755
rect 2560 -915 2565 -885
rect 2595 -915 2600 -885
rect 2400 -1035 2405 -1005
rect 2435 -1035 2440 -1005
rect 2400 -1165 2440 -1035
rect 2400 -1195 2405 -1165
rect 2435 -1195 2440 -1165
rect 2400 -1360 2440 -1195
rect 2480 -1005 2520 -960
rect 2480 -1035 2485 -1005
rect 2515 -1035 2520 -1005
rect 2480 -1165 2520 -1035
rect 2480 -1195 2485 -1165
rect 2515 -1195 2520 -1165
rect 2480 -1200 2520 -1195
rect 2560 -1005 2600 -915
rect 2560 -1035 2565 -1005
rect 2595 -1035 2600 -1005
rect 2560 -1165 2600 -1035
rect 2560 -1195 2565 -1165
rect 2595 -1195 2600 -1165
rect 2480 -1349 2520 -1320
rect 1200 -1440 1240 -1431
rect 2480 -1431 2484 -1349
rect 2516 -1431 2520 -1349
rect 2560 -1360 2600 -1195
rect 2640 -725 2680 -720
rect 2640 -755 2645 -725
rect 2675 -755 2680 -725
rect 2640 -885 2680 -755
rect 2640 -915 2645 -885
rect 2675 -915 2680 -885
rect 2640 -1005 2680 -915
rect 2640 -1035 2645 -1005
rect 2675 -1035 2680 -1005
rect 2640 -1165 2680 -1035
rect 2640 -1195 2645 -1165
rect 2675 -1195 2680 -1165
rect 2640 -1360 2680 -1195
rect 2720 -725 2760 -720
rect 2720 -755 2725 -725
rect 2755 -755 2760 -725
rect 2720 -885 2760 -755
rect 2720 -915 2725 -885
rect 2755 -915 2760 -885
rect 2720 -1005 2760 -915
rect 2720 -1035 2725 -1005
rect 2755 -1035 2760 -1005
rect 2720 -1165 2760 -1035
rect 2720 -1195 2725 -1165
rect 2755 -1195 2760 -1165
rect 2720 -1360 2760 -1195
rect 2800 -725 2840 -720
rect 2800 -755 2805 -725
rect 2835 -755 2840 -725
rect 2800 -885 2840 -755
rect 2800 -915 2805 -885
rect 2835 -915 2840 -885
rect 2800 -1005 2840 -915
rect 2800 -1035 2805 -1005
rect 2835 -1035 2840 -1005
rect 2800 -1165 2840 -1035
rect 2800 -1195 2805 -1165
rect 2835 -1195 2840 -1165
rect 2800 -1360 2840 -1195
rect 2880 -725 2920 -720
rect 2880 -755 2885 -725
rect 2915 -755 2920 -725
rect 2880 -885 2920 -755
rect 2880 -915 2885 -885
rect 2915 -915 2920 -885
rect 2880 -1005 2920 -915
rect 2880 -1035 2885 -1005
rect 2915 -1035 2920 -1005
rect 2880 -1165 2920 -1035
rect 2880 -1195 2885 -1165
rect 2915 -1195 2920 -1165
rect 2880 -1360 2920 -1195
rect 2960 -725 3000 -720
rect 2960 -755 2965 -725
rect 2995 -755 3000 -725
rect 2960 -885 3000 -755
rect 2960 -915 2965 -885
rect 2995 -915 3000 -885
rect 2960 -1005 3000 -915
rect 2960 -1035 2965 -1005
rect 2995 -1035 3000 -1005
rect 2960 -1165 3000 -1035
rect 2960 -1195 2965 -1165
rect 2995 -1195 3000 -1165
rect 2960 -1360 3000 -1195
rect 3040 -725 3080 -720
rect 3040 -755 3045 -725
rect 3075 -755 3080 -725
rect 3040 -885 3080 -755
rect 3040 -915 3045 -885
rect 3075 -915 3080 -885
rect 3040 -1005 3080 -915
rect 3120 -725 3160 -720
rect 3120 -755 3125 -725
rect 3155 -755 3160 -725
rect 3120 -885 3160 -755
rect 3120 -915 3125 -885
rect 3155 -915 3160 -885
rect 3120 -920 3160 -915
rect 3200 -725 3240 -720
rect 3200 -755 3205 -725
rect 3235 -755 3240 -725
rect 3200 -885 3240 -755
rect 3200 -915 3205 -885
rect 3235 -915 3240 -885
rect 3040 -1035 3045 -1005
rect 3075 -1035 3080 -1005
rect 3040 -1165 3080 -1035
rect 3040 -1195 3045 -1165
rect 3075 -1195 3080 -1165
rect 3040 -1360 3080 -1195
rect 3120 -1005 3160 -960
rect 3120 -1035 3125 -1005
rect 3155 -1035 3160 -1005
rect 3120 -1165 3160 -1035
rect 3120 -1195 3125 -1165
rect 3155 -1195 3160 -1165
rect 3120 -1200 3160 -1195
rect 3200 -1005 3240 -915
rect 3200 -1035 3205 -1005
rect 3235 -1035 3240 -1005
rect 3200 -1165 3240 -1035
rect 3200 -1195 3205 -1165
rect 3235 -1195 3240 -1165
rect 3200 -1360 3240 -1195
rect 3280 -725 3320 -720
rect 3280 -755 3285 -725
rect 3315 -755 3320 -725
rect 3280 -885 3320 -755
rect 3280 -915 3285 -885
rect 3315 -915 3320 -885
rect 3280 -1005 3320 -915
rect 3280 -1035 3285 -1005
rect 3315 -1035 3320 -1005
rect 3280 -1165 3320 -1035
rect 3280 -1195 3285 -1165
rect 3315 -1195 3320 -1165
rect 3280 -1360 3320 -1195
rect 3360 -725 3400 -720
rect 3360 -755 3365 -725
rect 3395 -755 3400 -725
rect 3360 -885 3400 -755
rect 3360 -915 3365 -885
rect 3395 -915 3400 -885
rect 3360 -1005 3400 -915
rect 3360 -1035 3365 -1005
rect 3395 -1035 3400 -1005
rect 3360 -1165 3400 -1035
rect 3360 -1195 3365 -1165
rect 3395 -1195 3400 -1165
rect 3360 -1360 3400 -1195
rect 3440 -725 3480 -720
rect 3440 -755 3445 -725
rect 3475 -755 3480 -725
rect 3440 -885 3480 -755
rect 3440 -915 3445 -885
rect 3475 -915 3480 -885
rect 3440 -1005 3480 -915
rect 3440 -1035 3445 -1005
rect 3475 -1035 3480 -1005
rect 3440 -1165 3480 -1035
rect 3440 -1195 3445 -1165
rect 3475 -1195 3480 -1165
rect 3440 -1360 3480 -1195
rect 3520 -725 3560 -720
rect 3520 -755 3525 -725
rect 3555 -755 3560 -725
rect 3520 -885 3560 -755
rect 3520 -915 3525 -885
rect 3555 -915 3560 -885
rect 3520 -1005 3560 -915
rect 3520 -1035 3525 -1005
rect 3555 -1035 3560 -1005
rect 3520 -1165 3560 -1035
rect 3520 -1195 3525 -1165
rect 3555 -1195 3560 -1165
rect 3520 -1360 3560 -1195
rect 3600 -725 3640 -720
rect 3600 -755 3605 -725
rect 3635 -755 3640 -725
rect 3600 -885 3640 -755
rect 3600 -915 3605 -885
rect 3635 -915 3640 -885
rect 3600 -1005 3640 -915
rect 3600 -1035 3605 -1005
rect 3635 -1035 3640 -1005
rect 3600 -1165 3640 -1035
rect 3600 -1195 3605 -1165
rect 3635 -1195 3640 -1165
rect 3600 -1360 3640 -1195
rect 3680 -725 3720 -720
rect 3680 -755 3685 -725
rect 3715 -755 3720 -725
rect 3680 -885 3720 -755
rect 3680 -915 3685 -885
rect 3715 -915 3720 -885
rect 3680 -1005 3720 -915
rect 3760 -725 3800 -720
rect 3760 -755 3765 -725
rect 3795 -755 3800 -725
rect 3760 -885 3800 -755
rect 3760 -915 3765 -885
rect 3795 -915 3800 -885
rect 3760 -920 3800 -915
rect 3840 -725 3880 -720
rect 3840 -755 3845 -725
rect 3875 -755 3880 -725
rect 3840 -885 3880 -755
rect 3840 -915 3845 -885
rect 3875 -915 3880 -885
rect 3680 -1035 3685 -1005
rect 3715 -1035 3720 -1005
rect 3680 -1165 3720 -1035
rect 3680 -1195 3685 -1165
rect 3715 -1195 3720 -1165
rect 3680 -1360 3720 -1195
rect 3760 -1005 3800 -960
rect 3760 -1035 3765 -1005
rect 3795 -1035 3800 -1005
rect 3760 -1165 3800 -1035
rect 3760 -1195 3765 -1165
rect 3795 -1195 3800 -1165
rect 3760 -1200 3800 -1195
rect 3840 -1005 3880 -915
rect 3840 -1035 3845 -1005
rect 3875 -1035 3880 -1005
rect 3840 -1165 3880 -1035
rect 3840 -1195 3845 -1165
rect 3875 -1195 3880 -1165
rect 3760 -1349 3800 -1320
rect 2480 -1440 2520 -1431
rect 3760 -1431 3764 -1349
rect 3796 -1431 3800 -1349
rect 3840 -1360 3880 -1195
rect 3920 -725 3960 -720
rect 3920 -755 3925 -725
rect 3955 -755 3960 -725
rect 3920 -885 3960 -755
rect 3920 -915 3925 -885
rect 3955 -915 3960 -885
rect 3920 -1005 3960 -915
rect 3920 -1035 3925 -1005
rect 3955 -1035 3960 -1005
rect 3920 -1165 3960 -1035
rect 3920 -1195 3925 -1165
rect 3955 -1195 3960 -1165
rect 3920 -1360 3960 -1195
rect 4000 -725 4040 -720
rect 4000 -755 4005 -725
rect 4035 -755 4040 -725
rect 4000 -885 4040 -755
rect 4000 -915 4005 -885
rect 4035 -915 4040 -885
rect 4000 -1005 4040 -915
rect 4000 -1035 4005 -1005
rect 4035 -1035 4040 -1005
rect 4000 -1165 4040 -1035
rect 4000 -1195 4005 -1165
rect 4035 -1195 4040 -1165
rect 4000 -1360 4040 -1195
rect 4080 -725 4120 -720
rect 4080 -755 4085 -725
rect 4115 -755 4120 -725
rect 4080 -885 4120 -755
rect 4080 -915 4085 -885
rect 4115 -915 4120 -885
rect 4080 -1005 4120 -915
rect 4080 -1035 4085 -1005
rect 4115 -1035 4120 -1005
rect 4080 -1165 4120 -1035
rect 4080 -1195 4085 -1165
rect 4115 -1195 4120 -1165
rect 4080 -1360 4120 -1195
rect 4160 -725 4200 -720
rect 4160 -755 4165 -725
rect 4195 -755 4200 -725
rect 4160 -885 4200 -755
rect 4160 -915 4165 -885
rect 4195 -915 4200 -885
rect 4160 -1005 4200 -915
rect 4160 -1035 4165 -1005
rect 4195 -1035 4200 -1005
rect 4160 -1165 4200 -1035
rect 4160 -1195 4165 -1165
rect 4195 -1195 4200 -1165
rect 4160 -1360 4200 -1195
rect 4240 -725 4280 -720
rect 4240 -755 4245 -725
rect 4275 -755 4280 -725
rect 4240 -885 4280 -755
rect 4240 -915 4245 -885
rect 4275 -915 4280 -885
rect 4240 -1005 4280 -915
rect 4240 -1035 4245 -1005
rect 4275 -1035 4280 -1005
rect 4240 -1165 4280 -1035
rect 4240 -1195 4245 -1165
rect 4275 -1195 4280 -1165
rect 4240 -1360 4280 -1195
rect 4320 -725 4360 -720
rect 4320 -755 4325 -725
rect 4355 -755 4360 -725
rect 4320 -885 4360 -755
rect 4320 -915 4325 -885
rect 4355 -915 4360 -885
rect 4320 -1005 4360 -915
rect 4400 -725 4440 -720
rect 4400 -755 4405 -725
rect 4435 -755 4440 -725
rect 4400 -885 4440 -755
rect 4400 -915 4405 -885
rect 4435 -915 4440 -885
rect 4400 -920 4440 -915
rect 4480 -725 4520 -720
rect 4480 -755 4485 -725
rect 4515 -755 4520 -725
rect 4480 -885 4520 -755
rect 4480 -915 4485 -885
rect 4515 -915 4520 -885
rect 4320 -1035 4325 -1005
rect 4355 -1035 4360 -1005
rect 4320 -1165 4360 -1035
rect 4320 -1195 4325 -1165
rect 4355 -1195 4360 -1165
rect 4320 -1360 4360 -1195
rect 4400 -1005 4440 -960
rect 4400 -1035 4405 -1005
rect 4435 -1035 4440 -1005
rect 4400 -1165 4440 -1035
rect 4400 -1195 4405 -1165
rect 4435 -1195 4440 -1165
rect 4400 -1200 4440 -1195
rect 4480 -1005 4520 -915
rect 4480 -1035 4485 -1005
rect 4515 -1035 4520 -1005
rect 4480 -1165 4520 -1035
rect 4480 -1195 4485 -1165
rect 4515 -1195 4520 -1165
rect 4480 -1360 4520 -1195
rect 4560 -725 4600 -720
rect 4560 -755 4565 -725
rect 4595 -755 4600 -725
rect 4560 -885 4600 -755
rect 4560 -915 4565 -885
rect 4595 -915 4600 -885
rect 4560 -1005 4600 -915
rect 4560 -1035 4565 -1005
rect 4595 -1035 4600 -1005
rect 4560 -1165 4600 -1035
rect 4560 -1195 4565 -1165
rect 4595 -1195 4600 -1165
rect 4560 -1360 4600 -1195
rect 4640 -725 4680 -720
rect 4640 -755 4645 -725
rect 4675 -755 4680 -725
rect 4640 -885 4680 -755
rect 4640 -915 4645 -885
rect 4675 -915 4680 -885
rect 4640 -1005 4680 -915
rect 4640 -1035 4645 -1005
rect 4675 -1035 4680 -1005
rect 4640 -1165 4680 -1035
rect 4640 -1195 4645 -1165
rect 4675 -1195 4680 -1165
rect 4640 -1360 4680 -1195
rect 4720 -725 4760 -720
rect 4720 -755 4725 -725
rect 4755 -755 4760 -725
rect 4720 -885 4760 -755
rect 4720 -915 4725 -885
rect 4755 -915 4760 -885
rect 4720 -1005 4760 -915
rect 4720 -1035 4725 -1005
rect 4755 -1035 4760 -1005
rect 4720 -1165 4760 -1035
rect 4720 -1195 4725 -1165
rect 4755 -1195 4760 -1165
rect 4720 -1360 4760 -1195
rect 4800 -725 4840 -720
rect 4800 -755 4805 -725
rect 4835 -755 4840 -725
rect 4800 -885 4840 -755
rect 4800 -915 4805 -885
rect 4835 -915 4840 -885
rect 4800 -1005 4840 -915
rect 4800 -1035 4805 -1005
rect 4835 -1035 4840 -1005
rect 4800 -1165 4840 -1035
rect 4800 -1195 4805 -1165
rect 4835 -1195 4840 -1165
rect 4800 -1360 4840 -1195
rect 4880 -725 4920 -720
rect 4880 -755 4885 -725
rect 4915 -755 4920 -725
rect 4880 -885 4920 -755
rect 4880 -915 4885 -885
rect 4915 -915 4920 -885
rect 4880 -1005 4920 -915
rect 4880 -1035 4885 -1005
rect 4915 -1035 4920 -1005
rect 4880 -1165 4920 -1035
rect 4880 -1195 4885 -1165
rect 4915 -1195 4920 -1165
rect 4880 -1360 4920 -1195
rect 4960 -725 5000 -720
rect 4960 -755 4965 -725
rect 4995 -755 5000 -725
rect 4960 -885 5000 -755
rect 4960 -915 4965 -885
rect 4995 -915 5000 -885
rect 4960 -1005 5000 -915
rect 4960 -1035 4965 -1005
rect 4995 -1035 5000 -1005
rect 4960 -1165 5000 -1035
rect 4960 -1195 4965 -1165
rect 4995 -1195 5000 -1165
rect 4960 -1360 5000 -1195
rect 5040 -725 5080 -720
rect 5040 -755 5045 -725
rect 5075 -755 5080 -725
rect 5040 -885 5080 -755
rect 5040 -915 5045 -885
rect 5075 -915 5080 -885
rect 5040 -1005 5080 -915
rect 5040 -1035 5045 -1005
rect 5075 -1035 5080 -1005
rect 5040 -1165 5080 -1035
rect 5040 -1195 5045 -1165
rect 5075 -1195 5080 -1165
rect 5040 -1349 5080 -1195
rect 3760 -1440 3800 -1431
rect 5040 -1431 5044 -1349
rect 5076 -1431 5080 -1349
rect 5120 -725 5160 -720
rect 5120 -755 5125 -725
rect 5155 -755 5160 -725
rect 5120 -885 5160 -755
rect 5120 -915 5125 -885
rect 5155 -915 5160 -885
rect 5120 -1005 5160 -915
rect 5120 -1035 5125 -1005
rect 5155 -1035 5160 -1005
rect 5120 -1165 5160 -1035
rect 5120 -1195 5125 -1165
rect 5155 -1195 5160 -1165
rect 5120 -1360 5160 -1195
rect 5200 -725 5240 -720
rect 5200 -755 5205 -725
rect 5235 -755 5240 -725
rect 5200 -885 5240 -755
rect 5200 -915 5205 -885
rect 5235 -915 5240 -885
rect 5200 -1165 5240 -915
rect 5200 -1195 5205 -1165
rect 5235 -1195 5240 -1165
rect 5200 -1360 5240 -1195
rect 5040 -1440 5080 -1431
<< via3 >>
rect -76 -1360 -44 -1349
rect -76 -1430 -75 -1360
rect -75 -1430 -45 -1360
rect -45 -1430 -44 -1360
rect -76 -1431 -44 -1430
rect 1204 -1360 1236 -1349
rect 1204 -1430 1205 -1360
rect 1205 -1430 1235 -1360
rect 1235 -1430 1236 -1360
rect 1204 -1431 1236 -1430
rect 2484 -1360 2516 -1349
rect 2484 -1430 2485 -1360
rect 2485 -1430 2515 -1360
rect 2515 -1430 2516 -1360
rect 2484 -1431 2516 -1430
rect 3764 -1360 3796 -1349
rect 3764 -1430 3765 -1360
rect 3765 -1430 3795 -1360
rect 3795 -1430 3796 -1360
rect 3764 -1431 3796 -1430
rect 5044 -1360 5076 -1349
rect 5044 -1430 5045 -1360
rect 5045 -1430 5075 -1360
rect 5075 -1430 5076 -1360
rect 5044 -1431 5076 -1430
<< metal4 >>
rect -240 -880 5240 -840
rect -240 -1000 -120 -880
rect 0 -1000 1160 -880
rect 1280 -1000 2440 -880
rect 2560 -1000 3720 -880
rect 3840 -1000 5000 -880
rect 5120 -1000 5240 -880
rect -240 -1040 5240 -1000
rect -240 -1349 5240 -1320
rect -240 -1431 -76 -1349
rect -44 -1360 1204 -1349
rect -44 -1431 520 -1360
rect -240 -1480 520 -1431
rect 640 -1431 1204 -1360
rect 1236 -1360 2484 -1349
rect 1236 -1431 1800 -1360
rect 640 -1480 1800 -1431
rect 1920 -1431 2484 -1360
rect 2516 -1360 3764 -1349
rect 2516 -1431 3080 -1360
rect 1920 -1480 3080 -1431
rect 3200 -1431 3764 -1360
rect 3796 -1360 5044 -1349
rect 3796 -1431 4360 -1360
rect 3200 -1480 4360 -1431
rect 4480 -1431 5044 -1360
rect 5076 -1431 5240 -1349
rect 4480 -1480 5240 -1431
rect -240 -1520 5240 -1480
<< via4 >>
rect -120 -1000 0 -880
rect 1160 -1000 1280 -880
rect 2440 -1000 2560 -880
rect 3720 -1000 3840 -880
rect 5000 -1000 5120 -880
rect 520 -1480 640 -1360
rect 1800 -1480 1920 -1360
rect 3080 -1480 3200 -1360
rect 4360 -1480 4480 -1360
<< metal5 >>
rect -160 -880 40 -720
rect -160 -1000 -120 -880
rect 0 -1000 40 -880
rect -160 -1520 40 -1000
rect 480 -1360 680 -720
rect 480 -1480 520 -1360
rect 640 -1480 680 -1360
rect 480 -1520 680 -1480
rect 1120 -880 1320 -720
rect 1120 -1000 1160 -880
rect 1280 -1000 1320 -880
rect 1120 -1520 1320 -1000
rect 1760 -1360 1960 -720
rect 1760 -1480 1800 -1360
rect 1920 -1480 1960 -1360
rect 1760 -1520 1960 -1480
rect 2400 -880 2600 -720
rect 2400 -1000 2440 -880
rect 2560 -1000 2600 -880
rect 2400 -1520 2600 -1000
rect 3040 -1360 3240 -720
rect 3040 -1480 3080 -1360
rect 3200 -1480 3240 -1360
rect 3040 -1520 3240 -1480
rect 3680 -880 3880 -720
rect 3680 -1000 3720 -880
rect 3840 -1000 3880 -880
rect 3680 -1520 3880 -1000
rect 4320 -1360 4520 -720
rect 4320 -1480 4360 -1360
rect 4480 -1480 4520 -1360
rect 4320 -1520 4520 -1480
rect 4960 -880 5160 -720
rect 4960 -1000 5000 -880
rect 5120 -1000 5160 -880
rect 4960 -1520 5160 -1000
<< labels >>
rlabel locali 2480 -1320 2520 -1280 0 xn
rlabel metal2 5200 -840 5240 -800 0 gnb
port 0 nsew
rlabel metal2 5200 -1120 5240 -1080 0 gna
port 1 nsew
rlabel metal5 -160 -760 40 -720 0 vdda
port 2 nsew
rlabel metal5 480 -760 680 -720 0 vssa
port 3 nsew
rlabel metal1 240 -1440 280 -1340 0 n1
rlabel metal1 880 -1440 920 -1340 0 n2
rlabel metal1 1520 -1440 1560 -1340 0 n3
rlabel metal1 2160 -1440 2200 -1340 0 n4
rlabel metal1 2800 -1440 2840 -1340 0 n5
rlabel metal1 3440 -1440 3480 -1340 0 n6
rlabel metal1 4080 -1440 4120 -1340 0 n7
rlabel metal1 4720 -1440 4760 -1340 0 n8
<< end >>
