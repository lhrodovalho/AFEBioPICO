* NGSPICE file created from opamp.ext - technology: sky130A

.subckt p1_8 D G S B SUB
X0 D G a7 B sky130_fd_pr__pfet_01v8_lvt ad=1.5e+12p pd=7e+06u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X1 a6 G a5 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X2 S G a1 B sky130_fd_pr__pfet_01v8_lvt ad=1.5e+12p pd=7e+06u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X3 a6 G a7 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X4 a2 G a3 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=3e+12p ps=1.4e+07u w=3e+06u l=8e+06u
X5 a2 G a1 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X6 a4 G a5 B sky130_fd_pr__pfet_01v8_lvt ad=3e+12p pd=1.4e+07u as=0p ps=0u w=3e+06u l=8e+06u
X7 a4 G a3 B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
.ends

.subckt n1_8 D G S B
X0 a5 G a6 B sky130_fd_pr__nfet_01v8_lvt ad=1e+12p pd=6e+06u as=1e+12p ps=6e+06u w=1e+06u l=8e+06u
X1 a1 G a2 B sky130_fd_pr__nfet_01v8_lvt ad=1e+12p pd=6e+06u as=1e+12p ps=6e+06u w=1e+06u l=8e+06u
X2 a1 G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=8e+06u
X3 a7 G D B sky130_fd_pr__nfet_01v8_lvt ad=1e+12p pd=6e+06u as=5e+11p ps=3e+06u w=1e+06u l=8e+06u
X4 a3 G a4 B sky130_fd_pr__nfet_01v8_lvt ad=1e+12p pd=6e+06u as=1e+12p ps=6e+06u w=1e+06u l=8e+06u
X5 a5 G a4 B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X6 a3 G a2 B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X7 a7 G a6 B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
.ends

.subckt n4_2 D G S B
X0 X G D B sky130_fd_pr__nfet_01v8_lvt ad=4e+12p pd=2.4e+07u as=2e+12p ps=1.2e+07u w=1e+06u l=8e+06u
X1 X G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2e+12p ps=1.2e+07u w=1e+06u l=8e+06u
X2 X G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X3 X G D B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X4 X G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X5 X G D B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X6 X G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X7 X G D B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
.ends

.subckt p8_1 D G S B SUB
X0 S G D B sky130_fd_pr__pfet_01v8_lvt ad=1.2e+13p pd=5.6e+07u as=1.2e+13p ps=5.6e+07u w=3e+06u l=8e+06u
X1 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X2 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X3 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X4 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X5 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X6 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X7 S G D B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
.ends

.subckt n8_1 D G S B
X0 D G S B sky130_fd_pr__nfet_01v8_lvt ad=4e+12p pd=2.4e+07u as=4e+12p ps=2.4e+07u w=1e+06u l=8e+06u
X1 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X2 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X3 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X4 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X5 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X6 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
X7 D G S B sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=8e+06u
.ends

.subckt p4_2 D G S B SUB
X0 D G X B sky130_fd_pr__pfet_01v8_lvt ad=6e+12p pd=2.8e+07u as=1.2e+13p ps=5.6e+07u w=3e+06u l=8e+06u
X1 D G X B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X2 S G X B sky130_fd_pr__pfet_01v8_lvt ad=6e+12p pd=2.8e+07u as=0p ps=0u w=3e+06u l=8e+06u
X3 D G X B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X4 S G X B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X5 S G X B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X6 D G X B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
X7 S G X B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
.ends

.subckt opamp inm inp out ib vdda gnda vssa
Xp1_8_31 x p1 vdda vdda vssa p1_8
Xp1_8_20 n2 p1 vdda vdda vssa p1_8
Xn1_8_40 n1 n1 vssa vssa n1_8
Xn4_2_6 out c vssa vssa n4_2
Xp1_8_5 b p1 vdda vdda vssa p1_8
Xp1_8_10 x p1 vdda vdda vssa p1_8
Xp1_8_32 n2 p1 vdda vdda vssa p1_8
Xp1_8_21 a p1 vdda vdda vssa p1_8
Xn4_2_7 out c vssa vssa n4_2
Xn1_8_41 xm a vssa vssa n1_8
Xn1_8_30 xp a vssa vssa n1_8
Xp1_8_6 p1 p1 vdda vdda vssa p1_8
Xp1_8_11 b p1 vdda vdda vssa p1_8
Xp1_8_33 a p1 vdda vdda vssa p1_8
Xp1_8_22 x p1 vdda vdda vssa p1_8
Xp1_8_7 x p1 vdda vdda vssa p1_8
Xn1_8_31 xm a vssa vssa n1_8
Xn1_8_20 xm a vssa vssa n1_8
Xpa2_1 ib ib p1 vdda vssa p8_1
Xp1_8_12 a p1 vdda vdda vssa p1_8
Xp1_8_34 x p1 vdda vdda vssa p1_8
Xp1_8_23 b p1 vdda vdda vssa p1_8
Xpd2_1 x inp xp vdda vssa p8_1
Xn1_8_10 xp a vssa vssa n1_8
Xn1_8_32 xp a vssa vssa n1_8
Xn1_8_21 n1 n1 vssa vssa n1_8
Xp1_8_8 n2 p1 vdda vdda vssa p1_8
Xp1_8_13 b p1 vdda vdda vssa p1_8
Xp1_8_35 b p1 vdda vdda vssa p1_8
Xp1_8_24 a p1 vdda vdda vssa p1_8
Xpd2_2 x inp xp vdda vssa p8_1
Xn1_8_11 xm a vssa vssa n1_8
Xp1_8_9 a p1 vdda vdda vssa p1_8
Xn1_8_33 xm a vssa vssa n1_8
Xn1_8_22 xm a vssa vssa n1_8
Xp1_8_14 x p1 vdda vdda vssa p1_8
Xp1_8_25 b p1 vdda vdda vssa p1_8
Xp1_8_36 a p1 vdda vdda vssa p1_8
Xn1_8_12 xp a vssa vssa n1_8
Xn1_8_34 xp a vssa vssa n1_8
Xn1_8_23 n1 n1 vssa vssa n1_8
Xn8_1_0 n2 n2 n1 vssa n8_1
Xp1_8_15 x p1 vdda vdda vssa p1_8
Xp1_8_26 x p1 vdda vdda vssa p1_8
Xp1_8_37 b p1 vdda vdda vssa p1_8
Xn8_1_1 a a xm vssa n8_1
Xn1_8_13 xm a vssa vssa n1_8
Xn1_8_35 xp a vssa vssa n1_8
Xn1_8_24 xp a vssa vssa n1_8
Xp1_8_16 p1 p1 vdda vdda vssa p1_8
Xp1_8_27 p1 p1 vdda vdda vssa p1_8
Xp1_8_38 x p1 vdda vdda vssa p1_8
Xn1_8_14 xp a vssa vssa n1_8
Xn1_8_36 vssa n1 vssa vssa n1_8
Xn1_8_25 xp a vssa vssa n1_8
Xn8_1_2 c a xp vssa n8_1
Xp4_2_0 out b vdda vdda vssa p4_2
Xp1_8_17 n2 p1 vdda vdda vssa p1_8
Xp1_8_28 n2 p1 vdda vdda vssa p1_8
Xp1_8_39 p1 p1 vdda vdda vssa p1_8
Xn1_8_15 xm a vssa vssa n1_8
Xn1_8_37 n1 n1 vssa vssa n1_8
Xn1_8_26 xp a vssa vssa n1_8
Xn8_1_3 c a xp vssa n8_1
Xp1_8_29 x p1 vdda vdda vssa p1_8
Xp1_8_18 p1 p1 vdda vdda vssa p1_8
Xp4_2_1 out b vdda vdda vssa p4_2
Xn1_8_16 vssa n1 vssa vssa n1_8
Xn1_8_38 xm a vssa vssa n1_8
Xn1_8_27 xp a vssa vssa n1_8
Xn8_1_4 a a xm vssa n8_1
Xp4_2_2 out b vdda vdda vssa p4_2
Xp1_8_19 x p1 vdda vdda vssa p1_8
Xn1_8_17 n1 n1 vssa vssa n1_8
Xn1_8_39 vssa n1 vssa vssa n1_8
Xn1_8_28 xm a vssa vssa n1_8
Xn8_1_5 c n2 b vssa n8_1
Xnf4_1 xp a vssa vssa n1_8
Xpc1_1 x p1 vdda vdda vssa p1_8
Xp4_2_3 out b vdda vdda vssa p4_2
Xn1_8_29 xm a vssa vssa n1_8
Xn1_8_18 vssa n1 vssa vssa n1_8
Xpf1_1 b p1 vdda vdda vssa p1_8
Xn8_1_6 vssa n1 vssa vssa n8_1
Xnf4_2 xp a vssa vssa n1_8
Xp4_2_4 out b vdda vdda vssa p4_2
Xn1_8_19 vssa n1 vssa vssa n1_8
Xn8_1_7 vssa n1 vssa vssa n8_1
Xp4_2_5 out b vdda vdda vssa p4_2
Xn8_1_8 vssa n1 vssa vssa n8_1
Xnf2_1 c n2 b vssa n8_1
Xp4_2_6 out b vdda vdda vssa p4_2
Xn8_1_9 a a xm vssa n8_1
Xp8_1_40 b ib c vdda vssa p8_1
Xp4_2_7 out b vdda vdda vssa p4_2
Xp8_1_41 x inm xm vdda vssa p8_1
Xp8_1_30 x inp xp vdda vssa p8_1
Xp8_1_20 ib ib p1 vdda vssa p8_1
Xp8_1_42 x inp xp vdda vssa p8_1
Xp8_1_31 x inm xm vdda vssa p8_1
Xn8_1_40 c a xp vssa n8_1
Xnb3_1 n2 n2 n1 vssa n8_1
Xp8_1_10 ib ib p1 vdda vssa p8_1
Xp8_1_21 vdda p1 vdda vdda vssa p8_1
Xp8_1_43 b ib c vdda vssa p8_1
Xp8_1_32 x inm xm vdda vssa p8_1
Xn1_8_0 n1 n1 vssa vssa n1_8
Xn8_1_41 a a xm vssa n8_1
Xn8_1_30 c n2 b vssa n8_1
Xne3_1 a a xm vssa n8_1
Xp8_1_11 x inp xp vdda vssa p8_1
Xp8_1_33 x inp xp vdda vssa p8_1
Xp8_1_22 vdda p1 vdda vdda vssa p8_1
Xp8_1_44 x inp xp vdda vssa p8_1
Xn1_8_1 vssa n1 vssa vssa n1_8
Xne3_2 a a xm vssa n8_1
Xn8_1_20 n2 n2 n1 vssa n8_1
Xn8_1_42 a a xm vssa n8_1
Xn8_1_31 a a xm vssa n8_1
Xp8_1_0 ib ib p1 vdda vssa p8_1
Xp8_1_12 x inp xp vdda vssa p8_1
Xp8_1_34 ib ib p1 vdda vssa p8_1
Xp8_1_23 ib ib p1 vdda vssa p8_1
Xp8_1_45 x inm xm vdda vssa p8_1
Xn1_8_2 xm a vssa vssa n1_8
Xn8_1_10 n2 n2 n1 vssa n8_1
Xn8_1_21 vssa n1 vssa vssa n8_1
Xn8_1_43 c a xp vssa n8_1
Xn8_1_32 c a xp vssa n8_1
Xp8_1_1 x inm xm vdda vssa p8_1
Xp8_1_13 b ib c vdda vssa p8_1
Xp8_1_35 vdda p1 vdda vdda vssa p8_1
Xp8_1_24 x inp xp vdda vssa p8_1
Xp8_1_46 x inm xm vdda vssa p8_1
Xn1_8_3 xp a vssa vssa n1_8
Xn8_1_11 c a xp vssa n8_1
Xn8_1_44 a a xm vssa n8_1
Xn8_1_33 c n2 b vssa n8_1
Xn8_1_22 vssa n1 vssa vssa n8_1
Xp8_1_2 x inp xp vdda vssa p8_1
Xp8_1_14 x inm xm vdda vssa p8_1
Xp8_1_36 vdda p1 vdda vdda vssa p8_1
Xp8_1_25 x inm xm vdda vssa p8_1
Xp8_1_47 x inp xp vdda vssa p8_1
Xn1_8_4 xp a vssa vssa n1_8
Xna4_1 vssa n1 vssa vssa n1_8
Xn8_1_12 c a xp vssa n8_1
Xn8_1_45 c a xp vssa n8_1
Xn8_1_34 a a xm vssa n8_1
Xn8_1_23 vssa n1 vssa vssa n8_1
Xpa1_1 p1 p1 vdda vdda vssa p1_8
Xp8_1_3 x inp xp vdda vssa p8_1
Xp8_1_15 x inm xm vdda vssa p8_1
Xp8_1_37 ib ib p1 vdda vssa p8_1
Xp8_1_26 b ib c vdda vssa p8_1
Xp8_1_48 ib ib p1 vdda vssa p8_1
Xn1_8_5 xm a vssa vssa n1_8
Xpd1_1 x p1 vdda vdda vssa p1_8
Xn8_1_13 c n2 b vssa n8_1
Xn8_1_46 n2 n2 n1 vssa n8_1
Xn8_1_35 c a xp vssa n8_1
Xn8_1_24 n2 n2 n1 vssa n8_1
Xp8_1_4 x inm xm vdda vssa p8_1
Xp8_1_16 b ib c vdda vssa p8_1
Xp8_1_38 x inp xp vdda vssa p8_1
Xp8_1_27 x inm xm vdda vssa p8_1
Xp8_1_49 vdda p1 vdda vdda vssa p8_1
Xn1_8_6 vssa n1 vssa vssa n1_8
Xn8_1_14 a a xm vssa n8_1
Xn8_1_47 n2 n2 n1 vssa n8_1
Xn8_1_36 c n2 b vssa n8_1
Xn8_1_25 n2 n2 n1 vssa n8_1
Xp8_1_5 b ib c vdda vssa p8_1
Xp8_1_17 x inp xp vdda vssa p8_1
Xp8_1_39 x inm xm vdda vssa p8_1
Xp8_1_28 x inp xp vdda vssa p8_1
Xn1_8_7 xm a vssa vssa n1_8
Xn8_1_15 c n2 b vssa n8_1
Xn8_1_48 vssa n1 vssa vssa n8_1
Xn8_1_37 c n2 b vssa n8_1
Xn8_1_26 c a xp vssa n8_1
Xp8_1_6 vdda p1 vdda vdda vssa p8_1
Xp8_1_18 x inm xm vdda vssa p8_1
Xp8_1_29 b ib c vdda vssa p8_1
Xn1_8_8 n1 n1 vssa vssa n1_8
Xn8_1_16 a a xm vssa n8_1
Xn8_1_49 vssa n1 vssa vssa n8_1
Xn8_1_38 c a xp vssa n8_1
Xn8_1_27 a a xm vssa n8_1
Xp8_1_7 vdda p1 vdda vdda vssa p8_1
Xp8_1_19 x inp xp vdda vssa p8_1
Xn1_8_9 xp a vssa vssa n1_8
Xn8_1_17 c a xp vssa n8_1
Xn8_1_39 a a xm vssa n8_1
Xn8_1_28 c a xp vssa n8_1
Xp8_1_8 vdda p1 vdda vdda vssa p8_1
Xpc2_1 x inm xm vdda vssa p8_1
Xpf2_1 b ib c vdda vssa p8_1
Xpc2_2 x inm xm vdda vssa p8_1
Xn8_1_18 a a xm vssa n8_1
Xn8_1_29 a a xm vssa n8_1
Xp8_1_9 x inm xm vdda vssa p8_1
Xn8_1_19 c a xp vssa n8_1
Xn4_2_0 out c vssa vssa n4_2
Xnf3_1 c a xp vssa n8_1
Xn4_2_1 out c vssa vssa n4_2
Xp1_8_0 p1 p1 vdda vdda vssa p1_8
Xnf3_2 c a xp vssa n8_1
Xn4_2_2 out c vssa vssa n4_2
Xp1_8_1 n2 p1 vdda vdda vssa p1_8
Xn4_2_3 out c vssa vssa n4_2
Xp1_8_2 x p1 vdda vdda vssa p1_8
Xnb4_1 n1 n1 vssa vssa n1_8
Xp1_8_40 n2 p1 vdda vdda vssa p1_8
Xn4_2_4 out c vssa vssa n4_2
Xp1_8_3 x p1 vdda vdda vssa p1_8
Xpb1_1 n2 p1 vdda vdda vssa p1_8
Xne4_1 xm a vssa vssa n1_8
Xp1_8_30 p1 p1 vdda vdda vssa p1_8
Xp1_8_41 x p1 vdda vdda vssa p1_8
Xpe1_1 a p1 vdda vdda vssa p1_8
Xn4_2_5 out c vssa vssa n4_2
Xp1_8_4 a p1 vdda vdda vssa p1_8
Xne4_2 xm a vssa vssa n1_8
X0 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X2 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X3 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X4 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X5 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X6 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X7 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X8 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X9 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X10 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X11 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X12 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X13 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X14 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X15 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X16 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X17 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X18 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X19 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X20 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X21 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X22 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X23 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X24 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X25 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X26 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X27 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X28 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X29 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X30 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X31 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X32 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X33 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X34 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X35 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X36 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X37 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X38 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X39 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X40 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X41 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X42 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X43 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X44 c out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X45 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X46 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X47 b out sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
C0 n1 gnda 701.66fF
C1 vdda gnda 118.61fF
C2 ib gnda 739.58fF
C3 out gnda 869.70fF
C4 a b 105.59fF
C5 p1 gnda 712.25fF
C6 c gnda 789.60fF
C7 out c 298.49fF
C8 inp gnda 748.76fF
C9 inm gnda 744.38fF
C10 gnda b 817.83fF
C11 out b 295.48fF
C12 n2 gnda 767.67fF
C13 x gnda 763.14fF
C14 gnda a 868.00fF
C15 xp gnda 776.34fF
C16 xm gnda 788.93fF
.ends

