magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< error_s >>
rect -952 70691 7432 70712
rect 11528 70691 19912 70712
rect 20160 70697 28472 70712
rect -952 70657 7417 70691
rect 11543 70657 19912 70691
rect -952 70640 7432 70657
rect -952 70560 -880 70640
rect -866 70600 7346 70626
rect -866 69480 -840 70600
rect -800 70534 7280 70560
rect -800 69592 -728 70534
rect 7254 69592 7280 70534
rect -800 69520 7280 69592
rect 7320 69480 7346 70600
rect 7360 69520 7432 70640
rect 11528 70640 19912 70657
rect 11528 70560 11600 70640
rect 11614 70600 19826 70626
rect -866 69454 7346 69480
rect 11614 69480 11640 70600
rect 11680 70534 19760 70560
rect 11680 69592 11752 70534
rect 19734 69592 19760 70534
rect 11680 69520 19760 69592
rect 19800 69480 19826 70600
rect 19840 69520 19912 70640
rect 20088 70691 28472 70697
rect 32568 70691 40952 70712
rect 20088 70657 28457 70691
rect 32583 70657 40952 70691
rect 20088 70640 28472 70657
rect 20088 70560 20160 70640
rect 20174 70600 28386 70626
rect 11614 69454 19826 69480
rect 20174 69480 20200 70600
rect 20240 70534 28320 70560
rect 20240 69592 20312 70534
rect 28294 69592 28320 70534
rect 20240 69520 28320 69592
rect 28360 69480 28386 70600
rect 28400 69520 28472 70640
rect 32568 70640 40952 70657
rect 32568 70560 32640 70640
rect 32654 70600 40866 70626
rect 20174 69454 28386 69480
rect 32654 69480 32680 70600
rect 32720 70534 40800 70560
rect 32720 69592 32792 70534
rect 40774 69592 40800 70534
rect 32720 69520 40800 69592
rect 40840 69480 40866 70600
rect 40880 69520 40952 70640
rect 32654 69454 40866 69480
rect -952 69200 7432 69272
rect -952 69120 -880 69200
rect -866 69160 7346 69186
rect -866 68040 -840 69160
rect -800 69094 7280 69120
rect -800 68152 -728 69094
rect 7254 68152 7280 69094
rect -800 68080 7280 68152
rect 7320 68040 7346 69160
rect 7360 68080 7432 69200
rect 11528 69200 19912 69272
rect 20160 69257 28472 69272
rect 11528 69120 11600 69200
rect 11614 69160 19826 69186
rect -866 68014 7346 68040
rect 11614 68040 11640 69160
rect 11680 69094 19760 69120
rect 11680 68152 11752 69094
rect 19734 68152 19760 69094
rect 11680 68080 19760 68152
rect 19800 68040 19826 69160
rect 19840 68080 19912 69200
rect 20088 69200 28472 69257
rect 20088 69120 20160 69200
rect 20174 69160 28386 69186
rect 11614 68014 19826 68040
rect 20174 68040 20200 69160
rect 20240 69094 28320 69120
rect 20240 68152 20312 69094
rect 28294 68152 28320 69094
rect 20240 68080 28320 68152
rect 28360 68040 28386 69160
rect 28400 68080 28472 69200
rect 32568 69200 40952 69272
rect 32568 69120 32640 69200
rect 32654 69160 40866 69186
rect 20174 68014 28386 68040
rect 32654 68040 32680 69160
rect 32720 69094 40800 69120
rect 32720 68152 32792 69094
rect 40774 68152 40800 69094
rect 32720 68080 40800 68152
rect 40840 68040 40866 69160
rect 40880 68080 40952 69200
rect 32654 68014 40866 68040
rect -952 67760 7432 67832
rect -952 67680 -880 67760
rect -866 67720 7346 67746
rect -866 66600 -840 67720
rect -800 67654 7280 67680
rect -800 66712 -728 67654
rect 7254 66712 7280 67654
rect -800 66640 7280 66712
rect 7320 66600 7346 67720
rect 7360 66640 7432 67760
rect 11528 67760 19912 67832
rect 20160 67817 28472 67832
rect 11528 67680 11600 67760
rect 11614 67720 19826 67746
rect -866 66574 7346 66600
rect 11614 66600 11640 67720
rect 11680 67654 19760 67680
rect 11680 66712 11752 67654
rect 19734 66712 19760 67654
rect 11680 66640 19760 66712
rect 19800 66600 19826 67720
rect 19840 66640 19912 67760
rect 20088 67760 28472 67817
rect 20088 67680 20160 67760
rect 20174 67720 28386 67746
rect 11614 66574 19826 66600
rect 20174 66600 20200 67720
rect 20240 67654 28320 67680
rect 20240 66712 20312 67654
rect 28294 66712 28320 67654
rect 20240 66640 28320 66712
rect 28360 66600 28386 67720
rect 28400 66640 28472 67760
rect 32568 67760 40952 67832
rect 32568 67680 32640 67760
rect 32654 67720 40866 67746
rect 20174 66574 28386 66600
rect 32654 66600 32680 67720
rect 32720 67654 40800 67680
rect 32720 66712 32792 67654
rect 40774 66712 40800 67654
rect 32720 66640 40800 66712
rect 40840 66600 40866 67720
rect 40880 66640 40952 67760
rect 32654 66574 40866 66600
rect -952 63120 7432 63192
rect -952 63040 -880 63120
rect -866 63080 7346 63106
rect -866 61960 -840 63080
rect -800 63014 7280 63040
rect -800 62072 -728 63014
rect 7254 62072 7280 63014
rect -800 62000 7280 62072
rect 7320 61960 7346 63080
rect 7360 62000 7432 63120
rect 11528 63120 19912 63192
rect 20160 63177 28472 63192
rect 11528 63040 11600 63120
rect 11614 63080 19826 63106
rect -866 61934 7346 61960
rect 11614 61960 11640 63080
rect 11680 63014 19760 63040
rect 11680 62072 11752 63014
rect 19734 62072 19760 63014
rect 11680 62000 19760 62072
rect 19800 61960 19826 63080
rect 19840 62000 19912 63120
rect 20088 63120 28472 63177
rect 20088 63040 20160 63120
rect 20174 63080 28386 63106
rect 11614 61934 19826 61960
rect 20174 61960 20200 63080
rect 20240 63014 28320 63040
rect 20240 62072 20312 63014
rect 28294 62072 28320 63014
rect 20240 62000 28320 62072
rect 28360 61960 28386 63080
rect 28400 62000 28472 63120
rect 32568 63120 40952 63192
rect 32568 63040 32640 63120
rect 32654 63080 40866 63106
rect 20174 61934 28386 61960
rect 32654 61960 32680 63080
rect 32720 63014 40800 63040
rect 32720 62072 32792 63014
rect 40774 62072 40800 63014
rect 32720 62000 40800 62072
rect 40840 61960 40866 63080
rect 40880 62000 40952 63120
rect 32654 61934 40866 61960
rect -952 60480 7432 60552
rect -952 60400 -880 60480
rect -866 60440 7346 60466
rect -866 59320 -840 60440
rect -800 60374 7280 60400
rect -800 59432 -728 60374
rect 7254 59432 7280 60374
rect -800 59360 7280 59432
rect 7320 59320 7346 60440
rect 7360 59360 7432 60480
rect 11528 60480 19912 60552
rect 20160 60537 28472 60552
rect 11528 60400 11600 60480
rect 11614 60440 19826 60466
rect -866 59294 7346 59320
rect 11614 59320 11640 60440
rect 11680 60374 19760 60400
rect 11680 59432 11752 60374
rect 19734 59432 19760 60374
rect 11680 59360 19760 59432
rect 19800 59320 19826 60440
rect 19840 59360 19912 60480
rect 20088 60480 28472 60537
rect 20088 60400 20160 60480
rect 20174 60440 28386 60466
rect 11614 59294 19826 59320
rect 20174 59320 20200 60440
rect 20240 60374 28320 60400
rect 20240 59432 20312 60374
rect 28294 59432 28320 60374
rect 20240 59360 28320 59432
rect 28360 59320 28386 60440
rect 28400 59360 28472 60480
rect 32568 60480 40952 60552
rect 32568 60400 32640 60480
rect 32654 60440 40866 60466
rect 20174 59294 28386 59320
rect 32654 59320 32680 60440
rect 32720 60374 40800 60400
rect 32720 59432 32792 60374
rect 40774 59432 40800 60374
rect 32720 59360 40800 59432
rect 40840 59320 40866 60440
rect 40880 59360 40952 60480
rect 32654 59294 40866 59320
rect -952 59040 7432 59112
rect -952 58960 -880 59040
rect -866 59000 7346 59026
rect -866 57880 -840 59000
rect -800 58934 7280 58960
rect -800 57992 -728 58934
rect 7254 57992 7280 58934
rect -800 57920 7280 57992
rect 7320 57880 7346 59000
rect 7360 57920 7432 59040
rect 11528 59040 19912 59112
rect 20160 59097 28472 59112
rect 11528 58960 11600 59040
rect 11614 59000 19826 59026
rect -866 57854 7346 57880
rect 11614 57880 11640 59000
rect 11680 58934 19760 58960
rect 11680 57992 11752 58934
rect 19734 57992 19760 58934
rect 11680 57920 19760 57992
rect 19800 57880 19826 59000
rect 19840 57920 19912 59040
rect 20088 59040 28472 59097
rect 20088 58960 20160 59040
rect 20174 59000 28386 59026
rect 11614 57854 19826 57880
rect 20174 57880 20200 59000
rect 20240 58934 28320 58960
rect 20240 57992 20312 58934
rect 28294 57992 28320 58934
rect 20240 57920 28320 57992
rect 28360 57880 28386 59000
rect 28400 57920 28472 59040
rect 32568 59040 40952 59112
rect 32568 58960 32640 59040
rect 32654 59000 40866 59026
rect 20174 57854 28386 57880
rect 32654 57880 32680 59000
rect 32720 58934 40800 58960
rect 32720 57992 32792 58934
rect 40774 57992 40800 58934
rect 32720 57920 40800 57992
rect 40840 57880 40866 59000
rect 40880 57920 40952 59040
rect 32654 57854 40866 57880
rect -952 57600 7432 57672
rect -952 57520 -880 57600
rect -866 57560 7346 57586
rect -866 56440 -840 57560
rect -800 57494 7280 57520
rect -800 56552 -728 57494
rect 7254 56552 7280 57494
rect -800 56480 7280 56552
rect 7320 56440 7346 57560
rect 7360 56480 7432 57600
rect 11528 57600 19912 57672
rect 20160 57657 28472 57672
rect 11528 57520 11600 57600
rect 11614 57560 19826 57586
rect -866 56414 7346 56440
rect 11614 56440 11640 57560
rect 11680 57494 19760 57520
rect 11680 56552 11752 57494
rect 19734 56552 19760 57494
rect 11680 56480 19760 56552
rect 19800 56440 19826 57560
rect 19840 56480 19912 57600
rect 20088 57600 28472 57657
rect 20088 57520 20160 57600
rect 20174 57560 28386 57586
rect 11614 56414 19826 56440
rect 20174 56440 20200 57560
rect 20240 57494 28320 57520
rect 20240 56552 20312 57494
rect 28294 56552 28320 57494
rect 20240 56480 28320 56552
rect 28360 56440 28386 57560
rect 28400 56480 28472 57600
rect 32568 57600 40952 57672
rect 32568 57520 32640 57600
rect 32654 57560 40866 57586
rect 20174 56414 28386 56440
rect 32654 56440 32680 57560
rect 32720 57494 40800 57520
rect 32720 56552 32792 57494
rect 40774 56552 40800 57494
rect 32720 56480 40800 56552
rect 40840 56440 40866 57560
rect 40880 56480 40952 57600
rect 32654 56414 40866 56440
rect -952 56160 7432 56232
rect -952 56080 -880 56160
rect -866 56120 7346 56146
rect -866 55000 -840 56120
rect -800 56054 7280 56080
rect -800 55112 -728 56054
rect 7254 55112 7280 56054
rect -800 55040 7280 55112
rect 7320 55000 7346 56120
rect 7360 55040 7432 56160
rect 11528 56160 19912 56232
rect 20160 56217 28472 56232
rect 11528 56080 11600 56160
rect 11614 56120 19826 56146
rect -866 54974 7346 55000
rect 11614 55000 11640 56120
rect 11680 56054 19760 56080
rect 11680 55112 11752 56054
rect 19734 55112 19760 56054
rect 11680 55040 19760 55112
rect 19800 55000 19826 56120
rect 19840 55040 19912 56160
rect 20088 56160 28472 56217
rect 20088 56080 20160 56160
rect 20174 56120 28386 56146
rect 11614 54974 19826 55000
rect 20174 55000 20200 56120
rect 20240 56054 28320 56080
rect 20240 55112 20312 56054
rect 28294 55112 28320 56054
rect 20240 55040 28320 55112
rect 28360 55000 28386 56120
rect 28400 55040 28472 56160
rect 32568 56160 40952 56232
rect 32568 56080 32640 56160
rect 32654 56120 40866 56146
rect 20174 54974 28386 55000
rect 32654 55000 32680 56120
rect 32720 56054 40800 56080
rect 32720 55112 32792 56054
rect 40774 55112 40800 56054
rect 32720 55040 40800 55112
rect 40840 55000 40866 56120
rect 40880 55040 40952 56160
rect 32654 54974 40866 55000
rect -952 52320 7432 52392
rect -952 52240 -880 52320
rect -866 52280 7346 52306
rect -866 51160 -840 52280
rect -800 52214 7280 52240
rect -800 51272 -728 52214
rect 7254 51272 7280 52214
rect -800 51200 7280 51272
rect 7320 51160 7346 52280
rect 7360 51200 7432 52320
rect 11528 52320 19912 52392
rect 20160 52377 28472 52392
rect 11528 52240 11600 52320
rect 11614 52280 19826 52306
rect -866 51134 7346 51160
rect 11614 51160 11640 52280
rect 11680 52214 19760 52240
rect 11680 51272 11752 52214
rect 19734 51272 19760 52214
rect 11680 51200 19760 51272
rect 19800 51160 19826 52280
rect 19840 51200 19912 52320
rect 20088 52320 28472 52377
rect 20088 52240 20160 52320
rect 20174 52280 28386 52306
rect 11614 51134 19826 51160
rect 20174 51160 20200 52280
rect 20240 52214 28320 52240
rect 20240 51272 20312 52214
rect 28294 51272 28320 52214
rect 20240 51200 28320 51272
rect 28360 51160 28386 52280
rect 28400 51200 28472 52320
rect 32568 52320 40952 52392
rect 32568 52240 32640 52320
rect 32654 52280 40866 52306
rect 20174 51134 28386 51160
rect 32654 51160 32680 52280
rect 32720 52214 40800 52240
rect 32720 51272 32792 52214
rect 40774 51272 40800 52214
rect 32720 51200 40800 51272
rect 40840 51160 40866 52280
rect 40880 51200 40952 52320
rect 32654 51134 40866 51160
rect -952 50880 7432 50952
rect -952 50800 -880 50880
rect -866 50840 7346 50866
rect -866 49720 -840 50840
rect -800 50774 7280 50800
rect -800 49832 -728 50774
rect 7254 49832 7280 50774
rect -800 49760 7280 49832
rect 7320 49720 7346 50840
rect 7360 49760 7432 50880
rect 11528 50880 19912 50952
rect 20160 50937 28472 50952
rect 11528 50800 11600 50880
rect 11614 50840 19826 50866
rect -866 49694 7346 49720
rect 11614 49720 11640 50840
rect 11680 50774 19760 50800
rect 11680 49832 11752 50774
rect 19734 49832 19760 50774
rect 11680 49760 19760 49832
rect 19800 49720 19826 50840
rect 19840 49760 19912 50880
rect 20088 50880 28472 50937
rect 20088 50800 20160 50880
rect 20174 50840 28386 50866
rect 11614 49694 19826 49720
rect 20174 49720 20200 50840
rect 20240 50774 28320 50800
rect 20240 49832 20312 50774
rect 28294 49832 28320 50774
rect 20240 49760 28320 49832
rect 28360 49720 28386 50840
rect 28400 49760 28472 50880
rect 32568 50880 40952 50952
rect 32568 50800 32640 50880
rect 32654 50840 40866 50866
rect 20174 49694 28386 49720
rect 32654 49720 32680 50840
rect 32720 50774 40800 50800
rect 32720 49832 32792 50774
rect 40774 49832 40800 50774
rect 32720 49760 40800 49832
rect 40840 49720 40866 50840
rect 40880 49760 40952 50880
rect 32654 49694 40866 49720
rect -952 49440 7432 49512
rect -952 49360 -880 49440
rect -866 49400 7346 49426
rect -866 48280 -840 49400
rect -800 49334 7280 49360
rect -800 48392 -728 49334
rect 7254 48392 7280 49334
rect -800 48320 7280 48392
rect 7320 48280 7346 49400
rect 7360 48320 7432 49440
rect 11528 49440 19912 49512
rect 20160 49497 28472 49512
rect 11528 49360 11600 49440
rect 11614 49400 19826 49426
rect -866 48254 7346 48280
rect 11614 48280 11640 49400
rect 11680 49334 19760 49360
rect 11680 48392 11752 49334
rect 19734 48392 19760 49334
rect 11680 48320 19760 48392
rect 19800 48280 19826 49400
rect 19840 48320 19912 49440
rect 20088 49440 28472 49497
rect 20088 49360 20160 49440
rect 20174 49400 28386 49426
rect 11614 48254 19826 48280
rect 20174 48280 20200 49400
rect 20240 49334 28320 49360
rect 20240 48392 20312 49334
rect 28294 48392 28320 49334
rect 20240 48320 28320 48392
rect 28360 48280 28386 49400
rect 28400 48320 28472 49440
rect 32568 49440 40952 49512
rect 32568 49360 32640 49440
rect 32654 49400 40866 49426
rect 20174 48254 28386 48280
rect 32654 48280 32680 49400
rect 32720 49334 40800 49360
rect 32720 48392 32792 49334
rect 40774 48392 40800 49334
rect 32720 48320 40800 48392
rect 40840 48280 40866 49400
rect 40880 48320 40952 49440
rect 32654 48254 40866 48280
rect -952 48000 7432 48072
rect -952 47920 -880 48000
rect -866 47960 7346 47986
rect -866 46840 -840 47960
rect -800 47894 7280 47920
rect -800 46952 -728 47894
rect 7254 46952 7280 47894
rect -800 46880 7280 46952
rect 7320 46840 7346 47960
rect 7360 46880 7432 48000
rect 11528 48000 19912 48072
rect 20160 48057 28472 48072
rect 11528 47920 11600 48000
rect 11614 47960 19826 47986
rect -866 46814 7346 46840
rect 11614 46840 11640 47960
rect 11680 47894 19760 47920
rect 11680 46952 11752 47894
rect 19734 46952 19760 47894
rect 11680 46880 19760 46952
rect 19800 46840 19826 47960
rect 19840 46880 19912 48000
rect 20088 48000 28472 48057
rect 20088 47920 20160 48000
rect 20174 47960 28386 47986
rect 11614 46814 19826 46840
rect 20174 46840 20200 47960
rect 20240 47894 28320 47920
rect 20240 46952 20312 47894
rect 28294 46952 28320 47894
rect 20240 46880 28320 46952
rect 28360 46840 28386 47960
rect 28400 46880 28472 48000
rect 32568 48000 40952 48072
rect 32568 47920 32640 48000
rect 32654 47960 40866 47986
rect 20174 46814 28386 46840
rect 32654 46840 32680 47960
rect 32720 47894 40800 47920
rect 32720 46952 32792 47894
rect 40774 46952 40800 47894
rect 32720 46880 40800 46952
rect 40840 46840 40866 47960
rect 40880 46880 40952 48000
rect 32654 46814 40866 46840
rect -952 44160 7432 44232
rect -952 44080 -880 44160
rect -866 44120 7346 44146
rect -866 43000 -840 44120
rect -800 44054 7280 44080
rect -800 43112 -728 44054
rect 7254 43112 7280 44054
rect -800 43040 7280 43112
rect 7320 43000 7346 44120
rect 7360 43040 7432 44160
rect 11528 44160 19912 44232
rect 20160 44217 28472 44232
rect 11528 44080 11600 44160
rect 11614 44120 19826 44146
rect -866 42974 7346 43000
rect 11614 43000 11640 44120
rect 11680 44054 19760 44080
rect 11680 43112 11752 44054
rect 19734 43112 19760 44054
rect 11680 43040 19760 43112
rect 19800 43000 19826 44120
rect 19840 43040 19912 44160
rect 20088 44160 28472 44217
rect 20088 44080 20160 44160
rect 20174 44120 28386 44146
rect 11614 42974 19826 43000
rect 20174 43000 20200 44120
rect 20240 44054 28320 44080
rect 20240 43112 20312 44054
rect 28294 43112 28320 44054
rect 20240 43040 28320 43112
rect 28360 43000 28386 44120
rect 28400 43040 28472 44160
rect 32568 44160 40952 44232
rect 32568 44080 32640 44160
rect 32654 44120 40866 44146
rect 20174 42974 28386 43000
rect 32654 43000 32680 44120
rect 32720 44054 40800 44080
rect 32720 43112 32792 44054
rect 40774 43112 40800 44054
rect 32720 43040 40800 43112
rect 40840 43000 40866 44120
rect 40880 43040 40952 44160
rect 32654 42974 40866 43000
rect -952 42720 7432 42792
rect -952 42640 -880 42720
rect -866 42680 7346 42706
rect -866 41560 -840 42680
rect -800 42614 7280 42640
rect -800 41672 -728 42614
rect 7254 41672 7280 42614
rect -800 41600 7280 41672
rect 7320 41560 7346 42680
rect 7360 41600 7432 42720
rect 11528 42720 19912 42792
rect 20160 42777 28472 42792
rect 11528 42640 11600 42720
rect 11614 42680 19826 42706
rect -866 41534 7346 41560
rect 11614 41560 11640 42680
rect 11680 42614 19760 42640
rect 11680 41672 11752 42614
rect 19734 41672 19760 42614
rect 11680 41600 19760 41672
rect 19800 41560 19826 42680
rect 19840 41600 19912 42720
rect 20088 42720 28472 42777
rect 20088 42640 20160 42720
rect 20174 42680 28386 42706
rect 11614 41534 19826 41560
rect 20174 41560 20200 42680
rect 20240 42614 28320 42640
rect 20240 41672 20312 42614
rect 28294 41672 28320 42614
rect 20240 41600 28320 41672
rect 28360 41560 28386 42680
rect 28400 41600 28472 42720
rect 32568 42720 40952 42792
rect 32568 42640 32640 42720
rect 32654 42680 40866 42706
rect 20174 41534 28386 41560
rect 32654 41560 32680 42680
rect 32720 42614 40800 42640
rect 32720 41672 32792 42614
rect 40774 41672 40800 42614
rect 32720 41600 40800 41672
rect 40840 41560 40866 42680
rect 40880 41600 40952 42720
rect 32654 41534 40866 41560
rect -17272 39840 -12248 39912
rect -17272 39760 -17200 39840
rect -17186 39800 -12334 39826
rect -17186 38840 -17160 39800
rect -17120 39734 -12400 39760
rect -17120 38952 -17048 39734
rect -12426 38952 -12400 39734
rect -17120 38880 -12400 38952
rect -12360 38840 -12334 39800
rect -12320 38880 -12248 39840
rect -8792 39840 -3768 39912
rect -8792 39760 -8720 39840
rect -8706 39800 -3854 39826
rect -17186 38814 -12334 38840
rect -8706 38840 -8680 39800
rect -8640 39734 -3920 39760
rect -8640 38952 -8568 39734
rect -3946 38952 -3920 39734
rect -8640 38880 -3920 38952
rect -3880 38840 -3854 39800
rect -3840 38880 -3768 39840
rect -8706 38814 -3854 38840
rect -17272 38560 -12248 38632
rect -17272 38480 -17200 38560
rect -17186 38520 -12334 38546
rect -17186 37560 -17160 38520
rect -17120 38454 -12400 38480
rect -17120 37672 -17048 38454
rect -12426 37672 -12400 38454
rect -17120 37600 -12400 37672
rect -12360 37560 -12334 38520
rect -12320 37600 -12248 38560
rect -8792 38560 -3768 38632
rect -8792 38480 -8720 38560
rect -8706 38520 -3854 38546
rect -17186 37534 -12334 37560
rect -8706 37560 -8680 38520
rect -8640 38454 -3920 38480
rect -8640 37672 -8568 38454
rect -3946 37672 -3920 38454
rect -8640 37600 -3920 37672
rect -3880 37560 -3854 38520
rect -3840 37600 -3768 38560
rect -8706 37534 -3854 37560
rect -17272 37280 -12248 37352
rect -17272 37200 -17200 37280
rect -17186 37240 -12334 37266
rect -17186 36280 -17160 37240
rect -17120 37174 -12400 37200
rect -17120 36392 -17048 37174
rect -12426 36392 -12400 37174
rect -17120 36320 -12400 36392
rect -12360 36280 -12334 37240
rect -12320 36320 -12248 37280
rect -8792 37280 -3768 37352
rect -8792 37200 -8720 37280
rect -8706 37240 -3854 37266
rect -17186 36254 -12334 36280
rect -8706 36280 -8680 37240
rect -8640 37174 -3920 37200
rect -8640 36392 -8568 37174
rect -3946 36392 -3920 37174
rect -8640 36320 -3920 36392
rect -3880 36280 -3854 37240
rect -3840 36320 -3768 37280
rect -8706 36254 -3854 36280
rect -17272 36000 -12248 36072
rect -17272 35920 -17200 36000
rect -17186 35960 -12334 35986
rect -17186 35000 -17160 35960
rect -17120 35894 -12400 35920
rect -17120 35112 -17048 35894
rect -12426 35112 -12400 35894
rect -17120 35040 -12400 35112
rect -12360 35000 -12334 35960
rect -12320 35040 -12248 36000
rect -8792 36000 -3768 36072
rect -8792 35920 -8720 36000
rect -8706 35960 -3854 35986
rect -17186 34974 -12334 35000
rect -8706 35000 -8680 35960
rect -8640 35894 -3920 35920
rect -8640 35112 -8568 35894
rect -3946 35112 -3920 35894
rect -8640 35040 -3920 35112
rect -3880 35000 -3854 35960
rect -3840 35040 -3768 36000
rect -8706 34974 -3854 35000
rect -952 33280 7432 33352
rect -952 33200 -880 33280
rect -866 33240 7346 33266
rect -866 32120 -840 33240
rect -800 33174 7280 33200
rect -800 32232 -728 33174
rect 7254 32232 7280 33174
rect -800 32160 7280 32232
rect 7320 32120 7346 33240
rect 7360 32160 7432 33280
rect 11528 33280 19912 33352
rect 20160 33337 28472 33352
rect 11528 33200 11600 33280
rect 11614 33240 19826 33266
rect -866 32094 7346 32120
rect 11614 32120 11640 33240
rect 11680 33174 19760 33200
rect 11680 32232 11752 33174
rect 19734 32232 19760 33174
rect 11680 32160 19760 32232
rect 19800 32120 19826 33240
rect 19840 32160 19912 33280
rect 20088 33280 28472 33337
rect 20088 33200 20160 33280
rect 20174 33240 28386 33266
rect 11614 32094 19826 32120
rect 20174 32120 20200 33240
rect 20240 33174 28320 33200
rect 20240 32232 20312 33174
rect 28294 32232 28320 33174
rect 20240 32160 28320 32232
rect 28360 32120 28386 33240
rect 28400 32160 28472 33280
rect 32568 33280 40952 33352
rect 32568 33200 32640 33280
rect 32654 33240 40866 33266
rect 20174 32094 28386 32120
rect 32654 32120 32680 33240
rect 32720 33174 40800 33200
rect 32720 32232 32792 33174
rect 40774 32232 40800 33174
rect 32720 32160 40800 32232
rect 40840 32120 40866 33240
rect 40880 32160 40952 33280
rect 32654 32094 40866 32120
rect -952 31840 7432 31912
rect -952 31760 -880 31840
rect -866 31800 7346 31826
rect -866 30680 -840 31800
rect -800 31734 7280 31760
rect -800 30792 -728 31734
rect 7254 30792 7280 31734
rect -800 30720 7280 30792
rect 7320 30680 7346 31800
rect 7360 30720 7432 31840
rect 11528 31840 19912 31912
rect 20160 31897 28472 31912
rect 11528 31760 11600 31840
rect 11614 31800 19826 31826
rect -866 30654 7346 30680
rect 11614 30680 11640 31800
rect 11680 31734 19760 31760
rect 11680 30792 11752 31734
rect 19734 30792 19760 31734
rect 11680 30720 19760 30792
rect 19800 30680 19826 31800
rect 19840 30720 19912 31840
rect 20088 31840 28472 31897
rect 20088 31760 20160 31840
rect 20174 31800 28386 31826
rect 11614 30654 19826 30680
rect 20174 30680 20200 31800
rect 20240 31734 28320 31760
rect 20240 30792 20312 31734
rect 28294 30792 28320 31734
rect 20240 30720 28320 30792
rect 28360 30680 28386 31800
rect 28400 30720 28472 31840
rect 32568 31840 40952 31912
rect 32568 31760 32640 31840
rect 32654 31800 40866 31826
rect 20174 30654 28386 30680
rect 32654 30680 32680 31800
rect 32720 31734 40800 31760
rect 32720 30792 32792 31734
rect 40774 30792 40800 31734
rect 32720 30720 40800 30792
rect 40840 30680 40866 31800
rect 40880 30720 40952 31840
rect 32654 30654 40866 30680
rect -952 28000 7432 28072
rect -952 27920 -880 28000
rect -866 27960 7346 27986
rect -866 26840 -840 27960
rect -800 27894 7280 27920
rect -800 26952 -728 27894
rect 7254 26952 7280 27894
rect -800 26880 7280 26952
rect 7320 26840 7346 27960
rect 7360 26880 7432 28000
rect 11528 28000 19912 28072
rect 20160 28057 28472 28072
rect 11528 27920 11600 28000
rect 11614 27960 19826 27986
rect -866 26814 7346 26840
rect 11614 26840 11640 27960
rect 11680 27894 19760 27920
rect 11680 26952 11752 27894
rect 19734 26952 19760 27894
rect 11680 26880 19760 26952
rect 19800 26840 19826 27960
rect 19840 26880 19912 28000
rect 20088 28000 28472 28057
rect 20088 27920 20160 28000
rect 20174 27960 28386 27986
rect 11614 26814 19826 26840
rect 20174 26840 20200 27960
rect 20240 27894 28320 27920
rect 20240 26952 20312 27894
rect 28294 26952 28320 27894
rect 20240 26880 28320 26952
rect 28360 26840 28386 27960
rect 28400 26880 28472 28000
rect 32568 28000 40952 28072
rect 32568 27920 32640 28000
rect 32654 27960 40866 27986
rect 20174 26814 28386 26840
rect 32654 26840 32680 27960
rect 32720 27894 40800 27920
rect 32720 26952 32792 27894
rect 40774 26952 40800 27894
rect 32720 26880 40800 26952
rect 40840 26840 40866 27960
rect 40880 26880 40952 28000
rect 32654 26814 40866 26840
rect -952 26560 7432 26632
rect -952 26480 -880 26560
rect -866 26520 7346 26546
rect -866 25400 -840 26520
rect -800 26454 7280 26480
rect -800 25512 -728 26454
rect 7254 25512 7280 26454
rect -800 25440 7280 25512
rect 7320 25400 7346 26520
rect 7360 25440 7432 26560
rect 11528 26560 19912 26632
rect 20160 26617 28472 26632
rect 11528 26480 11600 26560
rect 11614 26520 19826 26546
rect -866 25374 7346 25400
rect 11614 25400 11640 26520
rect 11680 26454 19760 26480
rect 11680 25512 11752 26454
rect 19734 25512 19760 26454
rect 11680 25440 19760 25512
rect 19800 25400 19826 26520
rect 19840 25440 19912 26560
rect 20088 26560 28472 26617
rect 20088 26480 20160 26560
rect 20174 26520 28386 26546
rect 11614 25374 19826 25400
rect 20174 25400 20200 26520
rect 20240 26454 28320 26480
rect 20240 25512 20312 26454
rect 28294 25512 28320 26454
rect 20240 25440 28320 25512
rect 28360 25400 28386 26520
rect 28400 25440 28472 26560
rect 32568 26560 40952 26632
rect 32568 26480 32640 26560
rect 32654 26520 40866 26546
rect 20174 25374 28386 25400
rect 32654 25400 32680 26520
rect 32720 26454 40800 26480
rect 32720 25512 32792 26454
rect 40774 25512 40800 26454
rect 32720 25440 40800 25512
rect 40840 25400 40866 26520
rect 40880 25440 40952 26560
rect 32654 25374 40866 25400
rect -952 25120 7432 25192
rect -952 25040 -880 25120
rect -866 25080 7346 25106
rect -866 23960 -840 25080
rect -800 25014 7280 25040
rect -800 24072 -728 25014
rect 7254 24072 7280 25014
rect -800 24000 7280 24072
rect 7320 23960 7346 25080
rect 7360 24000 7432 25120
rect 11528 25120 19912 25192
rect 20160 25177 28472 25192
rect 11528 25040 11600 25120
rect 11614 25080 19826 25106
rect -866 23934 7346 23960
rect 11614 23960 11640 25080
rect 11680 25014 19760 25040
rect 11680 24072 11752 25014
rect 19734 24072 19760 25014
rect 11680 24000 19760 24072
rect 19800 23960 19826 25080
rect 19840 24000 19912 25120
rect 20088 25120 28472 25177
rect 20088 25040 20160 25120
rect 20174 25080 28386 25106
rect 11614 23934 19826 23960
rect 20174 23960 20200 25080
rect 20240 25014 28320 25040
rect 20240 24072 20312 25014
rect 28294 24072 28320 25014
rect 20240 24000 28320 24072
rect 28360 23960 28386 25080
rect 28400 24000 28472 25120
rect 32568 25120 40952 25192
rect 32568 25040 32640 25120
rect 32654 25080 40866 25106
rect 20174 23934 28386 23960
rect 32654 23960 32680 25080
rect 32720 25014 40800 25040
rect 32720 24072 32792 25014
rect 40774 24072 40800 25014
rect 32720 24000 40800 24072
rect 40840 23960 40866 25080
rect 40880 24000 40952 25120
rect 32654 23934 40866 23960
rect -952 23680 7432 23752
rect -952 23600 -880 23680
rect -866 23640 7346 23666
rect -866 22520 -840 23640
rect -800 23574 7280 23600
rect -800 22632 -728 23574
rect 7254 22632 7280 23574
rect -800 22560 7280 22632
rect 7320 22520 7346 23640
rect 7360 22560 7432 23680
rect 11528 23680 19912 23752
rect 20160 23737 28472 23752
rect 11528 23600 11600 23680
rect 11614 23640 19826 23666
rect -866 22494 7346 22520
rect 11614 22520 11640 23640
rect 11680 23574 19760 23600
rect 11680 22632 11752 23574
rect 19734 22632 19760 23574
rect 11680 22560 19760 22632
rect 19800 22520 19826 23640
rect 19840 22560 19912 23680
rect 20088 23680 28472 23737
rect 20088 23600 20160 23680
rect 20174 23640 28386 23666
rect 11614 22494 19826 22520
rect 20174 22520 20200 23640
rect 20240 23574 28320 23600
rect 20240 22632 20312 23574
rect 28294 22632 28320 23574
rect 20240 22560 28320 22632
rect 28360 22520 28386 23640
rect 28400 22560 28472 23680
rect 32568 23680 40952 23752
rect 32568 23600 32640 23680
rect 32654 23640 40866 23666
rect 20174 22494 28386 22520
rect 32654 22520 32680 23640
rect 32720 23574 40800 23600
rect 32720 22632 32792 23574
rect 40774 22632 40800 23574
rect 32720 22560 40800 22632
rect 40840 22520 40866 23640
rect 40880 22560 40952 23680
rect 32654 22494 40866 22520
rect -952 19840 300 19912
rect 39700 19840 40952 19912
rect -952 19760 -880 19840
rect -866 19800 300 19826
rect 39700 19800 40866 19826
rect -866 18680 -840 19800
rect -800 19734 300 19760
rect 39700 19734 40800 19760
rect -800 18792 -728 19734
rect 40774 18792 40800 19734
rect -800 18720 300 18792
rect 39700 18720 40800 18792
rect 40840 18680 40866 19800
rect 40880 18720 40952 19840
rect -866 18654 300 18680
rect 39700 18654 40866 18680
rect -952 18400 300 18472
rect 39700 18400 40952 18472
rect -952 18320 -880 18400
rect -866 18360 300 18386
rect 39700 18360 40866 18386
rect -866 17240 -840 18360
rect -800 18294 300 18320
rect 39700 18294 40800 18320
rect -800 17352 -728 18294
rect 40774 17352 40800 18294
rect -800 17280 300 17352
rect 39700 17280 40800 17352
rect 40840 17240 40866 18360
rect 40880 17280 40952 18400
rect -866 17214 300 17240
rect 39700 17214 40866 17240
rect -952 16960 300 17032
rect 39700 16960 40952 17032
rect -952 16880 -880 16960
rect -866 16920 300 16946
rect 39700 16920 40866 16946
rect -866 15800 -840 16920
rect -800 16854 300 16880
rect 39700 16854 40800 16880
rect -800 15912 -728 16854
rect 40774 15912 40800 16854
rect -800 15840 300 15912
rect 39700 15840 40800 15912
rect 40840 15800 40866 16920
rect 40880 15840 40952 16960
rect -866 15774 300 15800
rect 39700 15774 40866 15800
rect -952 15520 300 15592
rect 39700 15520 40952 15592
rect -952 15440 -880 15520
rect -866 15480 300 15506
rect 39700 15480 40866 15506
rect -866 14360 -840 15480
rect -800 15414 300 15440
rect 39700 15414 40800 15440
rect -800 14472 -728 15414
rect 40774 14472 40800 15414
rect -800 14400 300 14472
rect 39700 14400 40800 14472
rect 40840 14360 40866 15480
rect 40880 14400 40952 15520
rect -866 14334 300 14360
rect 39700 14334 40866 14360
rect -952 12880 300 12952
rect 39700 12880 40952 12952
rect -952 12800 -880 12880
rect -866 12840 300 12866
rect 39700 12840 40866 12866
rect -866 11720 -840 12840
rect -800 12774 300 12800
rect 39700 12774 40800 12800
rect -800 11832 -728 12774
rect 40774 11832 40800 12774
rect -800 11760 300 11832
rect 39700 11760 40800 11832
rect 40840 11720 40866 12840
rect 40880 11760 40952 12880
rect -866 11694 300 11720
rect 39700 11694 40866 11720
rect -952 8240 300 8312
rect 39700 8240 40952 8312
rect -952 8160 -880 8240
rect -866 8200 300 8226
rect 39700 8200 40866 8226
rect -866 7080 -840 8200
rect -800 8134 300 8160
rect 39700 8134 40800 8160
rect -800 7192 -728 8134
rect 40774 7192 40800 8134
rect -800 7120 300 7192
rect 39700 7120 40800 7192
rect 40840 7080 40866 8200
rect 40880 7120 40952 8240
rect -866 7054 300 7080
rect 39700 7054 40866 7080
rect -952 6800 300 6872
rect 39700 6800 40952 6872
rect -952 6720 -880 6800
rect -866 6760 300 6786
rect 39700 6760 40866 6786
rect -866 5640 -840 6760
rect -800 6694 300 6720
rect 39700 6694 40800 6720
rect -800 5752 -728 6694
rect 40774 5752 40800 6694
rect -800 5680 300 5752
rect 39700 5680 40800 5752
rect 40840 5640 40866 6760
rect 40880 5680 40952 6800
rect -866 5614 300 5640
rect 39700 5614 40866 5640
rect -952 5360 300 5432
rect 39700 5360 40952 5432
rect -952 5280 -880 5360
rect -866 5320 300 5346
rect 39700 5320 40866 5346
rect -866 4200 -840 5320
rect -800 5254 300 5280
rect 39700 5254 40800 5280
rect -800 4312 -728 5254
rect 40774 4312 40800 5254
rect -800 4240 300 4312
rect 39700 4240 40800 4312
rect 40840 4200 40866 5320
rect 40880 4240 40952 5360
rect -866 4174 300 4200
rect 39700 4174 40866 4200
<< locali >>
rect -29920 42857 -29840 42880
rect -29920 42823 -29897 42857
rect -29863 42823 -29840 42857
rect -29920 42537 -29840 42823
rect -29920 42503 -29897 42537
rect -29863 42503 -29840 42537
rect -29920 42217 -29840 42503
rect -29920 42183 -29897 42217
rect -29863 42183 -29840 42217
rect -29920 41897 -29840 42183
rect -29920 41863 -29897 41897
rect -29863 41863 -29840 41897
rect -29920 41840 -29840 41863
rect -29760 42857 -29680 42880
rect -29760 42823 -29737 42857
rect -29703 42823 -29680 42857
rect -29760 42537 -29680 42823
rect -29760 42503 -29737 42537
rect -29703 42503 -29680 42537
rect -29760 42217 -29680 42503
rect -29760 42183 -29737 42217
rect -29703 42183 -29680 42217
rect -29760 41897 -29680 42183
rect -29760 41863 -29737 41897
rect -29703 41863 -29680 41897
rect -29760 41840 -29680 41863
rect -29600 42857 -29520 42880
rect -29600 42823 -29577 42857
rect -29543 42823 -29520 42857
rect -29600 42537 -29520 42823
rect -29600 42503 -29577 42537
rect -29543 42503 -29520 42537
rect -29600 42217 -29520 42503
rect -29600 42183 -29577 42217
rect -29543 42183 -29520 42217
rect -29600 41897 -29520 42183
rect -29600 41863 -29577 41897
rect -29543 41863 -29520 41897
rect -29600 41840 -29520 41863
rect -29440 42857 -29360 42880
rect -29440 42823 -29417 42857
rect -29383 42823 -29360 42857
rect -29440 42537 -29360 42823
rect -29440 42503 -29417 42537
rect -29383 42503 -29360 42537
rect -29440 42217 -29360 42503
rect -29440 42183 -29417 42217
rect -29383 42183 -29360 42217
rect -29440 41897 -29360 42183
rect -29440 41863 -29417 41897
rect -29383 41863 -29360 41897
rect -29440 41840 -29360 41863
rect -29280 42857 -29200 42880
rect -29280 42823 -29257 42857
rect -29223 42823 -29200 42857
rect -29280 42537 -29200 42823
rect -29280 42503 -29257 42537
rect -29223 42503 -29200 42537
rect -29280 42217 -29200 42503
rect -29280 42183 -29257 42217
rect -29223 42183 -29200 42217
rect -29280 41897 -29200 42183
rect -29280 41863 -29257 41897
rect -29223 41863 -29200 41897
rect -29280 41840 -29200 41863
rect -29120 42857 -29040 42880
rect -29120 42823 -29097 42857
rect -29063 42823 -29040 42857
rect -29120 42537 -29040 42823
rect -29120 42503 -29097 42537
rect -29063 42503 -29040 42537
rect -29120 42217 -29040 42503
rect -29120 42183 -29097 42217
rect -29063 42183 -29040 42217
rect -29120 41897 -29040 42183
rect -29120 41863 -29097 41897
rect -29063 41863 -29040 41897
rect -29120 41840 -29040 41863
rect -28960 42857 -28880 42880
rect -28960 42823 -28937 42857
rect -28903 42823 -28880 42857
rect -28960 42537 -28880 42823
rect -28960 42503 -28937 42537
rect -28903 42503 -28880 42537
rect -28960 42217 -28880 42503
rect -28960 42183 -28937 42217
rect -28903 42183 -28880 42217
rect -28960 41897 -28880 42183
rect -28960 41863 -28937 41897
rect -28903 41863 -28880 41897
rect -28960 41840 -28880 41863
rect -28800 42857 -28720 42880
rect -28800 42823 -28777 42857
rect -28743 42823 -28720 42857
rect -28800 42537 -28720 42823
rect -28800 42503 -28777 42537
rect -28743 42503 -28720 42537
rect -28800 42217 -28720 42503
rect -28800 42183 -28777 42217
rect -28743 42183 -28720 42217
rect -28800 41897 -28720 42183
rect -28800 41863 -28777 41897
rect -28743 41863 -28720 41897
rect -28800 41840 -28720 41863
rect -28640 42857 -28560 42880
rect -28640 42823 -28617 42857
rect -28583 42823 -28560 42857
rect -28640 42537 -28560 42823
rect -28640 42503 -28617 42537
rect -28583 42503 -28560 42537
rect -28640 42217 -28560 42503
rect -28640 42183 -28617 42217
rect -28583 42183 -28560 42217
rect -28640 41897 -28560 42183
rect -28640 41863 -28617 41897
rect -28583 41863 -28560 41897
rect -28640 41840 -28560 41863
rect -28480 42857 -28400 42880
rect -28480 42823 -28457 42857
rect -28423 42823 -28400 42857
rect -28480 42537 -28400 42823
rect -28480 42503 -28457 42537
rect -28423 42503 -28400 42537
rect -28480 42217 -28400 42503
rect -28480 42183 -28457 42217
rect -28423 42183 -28400 42217
rect -28480 41897 -28400 42183
rect -28480 41863 -28457 41897
rect -28423 41863 -28400 41897
rect -28480 41840 -28400 41863
rect -28320 42857 -28240 42880
rect -28320 42823 -28297 42857
rect -28263 42823 -28240 42857
rect -28320 42537 -28240 42823
rect -28320 42503 -28297 42537
rect -28263 42503 -28240 42537
rect -28320 42217 -28240 42503
rect -28320 42183 -28297 42217
rect -28263 42183 -28240 42217
rect -28320 41897 -28240 42183
rect -28320 41863 -28297 41897
rect -28263 41863 -28240 41897
rect -28320 41840 -28240 41863
rect -28160 42857 -28080 42880
rect -28160 42823 -28137 42857
rect -28103 42823 -28080 42857
rect -28160 42537 -28080 42823
rect -28160 42503 -28137 42537
rect -28103 42503 -28080 42537
rect -28160 42217 -28080 42503
rect -28160 42183 -28137 42217
rect -28103 42183 -28080 42217
rect -28160 41897 -28080 42183
rect -28160 41863 -28137 41897
rect -28103 41863 -28080 41897
rect -28160 41840 -28080 41863
rect -28000 42857 -27920 42880
rect -28000 42823 -27977 42857
rect -27943 42823 -27920 42857
rect -28000 42537 -27920 42823
rect -28000 42503 -27977 42537
rect -27943 42503 -27920 42537
rect -28000 42217 -27920 42503
rect -28000 42183 -27977 42217
rect -27943 42183 -27920 42217
rect -28000 41897 -27920 42183
rect -28000 41863 -27977 41897
rect -27943 41863 -27920 41897
rect -28000 41840 -27920 41863
rect -27840 42857 -27760 42880
rect -27840 42823 -27817 42857
rect -27783 42823 -27760 42857
rect -27840 42537 -27760 42823
rect -27840 42503 -27817 42537
rect -27783 42503 -27760 42537
rect -27840 42217 -27760 42503
rect -27840 42183 -27817 42217
rect -27783 42183 -27760 42217
rect -27840 41897 -27760 42183
rect -27840 41863 -27817 41897
rect -27783 41863 -27760 41897
rect -27840 41840 -27760 41863
rect -27680 42857 -27600 42880
rect -27680 42823 -27657 42857
rect -27623 42823 -27600 42857
rect -27680 42537 -27600 42823
rect -27680 42503 -27657 42537
rect -27623 42503 -27600 42537
rect -27680 42217 -27600 42503
rect -27680 42183 -27657 42217
rect -27623 42183 -27600 42217
rect -27680 41897 -27600 42183
rect -27680 41863 -27657 41897
rect -27623 41863 -27600 41897
rect -27680 41840 -27600 41863
rect -27520 42857 -27440 42880
rect -27520 42823 -27497 42857
rect -27463 42823 -27440 42857
rect -27520 42537 -27440 42823
rect -27520 42503 -27497 42537
rect -27463 42503 -27440 42537
rect -27520 42217 -27440 42503
rect -27520 42183 -27497 42217
rect -27463 42183 -27440 42217
rect -27520 41897 -27440 42183
rect -27520 41863 -27497 41897
rect -27463 41863 -27440 41897
rect -27520 41840 -27440 41863
rect -27360 42857 -27280 42880
rect -27360 42823 -27337 42857
rect -27303 42823 -27280 42857
rect -27360 42537 -27280 42823
rect -27360 42503 -27337 42537
rect -27303 42503 -27280 42537
rect -27360 42217 -27280 42503
rect -27360 42183 -27337 42217
rect -27303 42183 -27280 42217
rect -27360 41897 -27280 42183
rect -27360 41863 -27337 41897
rect -27303 41863 -27280 41897
rect -27360 41840 -27280 41863
rect -27200 42857 -27120 42880
rect -27200 42823 -27177 42857
rect -27143 42823 -27120 42857
rect -27200 42537 -27120 42823
rect -27200 42503 -27177 42537
rect -27143 42503 -27120 42537
rect -27200 42217 -27120 42503
rect -27200 42183 -27177 42217
rect -27143 42183 -27120 42217
rect -27200 41897 -27120 42183
rect -27200 41863 -27177 41897
rect -27143 41863 -27120 41897
rect -27200 41840 -27120 41863
rect -27040 42857 -26960 42880
rect -27040 42823 -27017 42857
rect -26983 42823 -26960 42857
rect -27040 42537 -26960 42823
rect -27040 42503 -27017 42537
rect -26983 42503 -26960 42537
rect -27040 42217 -26960 42503
rect -27040 42183 -27017 42217
rect -26983 42183 -26960 42217
rect -27040 41897 -26960 42183
rect -27040 41863 -27017 41897
rect -26983 41863 -26960 41897
rect -27040 41840 -26960 41863
rect -26880 42857 -26800 42880
rect -26880 42823 -26857 42857
rect -26823 42823 -26800 42857
rect -26880 42537 -26800 42823
rect -26880 42503 -26857 42537
rect -26823 42503 -26800 42537
rect -26880 42217 -26800 42503
rect -26880 42183 -26857 42217
rect -26823 42183 -26800 42217
rect -26880 41897 -26800 42183
rect -26880 41863 -26857 41897
rect -26823 41863 -26800 41897
rect -26880 41840 -26800 41863
rect -26720 42857 -26640 42880
rect -26720 42823 -26697 42857
rect -26663 42823 -26640 42857
rect -26720 42537 -26640 42823
rect -26720 42503 -26697 42537
rect -26663 42503 -26640 42537
rect -26720 42217 -26640 42503
rect -26720 42183 -26697 42217
rect -26663 42183 -26640 42217
rect -26720 41897 -26640 42183
rect -26720 41863 -26697 41897
rect -26663 41863 -26640 41897
rect -26720 41840 -26640 41863
rect -26560 42857 -26480 42880
rect -26560 42823 -26537 42857
rect -26503 42823 -26480 42857
rect -26560 42537 -26480 42823
rect -26560 42503 -26537 42537
rect -26503 42503 -26480 42537
rect -26560 42217 -26480 42503
rect -26560 42183 -26537 42217
rect -26503 42183 -26480 42217
rect -26560 41897 -26480 42183
rect -26560 41863 -26537 41897
rect -26503 41863 -26480 41897
rect -26560 41840 -26480 41863
rect -26400 42857 -26320 42880
rect -26400 42823 -26377 42857
rect -26343 42823 -26320 42857
rect -26400 42537 -26320 42823
rect -26400 42503 -26377 42537
rect -26343 42503 -26320 42537
rect -26400 42217 -26320 42503
rect -26400 42183 -26377 42217
rect -26343 42183 -26320 42217
rect -26400 41897 -26320 42183
rect -26400 41863 -26377 41897
rect -26343 41863 -26320 41897
rect -26400 41840 -26320 41863
rect -26240 42857 -26160 42880
rect -26240 42823 -26217 42857
rect -26183 42823 -26160 42857
rect -26240 42537 -26160 42823
rect -26240 42503 -26217 42537
rect -26183 42503 -26160 42537
rect -26240 42217 -26160 42503
rect -26240 42183 -26217 42217
rect -26183 42183 -26160 42217
rect -26240 41897 -26160 42183
rect -26240 41863 -26217 41897
rect -26183 41863 -26160 41897
rect -26240 41840 -26160 41863
rect -26080 42857 -26000 42880
rect -26080 42823 -26057 42857
rect -26023 42823 -26000 42857
rect -26080 42537 -26000 42823
rect -26080 42503 -26057 42537
rect -26023 42503 -26000 42537
rect -26080 42217 -26000 42503
rect -26080 42183 -26057 42217
rect -26023 42183 -26000 42217
rect -26080 41897 -26000 42183
rect -26080 41863 -26057 41897
rect -26023 41863 -26000 41897
rect -26080 41840 -26000 41863
rect -25920 42857 -25840 42880
rect -25920 42823 -25897 42857
rect -25863 42823 -25840 42857
rect -25920 42537 -25840 42823
rect -25920 42503 -25897 42537
rect -25863 42503 -25840 42537
rect -25920 42217 -25840 42503
rect -25920 42183 -25897 42217
rect -25863 42183 -25840 42217
rect -25920 41897 -25840 42183
rect -25920 41863 -25897 41897
rect -25863 41863 -25840 41897
rect -25920 41840 -25840 41863
rect -25760 42857 -25680 42880
rect -25760 42823 -25737 42857
rect -25703 42823 -25680 42857
rect -25760 42537 -25680 42823
rect -25760 42503 -25737 42537
rect -25703 42503 -25680 42537
rect -25760 42217 -25680 42503
rect -25760 42183 -25737 42217
rect -25703 42183 -25680 42217
rect -25760 41897 -25680 42183
rect -25760 41863 -25737 41897
rect -25703 41863 -25680 41897
rect -25760 41840 -25680 41863
rect -25600 42857 -25520 42880
rect -25600 42823 -25577 42857
rect -25543 42823 -25520 42857
rect -25600 42537 -25520 42823
rect -25600 42503 -25577 42537
rect -25543 42503 -25520 42537
rect -25600 42217 -25520 42503
rect -25600 42183 -25577 42217
rect -25543 42183 -25520 42217
rect -25600 41897 -25520 42183
rect -25600 41863 -25577 41897
rect -25543 41863 -25520 41897
rect -25600 41840 -25520 41863
rect -25440 42857 -25360 42880
rect -25440 42823 -25417 42857
rect -25383 42823 -25360 42857
rect -25440 42537 -25360 42823
rect -25440 42503 -25417 42537
rect -25383 42503 -25360 42537
rect -25440 42217 -25360 42503
rect -25440 42183 -25417 42217
rect -25383 42183 -25360 42217
rect -25440 41897 -25360 42183
rect -25440 41863 -25417 41897
rect -25383 41863 -25360 41897
rect -25440 41840 -25360 41863
rect -25280 42857 -25200 42880
rect -25280 42823 -25257 42857
rect -25223 42823 -25200 42857
rect -25280 42537 -25200 42823
rect -25280 42503 -25257 42537
rect -25223 42503 -25200 42537
rect -25280 42217 -25200 42503
rect -25280 42183 -25257 42217
rect -25223 42183 -25200 42217
rect -25280 41897 -25200 42183
rect -25280 41863 -25257 41897
rect -25223 41863 -25200 41897
rect -25280 41840 -25200 41863
rect -25120 42857 -25040 42880
rect -25120 42823 -25097 42857
rect -25063 42823 -25040 42857
rect -25120 42537 -25040 42823
rect -25120 42503 -25097 42537
rect -25063 42503 -25040 42537
rect -25120 42217 -25040 42503
rect -25120 42183 -25097 42217
rect -25063 42183 -25040 42217
rect -25120 41897 -25040 42183
rect -25120 41863 -25097 41897
rect -25063 41863 -25040 41897
rect -25120 41840 -25040 41863
rect -24960 42857 -24880 42880
rect -24960 42823 -24937 42857
rect -24903 42823 -24880 42857
rect -24960 42537 -24880 42823
rect -24960 42503 -24937 42537
rect -24903 42503 -24880 42537
rect -24960 42217 -24880 42503
rect -24960 42183 -24937 42217
rect -24903 42183 -24880 42217
rect -24960 41897 -24880 42183
rect -24960 41863 -24937 41897
rect -24903 41863 -24880 41897
rect -24960 41840 -24880 41863
rect -24800 42857 -24720 42880
rect -24800 42823 -24777 42857
rect -24743 42823 -24720 42857
rect -24800 42537 -24720 42823
rect -24800 42503 -24777 42537
rect -24743 42503 -24720 42537
rect -24800 42217 -24720 42503
rect -24800 42183 -24777 42217
rect -24743 42183 -24720 42217
rect -24800 41897 -24720 42183
rect -24800 41863 -24777 41897
rect -24743 41863 -24720 41897
rect -24800 41840 -24720 41863
rect -24640 42857 -24560 42880
rect -24640 42823 -24617 42857
rect -24583 42823 -24560 42857
rect -24640 42537 -24560 42823
rect -24640 42503 -24617 42537
rect -24583 42503 -24560 42537
rect -24640 42217 -24560 42503
rect -24640 42183 -24617 42217
rect -24583 42183 -24560 42217
rect -24640 41897 -24560 42183
rect -24640 41863 -24617 41897
rect -24583 41863 -24560 41897
rect -24640 41840 -24560 41863
rect -24480 42857 -24400 42880
rect -24480 42823 -24457 42857
rect -24423 42823 -24400 42857
rect -24480 42537 -24400 42823
rect -24480 42503 -24457 42537
rect -24423 42503 -24400 42537
rect -24480 42217 -24400 42503
rect -24480 42183 -24457 42217
rect -24423 42183 -24400 42217
rect -24480 41897 -24400 42183
rect -24480 41863 -24457 41897
rect -24423 41863 -24400 41897
rect -24480 41840 -24400 41863
rect -24320 42857 -24240 42880
rect -24320 42823 -24297 42857
rect -24263 42823 -24240 42857
rect -24320 42537 -24240 42823
rect -24320 42503 -24297 42537
rect -24263 42503 -24240 42537
rect -24320 42217 -24240 42503
rect -24320 42183 -24297 42217
rect -24263 42183 -24240 42217
rect -24320 41897 -24240 42183
rect -24320 41863 -24297 41897
rect -24263 41863 -24240 41897
rect -24320 41840 -24240 41863
rect -24160 42857 -24080 42880
rect -24160 42823 -24137 42857
rect -24103 42823 -24080 42857
rect -24160 42537 -24080 42823
rect -24160 42503 -24137 42537
rect -24103 42503 -24080 42537
rect -24160 42217 -24080 42503
rect -24160 42183 -24137 42217
rect -24103 42183 -24080 42217
rect -24160 41897 -24080 42183
rect -24160 41863 -24137 41897
rect -24103 41863 -24080 41897
rect -24160 41840 -24080 41863
rect -24000 42857 -23920 42880
rect -24000 42823 -23977 42857
rect -23943 42823 -23920 42857
rect -24000 42537 -23920 42823
rect -24000 42503 -23977 42537
rect -23943 42503 -23920 42537
rect -24000 42217 -23920 42503
rect -24000 42183 -23977 42217
rect -23943 42183 -23920 42217
rect -24000 41897 -23920 42183
rect -24000 41863 -23977 41897
rect -23943 41863 -23920 41897
rect -24000 41840 -23920 41863
rect -23840 42857 -23760 42880
rect -23840 42823 -23817 42857
rect -23783 42823 -23760 42857
rect -23840 42537 -23760 42823
rect -23840 42503 -23817 42537
rect -23783 42503 -23760 42537
rect -23840 42217 -23760 42503
rect -23840 42183 -23817 42217
rect -23783 42183 -23760 42217
rect -23840 41897 -23760 42183
rect -23840 41863 -23817 41897
rect -23783 41863 -23760 41897
rect -23840 41840 -23760 41863
rect -23680 42857 -23600 42880
rect -23680 42823 -23657 42857
rect -23623 42823 -23600 42857
rect -23680 42537 -23600 42823
rect -23680 42503 -23657 42537
rect -23623 42503 -23600 42537
rect -23680 42217 -23600 42503
rect -23680 42183 -23657 42217
rect -23623 42183 -23600 42217
rect -23680 41897 -23600 42183
rect -23680 41863 -23657 41897
rect -23623 41863 -23600 41897
rect -23680 41840 -23600 41863
rect -23520 42857 -23440 42880
rect -23520 42823 -23497 42857
rect -23463 42823 -23440 42857
rect -23520 42537 -23440 42823
rect -23520 42503 -23497 42537
rect -23463 42503 -23440 42537
rect -23520 42217 -23440 42503
rect -23520 42183 -23497 42217
rect -23463 42183 -23440 42217
rect -23520 41897 -23440 42183
rect -23520 41863 -23497 41897
rect -23463 41863 -23440 41897
rect -23520 41840 -23440 41863
rect -23360 42857 -23280 42880
rect -23360 42823 -23337 42857
rect -23303 42823 -23280 42857
rect -23360 42537 -23280 42823
rect -23360 42503 -23337 42537
rect -23303 42503 -23280 42537
rect -23360 42217 -23280 42503
rect -23360 42183 -23337 42217
rect -23303 42183 -23280 42217
rect -23360 41897 -23280 42183
rect -23360 41863 -23337 41897
rect -23303 41863 -23280 41897
rect -23360 41840 -23280 41863
rect -23200 42857 -23120 42880
rect -23200 42823 -23177 42857
rect -23143 42823 -23120 42857
rect -23200 42537 -23120 42823
rect -23200 42503 -23177 42537
rect -23143 42503 -23120 42537
rect -23200 42217 -23120 42503
rect -23200 42183 -23177 42217
rect -23143 42183 -23120 42217
rect -23200 41897 -23120 42183
rect -23200 41863 -23177 41897
rect -23143 41863 -23120 41897
rect -23200 41840 -23120 41863
rect -23040 42857 -22960 42880
rect -23040 42823 -23017 42857
rect -22983 42823 -22960 42857
rect -23040 42537 -22960 42823
rect -23040 42503 -23017 42537
rect -22983 42503 -22960 42537
rect -23040 42217 -22960 42503
rect -23040 42183 -23017 42217
rect -22983 42183 -22960 42217
rect -23040 41897 -22960 42183
rect -23040 41863 -23017 41897
rect -22983 41863 -22960 41897
rect -23040 41840 -22960 41863
rect -22880 42857 -22800 42880
rect -22880 42823 -22857 42857
rect -22823 42823 -22800 42857
rect -22880 42537 -22800 42823
rect -22880 42503 -22857 42537
rect -22823 42503 -22800 42537
rect -22880 42217 -22800 42503
rect -22880 42183 -22857 42217
rect -22823 42183 -22800 42217
rect -22880 41897 -22800 42183
rect -22880 41863 -22857 41897
rect -22823 41863 -22800 41897
rect -22880 41840 -22800 41863
rect -22720 42857 -22640 42880
rect -22720 42823 -22697 42857
rect -22663 42823 -22640 42857
rect -22720 42537 -22640 42823
rect -22720 42503 -22697 42537
rect -22663 42503 -22640 42537
rect -22720 42217 -22640 42503
rect -22720 42183 -22697 42217
rect -22663 42183 -22640 42217
rect -22720 41897 -22640 42183
rect -22720 41863 -22697 41897
rect -22663 41863 -22640 41897
rect -22720 41840 -22640 41863
rect -22560 42857 -22480 42880
rect -22560 42823 -22537 42857
rect -22503 42823 -22480 42857
rect -22560 42537 -22480 42823
rect -22560 42503 -22537 42537
rect -22503 42503 -22480 42537
rect -22560 42217 -22480 42503
rect -22560 42183 -22537 42217
rect -22503 42183 -22480 42217
rect -22560 41897 -22480 42183
rect -22560 41863 -22537 41897
rect -22503 41863 -22480 41897
rect -22560 41840 -22480 41863
rect -22400 42857 -22320 42880
rect -22400 42823 -22377 42857
rect -22343 42823 -22320 42857
rect -22400 42537 -22320 42823
rect -22400 42503 -22377 42537
rect -22343 42503 -22320 42537
rect -22400 42217 -22320 42503
rect -22400 42183 -22377 42217
rect -22343 42183 -22320 42217
rect -22400 41897 -22320 42183
rect -22400 41863 -22377 41897
rect -22343 41863 -22320 41897
rect -22400 41840 -22320 41863
rect -22240 42857 -22160 42880
rect -22240 42823 -22217 42857
rect -22183 42823 -22160 42857
rect -22240 42537 -22160 42823
rect -22240 42503 -22217 42537
rect -22183 42503 -22160 42537
rect -22240 42217 -22160 42503
rect -22240 42183 -22217 42217
rect -22183 42183 -22160 42217
rect -22240 41897 -22160 42183
rect -22240 41863 -22217 41897
rect -22183 41863 -22160 41897
rect -22240 41840 -22160 41863
rect -22080 42857 -22000 42880
rect -22080 42823 -22057 42857
rect -22023 42823 -22000 42857
rect -22080 42537 -22000 42823
rect -22080 42503 -22057 42537
rect -22023 42503 -22000 42537
rect -22080 42217 -22000 42503
rect -22080 42183 -22057 42217
rect -22023 42183 -22000 42217
rect -22080 41897 -22000 42183
rect -22080 41863 -22057 41897
rect -22023 41863 -22000 41897
rect -22080 41840 -22000 41863
rect -21920 42857 -21840 42880
rect -21920 42823 -21897 42857
rect -21863 42823 -21840 42857
rect -21920 42537 -21840 42823
rect -21920 42503 -21897 42537
rect -21863 42503 -21840 42537
rect -21920 42217 -21840 42503
rect -21920 42183 -21897 42217
rect -21863 42183 -21840 42217
rect -21920 41897 -21840 42183
rect -21920 41863 -21897 41897
rect -21863 41863 -21840 41897
rect -21920 41840 -21840 41863
rect -21760 42857 -21680 42880
rect -21760 42823 -21737 42857
rect -21703 42823 -21680 42857
rect -21760 42537 -21680 42823
rect -21760 42503 -21737 42537
rect -21703 42503 -21680 42537
rect -21760 42217 -21680 42503
rect -21760 42183 -21737 42217
rect -21703 42183 -21680 42217
rect -21760 41897 -21680 42183
rect -21760 41863 -21737 41897
rect -21703 41863 -21680 41897
rect -21760 41840 -21680 41863
rect -21600 42857 -21520 42880
rect -21600 42823 -21577 42857
rect -21543 42823 -21520 42857
rect -21600 42537 -21520 42823
rect -21600 42503 -21577 42537
rect -21543 42503 -21520 42537
rect -21600 42217 -21520 42503
rect -21600 42183 -21577 42217
rect -21543 42183 -21520 42217
rect -21600 41897 -21520 42183
rect -21600 41863 -21577 41897
rect -21543 41863 -21520 41897
rect -21600 41840 -21520 41863
rect -21440 42857 -21360 42880
rect -21440 42823 -21417 42857
rect -21383 42823 -21360 42857
rect -21440 42537 -21360 42823
rect -21440 42503 -21417 42537
rect -21383 42503 -21360 42537
rect -21440 42217 -21360 42503
rect -21440 42183 -21417 42217
rect -21383 42183 -21360 42217
rect -21440 41897 -21360 42183
rect -21440 41863 -21417 41897
rect -21383 41863 -21360 41897
rect -21440 41840 -21360 41863
rect -21280 42857 -21200 42880
rect -21280 42823 -21257 42857
rect -21223 42823 -21200 42857
rect -21280 42537 -21200 42823
rect -21280 42503 -21257 42537
rect -21223 42503 -21200 42537
rect -21280 42217 -21200 42503
rect -21280 42183 -21257 42217
rect -21223 42183 -21200 42217
rect -21280 41897 -21200 42183
rect -21280 41863 -21257 41897
rect -21223 41863 -21200 41897
rect -21280 41840 -21200 41863
rect -21120 42857 -21040 42880
rect -21120 42823 -21097 42857
rect -21063 42823 -21040 42857
rect -21120 42537 -21040 42823
rect -21120 42503 -21097 42537
rect -21063 42503 -21040 42537
rect -21120 42217 -21040 42503
rect -21120 42183 -21097 42217
rect -21063 42183 -21040 42217
rect -21120 41897 -21040 42183
rect -21120 41863 -21097 41897
rect -21063 41863 -21040 41897
rect -21120 41840 -21040 41863
rect -20960 42857 -20880 42880
rect -20960 42823 -20937 42857
rect -20903 42823 -20880 42857
rect -20960 42537 -20880 42823
rect -20960 42503 -20937 42537
rect -20903 42503 -20880 42537
rect -20960 42217 -20880 42503
rect -20960 42183 -20937 42217
rect -20903 42183 -20880 42217
rect -20960 41897 -20880 42183
rect -20960 41863 -20937 41897
rect -20903 41863 -20880 41897
rect -20960 41840 -20880 41863
rect -20800 42857 -20720 42880
rect -20800 42823 -20777 42857
rect -20743 42823 -20720 42857
rect -20800 42537 -20720 42823
rect -20800 42503 -20777 42537
rect -20743 42503 -20720 42537
rect -20800 42217 -20720 42503
rect -20800 42183 -20777 42217
rect -20743 42183 -20720 42217
rect -20800 41897 -20720 42183
rect -20800 41863 -20777 41897
rect -20743 41863 -20720 41897
rect -20800 41840 -20720 41863
rect -20640 42857 -20560 42880
rect -20640 42823 -20617 42857
rect -20583 42823 -20560 42857
rect -20640 42537 -20560 42823
rect -20640 42503 -20617 42537
rect -20583 42503 -20560 42537
rect -20640 42217 -20560 42503
rect -20640 42183 -20617 42217
rect -20583 42183 -20560 42217
rect -20640 41897 -20560 42183
rect -20640 41863 -20617 41897
rect -20583 41863 -20560 41897
rect -20640 41840 -20560 41863
rect -20480 42857 -20400 42880
rect -20480 42823 -20457 42857
rect -20423 42823 -20400 42857
rect -20480 42537 -20400 42823
rect -20480 42503 -20457 42537
rect -20423 42503 -20400 42537
rect -20480 42217 -20400 42503
rect -20480 42183 -20457 42217
rect -20423 42183 -20400 42217
rect -20480 41897 -20400 42183
rect -20480 41863 -20457 41897
rect -20423 41863 -20400 41897
rect -20480 41840 -20400 41863
rect -20320 42857 -20240 42880
rect -20320 42823 -20297 42857
rect -20263 42823 -20240 42857
rect -20320 42537 -20240 42823
rect -20320 42503 -20297 42537
rect -20263 42503 -20240 42537
rect -20320 42217 -20240 42503
rect -20320 42183 -20297 42217
rect -20263 42183 -20240 42217
rect -20320 41897 -20240 42183
rect -20320 41863 -20297 41897
rect -20263 41863 -20240 41897
rect -20320 41840 -20240 41863
rect -20160 42857 -20080 42880
rect -20160 42823 -20137 42857
rect -20103 42823 -20080 42857
rect -20160 42537 -20080 42823
rect -20160 42503 -20137 42537
rect -20103 42503 -20080 42537
rect -20160 42217 -20080 42503
rect -20160 42183 -20137 42217
rect -20103 42183 -20080 42217
rect -20160 41897 -20080 42183
rect -20160 41863 -20137 41897
rect -20103 41863 -20080 41897
rect -20160 41840 -20080 41863
rect -20000 42857 -19920 42880
rect -20000 42823 -19977 42857
rect -19943 42823 -19920 42857
rect -20000 42537 -19920 42823
rect -20000 42503 -19977 42537
rect -19943 42503 -19920 42537
rect -20000 42217 -19920 42503
rect -20000 42183 -19977 42217
rect -19943 42183 -19920 42217
rect -20000 41897 -19920 42183
rect -20000 41863 -19977 41897
rect -19943 41863 -19920 41897
rect -20000 41840 -19920 41863
rect -19840 42857 -19760 42880
rect -19840 42823 -19817 42857
rect -19783 42823 -19760 42857
rect -19840 42537 -19760 42823
rect -19840 42503 -19817 42537
rect -19783 42503 -19760 42537
rect -19840 42217 -19760 42503
rect -19840 42183 -19817 42217
rect -19783 42183 -19760 42217
rect -19840 41897 -19760 42183
rect -19840 41863 -19817 41897
rect -19783 41863 -19760 41897
rect -19840 41840 -19760 41863
rect -19680 42857 -19600 42880
rect -19680 42823 -19657 42857
rect -19623 42823 -19600 42857
rect -19680 42537 -19600 42823
rect -19680 42503 -19657 42537
rect -19623 42503 -19600 42537
rect -19680 42217 -19600 42503
rect -19680 42183 -19657 42217
rect -19623 42183 -19600 42217
rect -19680 41897 -19600 42183
rect -19680 41863 -19657 41897
rect -19623 41863 -19600 41897
rect -19680 41840 -19600 41863
rect -19520 42857 -19440 42880
rect -19520 42823 -19497 42857
rect -19463 42823 -19440 42857
rect -19520 42537 -19440 42823
rect -19520 42503 -19497 42537
rect -19463 42503 -19440 42537
rect -19520 42217 -19440 42503
rect -19520 42183 -19497 42217
rect -19463 42183 -19440 42217
rect -19520 41897 -19440 42183
rect -19520 41863 -19497 41897
rect -19463 41863 -19440 41897
rect -19520 41840 -19440 41863
rect -19360 42857 -19280 42880
rect -19360 42823 -19337 42857
rect -19303 42823 -19280 42857
rect -19360 42537 -19280 42823
rect -19360 42503 -19337 42537
rect -19303 42503 -19280 42537
rect -19360 42217 -19280 42503
rect -19360 42183 -19337 42217
rect -19303 42183 -19280 42217
rect -19360 41897 -19280 42183
rect -19360 41863 -19337 41897
rect -19303 41863 -19280 41897
rect -19360 41840 -19280 41863
rect -19200 42857 -19120 42880
rect -19200 42823 -19177 42857
rect -19143 42823 -19120 42857
rect -19200 42537 -19120 42823
rect -19200 42503 -19177 42537
rect -19143 42503 -19120 42537
rect -19200 42217 -19120 42503
rect -19200 42183 -19177 42217
rect -19143 42183 -19120 42217
rect -19200 41897 -19120 42183
rect -19200 41863 -19177 41897
rect -19143 41863 -19120 41897
rect -19200 41840 -19120 41863
rect -19040 42857 -18960 42880
rect -19040 42823 -19017 42857
rect -18983 42823 -18960 42857
rect -19040 42537 -18960 42823
rect -19040 42503 -19017 42537
rect -18983 42503 -18960 42537
rect -19040 42217 -18960 42503
rect -19040 42183 -19017 42217
rect -18983 42183 -18960 42217
rect -19040 41897 -18960 42183
rect -19040 41863 -19017 41897
rect -18983 41863 -18960 41897
rect -19040 41840 -18960 41863
rect -18880 42857 -18800 42880
rect -18880 42823 -18857 42857
rect -18823 42823 -18800 42857
rect -18880 42537 -18800 42823
rect -18880 42503 -18857 42537
rect -18823 42503 -18800 42537
rect -18880 42217 -18800 42503
rect -18880 42183 -18857 42217
rect -18823 42183 -18800 42217
rect -18880 41897 -18800 42183
rect -18880 41863 -18857 41897
rect -18823 41863 -18800 41897
rect -18880 41840 -18800 41863
rect -18720 42857 -18640 42880
rect -18720 42823 -18697 42857
rect -18663 42823 -18640 42857
rect -18720 42537 -18640 42823
rect -18720 42503 -18697 42537
rect -18663 42503 -18640 42537
rect -18720 42217 -18640 42503
rect -18720 42183 -18697 42217
rect -18663 42183 -18640 42217
rect -18720 41897 -18640 42183
rect -18720 41863 -18697 41897
rect -18663 41863 -18640 41897
rect -18720 41840 -18640 41863
rect -18560 42857 -18480 42880
rect -18560 42823 -18537 42857
rect -18503 42823 -18480 42857
rect -18560 42537 -18480 42823
rect -18560 42503 -18537 42537
rect -18503 42503 -18480 42537
rect -18560 42217 -18480 42503
rect -18560 42183 -18537 42217
rect -18503 42183 -18480 42217
rect -18560 41897 -18480 42183
rect -18560 41863 -18537 41897
rect -18503 41863 -18480 41897
rect -18560 41840 -18480 41863
rect -18400 42857 -18320 42880
rect -18400 42823 -18377 42857
rect -18343 42823 -18320 42857
rect -18400 42537 -18320 42823
rect -18400 42503 -18377 42537
rect -18343 42503 -18320 42537
rect -18400 42217 -18320 42503
rect -18400 42183 -18377 42217
rect -18343 42183 -18320 42217
rect -18400 41897 -18320 42183
rect -18400 41863 -18377 41897
rect -18343 41863 -18320 41897
rect -18400 41840 -18320 41863
rect -18240 42857 -18160 42880
rect -18240 42823 -18217 42857
rect -18183 42823 -18160 42857
rect -18240 42537 -18160 42823
rect -18240 42503 -18217 42537
rect -18183 42503 -18160 42537
rect -18240 42217 -18160 42503
rect -18240 42183 -18217 42217
rect -18183 42183 -18160 42217
rect -18240 41897 -18160 42183
rect -18240 41863 -18217 41897
rect -18183 41863 -18160 41897
rect -18240 41840 -18160 41863
rect -18080 42857 -18000 42880
rect -18080 42823 -18057 42857
rect -18023 42823 -18000 42857
rect -18080 42537 -18000 42823
rect -18080 42503 -18057 42537
rect -18023 42503 -18000 42537
rect -18080 42217 -18000 42503
rect -18080 42183 -18057 42217
rect -18023 42183 -18000 42217
rect -18080 41897 -18000 42183
rect -18080 41863 -18057 41897
rect -18023 41863 -18000 41897
rect -18080 41840 -18000 41863
rect -17920 42857 -17840 42880
rect -17920 42823 -17897 42857
rect -17863 42823 -17840 42857
rect -17920 42537 -17840 42823
rect -17920 42503 -17897 42537
rect -17863 42503 -17840 42537
rect -17920 42217 -17840 42503
rect -17920 42183 -17897 42217
rect -17863 42183 -17840 42217
rect -17920 41897 -17840 42183
rect -17920 41863 -17897 41897
rect -17863 41863 -17840 41897
rect -17920 41840 -17840 41863
rect -17760 42857 -17680 42880
rect -17760 42823 -17737 42857
rect -17703 42823 -17680 42857
rect -17760 42537 -17680 42823
rect -17760 42503 -17737 42537
rect -17703 42503 -17680 42537
rect -17760 42217 -17680 42503
rect -17760 42183 -17737 42217
rect -17703 42183 -17680 42217
rect -17760 41897 -17680 42183
rect -17760 41863 -17737 41897
rect -17703 41863 -17680 41897
rect -17760 41840 -17680 41863
rect -17600 42857 -17520 42880
rect -17600 42823 -17577 42857
rect -17543 42823 -17520 42857
rect -17600 42537 -17520 42823
rect -17600 42503 -17577 42537
rect -17543 42503 -17520 42537
rect -17600 42217 -17520 42503
rect -17600 42183 -17577 42217
rect -17543 42183 -17520 42217
rect -17600 41897 -17520 42183
rect -17600 41863 -17577 41897
rect -17543 41863 -17520 41897
rect -17600 41840 -17520 41863
rect -17440 42857 -17360 42880
rect -17440 42823 -17417 42857
rect -17383 42823 -17360 42857
rect -17440 42537 -17360 42823
rect -17440 42503 -17417 42537
rect -17383 42503 -17360 42537
rect -17440 42217 -17360 42503
rect -17440 42183 -17417 42217
rect -17383 42183 -17360 42217
rect -17440 41897 -17360 42183
rect -17440 41863 -17417 41897
rect -17383 41863 -17360 41897
rect -17440 41840 -17360 41863
rect -17280 42857 -17200 42880
rect -17280 42823 -17257 42857
rect -17223 42823 -17200 42857
rect -17280 42537 -17200 42823
rect -17280 42503 -17257 42537
rect -17223 42503 -17200 42537
rect -17280 42217 -17200 42503
rect -17280 42183 -17257 42217
rect -17223 42183 -17200 42217
rect -17280 41897 -17200 42183
rect -17280 41863 -17257 41897
rect -17223 41863 -17200 41897
rect -17280 41840 -17200 41863
rect -17120 42857 -17040 42880
rect -17120 42823 -17097 42857
rect -17063 42823 -17040 42857
rect -17120 42537 -17040 42823
rect -17120 42503 -17097 42537
rect -17063 42503 -17040 42537
rect -17120 42217 -17040 42503
rect -17120 42183 -17097 42217
rect -17063 42183 -17040 42217
rect -17120 41897 -17040 42183
rect -17120 41863 -17097 41897
rect -17063 41863 -17040 41897
rect -17120 41840 -17040 41863
rect -16960 42857 -16880 42880
rect -16960 42823 -16937 42857
rect -16903 42823 -16880 42857
rect -16960 42537 -16880 42823
rect -16960 42503 -16937 42537
rect -16903 42503 -16880 42537
rect -16960 42217 -16880 42503
rect -16960 42183 -16937 42217
rect -16903 42183 -16880 42217
rect -16960 41897 -16880 42183
rect -16960 41863 -16937 41897
rect -16903 41863 -16880 41897
rect -16960 41840 -16880 41863
rect -16800 42857 -16720 42880
rect -16800 42823 -16777 42857
rect -16743 42823 -16720 42857
rect -16800 42537 -16720 42823
rect -16800 42503 -16777 42537
rect -16743 42503 -16720 42537
rect -16800 42217 -16720 42503
rect -16800 42183 -16777 42217
rect -16743 42183 -16720 42217
rect -16800 41897 -16720 42183
rect -16800 41863 -16777 41897
rect -16743 41863 -16720 41897
rect -16800 41840 -16720 41863
rect -16640 42857 -16560 42880
rect -16640 42823 -16617 42857
rect -16583 42823 -16560 42857
rect -16640 42537 -16560 42823
rect -16640 42503 -16617 42537
rect -16583 42503 -16560 42537
rect -16640 42217 -16560 42503
rect -16640 42183 -16617 42217
rect -16583 42183 -16560 42217
rect -16640 41897 -16560 42183
rect -16640 41863 -16617 41897
rect -16583 41863 -16560 41897
rect -16640 41840 -16560 41863
rect -16480 42857 -16400 42880
rect -16480 42823 -16457 42857
rect -16423 42823 -16400 42857
rect -16480 42537 -16400 42823
rect -16480 42503 -16457 42537
rect -16423 42503 -16400 42537
rect -16480 42217 -16400 42503
rect -16480 42183 -16457 42217
rect -16423 42183 -16400 42217
rect -16480 41897 -16400 42183
rect -16480 41863 -16457 41897
rect -16423 41863 -16400 41897
rect -16480 41840 -16400 41863
rect -16320 42857 -16240 42880
rect -16320 42823 -16297 42857
rect -16263 42823 -16240 42857
rect -16320 42537 -16240 42823
rect -16320 42503 -16297 42537
rect -16263 42503 -16240 42537
rect -16320 42217 -16240 42503
rect -16320 42183 -16297 42217
rect -16263 42183 -16240 42217
rect -16320 41897 -16240 42183
rect -16320 41863 -16297 41897
rect -16263 41863 -16240 41897
rect -16320 41840 -16240 41863
rect -16160 42857 -16080 42880
rect -16160 42823 -16137 42857
rect -16103 42823 -16080 42857
rect -16160 42537 -16080 42823
rect -16160 42503 -16137 42537
rect -16103 42503 -16080 42537
rect -16160 42217 -16080 42503
rect -16160 42183 -16137 42217
rect -16103 42183 -16080 42217
rect -16160 41897 -16080 42183
rect -16160 41863 -16137 41897
rect -16103 41863 -16080 41897
rect -16160 41840 -16080 41863
rect -16000 42857 -15920 42880
rect -16000 42823 -15977 42857
rect -15943 42823 -15920 42857
rect -16000 42537 -15920 42823
rect -16000 42503 -15977 42537
rect -15943 42503 -15920 42537
rect -16000 42217 -15920 42503
rect -16000 42183 -15977 42217
rect -15943 42183 -15920 42217
rect -16000 41897 -15920 42183
rect -16000 41863 -15977 41897
rect -15943 41863 -15920 41897
rect -16000 41840 -15920 41863
rect -15840 42857 -15760 42880
rect -15840 42823 -15817 42857
rect -15783 42823 -15760 42857
rect -15840 42537 -15760 42823
rect -15840 42503 -15817 42537
rect -15783 42503 -15760 42537
rect -15840 42217 -15760 42503
rect -15840 42183 -15817 42217
rect -15783 42183 -15760 42217
rect -15840 41897 -15760 42183
rect -15840 41863 -15817 41897
rect -15783 41863 -15760 41897
rect -15840 41840 -15760 41863
rect -15680 42857 -15600 42880
rect -15680 42823 -15657 42857
rect -15623 42823 -15600 42857
rect -15680 42537 -15600 42823
rect -15680 42503 -15657 42537
rect -15623 42503 -15600 42537
rect -15680 42217 -15600 42503
rect -15680 42183 -15657 42217
rect -15623 42183 -15600 42217
rect -15680 41897 -15600 42183
rect -15680 41863 -15657 41897
rect -15623 41863 -15600 41897
rect -15680 41840 -15600 41863
rect -15520 42857 -15440 42880
rect -15520 42823 -15497 42857
rect -15463 42823 -15440 42857
rect -15520 42537 -15440 42823
rect -15520 42503 -15497 42537
rect -15463 42503 -15440 42537
rect -15520 42217 -15440 42503
rect -15520 42183 -15497 42217
rect -15463 42183 -15440 42217
rect -15520 41897 -15440 42183
rect -15520 41863 -15497 41897
rect -15463 41863 -15440 41897
rect -15520 41840 -15440 41863
rect -15360 42857 -15280 42880
rect -15360 42823 -15337 42857
rect -15303 42823 -15280 42857
rect -15360 42537 -15280 42823
rect -15360 42503 -15337 42537
rect -15303 42503 -15280 42537
rect -15360 42217 -15280 42503
rect -15360 42183 -15337 42217
rect -15303 42183 -15280 42217
rect -15360 41897 -15280 42183
rect -15360 41863 -15337 41897
rect -15303 41863 -15280 41897
rect -15360 41840 -15280 41863
rect -15200 42857 -15120 42880
rect -15200 42823 -15177 42857
rect -15143 42823 -15120 42857
rect -15200 42537 -15120 42823
rect -15200 42503 -15177 42537
rect -15143 42503 -15120 42537
rect -15200 42217 -15120 42503
rect -15200 42183 -15177 42217
rect -15143 42183 -15120 42217
rect -15200 41897 -15120 42183
rect -15200 41863 -15177 41897
rect -15143 41863 -15120 41897
rect -15200 41840 -15120 41863
rect -15040 42857 -14960 42880
rect -15040 42823 -15017 42857
rect -14983 42823 -14960 42857
rect -15040 42537 -14960 42823
rect -15040 42503 -15017 42537
rect -14983 42503 -14960 42537
rect -15040 42217 -14960 42503
rect -15040 42183 -15017 42217
rect -14983 42183 -14960 42217
rect -15040 41897 -14960 42183
rect -15040 41863 -15017 41897
rect -14983 41863 -14960 41897
rect -15040 41840 -14960 41863
rect -14880 42857 -14800 42880
rect -14880 42823 -14857 42857
rect -14823 42823 -14800 42857
rect -14880 42537 -14800 42823
rect -14880 42503 -14857 42537
rect -14823 42503 -14800 42537
rect -14880 42217 -14800 42503
rect -14880 42183 -14857 42217
rect -14823 42183 -14800 42217
rect -14880 41897 -14800 42183
rect -14880 41863 -14857 41897
rect -14823 41863 -14800 41897
rect -14880 41840 -14800 41863
rect -14720 42857 -14640 42880
rect -14720 42823 -14697 42857
rect -14663 42823 -14640 42857
rect -14720 42537 -14640 42823
rect -14720 42503 -14697 42537
rect -14663 42503 -14640 42537
rect -14720 42217 -14640 42503
rect -14720 42183 -14697 42217
rect -14663 42183 -14640 42217
rect -14720 41897 -14640 42183
rect -14720 41863 -14697 41897
rect -14663 41863 -14640 41897
rect -14720 41840 -14640 41863
rect -14560 42857 -14480 42880
rect -14560 42823 -14537 42857
rect -14503 42823 -14480 42857
rect -14560 42537 -14480 42823
rect -14560 42503 -14537 42537
rect -14503 42503 -14480 42537
rect -14560 42217 -14480 42503
rect -14560 42183 -14537 42217
rect -14503 42183 -14480 42217
rect -14560 41897 -14480 42183
rect -14560 41863 -14537 41897
rect -14503 41863 -14480 41897
rect -14560 41840 -14480 41863
rect -14400 42857 -14320 42880
rect -14400 42823 -14377 42857
rect -14343 42823 -14320 42857
rect -14400 42537 -14320 42823
rect -14400 42503 -14377 42537
rect -14343 42503 -14320 42537
rect -14400 42217 -14320 42503
rect -14400 42183 -14377 42217
rect -14343 42183 -14320 42217
rect -14400 41897 -14320 42183
rect -14400 41863 -14377 41897
rect -14343 41863 -14320 41897
rect -14400 41840 -14320 41863
rect -14240 42857 -14160 42880
rect -14240 42823 -14217 42857
rect -14183 42823 -14160 42857
rect -14240 42537 -14160 42823
rect -14240 42503 -14217 42537
rect -14183 42503 -14160 42537
rect -14240 42217 -14160 42503
rect -14240 42183 -14217 42217
rect -14183 42183 -14160 42217
rect -14240 41897 -14160 42183
rect -14240 41863 -14217 41897
rect -14183 41863 -14160 41897
rect -14240 41840 -14160 41863
rect -14080 42857 -14000 42880
rect -14080 42823 -14057 42857
rect -14023 42823 -14000 42857
rect -14080 42537 -14000 42823
rect -14080 42503 -14057 42537
rect -14023 42503 -14000 42537
rect -14080 42217 -14000 42503
rect -14080 42183 -14057 42217
rect -14023 42183 -14000 42217
rect -14080 41897 -14000 42183
rect -14080 41863 -14057 41897
rect -14023 41863 -14000 41897
rect -14080 41840 -14000 41863
rect -13920 42857 -13840 42880
rect -13920 42823 -13897 42857
rect -13863 42823 -13840 42857
rect -13920 42537 -13840 42823
rect -13920 42503 -13897 42537
rect -13863 42503 -13840 42537
rect -13920 42217 -13840 42503
rect -13920 42183 -13897 42217
rect -13863 42183 -13840 42217
rect -13920 41897 -13840 42183
rect -13920 41863 -13897 41897
rect -13863 41863 -13840 41897
rect -13920 41840 -13840 41863
rect -13760 42857 -13680 42880
rect -13760 42823 -13737 42857
rect -13703 42823 -13680 42857
rect -13760 42537 -13680 42823
rect -13760 42503 -13737 42537
rect -13703 42503 -13680 42537
rect -13760 42217 -13680 42503
rect -13760 42183 -13737 42217
rect -13703 42183 -13680 42217
rect -13760 41897 -13680 42183
rect -13760 41863 -13737 41897
rect -13703 41863 -13680 41897
rect -13760 41840 -13680 41863
rect -13600 42857 -13520 42880
rect -13600 42823 -13577 42857
rect -13543 42823 -13520 42857
rect -13600 42537 -13520 42823
rect -13600 42503 -13577 42537
rect -13543 42503 -13520 42537
rect -13600 42217 -13520 42503
rect -13600 42183 -13577 42217
rect -13543 42183 -13520 42217
rect -13600 41897 -13520 42183
rect -13600 41863 -13577 41897
rect -13543 41863 -13520 41897
rect -13600 41840 -13520 41863
rect -13440 42857 -13360 42880
rect -13440 42823 -13417 42857
rect -13383 42823 -13360 42857
rect -13440 42537 -13360 42823
rect -13440 42503 -13417 42537
rect -13383 42503 -13360 42537
rect -13440 42217 -13360 42503
rect -13440 42183 -13417 42217
rect -13383 42183 -13360 42217
rect -13440 41897 -13360 42183
rect -13440 41863 -13417 41897
rect -13383 41863 -13360 41897
rect -13440 41840 -13360 41863
rect -13280 42857 -13200 42880
rect -13280 42823 -13257 42857
rect -13223 42823 -13200 42857
rect -13280 42537 -13200 42823
rect -13280 42503 -13257 42537
rect -13223 42503 -13200 42537
rect -13280 42217 -13200 42503
rect -13280 42183 -13257 42217
rect -13223 42183 -13200 42217
rect -13280 41897 -13200 42183
rect -13280 41863 -13257 41897
rect -13223 41863 -13200 41897
rect -13280 41840 -13200 41863
rect -13120 42857 -13040 42880
rect -13120 42823 -13097 42857
rect -13063 42823 -13040 42857
rect -13120 42537 -13040 42823
rect -13120 42503 -13097 42537
rect -13063 42503 -13040 42537
rect -13120 42217 -13040 42503
rect -13120 42183 -13097 42217
rect -13063 42183 -13040 42217
rect -13120 41897 -13040 42183
rect -13120 41863 -13097 41897
rect -13063 41863 -13040 41897
rect -13120 41840 -13040 41863
rect -12960 42857 -12880 42880
rect -12960 42823 -12937 42857
rect -12903 42823 -12880 42857
rect -12960 42537 -12880 42823
rect -12960 42503 -12937 42537
rect -12903 42503 -12880 42537
rect -12960 42217 -12880 42503
rect -12960 42183 -12937 42217
rect -12903 42183 -12880 42217
rect -12960 41897 -12880 42183
rect -12960 41863 -12937 41897
rect -12903 41863 -12880 41897
rect -12960 41840 -12880 41863
rect -12800 42857 -12720 42880
rect -12800 42823 -12777 42857
rect -12743 42823 -12720 42857
rect -12800 42537 -12720 42823
rect -12800 42503 -12777 42537
rect -12743 42503 -12720 42537
rect -12800 42217 -12720 42503
rect -12800 42183 -12777 42217
rect -12743 42183 -12720 42217
rect -12800 41897 -12720 42183
rect -12800 41863 -12777 41897
rect -12743 41863 -12720 41897
rect -12800 41840 -12720 41863
rect -12640 42857 -12560 42880
rect -12640 42823 -12617 42857
rect -12583 42823 -12560 42857
rect -12640 42537 -12560 42823
rect -12640 42503 -12617 42537
rect -12583 42503 -12560 42537
rect -12640 42217 -12560 42503
rect -12640 42183 -12617 42217
rect -12583 42183 -12560 42217
rect -12640 41897 -12560 42183
rect -12640 41863 -12617 41897
rect -12583 41863 -12560 41897
rect -12640 41840 -12560 41863
rect -12480 42857 -12400 42880
rect -12480 42823 -12457 42857
rect -12423 42823 -12400 42857
rect -12480 42537 -12400 42823
rect -12480 42503 -12457 42537
rect -12423 42503 -12400 42537
rect -12480 42217 -12400 42503
rect -12480 42183 -12457 42217
rect -12423 42183 -12400 42217
rect -12480 41897 -12400 42183
rect -12480 41863 -12457 41897
rect -12423 41863 -12400 41897
rect -12480 41840 -12400 41863
rect -12320 42857 -12240 42880
rect -12320 42823 -12297 42857
rect -12263 42823 -12240 42857
rect -12320 42537 -12240 42823
rect -12320 42503 -12297 42537
rect -12263 42503 -12240 42537
rect -12320 42217 -12240 42503
rect -12320 42183 -12297 42217
rect -12263 42183 -12240 42217
rect -12320 41897 -12240 42183
rect -12320 41863 -12297 41897
rect -12263 41863 -12240 41897
rect -12320 41840 -12240 41863
rect -11360 42857 -11280 42880
rect -11360 42823 -11337 42857
rect -11303 42823 -11280 42857
rect -11360 42537 -11280 42823
rect -11360 42503 -11337 42537
rect -11303 42503 -11280 42537
rect -11360 42217 -11280 42503
rect -11360 42183 -11337 42217
rect -11303 42183 -11280 42217
rect -11360 41897 -11280 42183
rect -11360 41863 -11337 41897
rect -11303 41863 -11280 41897
rect -11360 41840 -11280 41863
rect -11200 42857 -11120 42880
rect -11200 42823 -11177 42857
rect -11143 42823 -11120 42857
rect -11200 42537 -11120 42823
rect -11200 42503 -11177 42537
rect -11143 42503 -11120 42537
rect -11200 42217 -11120 42503
rect -11200 42183 -11177 42217
rect -11143 42183 -11120 42217
rect -11200 41897 -11120 42183
rect -11200 41863 -11177 41897
rect -11143 41863 -11120 41897
rect -11200 41840 -11120 41863
rect -11040 42857 -10960 42880
rect -11040 42823 -11017 42857
rect -10983 42823 -10960 42857
rect -11040 42537 -10960 42823
rect -11040 42503 -11017 42537
rect -10983 42503 -10960 42537
rect -11040 42217 -10960 42503
rect -11040 42183 -11017 42217
rect -10983 42183 -10960 42217
rect -11040 41897 -10960 42183
rect -11040 41863 -11017 41897
rect -10983 41863 -10960 41897
rect -11040 41840 -10960 41863
rect -10880 42857 -10800 42880
rect -10880 42823 -10857 42857
rect -10823 42823 -10800 42857
rect -10880 42537 -10800 42823
rect -10880 42503 -10857 42537
rect -10823 42503 -10800 42537
rect -10880 42217 -10800 42503
rect -10880 42183 -10857 42217
rect -10823 42183 -10800 42217
rect -10880 41897 -10800 42183
rect -10880 41863 -10857 41897
rect -10823 41863 -10800 41897
rect -10880 41840 -10800 41863
rect -10720 42857 -10640 42880
rect -10720 42823 -10697 42857
rect -10663 42823 -10640 42857
rect -10720 42537 -10640 42823
rect -10720 42503 -10697 42537
rect -10663 42503 -10640 42537
rect -10720 42217 -10640 42503
rect -10720 42183 -10697 42217
rect -10663 42183 -10640 42217
rect -10720 41897 -10640 42183
rect -10720 41863 -10697 41897
rect -10663 41863 -10640 41897
rect -10720 41840 -10640 41863
rect -10560 42857 -10480 42880
rect -10560 42823 -10537 42857
rect -10503 42823 -10480 42857
rect -10560 42537 -10480 42823
rect -10560 42503 -10537 42537
rect -10503 42503 -10480 42537
rect -10560 42217 -10480 42503
rect -10560 42183 -10537 42217
rect -10503 42183 -10480 42217
rect -10560 41897 -10480 42183
rect -10560 41863 -10537 41897
rect -10503 41863 -10480 41897
rect -10560 41840 -10480 41863
rect -10400 42857 -10320 42880
rect -10400 42823 -10377 42857
rect -10343 42823 -10320 42857
rect -10400 42537 -10320 42823
rect -10400 42503 -10377 42537
rect -10343 42503 -10320 42537
rect -10400 42217 -10320 42503
rect -10400 42183 -10377 42217
rect -10343 42183 -10320 42217
rect -10400 41897 -10320 42183
rect -10400 41863 -10377 41897
rect -10343 41863 -10320 41897
rect -10400 41840 -10320 41863
rect -10240 42857 -10160 42880
rect -10240 42823 -10217 42857
rect -10183 42823 -10160 42857
rect -10240 42537 -10160 42823
rect -10240 42503 -10217 42537
rect -10183 42503 -10160 42537
rect -10240 42217 -10160 42503
rect -10240 42183 -10217 42217
rect -10183 42183 -10160 42217
rect -10240 41897 -10160 42183
rect -10240 41863 -10217 41897
rect -10183 41863 -10160 41897
rect -10240 41840 -10160 41863
rect -10080 42857 -10000 42880
rect -10080 42823 -10057 42857
rect -10023 42823 -10000 42857
rect -10080 42537 -10000 42823
rect -10080 42503 -10057 42537
rect -10023 42503 -10000 42537
rect -10080 42217 -10000 42503
rect -10080 42183 -10057 42217
rect -10023 42183 -10000 42217
rect -10080 41897 -10000 42183
rect -10080 41863 -10057 41897
rect -10023 41863 -10000 41897
rect -10080 41840 -10000 41863
rect -9920 42857 -9840 42880
rect -9920 42823 -9897 42857
rect -9863 42823 -9840 42857
rect -9920 42537 -9840 42823
rect -9920 42503 -9897 42537
rect -9863 42503 -9840 42537
rect -9920 42217 -9840 42503
rect -9920 42183 -9897 42217
rect -9863 42183 -9840 42217
rect -9920 41897 -9840 42183
rect -9920 41863 -9897 41897
rect -9863 41863 -9840 41897
rect -9920 41840 -9840 41863
rect -9760 42857 -9680 42880
rect -9760 42823 -9737 42857
rect -9703 42823 -9680 42857
rect -9760 42537 -9680 42823
rect -9760 42503 -9737 42537
rect -9703 42503 -9680 42537
rect -9760 42217 -9680 42503
rect -9760 42183 -9737 42217
rect -9703 42183 -9680 42217
rect -9760 41897 -9680 42183
rect -9760 41863 -9737 41897
rect -9703 41863 -9680 41897
rect -9760 41840 -9680 41863
rect -9600 42857 -9520 42880
rect -9600 42823 -9577 42857
rect -9543 42823 -9520 42857
rect -9600 42537 -9520 42823
rect -9600 42503 -9577 42537
rect -9543 42503 -9520 42537
rect -9600 42217 -9520 42503
rect -9600 42183 -9577 42217
rect -9543 42183 -9520 42217
rect -9600 41897 -9520 42183
rect -9600 41863 -9577 41897
rect -9543 41863 -9520 41897
rect -9600 41840 -9520 41863
rect -9440 42857 -9360 42880
rect -9440 42823 -9417 42857
rect -9383 42823 -9360 42857
rect -9440 42537 -9360 42823
rect -9440 42503 -9417 42537
rect -9383 42503 -9360 42537
rect -9440 42217 -9360 42503
rect -9440 42183 -9417 42217
rect -9383 42183 -9360 42217
rect -9440 41897 -9360 42183
rect -9440 41863 -9417 41897
rect -9383 41863 -9360 41897
rect -9440 41840 -9360 41863
rect -9280 42857 -9200 42880
rect -9280 42823 -9257 42857
rect -9223 42823 -9200 42857
rect -9280 42537 -9200 42823
rect -9280 42503 -9257 42537
rect -9223 42503 -9200 42537
rect -9280 42217 -9200 42503
rect -9280 42183 -9257 42217
rect -9223 42183 -9200 42217
rect -9280 41897 -9200 42183
rect -9280 41863 -9257 41897
rect -9223 41863 -9200 41897
rect -9280 41840 -9200 41863
rect -9120 42857 -9040 42880
rect -9120 42823 -9097 42857
rect -9063 42823 -9040 42857
rect -9120 42537 -9040 42823
rect -9120 42503 -9097 42537
rect -9063 42503 -9040 42537
rect -9120 42217 -9040 42503
rect -9120 42183 -9097 42217
rect -9063 42183 -9040 42217
rect -9120 41897 -9040 42183
rect -9120 41863 -9097 41897
rect -9063 41863 -9040 41897
rect -9120 41840 -9040 41863
rect -8960 42857 -8880 42880
rect -8960 42823 -8937 42857
rect -8903 42823 -8880 42857
rect -8960 42537 -8880 42823
rect -8960 42503 -8937 42537
rect -8903 42503 -8880 42537
rect -8960 42217 -8880 42503
rect -8960 42183 -8937 42217
rect -8903 42183 -8880 42217
rect -8960 41897 -8880 42183
rect -8960 41863 -8937 41897
rect -8903 41863 -8880 41897
rect -8960 41840 -8880 41863
rect -8800 42857 -8720 42880
rect -8800 42823 -8777 42857
rect -8743 42823 -8720 42857
rect -8800 42537 -8720 42823
rect -8800 42503 -8777 42537
rect -8743 42503 -8720 42537
rect -8800 42217 -8720 42503
rect -8800 42183 -8777 42217
rect -8743 42183 -8720 42217
rect -8800 41897 -8720 42183
rect -8800 41863 -8777 41897
rect -8743 41863 -8720 41897
rect -8800 41840 -8720 41863
rect -8640 42857 -8560 42880
rect -8640 42823 -8617 42857
rect -8583 42823 -8560 42857
rect -8640 42537 -8560 42823
rect -8640 42503 -8617 42537
rect -8583 42503 -8560 42537
rect -8640 42217 -8560 42503
rect -8640 42183 -8617 42217
rect -8583 42183 -8560 42217
rect -8640 41897 -8560 42183
rect -8640 41863 -8617 41897
rect -8583 41863 -8560 41897
rect -8640 41840 -8560 41863
rect -8480 42857 -8400 42880
rect -8480 42823 -8457 42857
rect -8423 42823 -8400 42857
rect -8480 42537 -8400 42823
rect -8480 42503 -8457 42537
rect -8423 42503 -8400 42537
rect -8480 42217 -8400 42503
rect -8480 42183 -8457 42217
rect -8423 42183 -8400 42217
rect -8480 41897 -8400 42183
rect -8480 41863 -8457 41897
rect -8423 41863 -8400 41897
rect -8480 41840 -8400 41863
rect -8320 42857 -8240 42880
rect -8320 42823 -8297 42857
rect -8263 42823 -8240 42857
rect -8320 42537 -8240 42823
rect -8320 42503 -8297 42537
rect -8263 42503 -8240 42537
rect -8320 42217 -8240 42503
rect -8320 42183 -8297 42217
rect -8263 42183 -8240 42217
rect -8320 41897 -8240 42183
rect -8320 41863 -8297 41897
rect -8263 41863 -8240 41897
rect -8320 41840 -8240 41863
rect -8160 42857 -8080 42880
rect -8160 42823 -8137 42857
rect -8103 42823 -8080 42857
rect -8160 42537 -8080 42823
rect -8160 42503 -8137 42537
rect -8103 42503 -8080 42537
rect -8160 42217 -8080 42503
rect -8160 42183 -8137 42217
rect -8103 42183 -8080 42217
rect -8160 41897 -8080 42183
rect -8160 41863 -8137 41897
rect -8103 41863 -8080 41897
rect -8160 41840 -8080 41863
rect -8000 42857 -7920 42880
rect -8000 42823 -7977 42857
rect -7943 42823 -7920 42857
rect -8000 42537 -7920 42823
rect -8000 42503 -7977 42537
rect -7943 42503 -7920 42537
rect -8000 42217 -7920 42503
rect -8000 42183 -7977 42217
rect -7943 42183 -7920 42217
rect -8000 41897 -7920 42183
rect -8000 41863 -7977 41897
rect -7943 41863 -7920 41897
rect -8000 41840 -7920 41863
rect -7840 42857 -7760 42880
rect -7840 42823 -7817 42857
rect -7783 42823 -7760 42857
rect -7840 42537 -7760 42823
rect -7840 42503 -7817 42537
rect -7783 42503 -7760 42537
rect -7840 42217 -7760 42503
rect -7840 42183 -7817 42217
rect -7783 42183 -7760 42217
rect -7840 41897 -7760 42183
rect -7840 41863 -7817 41897
rect -7783 41863 -7760 41897
rect -7840 41840 -7760 41863
rect -7680 42857 -7600 42880
rect -7680 42823 -7657 42857
rect -7623 42823 -7600 42857
rect -7680 42537 -7600 42823
rect -7680 42503 -7657 42537
rect -7623 42503 -7600 42537
rect -7680 42217 -7600 42503
rect -7680 42183 -7657 42217
rect -7623 42183 -7600 42217
rect -7680 41897 -7600 42183
rect -7680 41863 -7657 41897
rect -7623 41863 -7600 41897
rect -7680 41840 -7600 41863
rect -7520 42857 -7440 42880
rect -7520 42823 -7497 42857
rect -7463 42823 -7440 42857
rect -7520 42537 -7440 42823
rect -7520 42503 -7497 42537
rect -7463 42503 -7440 42537
rect -7520 42217 -7440 42503
rect -7520 42183 -7497 42217
rect -7463 42183 -7440 42217
rect -7520 41897 -7440 42183
rect -7520 41863 -7497 41897
rect -7463 41863 -7440 41897
rect -7520 41840 -7440 41863
rect -7360 42857 -7280 42880
rect -7360 42823 -7337 42857
rect -7303 42823 -7280 42857
rect -7360 42537 -7280 42823
rect -7360 42503 -7337 42537
rect -7303 42503 -7280 42537
rect -7360 42217 -7280 42503
rect -7360 42183 -7337 42217
rect -7303 42183 -7280 42217
rect -7360 41897 -7280 42183
rect -7360 41863 -7337 41897
rect -7303 41863 -7280 41897
rect -7360 41840 -7280 41863
rect -7200 42857 -7120 42880
rect -7200 42823 -7177 42857
rect -7143 42823 -7120 42857
rect -7200 42537 -7120 42823
rect -7200 42503 -7177 42537
rect -7143 42503 -7120 42537
rect -7200 42217 -7120 42503
rect -7200 42183 -7177 42217
rect -7143 42183 -7120 42217
rect -7200 41897 -7120 42183
rect -7200 41863 -7177 41897
rect -7143 41863 -7120 41897
rect -7200 41840 -7120 41863
rect -7040 42857 -6960 42880
rect -7040 42823 -7017 42857
rect -6983 42823 -6960 42857
rect -7040 42537 -6960 42823
rect -7040 42503 -7017 42537
rect -6983 42503 -6960 42537
rect -7040 42217 -6960 42503
rect -7040 42183 -7017 42217
rect -6983 42183 -6960 42217
rect -7040 41897 -6960 42183
rect -7040 41863 -7017 41897
rect -6983 41863 -6960 41897
rect -7040 41840 -6960 41863
rect -6880 42857 -6800 42880
rect -6880 42823 -6857 42857
rect -6823 42823 -6800 42857
rect -6880 42537 -6800 42823
rect -6880 42503 -6857 42537
rect -6823 42503 -6800 42537
rect -6880 42217 -6800 42503
rect -6880 42183 -6857 42217
rect -6823 42183 -6800 42217
rect -6880 41897 -6800 42183
rect -6880 41863 -6857 41897
rect -6823 41863 -6800 41897
rect -6880 41840 -6800 41863
rect -6720 42857 -6640 42880
rect -6720 42823 -6697 42857
rect -6663 42823 -6640 42857
rect -6720 42537 -6640 42823
rect -6720 42503 -6697 42537
rect -6663 42503 -6640 42537
rect -6720 42217 -6640 42503
rect -6720 42183 -6697 42217
rect -6663 42183 -6640 42217
rect -6720 41897 -6640 42183
rect -6720 41863 -6697 41897
rect -6663 41863 -6640 41897
rect -6720 41840 -6640 41863
rect -6560 42857 -6480 42880
rect -6560 42823 -6537 42857
rect -6503 42823 -6480 42857
rect -6560 42537 -6480 42823
rect -6560 42503 -6537 42537
rect -6503 42503 -6480 42537
rect -6560 42217 -6480 42503
rect -6560 42183 -6537 42217
rect -6503 42183 -6480 42217
rect -6560 41897 -6480 42183
rect -6560 41863 -6537 41897
rect -6503 41863 -6480 41897
rect -6560 41840 -6480 41863
rect -6400 42857 -6320 42880
rect -6400 42823 -6377 42857
rect -6343 42823 -6320 42857
rect -6400 42537 -6320 42823
rect -6400 42503 -6377 42537
rect -6343 42503 -6320 42537
rect -6400 42217 -6320 42503
rect -6400 42183 -6377 42217
rect -6343 42183 -6320 42217
rect -6400 41897 -6320 42183
rect -6400 41863 -6377 41897
rect -6343 41863 -6320 41897
rect -6400 41840 -6320 41863
rect -6240 42857 -6160 42880
rect -6240 42823 -6217 42857
rect -6183 42823 -6160 42857
rect -6240 42537 -6160 42823
rect -6240 42503 -6217 42537
rect -6183 42503 -6160 42537
rect -6240 42217 -6160 42503
rect -6240 42183 -6217 42217
rect -6183 42183 -6160 42217
rect -6240 41897 -6160 42183
rect -6240 41863 -6217 41897
rect -6183 41863 -6160 41897
rect -6240 41840 -6160 41863
rect -6080 42857 -6000 42880
rect -6080 42823 -6057 42857
rect -6023 42823 -6000 42857
rect -6080 42537 -6000 42823
rect -6080 42503 -6057 42537
rect -6023 42503 -6000 42537
rect -6080 42217 -6000 42503
rect -6080 42183 -6057 42217
rect -6023 42183 -6000 42217
rect -6080 41897 -6000 42183
rect -6080 41863 -6057 41897
rect -6023 41863 -6000 41897
rect -6080 41840 -6000 41863
rect -5920 42857 -5840 42880
rect -5920 42823 -5897 42857
rect -5863 42823 -5840 42857
rect -5920 42537 -5840 42823
rect -5920 42503 -5897 42537
rect -5863 42503 -5840 42537
rect -5920 42217 -5840 42503
rect -5920 42183 -5897 42217
rect -5863 42183 -5840 42217
rect -5920 41897 -5840 42183
rect -5920 41863 -5897 41897
rect -5863 41863 -5840 41897
rect -5920 41840 -5840 41863
rect -5760 42857 -5680 42880
rect -5760 42823 -5737 42857
rect -5703 42823 -5680 42857
rect -5760 42537 -5680 42823
rect -5760 42503 -5737 42537
rect -5703 42503 -5680 42537
rect -5760 42217 -5680 42503
rect -5760 42183 -5737 42217
rect -5703 42183 -5680 42217
rect -5760 41897 -5680 42183
rect -5760 41863 -5737 41897
rect -5703 41863 -5680 41897
rect -5760 41840 -5680 41863
rect -5600 42857 -5520 42880
rect -5600 42823 -5577 42857
rect -5543 42823 -5520 42857
rect -5600 42537 -5520 42823
rect -5600 42503 -5577 42537
rect -5543 42503 -5520 42537
rect -5600 42217 -5520 42503
rect -5600 42183 -5577 42217
rect -5543 42183 -5520 42217
rect -5600 41897 -5520 42183
rect -5600 41863 -5577 41897
rect -5543 41863 -5520 41897
rect -5600 41840 -5520 41863
rect -5440 42857 -5360 42880
rect -5440 42823 -5417 42857
rect -5383 42823 -5360 42857
rect -5440 42537 -5360 42823
rect -5440 42503 -5417 42537
rect -5383 42503 -5360 42537
rect -5440 42217 -5360 42503
rect -5440 42183 -5417 42217
rect -5383 42183 -5360 42217
rect -5440 41897 -5360 42183
rect -5440 41863 -5417 41897
rect -5383 41863 -5360 41897
rect -5440 41840 -5360 41863
rect -5280 42857 -5200 42880
rect -5280 42823 -5257 42857
rect -5223 42823 -5200 42857
rect -5280 42537 -5200 42823
rect -5280 42503 -5257 42537
rect -5223 42503 -5200 42537
rect -5280 42217 -5200 42503
rect -5280 42183 -5257 42217
rect -5223 42183 -5200 42217
rect -5280 41897 -5200 42183
rect -5280 41863 -5257 41897
rect -5223 41863 -5200 41897
rect -5280 41840 -5200 41863
rect -5120 42857 -5040 42880
rect -5120 42823 -5097 42857
rect -5063 42823 -5040 42857
rect -5120 42537 -5040 42823
rect -5120 42503 -5097 42537
rect -5063 42503 -5040 42537
rect -5120 42217 -5040 42503
rect -5120 42183 -5097 42217
rect -5063 42183 -5040 42217
rect -5120 41897 -5040 42183
rect -5120 41863 -5097 41897
rect -5063 41863 -5040 41897
rect -5120 41840 -5040 41863
rect -4960 42857 -4880 42880
rect -4960 42823 -4937 42857
rect -4903 42823 -4880 42857
rect -4960 42537 -4880 42823
rect -4960 42503 -4937 42537
rect -4903 42503 -4880 42537
rect -4960 42217 -4880 42503
rect -4960 42183 -4937 42217
rect -4903 42183 -4880 42217
rect -4960 41897 -4880 42183
rect -4960 41863 -4937 41897
rect -4903 41863 -4880 41897
rect -4960 41840 -4880 41863
rect -4800 42857 -4720 42880
rect -4800 42823 -4777 42857
rect -4743 42823 -4720 42857
rect -4800 42537 -4720 42823
rect -4800 42503 -4777 42537
rect -4743 42503 -4720 42537
rect -4800 42217 -4720 42503
rect -4800 42183 -4777 42217
rect -4743 42183 -4720 42217
rect -4800 41897 -4720 42183
rect -4800 41863 -4777 41897
rect -4743 41863 -4720 41897
rect -4800 41840 -4720 41863
rect -4640 42857 -4560 42880
rect -4640 42823 -4617 42857
rect -4583 42823 -4560 42857
rect -4640 42537 -4560 42823
rect -4640 42503 -4617 42537
rect -4583 42503 -4560 42537
rect -4640 42217 -4560 42503
rect -4640 42183 -4617 42217
rect -4583 42183 -4560 42217
rect -4640 41897 -4560 42183
rect -4640 41863 -4617 41897
rect -4583 41863 -4560 41897
rect -4640 41840 -4560 41863
rect -4480 42857 -4400 42880
rect -4480 42823 -4457 42857
rect -4423 42823 -4400 42857
rect -4480 42537 -4400 42823
rect -4480 42503 -4457 42537
rect -4423 42503 -4400 42537
rect -4480 42217 -4400 42503
rect -4480 42183 -4457 42217
rect -4423 42183 -4400 42217
rect -4480 41897 -4400 42183
rect -4480 41863 -4457 41897
rect -4423 41863 -4400 41897
rect -4480 41840 -4400 41863
rect -4320 42857 -4240 42880
rect -4320 42823 -4297 42857
rect -4263 42823 -4240 42857
rect -4320 42537 -4240 42823
rect -4320 42503 -4297 42537
rect -4263 42503 -4240 42537
rect -4320 42217 -4240 42503
rect -4320 42183 -4297 42217
rect -4263 42183 -4240 42217
rect -4320 41897 -4240 42183
rect -4320 41863 -4297 41897
rect -4263 41863 -4240 41897
rect -4320 41840 -4240 41863
rect -4160 42857 -4080 42880
rect -4160 42823 -4137 42857
rect -4103 42823 -4080 42857
rect -4160 42537 -4080 42823
rect -4160 42503 -4137 42537
rect -4103 42503 -4080 42537
rect -4160 42217 -4080 42503
rect -4160 42183 -4137 42217
rect -4103 42183 -4080 42217
rect -4160 41897 -4080 42183
rect -4160 41863 -4137 41897
rect -4103 41863 -4080 41897
rect -4160 41840 -4080 41863
rect -4000 42857 -3920 42880
rect -4000 42823 -3977 42857
rect -3943 42823 -3920 42857
rect -4000 42537 -3920 42823
rect -4000 42503 -3977 42537
rect -3943 42503 -3920 42537
rect -4000 42217 -3920 42503
rect -4000 42183 -3977 42217
rect -3943 42183 -3920 42217
rect -4000 41897 -3920 42183
rect -4000 41863 -3977 41897
rect -3943 41863 -3920 41897
rect -4000 41840 -3920 41863
rect -33120 41337 -33040 41360
rect -33120 41303 -33097 41337
rect -33063 41303 -33040 41337
rect -33120 41017 -33040 41303
rect -33120 40983 -33097 41017
rect -33063 40983 -33040 41017
rect -33120 40960 -33040 40983
rect -32960 41337 -32880 41360
rect -32960 41303 -32937 41337
rect -32903 41303 -32880 41337
rect -32960 41017 -32880 41303
rect -32960 40983 -32937 41017
rect -32903 40983 -32880 41017
rect -32960 40960 -32880 40983
rect -32800 41337 -32720 41360
rect -32800 41303 -32777 41337
rect -32743 41303 -32720 41337
rect -32800 41017 -32720 41303
rect -32800 40983 -32777 41017
rect -32743 40983 -32720 41017
rect -32800 40960 -32720 40983
rect -32640 41337 -32560 41360
rect -32640 41303 -32617 41337
rect -32583 41303 -32560 41337
rect -32640 41017 -32560 41303
rect -32640 40983 -32617 41017
rect -32583 40983 -32560 41017
rect -32640 40960 -32560 40983
rect -32480 41337 -32400 41360
rect -32480 41303 -32457 41337
rect -32423 41303 -32400 41337
rect -32480 41017 -32400 41303
rect -32480 40983 -32457 41017
rect -32423 40983 -32400 41017
rect -32480 40960 -32400 40983
rect -32320 41337 -32240 41360
rect -32320 41303 -32297 41337
rect -32263 41303 -32240 41337
rect -32320 41017 -32240 41303
rect -32320 40983 -32297 41017
rect -32263 40983 -32240 41017
rect -32320 40960 -32240 40983
rect -32160 41337 -32080 41360
rect -32160 41303 -32137 41337
rect -32103 41303 -32080 41337
rect -32160 41017 -32080 41303
rect -32160 40983 -32137 41017
rect -32103 40983 -32080 41017
rect -32160 40960 -32080 40983
rect -32000 41337 -31920 41360
rect -32000 41303 -31977 41337
rect -31943 41303 -31920 41337
rect -32000 41017 -31920 41303
rect -32000 40983 -31977 41017
rect -31943 40983 -31920 41017
rect -32000 40960 -31920 40983
rect -31840 41337 -31760 41360
rect -31840 41303 -31817 41337
rect -31783 41303 -31760 41337
rect -31840 41017 -31760 41303
rect -31840 40983 -31817 41017
rect -31783 40983 -31760 41017
rect -31840 40960 -31760 40983
rect -31680 41337 -31600 41360
rect -31680 41303 -31657 41337
rect -31623 41303 -31600 41337
rect -31680 41017 -31600 41303
rect -31680 40983 -31657 41017
rect -31623 40983 -31600 41017
rect -31680 40960 -31600 40983
rect -31520 41337 -31440 41360
rect -31520 41303 -31497 41337
rect -31463 41303 -31440 41337
rect -31520 41017 -31440 41303
rect -31520 40983 -31497 41017
rect -31463 40983 -31440 41017
rect -31520 40960 -31440 40983
rect -31360 41337 -31280 41360
rect -31360 41303 -31337 41337
rect -31303 41303 -31280 41337
rect -31360 41017 -31280 41303
rect -31360 40983 -31337 41017
rect -31303 40983 -31280 41017
rect -31360 40960 -31280 40983
rect -31200 41337 -31120 41360
rect -31200 41303 -31177 41337
rect -31143 41303 -31120 41337
rect -31200 41017 -31120 41303
rect -31200 40983 -31177 41017
rect -31143 40983 -31120 41017
rect -31200 40960 -31120 40983
rect -29920 41337 -29840 41360
rect -29920 41303 -29897 41337
rect -29863 41303 -29840 41337
rect -29920 41017 -29840 41303
rect -29920 40983 -29897 41017
rect -29863 40983 -29840 41017
rect -29920 40960 -29840 40983
rect -29760 41337 -29680 41360
rect -29760 41303 -29737 41337
rect -29703 41303 -29680 41337
rect -29760 41017 -29680 41303
rect -29760 40983 -29737 41017
rect -29703 40983 -29680 41017
rect -29760 40960 -29680 40983
rect -29600 41337 -29520 41360
rect -29600 41303 -29577 41337
rect -29543 41303 -29520 41337
rect -29600 41017 -29520 41303
rect -29600 40983 -29577 41017
rect -29543 40983 -29520 41017
rect -29600 40960 -29520 40983
rect -29440 41337 -29360 41360
rect -29440 41303 -29417 41337
rect -29383 41303 -29360 41337
rect -29440 41017 -29360 41303
rect -29440 40983 -29417 41017
rect -29383 40983 -29360 41017
rect -29440 40960 -29360 40983
rect -29280 41337 -29200 41360
rect -29280 41303 -29257 41337
rect -29223 41303 -29200 41337
rect -29280 41017 -29200 41303
rect -29280 40983 -29257 41017
rect -29223 40983 -29200 41017
rect -29280 40960 -29200 40983
rect -29120 41337 -29040 41360
rect -29120 41303 -29097 41337
rect -29063 41303 -29040 41337
rect -29120 41017 -29040 41303
rect -29120 40983 -29097 41017
rect -29063 40983 -29040 41017
rect -29120 40960 -29040 40983
rect -28960 41337 -28880 41360
rect -28960 41303 -28937 41337
rect -28903 41303 -28880 41337
rect -28960 41017 -28880 41303
rect -28960 40983 -28937 41017
rect -28903 40983 -28880 41017
rect -28960 40960 -28880 40983
rect -28800 41337 -28720 41360
rect -28800 41303 -28777 41337
rect -28743 41303 -28720 41337
rect -28800 41017 -28720 41303
rect -28800 40983 -28777 41017
rect -28743 40983 -28720 41017
rect -28800 40960 -28720 40983
rect -28640 41337 -28560 41360
rect -28640 41303 -28617 41337
rect -28583 41303 -28560 41337
rect -28640 41017 -28560 41303
rect -28640 40983 -28617 41017
rect -28583 40983 -28560 41017
rect -28640 40960 -28560 40983
rect -28480 41337 -28400 41360
rect -28480 41303 -28457 41337
rect -28423 41303 -28400 41337
rect -28480 41017 -28400 41303
rect -28480 40983 -28457 41017
rect -28423 40983 -28400 41017
rect -28480 40960 -28400 40983
rect -28320 41337 -28240 41360
rect -28320 41303 -28297 41337
rect -28263 41303 -28240 41337
rect -28320 41017 -28240 41303
rect -28320 40983 -28297 41017
rect -28263 40983 -28240 41017
rect -28320 40960 -28240 40983
rect -28160 41337 -28080 41360
rect -28160 41303 -28137 41337
rect -28103 41303 -28080 41337
rect -28160 41017 -28080 41303
rect -28160 40983 -28137 41017
rect -28103 40983 -28080 41017
rect -28160 40960 -28080 40983
rect -28000 41337 -27920 41360
rect -28000 41303 -27977 41337
rect -27943 41303 -27920 41337
rect -28000 41017 -27920 41303
rect -28000 40983 -27977 41017
rect -27943 40983 -27920 41017
rect -28000 40960 -27920 40983
rect -27840 41337 -27760 41360
rect -27840 41303 -27817 41337
rect -27783 41303 -27760 41337
rect -27840 41017 -27760 41303
rect -27840 40983 -27817 41017
rect -27783 40983 -27760 41017
rect -27840 40960 -27760 40983
rect -27680 41337 -27600 41360
rect -27680 41303 -27657 41337
rect -27623 41303 -27600 41337
rect -27680 41017 -27600 41303
rect -27680 40983 -27657 41017
rect -27623 40983 -27600 41017
rect -27680 40960 -27600 40983
rect -27520 41337 -27440 41360
rect -27520 41303 -27497 41337
rect -27463 41303 -27440 41337
rect -27520 41017 -27440 41303
rect -27520 40983 -27497 41017
rect -27463 40983 -27440 41017
rect -27520 40960 -27440 40983
rect -27360 41337 -27280 41360
rect -27360 41303 -27337 41337
rect -27303 41303 -27280 41337
rect -27360 41017 -27280 41303
rect -27360 40983 -27337 41017
rect -27303 40983 -27280 41017
rect -27360 40960 -27280 40983
rect -27200 41337 -27120 41360
rect -27200 41303 -27177 41337
rect -27143 41303 -27120 41337
rect -27200 41017 -27120 41303
rect -27200 40983 -27177 41017
rect -27143 40983 -27120 41017
rect -27200 40960 -27120 40983
rect -27040 41337 -26960 41360
rect -27040 41303 -27017 41337
rect -26983 41303 -26960 41337
rect -27040 41017 -26960 41303
rect -27040 40983 -27017 41017
rect -26983 40983 -26960 41017
rect -27040 40960 -26960 40983
rect -26880 41337 -26800 41360
rect -26880 41303 -26857 41337
rect -26823 41303 -26800 41337
rect -26880 41017 -26800 41303
rect -26880 40983 -26857 41017
rect -26823 40983 -26800 41017
rect -26880 40960 -26800 40983
rect -26720 41337 -26640 41360
rect -26720 41303 -26697 41337
rect -26663 41303 -26640 41337
rect -26720 41017 -26640 41303
rect -26720 40983 -26697 41017
rect -26663 40983 -26640 41017
rect -26720 40960 -26640 40983
rect -26560 41337 -26480 41360
rect -26560 41303 -26537 41337
rect -26503 41303 -26480 41337
rect -26560 41017 -26480 41303
rect -26560 40983 -26537 41017
rect -26503 40983 -26480 41017
rect -26560 40960 -26480 40983
rect -26400 41337 -26320 41360
rect -26400 41303 -26377 41337
rect -26343 41303 -26320 41337
rect -26400 41017 -26320 41303
rect -26400 40983 -26377 41017
rect -26343 40983 -26320 41017
rect -26400 40960 -26320 40983
rect -26240 41337 -26160 41360
rect -26240 41303 -26217 41337
rect -26183 41303 -26160 41337
rect -26240 41017 -26160 41303
rect -26240 40983 -26217 41017
rect -26183 40983 -26160 41017
rect -26240 40960 -26160 40983
rect -26080 41337 -26000 41360
rect -26080 41303 -26057 41337
rect -26023 41303 -26000 41337
rect -26080 41017 -26000 41303
rect -26080 40983 -26057 41017
rect -26023 40983 -26000 41017
rect -26080 40960 -26000 40983
rect -25920 41337 -25840 41360
rect -25920 41303 -25897 41337
rect -25863 41303 -25840 41337
rect -25920 41017 -25840 41303
rect -25920 40983 -25897 41017
rect -25863 40983 -25840 41017
rect -25920 40960 -25840 40983
rect -25760 41337 -25680 41360
rect -25760 41303 -25737 41337
rect -25703 41303 -25680 41337
rect -25760 41017 -25680 41303
rect -25760 40983 -25737 41017
rect -25703 40983 -25680 41017
rect -25760 40960 -25680 40983
rect -25600 41337 -25520 41360
rect -25600 41303 -25577 41337
rect -25543 41303 -25520 41337
rect -25600 41017 -25520 41303
rect -25600 40983 -25577 41017
rect -25543 40983 -25520 41017
rect -25600 40960 -25520 40983
rect -25440 41337 -25360 41360
rect -25440 41303 -25417 41337
rect -25383 41303 -25360 41337
rect -25440 41017 -25360 41303
rect -25440 40983 -25417 41017
rect -25383 40983 -25360 41017
rect -25440 40960 -25360 40983
rect -25280 41337 -25200 41360
rect -25280 41303 -25257 41337
rect -25223 41303 -25200 41337
rect -25280 41017 -25200 41303
rect -25280 40983 -25257 41017
rect -25223 40983 -25200 41017
rect -25280 40960 -25200 40983
rect -25120 41337 -25040 41360
rect -25120 41303 -25097 41337
rect -25063 41303 -25040 41337
rect -25120 41017 -25040 41303
rect -25120 40983 -25097 41017
rect -25063 40983 -25040 41017
rect -25120 40960 -25040 40983
rect -24960 41337 -24880 41360
rect -24960 41303 -24937 41337
rect -24903 41303 -24880 41337
rect -24960 41017 -24880 41303
rect -24960 40983 -24937 41017
rect -24903 40983 -24880 41017
rect -24960 40960 -24880 40983
rect -24800 41337 -24720 41360
rect -24800 41303 -24777 41337
rect -24743 41303 -24720 41337
rect -24800 41017 -24720 41303
rect -24800 40983 -24777 41017
rect -24743 40983 -24720 41017
rect -24800 40960 -24720 40983
rect -24640 41337 -24560 41360
rect -24640 41303 -24617 41337
rect -24583 41303 -24560 41337
rect -24640 41017 -24560 41303
rect -24640 40983 -24617 41017
rect -24583 40983 -24560 41017
rect -24640 40960 -24560 40983
rect -24480 41337 -24400 41360
rect -24480 41303 -24457 41337
rect -24423 41303 -24400 41337
rect -24480 41017 -24400 41303
rect -24480 40983 -24457 41017
rect -24423 40983 -24400 41017
rect -24480 40960 -24400 40983
rect -24320 41337 -24240 41360
rect -24320 41303 -24297 41337
rect -24263 41303 -24240 41337
rect -24320 41017 -24240 41303
rect -24320 40983 -24297 41017
rect -24263 40983 -24240 41017
rect -24320 40960 -24240 40983
rect -24160 41337 -24080 41360
rect -24160 41303 -24137 41337
rect -24103 41303 -24080 41337
rect -24160 41017 -24080 41303
rect -24160 40983 -24137 41017
rect -24103 40983 -24080 41017
rect -24160 40960 -24080 40983
rect -24000 41337 -23920 41360
rect -24000 41303 -23977 41337
rect -23943 41303 -23920 41337
rect -24000 41017 -23920 41303
rect -24000 40983 -23977 41017
rect -23943 40983 -23920 41017
rect -24000 40960 -23920 40983
rect -23840 41337 -23760 41360
rect -23840 41303 -23817 41337
rect -23783 41303 -23760 41337
rect -23840 41017 -23760 41303
rect -23840 40983 -23817 41017
rect -23783 40983 -23760 41017
rect -23840 40960 -23760 40983
rect -23680 41337 -23600 41360
rect -23680 41303 -23657 41337
rect -23623 41303 -23600 41337
rect -23680 41017 -23600 41303
rect -23680 40983 -23657 41017
rect -23623 40983 -23600 41017
rect -23680 40960 -23600 40983
rect -23520 41337 -23440 41360
rect -23520 41303 -23497 41337
rect -23463 41303 -23440 41337
rect -23520 41017 -23440 41303
rect -23520 40983 -23497 41017
rect -23463 40983 -23440 41017
rect -23520 40960 -23440 40983
rect -23360 41337 -23280 41360
rect -23360 41303 -23337 41337
rect -23303 41303 -23280 41337
rect -23360 41017 -23280 41303
rect -23360 40983 -23337 41017
rect -23303 40983 -23280 41017
rect -23360 40960 -23280 40983
rect -23200 41337 -23120 41360
rect -23200 41303 -23177 41337
rect -23143 41303 -23120 41337
rect -23200 41017 -23120 41303
rect -23200 40983 -23177 41017
rect -23143 40983 -23120 41017
rect -23200 40960 -23120 40983
rect -23040 41337 -22960 41360
rect -23040 41303 -23017 41337
rect -22983 41303 -22960 41337
rect -23040 41017 -22960 41303
rect -23040 40983 -23017 41017
rect -22983 40983 -22960 41017
rect -23040 40960 -22960 40983
rect -22880 41337 -22800 41360
rect -22880 41303 -22857 41337
rect -22823 41303 -22800 41337
rect -22880 41017 -22800 41303
rect -22880 40983 -22857 41017
rect -22823 40983 -22800 41017
rect -22880 40960 -22800 40983
rect -22720 41337 -22640 41360
rect -22720 41303 -22697 41337
rect -22663 41303 -22640 41337
rect -22720 41017 -22640 41303
rect -22720 40983 -22697 41017
rect -22663 40983 -22640 41017
rect -22720 40960 -22640 40983
rect -22560 41337 -22480 41360
rect -22560 41303 -22537 41337
rect -22503 41303 -22480 41337
rect -22560 41017 -22480 41303
rect -22560 40983 -22537 41017
rect -22503 40983 -22480 41017
rect -22560 40960 -22480 40983
rect -22400 41337 -22320 41360
rect -22400 41303 -22377 41337
rect -22343 41303 -22320 41337
rect -22400 41017 -22320 41303
rect -22400 40983 -22377 41017
rect -22343 40983 -22320 41017
rect -22400 40960 -22320 40983
rect -22240 41337 -22160 41360
rect -22240 41303 -22217 41337
rect -22183 41303 -22160 41337
rect -22240 41017 -22160 41303
rect -22240 40983 -22217 41017
rect -22183 40983 -22160 41017
rect -22240 40960 -22160 40983
rect -22080 41337 -22000 41360
rect -22080 41303 -22057 41337
rect -22023 41303 -22000 41337
rect -22080 41017 -22000 41303
rect -22080 40983 -22057 41017
rect -22023 40983 -22000 41017
rect -22080 40960 -22000 40983
rect -21920 41337 -21840 41360
rect -21920 41303 -21897 41337
rect -21863 41303 -21840 41337
rect -21920 41017 -21840 41303
rect -21920 40983 -21897 41017
rect -21863 40983 -21840 41017
rect -21920 40960 -21840 40983
rect -21760 41337 -21680 41360
rect -21760 41303 -21737 41337
rect -21703 41303 -21680 41337
rect -21760 41017 -21680 41303
rect -21760 40983 -21737 41017
rect -21703 40983 -21680 41017
rect -21760 40960 -21680 40983
rect -21600 41337 -21520 41360
rect -21600 41303 -21577 41337
rect -21543 41303 -21520 41337
rect -21600 41017 -21520 41303
rect -21600 40983 -21577 41017
rect -21543 40983 -21520 41017
rect -21600 40960 -21520 40983
rect -21440 41337 -21360 41360
rect -21440 41303 -21417 41337
rect -21383 41303 -21360 41337
rect -21440 41017 -21360 41303
rect -21440 40983 -21417 41017
rect -21383 40983 -21360 41017
rect -21440 40960 -21360 40983
rect -21280 41337 -21200 41360
rect -21280 41303 -21257 41337
rect -21223 41303 -21200 41337
rect -21280 41017 -21200 41303
rect -21280 40983 -21257 41017
rect -21223 40983 -21200 41017
rect -21280 40960 -21200 40983
rect -21120 41337 -21040 41360
rect -21120 41303 -21097 41337
rect -21063 41303 -21040 41337
rect -21120 41017 -21040 41303
rect -21120 40983 -21097 41017
rect -21063 40983 -21040 41017
rect -21120 40960 -21040 40983
rect -20960 41337 -20880 41360
rect -20960 41303 -20937 41337
rect -20903 41303 -20880 41337
rect -20960 41017 -20880 41303
rect -20960 40983 -20937 41017
rect -20903 40983 -20880 41017
rect -20960 40960 -20880 40983
rect -20800 41337 -20720 41360
rect -20800 41303 -20777 41337
rect -20743 41303 -20720 41337
rect -20800 41017 -20720 41303
rect -20800 40983 -20777 41017
rect -20743 40983 -20720 41017
rect -20800 40960 -20720 40983
rect -20640 41337 -20560 41360
rect -20640 41303 -20617 41337
rect -20583 41303 -20560 41337
rect -20640 41017 -20560 41303
rect -20640 40983 -20617 41017
rect -20583 40983 -20560 41017
rect -20640 40960 -20560 40983
rect -20480 41337 -20400 41360
rect -20480 41303 -20457 41337
rect -20423 41303 -20400 41337
rect -20480 41017 -20400 41303
rect -20480 40983 -20457 41017
rect -20423 40983 -20400 41017
rect -20480 40960 -20400 40983
rect -20320 41337 -20240 41360
rect -20320 41303 -20297 41337
rect -20263 41303 -20240 41337
rect -20320 41017 -20240 41303
rect -20320 40983 -20297 41017
rect -20263 40983 -20240 41017
rect -20320 40960 -20240 40983
rect -20160 41337 -20080 41360
rect -20160 41303 -20137 41337
rect -20103 41303 -20080 41337
rect -20160 41017 -20080 41303
rect -20160 40983 -20137 41017
rect -20103 40983 -20080 41017
rect -20160 40960 -20080 40983
rect -20000 41337 -19920 41360
rect -20000 41303 -19977 41337
rect -19943 41303 -19920 41337
rect -20000 41017 -19920 41303
rect -20000 40983 -19977 41017
rect -19943 40983 -19920 41017
rect -20000 40960 -19920 40983
rect -19840 41337 -19760 41360
rect -19840 41303 -19817 41337
rect -19783 41303 -19760 41337
rect -19840 41017 -19760 41303
rect -19840 40983 -19817 41017
rect -19783 40983 -19760 41017
rect -19840 40960 -19760 40983
rect -19680 41337 -19600 41360
rect -19680 41303 -19657 41337
rect -19623 41303 -19600 41337
rect -19680 41017 -19600 41303
rect -19680 40983 -19657 41017
rect -19623 40983 -19600 41017
rect -19680 40960 -19600 40983
rect -19520 41337 -19440 41360
rect -19520 41303 -19497 41337
rect -19463 41303 -19440 41337
rect -19520 41017 -19440 41303
rect -19520 40983 -19497 41017
rect -19463 40983 -19440 41017
rect -19520 40960 -19440 40983
rect -19360 41337 -19280 41360
rect -19360 41303 -19337 41337
rect -19303 41303 -19280 41337
rect -19360 41017 -19280 41303
rect -19360 40983 -19337 41017
rect -19303 40983 -19280 41017
rect -19360 40960 -19280 40983
rect -19200 41337 -19120 41360
rect -19200 41303 -19177 41337
rect -19143 41303 -19120 41337
rect -19200 41017 -19120 41303
rect -19200 40983 -19177 41017
rect -19143 40983 -19120 41017
rect -19200 40960 -19120 40983
rect -19040 41337 -18960 41360
rect -19040 41303 -19017 41337
rect -18983 41303 -18960 41337
rect -19040 41017 -18960 41303
rect -19040 40983 -19017 41017
rect -18983 40983 -18960 41017
rect -19040 40960 -18960 40983
rect -18880 41337 -18800 41360
rect -18880 41303 -18857 41337
rect -18823 41303 -18800 41337
rect -18880 41017 -18800 41303
rect -18880 40983 -18857 41017
rect -18823 40983 -18800 41017
rect -18880 40960 -18800 40983
rect -18720 41337 -18640 41360
rect -18720 41303 -18697 41337
rect -18663 41303 -18640 41337
rect -18720 41017 -18640 41303
rect -18720 40983 -18697 41017
rect -18663 40983 -18640 41017
rect -18720 40960 -18640 40983
rect -18560 41337 -18480 41360
rect -18560 41303 -18537 41337
rect -18503 41303 -18480 41337
rect -18560 41017 -18480 41303
rect -18560 40983 -18537 41017
rect -18503 40983 -18480 41017
rect -18560 40960 -18480 40983
rect -18400 41337 -18320 41360
rect -18400 41303 -18377 41337
rect -18343 41303 -18320 41337
rect -18400 41017 -18320 41303
rect -18400 40983 -18377 41017
rect -18343 40983 -18320 41017
rect -18400 40960 -18320 40983
rect -18240 41337 -18160 41360
rect -18240 41303 -18217 41337
rect -18183 41303 -18160 41337
rect -18240 41017 -18160 41303
rect -18240 40983 -18217 41017
rect -18183 40983 -18160 41017
rect -18240 40960 -18160 40983
rect -18080 41337 -18000 41360
rect -18080 41303 -18057 41337
rect -18023 41303 -18000 41337
rect -18080 41017 -18000 41303
rect -18080 40983 -18057 41017
rect -18023 40983 -18000 41017
rect -18080 40960 -18000 40983
rect -17920 41337 -17840 41360
rect -17920 41303 -17897 41337
rect -17863 41303 -17840 41337
rect -17920 41017 -17840 41303
rect -17920 40983 -17897 41017
rect -17863 40983 -17840 41017
rect -17920 40960 -17840 40983
rect -17760 41337 -17680 41360
rect -17760 41303 -17737 41337
rect -17703 41303 -17680 41337
rect -17760 41017 -17680 41303
rect -17760 40983 -17737 41017
rect -17703 40983 -17680 41017
rect -17760 40960 -17680 40983
rect -17600 41337 -17520 41360
rect -17600 41303 -17577 41337
rect -17543 41303 -17520 41337
rect -17600 41017 -17520 41303
rect -17600 40983 -17577 41017
rect -17543 40983 -17520 41017
rect -17600 40960 -17520 40983
rect -17440 41337 -17360 41360
rect -17440 41303 -17417 41337
rect -17383 41303 -17360 41337
rect -17440 41017 -17360 41303
rect -17440 40983 -17417 41017
rect -17383 40983 -17360 41017
rect -17440 40960 -17360 40983
rect -17280 41337 -17200 41360
rect -17280 41303 -17257 41337
rect -17223 41303 -17200 41337
rect -17280 41017 -17200 41303
rect -17280 40983 -17257 41017
rect -17223 40983 -17200 41017
rect -17280 40960 -17200 40983
rect -17120 41337 -17040 41360
rect -17120 41303 -17097 41337
rect -17063 41303 -17040 41337
rect -17120 41017 -17040 41303
rect -17120 40983 -17097 41017
rect -17063 40983 -17040 41017
rect -17120 40960 -17040 40983
rect -16960 41337 -16880 41360
rect -16960 41303 -16937 41337
rect -16903 41303 -16880 41337
rect -16960 41017 -16880 41303
rect -16960 40983 -16937 41017
rect -16903 40983 -16880 41017
rect -16960 40960 -16880 40983
rect -16800 41337 -16720 41360
rect -16800 41303 -16777 41337
rect -16743 41303 -16720 41337
rect -16800 41017 -16720 41303
rect -16800 40983 -16777 41017
rect -16743 40983 -16720 41017
rect -16800 40960 -16720 40983
rect -16640 41337 -16560 41360
rect -16640 41303 -16617 41337
rect -16583 41303 -16560 41337
rect -16640 41017 -16560 41303
rect -16640 40983 -16617 41017
rect -16583 40983 -16560 41017
rect -16640 40960 -16560 40983
rect -16480 41337 -16400 41360
rect -16480 41303 -16457 41337
rect -16423 41303 -16400 41337
rect -16480 41017 -16400 41303
rect -16480 40983 -16457 41017
rect -16423 40983 -16400 41017
rect -16480 40960 -16400 40983
rect -16320 41337 -16240 41360
rect -16320 41303 -16297 41337
rect -16263 41303 -16240 41337
rect -16320 41017 -16240 41303
rect -16320 40983 -16297 41017
rect -16263 40983 -16240 41017
rect -16320 40960 -16240 40983
rect -16160 41337 -16080 41360
rect -16160 41303 -16137 41337
rect -16103 41303 -16080 41337
rect -16160 41017 -16080 41303
rect -16160 40983 -16137 41017
rect -16103 40983 -16080 41017
rect -16160 40960 -16080 40983
rect -16000 41337 -15920 41360
rect -16000 41303 -15977 41337
rect -15943 41303 -15920 41337
rect -16000 41017 -15920 41303
rect -16000 40983 -15977 41017
rect -15943 40983 -15920 41017
rect -16000 40960 -15920 40983
rect -15840 41337 -15760 41360
rect -15840 41303 -15817 41337
rect -15783 41303 -15760 41337
rect -15840 41017 -15760 41303
rect -15840 40983 -15817 41017
rect -15783 40983 -15760 41017
rect -15840 40960 -15760 40983
rect -15680 41337 -15600 41360
rect -15680 41303 -15657 41337
rect -15623 41303 -15600 41337
rect -15680 41017 -15600 41303
rect -15680 40983 -15657 41017
rect -15623 40983 -15600 41017
rect -15680 40960 -15600 40983
rect -15520 41337 -15440 41360
rect -15520 41303 -15497 41337
rect -15463 41303 -15440 41337
rect -15520 41017 -15440 41303
rect -15520 40983 -15497 41017
rect -15463 40983 -15440 41017
rect -15520 40960 -15440 40983
rect -15360 41337 -15280 41360
rect -15360 41303 -15337 41337
rect -15303 41303 -15280 41337
rect -15360 41017 -15280 41303
rect -15360 40983 -15337 41017
rect -15303 40983 -15280 41017
rect -15360 40960 -15280 40983
rect -15200 41337 -15120 41360
rect -15200 41303 -15177 41337
rect -15143 41303 -15120 41337
rect -15200 41017 -15120 41303
rect -15200 40983 -15177 41017
rect -15143 40983 -15120 41017
rect -15200 40960 -15120 40983
rect -15040 41337 -14960 41360
rect -15040 41303 -15017 41337
rect -14983 41303 -14960 41337
rect -15040 41017 -14960 41303
rect -15040 40983 -15017 41017
rect -14983 40983 -14960 41017
rect -15040 40960 -14960 40983
rect -14880 41337 -14800 41360
rect -14880 41303 -14857 41337
rect -14823 41303 -14800 41337
rect -14880 41017 -14800 41303
rect -14880 40983 -14857 41017
rect -14823 40983 -14800 41017
rect -14880 40960 -14800 40983
rect -14720 41337 -14640 41360
rect -14720 41303 -14697 41337
rect -14663 41303 -14640 41337
rect -14720 41017 -14640 41303
rect -14720 40983 -14697 41017
rect -14663 40983 -14640 41017
rect -14720 40960 -14640 40983
rect -14560 41337 -14480 41360
rect -14560 41303 -14537 41337
rect -14503 41303 -14480 41337
rect -14560 41017 -14480 41303
rect -14560 40983 -14537 41017
rect -14503 40983 -14480 41017
rect -14560 40960 -14480 40983
rect -14400 41337 -14320 41360
rect -14400 41303 -14377 41337
rect -14343 41303 -14320 41337
rect -14400 41017 -14320 41303
rect -14400 40983 -14377 41017
rect -14343 40983 -14320 41017
rect -14400 40960 -14320 40983
rect -14240 41337 -14160 41360
rect -14240 41303 -14217 41337
rect -14183 41303 -14160 41337
rect -14240 41017 -14160 41303
rect -14240 40983 -14217 41017
rect -14183 40983 -14160 41017
rect -14240 40960 -14160 40983
rect -14080 41337 -14000 41360
rect -14080 41303 -14057 41337
rect -14023 41303 -14000 41337
rect -14080 41017 -14000 41303
rect -14080 40983 -14057 41017
rect -14023 40983 -14000 41017
rect -14080 40960 -14000 40983
rect -13920 41337 -13840 41360
rect -13920 41303 -13897 41337
rect -13863 41303 -13840 41337
rect -13920 41017 -13840 41303
rect -13920 40983 -13897 41017
rect -13863 40983 -13840 41017
rect -13920 40960 -13840 40983
rect -13760 41337 -13680 41360
rect -13760 41303 -13737 41337
rect -13703 41303 -13680 41337
rect -13760 41017 -13680 41303
rect -13760 40983 -13737 41017
rect -13703 40983 -13680 41017
rect -13760 40960 -13680 40983
rect -13600 41337 -13520 41360
rect -13600 41303 -13577 41337
rect -13543 41303 -13520 41337
rect -13600 41017 -13520 41303
rect -13600 40983 -13577 41017
rect -13543 40983 -13520 41017
rect -13600 40960 -13520 40983
rect -13440 41337 -13360 41360
rect -13440 41303 -13417 41337
rect -13383 41303 -13360 41337
rect -13440 41017 -13360 41303
rect -13440 40983 -13417 41017
rect -13383 40983 -13360 41017
rect -13440 40960 -13360 40983
rect -13280 41337 -13200 41360
rect -13280 41303 -13257 41337
rect -13223 41303 -13200 41337
rect -13280 41017 -13200 41303
rect -13280 40983 -13257 41017
rect -13223 40983 -13200 41017
rect -13280 40960 -13200 40983
rect -13120 41337 -13040 41360
rect -13120 41303 -13097 41337
rect -13063 41303 -13040 41337
rect -13120 41017 -13040 41303
rect -13120 40983 -13097 41017
rect -13063 40983 -13040 41017
rect -13120 40960 -13040 40983
rect -12960 41337 -12880 41360
rect -12960 41303 -12937 41337
rect -12903 41303 -12880 41337
rect -12960 41017 -12880 41303
rect -12960 40983 -12937 41017
rect -12903 40983 -12880 41017
rect -12960 40960 -12880 40983
rect -12800 41337 -12720 41360
rect -12800 41303 -12777 41337
rect -12743 41303 -12720 41337
rect -12800 41017 -12720 41303
rect -12800 40983 -12777 41017
rect -12743 40983 -12720 41017
rect -12800 40960 -12720 40983
rect -12640 41337 -12560 41360
rect -12640 41303 -12617 41337
rect -12583 41303 -12560 41337
rect -12640 41017 -12560 41303
rect -12640 40983 -12617 41017
rect -12583 40983 -12560 41017
rect -12640 40960 -12560 40983
rect -12480 41337 -12400 41360
rect -12480 41303 -12457 41337
rect -12423 41303 -12400 41337
rect -12480 41017 -12400 41303
rect -12480 40983 -12457 41017
rect -12423 40983 -12400 41017
rect -12480 40960 -12400 40983
rect -12320 41337 -12240 41360
rect -12320 41303 -12297 41337
rect -12263 41303 -12240 41337
rect -12320 41017 -12240 41303
rect -12320 40983 -12297 41017
rect -12263 40983 -12240 41017
rect -12320 40960 -12240 40983
rect -11360 41337 -11280 41360
rect -11360 41303 -11337 41337
rect -11303 41303 -11280 41337
rect -11360 41017 -11280 41303
rect -11360 40983 -11337 41017
rect -11303 40983 -11280 41017
rect -11360 40960 -11280 40983
rect -11200 41337 -11120 41360
rect -11200 41303 -11177 41337
rect -11143 41303 -11120 41337
rect -11200 41017 -11120 41303
rect -11200 40983 -11177 41017
rect -11143 40983 -11120 41017
rect -11200 40960 -11120 40983
rect -11040 41337 -10960 41360
rect -11040 41303 -11017 41337
rect -10983 41303 -10960 41337
rect -11040 41017 -10960 41303
rect -11040 40983 -11017 41017
rect -10983 40983 -10960 41017
rect -11040 40960 -10960 40983
rect -10880 41337 -10800 41360
rect -10880 41303 -10857 41337
rect -10823 41303 -10800 41337
rect -10880 41017 -10800 41303
rect -10880 40983 -10857 41017
rect -10823 40983 -10800 41017
rect -10880 40960 -10800 40983
rect -10720 41337 -10640 41360
rect -10720 41303 -10697 41337
rect -10663 41303 -10640 41337
rect -10720 41017 -10640 41303
rect -10720 40983 -10697 41017
rect -10663 40983 -10640 41017
rect -10720 40960 -10640 40983
rect -10560 41337 -10480 41360
rect -10560 41303 -10537 41337
rect -10503 41303 -10480 41337
rect -10560 41017 -10480 41303
rect -10560 40983 -10537 41017
rect -10503 40983 -10480 41017
rect -10560 40960 -10480 40983
rect -10400 41337 -10320 41360
rect -10400 41303 -10377 41337
rect -10343 41303 -10320 41337
rect -10400 41017 -10320 41303
rect -10400 40983 -10377 41017
rect -10343 40983 -10320 41017
rect -10400 40960 -10320 40983
rect -10240 41337 -10160 41360
rect -10240 41303 -10217 41337
rect -10183 41303 -10160 41337
rect -10240 41017 -10160 41303
rect -10240 40983 -10217 41017
rect -10183 40983 -10160 41017
rect -10240 40960 -10160 40983
rect -10080 41337 -10000 41360
rect -10080 41303 -10057 41337
rect -10023 41303 -10000 41337
rect -10080 41017 -10000 41303
rect -10080 40983 -10057 41017
rect -10023 40983 -10000 41017
rect -10080 40960 -10000 40983
rect -9920 41337 -9840 41360
rect -9920 41303 -9897 41337
rect -9863 41303 -9840 41337
rect -9920 41017 -9840 41303
rect -9920 40983 -9897 41017
rect -9863 40983 -9840 41017
rect -9920 40960 -9840 40983
rect -9760 41337 -9680 41360
rect -9760 41303 -9737 41337
rect -9703 41303 -9680 41337
rect -9760 41017 -9680 41303
rect -9760 40983 -9737 41017
rect -9703 40983 -9680 41017
rect -9760 40960 -9680 40983
rect -9600 41337 -9520 41360
rect -9600 41303 -9577 41337
rect -9543 41303 -9520 41337
rect -9600 41017 -9520 41303
rect -9600 40983 -9577 41017
rect -9543 40983 -9520 41017
rect -9600 40960 -9520 40983
rect -9440 41337 -9360 41360
rect -9440 41303 -9417 41337
rect -9383 41303 -9360 41337
rect -9440 41017 -9360 41303
rect -9440 40983 -9417 41017
rect -9383 40983 -9360 41017
rect -9440 40960 -9360 40983
rect -9280 41337 -9200 41360
rect -9280 41303 -9257 41337
rect -9223 41303 -9200 41337
rect -9280 41017 -9200 41303
rect -9280 40983 -9257 41017
rect -9223 40983 -9200 41017
rect -9280 40960 -9200 40983
rect -9120 41337 -9040 41360
rect -9120 41303 -9097 41337
rect -9063 41303 -9040 41337
rect -9120 41017 -9040 41303
rect -9120 40983 -9097 41017
rect -9063 40983 -9040 41017
rect -9120 40960 -9040 40983
rect -8960 41337 -8880 41360
rect -8960 41303 -8937 41337
rect -8903 41303 -8880 41337
rect -8960 41017 -8880 41303
rect -8960 40983 -8937 41017
rect -8903 40983 -8880 41017
rect -8960 40960 -8880 40983
rect -8800 41337 -8720 41360
rect -8800 41303 -8777 41337
rect -8743 41303 -8720 41337
rect -8800 41017 -8720 41303
rect -8800 40983 -8777 41017
rect -8743 40983 -8720 41017
rect -8800 40960 -8720 40983
rect -8640 41337 -8560 41360
rect -8640 41303 -8617 41337
rect -8583 41303 -8560 41337
rect -8640 41017 -8560 41303
rect -8640 40983 -8617 41017
rect -8583 40983 -8560 41017
rect -8640 40960 -8560 40983
rect -8480 41337 -8400 41360
rect -8480 41303 -8457 41337
rect -8423 41303 -8400 41337
rect -8480 41017 -8400 41303
rect -8480 40983 -8457 41017
rect -8423 40983 -8400 41017
rect -8480 40960 -8400 40983
rect -8320 41337 -8240 41360
rect -8320 41303 -8297 41337
rect -8263 41303 -8240 41337
rect -8320 41017 -8240 41303
rect -8320 40983 -8297 41017
rect -8263 40983 -8240 41017
rect -8320 40960 -8240 40983
rect -8160 41337 -8080 41360
rect -8160 41303 -8137 41337
rect -8103 41303 -8080 41337
rect -8160 41017 -8080 41303
rect -8160 40983 -8137 41017
rect -8103 40983 -8080 41017
rect -8160 40960 -8080 40983
rect -8000 41337 -7920 41360
rect -8000 41303 -7977 41337
rect -7943 41303 -7920 41337
rect -8000 41017 -7920 41303
rect -8000 40983 -7977 41017
rect -7943 40983 -7920 41017
rect -8000 40960 -7920 40983
rect -7840 41337 -7760 41360
rect -7840 41303 -7817 41337
rect -7783 41303 -7760 41337
rect -7840 41017 -7760 41303
rect -7840 40983 -7817 41017
rect -7783 40983 -7760 41017
rect -7840 40960 -7760 40983
rect -7680 41337 -7600 41360
rect -7680 41303 -7657 41337
rect -7623 41303 -7600 41337
rect -7680 41017 -7600 41303
rect -7680 40983 -7657 41017
rect -7623 40983 -7600 41017
rect -7680 40960 -7600 40983
rect -7520 41337 -7440 41360
rect -7520 41303 -7497 41337
rect -7463 41303 -7440 41337
rect -7520 41017 -7440 41303
rect -7520 40983 -7497 41017
rect -7463 40983 -7440 41017
rect -7520 40960 -7440 40983
rect -7360 41337 -7280 41360
rect -7360 41303 -7337 41337
rect -7303 41303 -7280 41337
rect -7360 41017 -7280 41303
rect -7360 40983 -7337 41017
rect -7303 40983 -7280 41017
rect -7360 40960 -7280 40983
rect -7200 41337 -7120 41360
rect -7200 41303 -7177 41337
rect -7143 41303 -7120 41337
rect -7200 41017 -7120 41303
rect -7200 40983 -7177 41017
rect -7143 40983 -7120 41017
rect -7200 40960 -7120 40983
rect -7040 41337 -6960 41360
rect -7040 41303 -7017 41337
rect -6983 41303 -6960 41337
rect -7040 41017 -6960 41303
rect -7040 40983 -7017 41017
rect -6983 40983 -6960 41017
rect -7040 40960 -6960 40983
rect -6880 41337 -6800 41360
rect -6880 41303 -6857 41337
rect -6823 41303 -6800 41337
rect -6880 41017 -6800 41303
rect -6880 40983 -6857 41017
rect -6823 40983 -6800 41017
rect -6880 40960 -6800 40983
rect -6720 41337 -6640 41360
rect -6720 41303 -6697 41337
rect -6663 41303 -6640 41337
rect -6720 41017 -6640 41303
rect -6720 40983 -6697 41017
rect -6663 40983 -6640 41017
rect -6720 40960 -6640 40983
rect -6560 41337 -6480 41360
rect -6560 41303 -6537 41337
rect -6503 41303 -6480 41337
rect -6560 41017 -6480 41303
rect -6560 40983 -6537 41017
rect -6503 40983 -6480 41017
rect -6560 40960 -6480 40983
rect -6400 41337 -6320 41360
rect -6400 41303 -6377 41337
rect -6343 41303 -6320 41337
rect -6400 41017 -6320 41303
rect -6400 40983 -6377 41017
rect -6343 40983 -6320 41017
rect -6400 40960 -6320 40983
rect -6240 41337 -6160 41360
rect -6240 41303 -6217 41337
rect -6183 41303 -6160 41337
rect -6240 41017 -6160 41303
rect -6240 40983 -6217 41017
rect -6183 40983 -6160 41017
rect -6240 40960 -6160 40983
rect -6080 41337 -6000 41360
rect -6080 41303 -6057 41337
rect -6023 41303 -6000 41337
rect -6080 41017 -6000 41303
rect -6080 40983 -6057 41017
rect -6023 40983 -6000 41017
rect -6080 40960 -6000 40983
rect -5920 41337 -5840 41360
rect -5920 41303 -5897 41337
rect -5863 41303 -5840 41337
rect -5920 41017 -5840 41303
rect -5920 40983 -5897 41017
rect -5863 40983 -5840 41017
rect -5920 40960 -5840 40983
rect -5760 41337 -5680 41360
rect -5760 41303 -5737 41337
rect -5703 41303 -5680 41337
rect -5760 41017 -5680 41303
rect -5760 40983 -5737 41017
rect -5703 40983 -5680 41017
rect -5760 40960 -5680 40983
rect -5600 41337 -5520 41360
rect -5600 41303 -5577 41337
rect -5543 41303 -5520 41337
rect -5600 41017 -5520 41303
rect -5600 40983 -5577 41017
rect -5543 40983 -5520 41017
rect -5600 40960 -5520 40983
rect -5440 41337 -5360 41360
rect -5440 41303 -5417 41337
rect -5383 41303 -5360 41337
rect -5440 41017 -5360 41303
rect -5440 40983 -5417 41017
rect -5383 40983 -5360 41017
rect -5440 40960 -5360 40983
rect -5280 41337 -5200 41360
rect -5280 41303 -5257 41337
rect -5223 41303 -5200 41337
rect -5280 41017 -5200 41303
rect -5280 40983 -5257 41017
rect -5223 40983 -5200 41017
rect -5280 40960 -5200 40983
rect -5120 41337 -5040 41360
rect -5120 41303 -5097 41337
rect -5063 41303 -5040 41337
rect -5120 41017 -5040 41303
rect -5120 40983 -5097 41017
rect -5063 40983 -5040 41017
rect -5120 40960 -5040 40983
rect -4960 41337 -4880 41360
rect -4960 41303 -4937 41337
rect -4903 41303 -4880 41337
rect -4960 41017 -4880 41303
rect -4960 40983 -4937 41017
rect -4903 40983 -4880 41017
rect -4960 40960 -4880 40983
rect -4800 41337 -4720 41360
rect -4800 41303 -4777 41337
rect -4743 41303 -4720 41337
rect -4800 41017 -4720 41303
rect -4800 40983 -4777 41017
rect -4743 40983 -4720 41017
rect -4800 40960 -4720 40983
rect -4640 41337 -4560 41360
rect -4640 41303 -4617 41337
rect -4583 41303 -4560 41337
rect -4640 41017 -4560 41303
rect -4640 40983 -4617 41017
rect -4583 40983 -4560 41017
rect -4640 40960 -4560 40983
rect -4480 41337 -4400 41360
rect -4480 41303 -4457 41337
rect -4423 41303 -4400 41337
rect -4480 41017 -4400 41303
rect -4480 40983 -4457 41017
rect -4423 40983 -4400 41017
rect -4480 40960 -4400 40983
rect -4320 41337 -4240 41360
rect -4320 41303 -4297 41337
rect -4263 41303 -4240 41337
rect -4320 41017 -4240 41303
rect -4320 40983 -4297 41017
rect -4263 40983 -4240 41017
rect -4320 40960 -4240 40983
rect -4160 41337 -4080 41360
rect -4160 41303 -4137 41337
rect -4103 41303 -4080 41337
rect -4160 41017 -4080 41303
rect -4160 40983 -4137 41017
rect -4103 40983 -4080 41017
rect -4160 40960 -4080 40983
rect -4000 41337 -3920 41360
rect -4000 41303 -3977 41337
rect -3943 41303 -3920 41337
rect -4000 41017 -3920 41303
rect -4000 40983 -3977 41017
rect -3943 40983 -3920 41017
rect -4000 40960 -3920 40983
rect -3840 41337 -3760 42960
rect -3680 42857 -3600 42880
rect -3680 42823 -3657 42857
rect -3623 42823 -3600 42857
rect -3680 42537 -3600 42823
rect -3680 42503 -3657 42537
rect -3623 42503 -3600 42537
rect -3680 42217 -3600 42503
rect -3680 42183 -3657 42217
rect -3623 42183 -3600 42217
rect -3680 41897 -3600 42183
rect -3680 41863 -3657 41897
rect -3623 41863 -3600 41897
rect -3680 41840 -3600 41863
rect -3520 42857 -3440 42880
rect -3520 42823 -3497 42857
rect -3463 42823 -3440 42857
rect -3520 42537 -3440 42823
rect -3520 42503 -3497 42537
rect -3463 42503 -3440 42537
rect -3520 42217 -3440 42503
rect -3520 42183 -3497 42217
rect -3463 42183 -3440 42217
rect -3520 41897 -3440 42183
rect -3520 41863 -3497 41897
rect -3463 41863 -3440 41897
rect -3520 41840 -3440 41863
rect -3360 42857 -3280 42880
rect -3360 42823 -3337 42857
rect -3303 42823 -3280 42857
rect -3360 42537 -3280 42823
rect -3360 42503 -3337 42537
rect -3303 42503 -3280 42537
rect -3360 42217 -3280 42503
rect -3360 42183 -3337 42217
rect -3303 42183 -3280 42217
rect -3360 41897 -3280 42183
rect -3360 41863 -3337 41897
rect -3303 41863 -3280 41897
rect -3360 41840 -3280 41863
rect -3040 42857 -2960 42880
rect -3040 42823 -3017 42857
rect -2983 42823 -2960 42857
rect -3040 42537 -2960 42823
rect -3040 42503 -3017 42537
rect -2983 42503 -2960 42537
rect -3040 42217 -2960 42503
rect -3040 42183 -3017 42217
rect -2983 42183 -2960 42217
rect -3040 41897 -2960 42183
rect -3040 41863 -3017 41897
rect -2983 41863 -2960 41897
rect -3040 41840 -2960 41863
rect -2720 42857 -2640 42880
rect -2720 42823 -2697 42857
rect -2663 42823 -2640 42857
rect -2720 42537 -2640 42823
rect -2720 42503 -2697 42537
rect -2663 42503 -2640 42537
rect -2720 42217 -2640 42503
rect -2720 42183 -2697 42217
rect -2663 42183 -2640 42217
rect -2720 41897 -2640 42183
rect -2720 41863 -2697 41897
rect -2663 41863 -2640 41897
rect -2720 41840 -2640 41863
rect -2560 42857 -2480 42880
rect -2560 42823 -2537 42857
rect -2503 42823 -2480 42857
rect -2560 42537 -2480 42823
rect -2560 42503 -2537 42537
rect -2503 42503 -2480 42537
rect -2560 42217 -2480 42503
rect -2560 42183 -2537 42217
rect -2503 42183 -2480 42217
rect -2560 41897 -2480 42183
rect -2560 41863 -2537 41897
rect -2503 41863 -2480 41897
rect -2560 41840 -2480 41863
rect -2400 42857 -2320 42880
rect -2400 42823 -2377 42857
rect -2343 42823 -2320 42857
rect -2400 42537 -2320 42823
rect -2400 42503 -2377 42537
rect -2343 42503 -2320 42537
rect -2400 42217 -2320 42503
rect -2400 42183 -2377 42217
rect -2343 42183 -2320 42217
rect -2400 41897 -2320 42183
rect -2400 41863 -2377 41897
rect -2343 41863 -2320 41897
rect -2400 41840 -2320 41863
rect -2240 42857 -2160 42880
rect -2240 42823 -2217 42857
rect -2183 42823 -2160 42857
rect -2240 42537 -2160 42823
rect -2240 42503 -2217 42537
rect -2183 42503 -2160 42537
rect -2240 42217 -2160 42503
rect -2240 42183 -2217 42217
rect -2183 42183 -2160 42217
rect -2240 41897 -2160 42183
rect -2240 41863 -2217 41897
rect -2183 41863 -2160 41897
rect -2240 41840 -2160 41863
rect -2080 42857 -2000 42880
rect -2080 42823 -2057 42857
rect -2023 42823 -2000 42857
rect -2080 42537 -2000 42823
rect -2080 42503 -2057 42537
rect -2023 42503 -2000 42537
rect -2080 42217 -2000 42503
rect -2080 42183 -2057 42217
rect -2023 42183 -2000 42217
rect -2080 41897 -2000 42183
rect -2080 41863 -2057 41897
rect -2023 41863 -2000 41897
rect -2080 41840 -2000 41863
rect -1760 42857 -1680 42880
rect -1760 42823 -1737 42857
rect -1703 42823 -1680 42857
rect -1760 42537 -1680 42823
rect -1760 42503 -1737 42537
rect -1703 42503 -1680 42537
rect -1760 42217 -1680 42503
rect -1760 42183 -1737 42217
rect -1703 42183 -1680 42217
rect -1760 41897 -1680 42183
rect -1760 41863 -1737 41897
rect -1703 41863 -1680 41897
rect -1760 41840 -1680 41863
rect -1440 42857 -1360 42880
rect -1440 42823 -1417 42857
rect -1383 42823 -1360 42857
rect -1440 42537 -1360 42823
rect -1440 42503 -1417 42537
rect -1383 42503 -1360 42537
rect -1440 42217 -1360 42503
rect -1440 42183 -1417 42217
rect -1383 42183 -1360 42217
rect -1440 41897 -1360 42183
rect -1440 41863 -1417 41897
rect -1383 41863 -1360 41897
rect -1440 41840 -1360 41863
rect -1120 42857 -1040 42880
rect -1120 42823 -1097 42857
rect -1063 42823 -1040 42857
rect -1120 42537 -1040 42823
rect -1120 42503 -1097 42537
rect -1063 42503 -1040 42537
rect -1120 42217 -1040 42503
rect -1120 42183 -1097 42217
rect -1063 42183 -1040 42217
rect -1120 41897 -1040 42183
rect -1120 41863 -1097 41897
rect -1063 41863 -1040 41897
rect -1120 41840 -1040 41863
rect -3840 41303 -3817 41337
rect -3783 41303 -3760 41337
rect -3840 41017 -3760 41303
rect -3840 40983 -3817 41017
rect -3783 40983 -3760 41017
rect -10560 40697 -10480 40720
rect -10560 40663 -10537 40697
rect -10503 40663 -10480 40697
rect -10560 40377 -10480 40663
rect -10560 40343 -10537 40377
rect -10503 40343 -10480 40377
rect -10560 40320 -10480 40343
rect -10240 40697 -10160 40720
rect -10240 40663 -10217 40697
rect -10183 40663 -10160 40697
rect -10240 40377 -10160 40663
rect -10240 40343 -10217 40377
rect -10183 40343 -10160 40377
rect -10240 40320 -10160 40343
rect -10080 40697 -10000 40720
rect -10080 40663 -10057 40697
rect -10023 40663 -10000 40697
rect -10080 40377 -10000 40663
rect -10080 40343 -10057 40377
rect -10023 40343 -10000 40377
rect -10080 40320 -10000 40343
rect -9920 40697 -9840 40720
rect -9920 40663 -9897 40697
rect -9863 40663 -9840 40697
rect -9920 40377 -9840 40663
rect -9920 40343 -9897 40377
rect -9863 40343 -9840 40377
rect -9920 40320 -9840 40343
rect -9760 40697 -9680 40720
rect -9760 40663 -9737 40697
rect -9703 40663 -9680 40697
rect -9760 40377 -9680 40663
rect -9760 40343 -9737 40377
rect -9703 40343 -9680 40377
rect -9760 40320 -9680 40343
rect -9600 40697 -9520 40720
rect -9600 40663 -9577 40697
rect -9543 40663 -9520 40697
rect -9600 40377 -9520 40663
rect -9600 40343 -9577 40377
rect -9543 40343 -9520 40377
rect -9600 40320 -9520 40343
rect -9440 40697 -9360 40720
rect -9440 40663 -9417 40697
rect -9383 40663 -9360 40697
rect -9440 40377 -9360 40663
rect -9440 40343 -9417 40377
rect -9383 40343 -9360 40377
rect -9440 40320 -9360 40343
rect -9280 40697 -9200 40720
rect -9280 40663 -9257 40697
rect -9223 40663 -9200 40697
rect -9280 40377 -9200 40663
rect -9280 40343 -9257 40377
rect -9223 40343 -9200 40377
rect -9280 40320 -9200 40343
rect -9120 40697 -9040 40720
rect -9120 40663 -9097 40697
rect -9063 40663 -9040 40697
rect -9120 40377 -9040 40663
rect -9120 40343 -9097 40377
rect -9063 40343 -9040 40377
rect -9120 40320 -9040 40343
rect -8960 40697 -8880 40720
rect -8960 40663 -8937 40697
rect -8903 40663 -8880 40697
rect -8960 40377 -8880 40663
rect -8960 40343 -8937 40377
rect -8903 40343 -8880 40377
rect -8960 40320 -8880 40343
rect -8800 40697 -8720 40720
rect -8800 40663 -8777 40697
rect -8743 40663 -8720 40697
rect -8800 40377 -8720 40663
rect -8800 40343 -8777 40377
rect -8743 40343 -8720 40377
rect -8800 40320 -8720 40343
rect -8640 40697 -8560 40720
rect -8640 40663 -8617 40697
rect -8583 40663 -8560 40697
rect -8640 40377 -8560 40663
rect -8640 40343 -8617 40377
rect -8583 40343 -8560 40377
rect -8640 40320 -8560 40343
rect -8480 40697 -8400 40720
rect -8480 40663 -8457 40697
rect -8423 40663 -8400 40697
rect -8480 40377 -8400 40663
rect -8480 40343 -8457 40377
rect -8423 40343 -8400 40377
rect -8480 40320 -8400 40343
rect -8320 40697 -8240 40720
rect -8320 40663 -8297 40697
rect -8263 40663 -8240 40697
rect -8320 40377 -8240 40663
rect -8320 40343 -8297 40377
rect -8263 40343 -8240 40377
rect -8320 40320 -8240 40343
rect -8160 40697 -8080 40720
rect -8160 40663 -8137 40697
rect -8103 40663 -8080 40697
rect -8160 40377 -8080 40663
rect -8160 40343 -8137 40377
rect -8103 40343 -8080 40377
rect -8160 40320 -8080 40343
rect -8000 40697 -7920 40720
rect -8000 40663 -7977 40697
rect -7943 40663 -7920 40697
rect -8000 40377 -7920 40663
rect -8000 40343 -7977 40377
rect -7943 40343 -7920 40377
rect -8000 40320 -7920 40343
rect -7840 40697 -7760 40720
rect -7840 40663 -7817 40697
rect -7783 40663 -7760 40697
rect -7840 40377 -7760 40663
rect -7840 40343 -7817 40377
rect -7783 40343 -7760 40377
rect -7840 40320 -7760 40343
rect -7680 40697 -7600 40720
rect -7680 40663 -7657 40697
rect -7623 40663 -7600 40697
rect -7680 40377 -7600 40663
rect -7680 40343 -7657 40377
rect -7623 40343 -7600 40377
rect -7680 40320 -7600 40343
rect -7520 40697 -7440 40720
rect -7520 40663 -7497 40697
rect -7463 40663 -7440 40697
rect -7520 40377 -7440 40663
rect -7520 40343 -7497 40377
rect -7463 40343 -7440 40377
rect -7520 40320 -7440 40343
rect -7360 40697 -7280 40720
rect -7360 40663 -7337 40697
rect -7303 40663 -7280 40697
rect -7360 40377 -7280 40663
rect -7360 40343 -7337 40377
rect -7303 40343 -7280 40377
rect -7360 40320 -7280 40343
rect -7200 40697 -7120 40720
rect -7200 40663 -7177 40697
rect -7143 40663 -7120 40697
rect -7200 40377 -7120 40663
rect -7200 40343 -7177 40377
rect -7143 40343 -7120 40377
rect -7200 40320 -7120 40343
rect -7040 40697 -6960 40720
rect -7040 40663 -7017 40697
rect -6983 40663 -6960 40697
rect -7040 40377 -6960 40663
rect -7040 40343 -7017 40377
rect -6983 40343 -6960 40377
rect -7040 40320 -6960 40343
rect -6880 40697 -6800 40720
rect -6880 40663 -6857 40697
rect -6823 40663 -6800 40697
rect -6880 40377 -6800 40663
rect -6880 40343 -6857 40377
rect -6823 40343 -6800 40377
rect -6880 40320 -6800 40343
rect -6720 40697 -6640 40720
rect -6720 40663 -6697 40697
rect -6663 40663 -6640 40697
rect -6720 40377 -6640 40663
rect -6720 40343 -6697 40377
rect -6663 40343 -6640 40377
rect -6720 40320 -6640 40343
rect -6560 40697 -6480 40720
rect -6560 40663 -6537 40697
rect -6503 40663 -6480 40697
rect -6560 40377 -6480 40663
rect -6560 40343 -6537 40377
rect -6503 40343 -6480 40377
rect -6560 40320 -6480 40343
rect -6400 40697 -6320 40720
rect -6400 40663 -6377 40697
rect -6343 40663 -6320 40697
rect -6400 40377 -6320 40663
rect -6400 40343 -6377 40377
rect -6343 40343 -6320 40377
rect -6400 40320 -6320 40343
rect -6240 40697 -6160 40720
rect -6240 40663 -6217 40697
rect -6183 40663 -6160 40697
rect -6240 40377 -6160 40663
rect -6240 40343 -6217 40377
rect -6183 40343 -6160 40377
rect -6240 40320 -6160 40343
rect -6080 40697 -6000 40720
rect -6080 40663 -6057 40697
rect -6023 40663 -6000 40697
rect -6080 40377 -6000 40663
rect -6080 40343 -6057 40377
rect -6023 40343 -6000 40377
rect -6080 40320 -6000 40343
rect -5920 40697 -5840 40720
rect -5920 40663 -5897 40697
rect -5863 40663 -5840 40697
rect -5920 40377 -5840 40663
rect -5920 40343 -5897 40377
rect -5863 40343 -5840 40377
rect -5920 40320 -5840 40343
rect -5760 40697 -5680 40720
rect -5760 40663 -5737 40697
rect -5703 40663 -5680 40697
rect -5760 40377 -5680 40663
rect -5760 40343 -5737 40377
rect -5703 40343 -5680 40377
rect -5760 40320 -5680 40343
rect -5600 40697 -5520 40720
rect -5600 40663 -5577 40697
rect -5543 40663 -5520 40697
rect -5600 40377 -5520 40663
rect -5600 40343 -5577 40377
rect -5543 40343 -5520 40377
rect -5600 40320 -5520 40343
rect -5440 40697 -5360 40720
rect -5440 40663 -5417 40697
rect -5383 40663 -5360 40697
rect -5440 40377 -5360 40663
rect -5440 40343 -5417 40377
rect -5383 40343 -5360 40377
rect -5440 40320 -5360 40343
rect -5280 40697 -5200 40720
rect -5280 40663 -5257 40697
rect -5223 40663 -5200 40697
rect -5280 40377 -5200 40663
rect -5280 40343 -5257 40377
rect -5223 40343 -5200 40377
rect -5280 40320 -5200 40343
rect -5120 40697 -5040 40720
rect -5120 40663 -5097 40697
rect -5063 40663 -5040 40697
rect -5120 40377 -5040 40663
rect -5120 40343 -5097 40377
rect -5063 40343 -5040 40377
rect -5120 40320 -5040 40343
rect -4960 40697 -4880 40720
rect -4960 40663 -4937 40697
rect -4903 40663 -4880 40697
rect -4960 40377 -4880 40663
rect -4960 40343 -4937 40377
rect -4903 40343 -4880 40377
rect -4960 40320 -4880 40343
rect -4800 40697 -4720 40720
rect -4800 40663 -4777 40697
rect -4743 40663 -4720 40697
rect -4800 40377 -4720 40663
rect -4800 40343 -4777 40377
rect -4743 40343 -4720 40377
rect -4800 40320 -4720 40343
rect -4640 40697 -4560 40720
rect -4640 40663 -4617 40697
rect -4583 40663 -4560 40697
rect -4640 40377 -4560 40663
rect -4640 40343 -4617 40377
rect -4583 40343 -4560 40377
rect -4640 40320 -4560 40343
rect -4480 40697 -4400 40720
rect -4480 40663 -4457 40697
rect -4423 40663 -4400 40697
rect -4480 40377 -4400 40663
rect -4480 40343 -4457 40377
rect -4423 40343 -4400 40377
rect -4480 40320 -4400 40343
rect -4320 40697 -4240 40720
rect -4320 40663 -4297 40697
rect -4263 40663 -4240 40697
rect -4320 40377 -4240 40663
rect -4320 40343 -4297 40377
rect -4263 40343 -4240 40377
rect -4320 40320 -4240 40343
rect -4160 40697 -4080 40720
rect -4160 40663 -4137 40697
rect -4103 40663 -4080 40697
rect -4160 40377 -4080 40663
rect -4160 40343 -4137 40377
rect -4103 40343 -4080 40377
rect -4160 40320 -4080 40343
rect -4000 40697 -3920 40720
rect -4000 40663 -3977 40697
rect -3943 40663 -3920 40697
rect -4000 40377 -3920 40663
rect -4000 40343 -3977 40377
rect -3943 40343 -3920 40377
rect -4000 40320 -3920 40343
rect -3840 39920 -3760 40983
rect -3680 41337 -3600 41360
rect -3680 41303 -3657 41337
rect -3623 41303 -3600 41337
rect -3680 41017 -3600 41303
rect -3680 40983 -3657 41017
rect -3623 40983 -3600 41017
rect -3680 40960 -3600 40983
rect -3520 41337 -3440 41360
rect -3520 41303 -3497 41337
rect -3463 41303 -3440 41337
rect -3520 41017 -3440 41303
rect -3520 40983 -3497 41017
rect -3463 40983 -3440 41017
rect -3520 40960 -3440 40983
rect 41040 41337 41120 41360
rect 41040 41303 41063 41337
rect 41097 41303 41120 41337
rect 41040 41017 41120 41303
rect 41040 40983 41063 41017
rect 41097 40983 41120 41017
rect 41040 40960 41120 40983
rect 41200 41337 41280 41360
rect 41200 41303 41223 41337
rect 41257 41303 41280 41337
rect 41200 41017 41280 41303
rect 41200 40983 41223 41017
rect 41257 40983 41280 41017
rect 41200 40960 41280 40983
rect 41360 41337 41440 41360
rect 41360 41303 41383 41337
rect 41417 41303 41440 41337
rect 41360 41017 41440 41303
rect 41360 40983 41383 41017
rect 41417 40983 41440 41017
rect 41360 40960 41440 40983
rect 41520 41337 41600 41360
rect 41520 41303 41543 41337
rect 41577 41303 41600 41337
rect 41520 41017 41600 41303
rect 41520 40983 41543 41017
rect 41577 40983 41600 41017
rect 41520 40960 41600 40983
rect 41680 41337 41760 41360
rect 41680 41303 41703 41337
rect 41737 41303 41760 41337
rect 41680 41017 41760 41303
rect 41680 40983 41703 41017
rect 41737 40983 41760 41017
rect 41680 40960 41760 40983
rect 41840 41337 41920 41360
rect 41840 41303 41863 41337
rect 41897 41303 41920 41337
rect 41840 41017 41920 41303
rect 41840 40983 41863 41017
rect 41897 40983 41920 41017
rect 41840 40960 41920 40983
rect 42000 41337 42080 41360
rect 42000 41303 42023 41337
rect 42057 41303 42080 41337
rect 42000 41017 42080 41303
rect 42000 40983 42023 41017
rect 42057 40983 42080 41017
rect 42000 40960 42080 40983
rect 42160 41337 42240 41360
rect 42160 41303 42183 41337
rect 42217 41303 42240 41337
rect 42160 41017 42240 41303
rect 42160 40983 42183 41017
rect 42217 40983 42240 41017
rect 42160 40960 42240 40983
rect 42320 41337 42400 41360
rect 42320 41303 42343 41337
rect 42377 41303 42400 41337
rect 42320 41017 42400 41303
rect 42320 40983 42343 41017
rect 42377 40983 42400 41017
rect 42320 40960 42400 40983
rect 42480 41337 42560 41360
rect 42480 41303 42503 41337
rect 42537 41303 42560 41337
rect 42480 41017 42560 41303
rect 42480 40983 42503 41017
rect 42537 40983 42560 41017
rect 42480 40960 42560 40983
rect 42640 41337 42720 41360
rect 42640 41303 42663 41337
rect 42697 41303 42720 41337
rect 42640 41017 42720 41303
rect 42640 40983 42663 41017
rect 42697 40983 42720 41017
rect 42640 40960 42720 40983
rect 42800 41337 42880 41360
rect 42800 41303 42823 41337
rect 42857 41303 42880 41337
rect 42800 41017 42880 41303
rect 42800 40983 42823 41017
rect 42857 40983 42880 41017
rect 42800 40960 42880 40983
rect 42960 41337 43040 41360
rect 42960 41303 42983 41337
rect 43017 41303 43040 41337
rect 42960 41017 43040 41303
rect 42960 40983 42983 41017
rect 43017 40983 43040 41017
rect 42960 40960 43040 40983
rect 43120 41337 43200 41360
rect 43120 41303 43143 41337
rect 43177 41303 43200 41337
rect 43120 41017 43200 41303
rect 43120 40983 43143 41017
rect 43177 40983 43200 41017
rect 43120 40960 43200 40983
rect -3680 40697 -3600 40720
rect -3680 40663 -3657 40697
rect -3623 40663 -3600 40697
rect -3680 40377 -3600 40663
rect -3680 40343 -3657 40377
rect -3623 40343 -3600 40377
rect -3680 40320 -3600 40343
rect -3520 40697 -3440 40720
rect -3520 40663 -3497 40697
rect -3463 40663 -3440 40697
rect -3520 40377 -3440 40663
rect -3520 40343 -3497 40377
rect -3463 40343 -3440 40377
rect -3520 40320 -3440 40343
rect 41040 40057 41120 40080
rect 41040 40023 41063 40057
rect 41097 40023 41120 40057
rect 41040 39737 41120 40023
rect 41040 39703 41063 39737
rect 41097 39703 41120 39737
rect 41040 39680 41120 39703
rect 41200 40057 41280 40080
rect 41200 40023 41223 40057
rect 41257 40023 41280 40057
rect 41200 39737 41280 40023
rect 41200 39703 41223 39737
rect 41257 39703 41280 39737
rect 41200 39680 41280 39703
rect 41360 40057 41440 40080
rect 41360 40023 41383 40057
rect 41417 40023 41440 40057
rect 41360 39737 41440 40023
rect 41360 39703 41383 39737
rect 41417 39703 41440 39737
rect 41360 39680 41440 39703
rect 41520 40057 41600 40080
rect 41520 40023 41543 40057
rect 41577 40023 41600 40057
rect 41520 39737 41600 40023
rect 41520 39703 41543 39737
rect 41577 39703 41600 39737
rect 41520 39680 41600 39703
rect 41680 40057 41760 40080
rect 41680 40023 41703 40057
rect 41737 40023 41760 40057
rect 41680 39737 41760 40023
rect 41680 39703 41703 39737
rect 41737 39703 41760 39737
rect 41680 39680 41760 39703
rect 41840 40057 41920 40080
rect 41840 40023 41863 40057
rect 41897 40023 41920 40057
rect 41840 39737 41920 40023
rect 41840 39703 41863 39737
rect 41897 39703 41920 39737
rect 41840 39680 41920 39703
rect 42000 40057 42080 40080
rect 42000 40023 42023 40057
rect 42057 40023 42080 40057
rect 42000 39737 42080 40023
rect 42000 39703 42023 39737
rect 42057 39703 42080 39737
rect 42000 39680 42080 39703
rect 42160 40057 42240 40080
rect 42160 40023 42183 40057
rect 42217 40023 42240 40057
rect 42160 39737 42240 40023
rect 42160 39703 42183 39737
rect 42217 39703 42240 39737
rect 42160 39680 42240 39703
rect 42320 40057 42400 40080
rect 42320 40023 42343 40057
rect 42377 40023 42400 40057
rect 42320 39737 42400 40023
rect 42320 39703 42343 39737
rect 42377 39703 42400 39737
rect 42320 39680 42400 39703
rect 42480 40057 42560 40080
rect 42480 40023 42503 40057
rect 42537 40023 42560 40057
rect 42480 39737 42560 40023
rect 42480 39703 42503 39737
rect 42537 39703 42560 39737
rect 42480 39680 42560 39703
rect 42640 40057 42720 40080
rect 42640 40023 42663 40057
rect 42697 40023 42720 40057
rect 42640 39737 42720 40023
rect 42640 39703 42663 39737
rect 42697 39703 42720 39737
rect 42640 39680 42720 39703
rect 42800 40057 42880 40080
rect 42800 40023 42823 40057
rect 42857 40023 42880 40057
rect 42800 39737 42880 40023
rect 42800 39703 42823 39737
rect 42857 39703 42880 39737
rect 42800 39680 42880 39703
rect 42960 40057 43040 40080
rect 42960 40023 42983 40057
rect 43017 40023 43040 40057
rect 42960 39737 43040 40023
rect 42960 39703 42983 39737
rect 43017 39703 43040 39737
rect 42960 39680 43040 39703
rect 43120 40057 43200 40080
rect 43120 40023 43143 40057
rect 43177 40023 43200 40057
rect 43120 39737 43200 40023
rect 43120 39703 43143 39737
rect 43177 39703 43200 39737
rect 43120 39680 43200 39703
rect -33120 37737 -33040 37760
rect -33120 37703 -33097 37737
rect -33063 37703 -33040 37737
rect -33120 37417 -33040 37703
rect -33120 37383 -33097 37417
rect -33063 37383 -33040 37417
rect -33120 37097 -33040 37383
rect -33120 37063 -33097 37097
rect -33063 37063 -33040 37097
rect -33120 37040 -33040 37063
rect -32960 37737 -32880 37760
rect -32960 37703 -32937 37737
rect -32903 37703 -32880 37737
rect -32960 37417 -32880 37703
rect -32960 37383 -32937 37417
rect -32903 37383 -32880 37417
rect -32960 37097 -32880 37383
rect -32960 37063 -32937 37097
rect -32903 37063 -32880 37097
rect -32960 37040 -32880 37063
rect -32800 37737 -32720 37760
rect -32800 37703 -32777 37737
rect -32743 37703 -32720 37737
rect -32800 37417 -32720 37703
rect -32800 37383 -32777 37417
rect -32743 37383 -32720 37417
rect -32800 37097 -32720 37383
rect -32800 37063 -32777 37097
rect -32743 37063 -32720 37097
rect -32800 37040 -32720 37063
rect -32640 37737 -32560 37760
rect -32640 37703 -32617 37737
rect -32583 37703 -32560 37737
rect -32640 37417 -32560 37703
rect -32640 37383 -32617 37417
rect -32583 37383 -32560 37417
rect -32640 37097 -32560 37383
rect -32640 37063 -32617 37097
rect -32583 37063 -32560 37097
rect -32640 37040 -32560 37063
rect -32480 37737 -32400 37760
rect -32480 37703 -32457 37737
rect -32423 37703 -32400 37737
rect -32480 37417 -32400 37703
rect -32480 37383 -32457 37417
rect -32423 37383 -32400 37417
rect -32480 37097 -32400 37383
rect -32480 37063 -32457 37097
rect -32423 37063 -32400 37097
rect -32480 37040 -32400 37063
rect -32320 37737 -32240 37760
rect -32320 37703 -32297 37737
rect -32263 37703 -32240 37737
rect -32320 37417 -32240 37703
rect -32320 37383 -32297 37417
rect -32263 37383 -32240 37417
rect -32320 37097 -32240 37383
rect -32320 37063 -32297 37097
rect -32263 37063 -32240 37097
rect -32320 37040 -32240 37063
rect -32160 37737 -32080 37760
rect -32160 37703 -32137 37737
rect -32103 37703 -32080 37737
rect -32160 37417 -32080 37703
rect -32160 37383 -32137 37417
rect -32103 37383 -32080 37417
rect -32160 37097 -32080 37383
rect -32160 37063 -32137 37097
rect -32103 37063 -32080 37097
rect -32160 37040 -32080 37063
rect -32000 37737 -31920 37760
rect -32000 37703 -31977 37737
rect -31943 37703 -31920 37737
rect -32000 37417 -31920 37703
rect -32000 37383 -31977 37417
rect -31943 37383 -31920 37417
rect -32000 37097 -31920 37383
rect -32000 37063 -31977 37097
rect -31943 37063 -31920 37097
rect -32000 37040 -31920 37063
rect -31840 37737 -31760 37760
rect -31840 37703 -31817 37737
rect -31783 37703 -31760 37737
rect -31840 37417 -31760 37703
rect -31840 37383 -31817 37417
rect -31783 37383 -31760 37417
rect -31840 37097 -31760 37383
rect -31840 37063 -31817 37097
rect -31783 37063 -31760 37097
rect -31840 37040 -31760 37063
rect -31680 37737 -31600 37760
rect -31680 37703 -31657 37737
rect -31623 37703 -31600 37737
rect -31680 37417 -31600 37703
rect -31680 37383 -31657 37417
rect -31623 37383 -31600 37417
rect -31680 37097 -31600 37383
rect -31680 37063 -31657 37097
rect -31623 37063 -31600 37097
rect -31680 37040 -31600 37063
rect -31520 37737 -31440 37760
rect -31520 37703 -31497 37737
rect -31463 37703 -31440 37737
rect -31520 37417 -31440 37703
rect -31520 37383 -31497 37417
rect -31463 37383 -31440 37417
rect -31520 37097 -31440 37383
rect -31520 37063 -31497 37097
rect -31463 37063 -31440 37097
rect -31520 37040 -31440 37063
rect -31360 37737 -31280 37760
rect -31360 37703 -31337 37737
rect -31303 37703 -31280 37737
rect -31360 37417 -31280 37703
rect -31360 37383 -31337 37417
rect -31303 37383 -31280 37417
rect -31360 37097 -31280 37383
rect -31360 37063 -31337 37097
rect -31303 37063 -31280 37097
rect -31360 37040 -31280 37063
rect -31200 37737 -31120 37760
rect -31200 37703 -31177 37737
rect -31143 37703 -31120 37737
rect -31200 37417 -31120 37703
rect -31200 37383 -31177 37417
rect -31143 37383 -31120 37417
rect -31200 37097 -31120 37383
rect -31200 37063 -31177 37097
rect -31143 37063 -31120 37097
rect -31200 37040 -31120 37063
rect 41040 36057 41120 36080
rect 41040 36023 41063 36057
rect 41097 36023 41120 36057
rect 41040 35737 41120 36023
rect 41040 35703 41063 35737
rect 41097 35703 41120 35737
rect 41040 35680 41120 35703
rect 41200 36057 41280 36080
rect 41200 36023 41223 36057
rect 41257 36023 41280 36057
rect 41200 35737 41280 36023
rect 41200 35703 41223 35737
rect 41257 35703 41280 35737
rect 41200 35680 41280 35703
rect 41360 36057 41440 36080
rect 41360 36023 41383 36057
rect 41417 36023 41440 36057
rect 41360 35737 41440 36023
rect 41360 35703 41383 35737
rect 41417 35703 41440 35737
rect 41360 35680 41440 35703
rect 41520 36057 41600 36080
rect 41520 36023 41543 36057
rect 41577 36023 41600 36057
rect 41520 35737 41600 36023
rect 41520 35703 41543 35737
rect 41577 35703 41600 35737
rect 41520 35680 41600 35703
rect 41680 36057 41760 36080
rect 41680 36023 41703 36057
rect 41737 36023 41760 36057
rect 41680 35737 41760 36023
rect 41680 35703 41703 35737
rect 41737 35703 41760 35737
rect 41680 35680 41760 35703
rect 41840 36057 41920 36080
rect 41840 36023 41863 36057
rect 41897 36023 41920 36057
rect 41840 35737 41920 36023
rect 41840 35703 41863 35737
rect 41897 35703 41920 35737
rect 41840 35680 41920 35703
rect 42000 36057 42080 36080
rect 42000 36023 42023 36057
rect 42057 36023 42080 36057
rect 42000 35737 42080 36023
rect 42000 35703 42023 35737
rect 42057 35703 42080 35737
rect 42000 35680 42080 35703
rect 42160 36057 42240 36080
rect 42160 36023 42183 36057
rect 42217 36023 42240 36057
rect 42160 35737 42240 36023
rect 42160 35703 42183 35737
rect 42217 35703 42240 35737
rect 42160 35680 42240 35703
rect 42320 36057 42400 36080
rect 42320 36023 42343 36057
rect 42377 36023 42400 36057
rect 42320 35737 42400 36023
rect 42320 35703 42343 35737
rect 42377 35703 42400 35737
rect 42320 35680 42400 35703
rect 42480 36057 42560 36080
rect 42480 36023 42503 36057
rect 42537 36023 42560 36057
rect 42480 35737 42560 36023
rect 42480 35703 42503 35737
rect 42537 35703 42560 35737
rect 42480 35680 42560 35703
rect 42640 36057 42720 36080
rect 42640 36023 42663 36057
rect 42697 36023 42720 36057
rect 42640 35737 42720 36023
rect 42640 35703 42663 35737
rect 42697 35703 42720 35737
rect 42640 35680 42720 35703
rect 42800 36057 42880 36080
rect 42800 36023 42823 36057
rect 42857 36023 42880 36057
rect 42800 35737 42880 36023
rect 42800 35703 42823 35737
rect 42857 35703 42880 35737
rect 42800 35680 42880 35703
rect 42960 36057 43040 36080
rect 42960 36023 42983 36057
rect 43017 36023 43040 36057
rect 42960 35737 43040 36023
rect 42960 35703 42983 35737
rect 43017 35703 43040 35737
rect 42960 35680 43040 35703
rect 43120 36057 43200 36080
rect 43120 36023 43143 36057
rect 43177 36023 43200 36057
rect 43120 35737 43200 36023
rect 43120 35703 43143 35737
rect 43177 35703 43200 35737
rect 43120 35680 43200 35703
rect -33120 34697 -33040 34720
rect -33120 34663 -33097 34697
rect -33063 34663 -33040 34697
rect -33120 34377 -33040 34663
rect -33120 34343 -33097 34377
rect -33063 34343 -33040 34377
rect -33120 34320 -33040 34343
rect -32960 34697 -32880 34720
rect -32960 34663 -32937 34697
rect -32903 34663 -32880 34697
rect -32960 34377 -32880 34663
rect -32960 34343 -32937 34377
rect -32903 34343 -32880 34377
rect -32960 34320 -32880 34343
rect -32800 34697 -32720 34720
rect -32800 34663 -32777 34697
rect -32743 34663 -32720 34697
rect -32800 34377 -32720 34663
rect -32800 34343 -32777 34377
rect -32743 34343 -32720 34377
rect -32800 34320 -32720 34343
rect -32640 34697 -32560 34720
rect -32640 34663 -32617 34697
rect -32583 34663 -32560 34697
rect -32640 34377 -32560 34663
rect -32640 34343 -32617 34377
rect -32583 34343 -32560 34377
rect -32640 34320 -32560 34343
rect -32480 34697 -32400 34720
rect -32480 34663 -32457 34697
rect -32423 34663 -32400 34697
rect -32480 34377 -32400 34663
rect -32480 34343 -32457 34377
rect -32423 34343 -32400 34377
rect -32480 34320 -32400 34343
rect -32320 34697 -32240 34720
rect -32320 34663 -32297 34697
rect -32263 34663 -32240 34697
rect -32320 34377 -32240 34663
rect -32320 34343 -32297 34377
rect -32263 34343 -32240 34377
rect -32320 34320 -32240 34343
rect -32160 34697 -32080 34720
rect -32160 34663 -32137 34697
rect -32103 34663 -32080 34697
rect -32160 34377 -32080 34663
rect -32160 34343 -32137 34377
rect -32103 34343 -32080 34377
rect -32160 34320 -32080 34343
rect -32000 34697 -31920 34720
rect -32000 34663 -31977 34697
rect -31943 34663 -31920 34697
rect -32000 34377 -31920 34663
rect -32000 34343 -31977 34377
rect -31943 34343 -31920 34377
rect -32000 34320 -31920 34343
rect -31840 34697 -31760 34720
rect -31840 34663 -31817 34697
rect -31783 34663 -31760 34697
rect -31840 34377 -31760 34663
rect -31840 34343 -31817 34377
rect -31783 34343 -31760 34377
rect -31840 34320 -31760 34343
rect -31680 34697 -31600 34720
rect -31680 34663 -31657 34697
rect -31623 34663 -31600 34697
rect -31680 34377 -31600 34663
rect -31680 34343 -31657 34377
rect -31623 34343 -31600 34377
rect -31680 34320 -31600 34343
rect -31520 34697 -31440 34720
rect -31520 34663 -31497 34697
rect -31463 34663 -31440 34697
rect -31520 34377 -31440 34663
rect -31520 34343 -31497 34377
rect -31463 34343 -31440 34377
rect -31520 34320 -31440 34343
rect -31360 34697 -31280 34720
rect -31360 34663 -31337 34697
rect -31303 34663 -31280 34697
rect -31360 34377 -31280 34663
rect -31360 34343 -31337 34377
rect -31303 34343 -31280 34377
rect -31360 34320 -31280 34343
rect -31200 34697 -31120 34720
rect -31200 34663 -31177 34697
rect -31143 34663 -31120 34697
rect -31200 34377 -31120 34663
rect -31200 34343 -31177 34377
rect -31143 34343 -31120 34377
rect -31200 34320 -31120 34343
rect -29920 34697 -29840 34720
rect -29920 34663 -29897 34697
rect -29863 34663 -29840 34697
rect -29920 34377 -29840 34663
rect -29920 34343 -29897 34377
rect -29863 34343 -29840 34377
rect -29920 34320 -29840 34343
rect -29760 34697 -29680 34720
rect -29760 34663 -29737 34697
rect -29703 34663 -29680 34697
rect -29760 34377 -29680 34663
rect -29760 34343 -29737 34377
rect -29703 34343 -29680 34377
rect -29760 34320 -29680 34343
rect -29600 34697 -29520 34720
rect -29600 34663 -29577 34697
rect -29543 34663 -29520 34697
rect -29600 34377 -29520 34663
rect -29600 34343 -29577 34377
rect -29543 34343 -29520 34377
rect -29600 34320 -29520 34343
rect -29440 34697 -29360 34720
rect -29440 34663 -29417 34697
rect -29383 34663 -29360 34697
rect -29440 34377 -29360 34663
rect -29440 34343 -29417 34377
rect -29383 34343 -29360 34377
rect -29440 34320 -29360 34343
rect -29280 34697 -29200 34720
rect -29280 34663 -29257 34697
rect -29223 34663 -29200 34697
rect -29280 34377 -29200 34663
rect -29280 34343 -29257 34377
rect -29223 34343 -29200 34377
rect -29280 34320 -29200 34343
rect -29120 34697 -29040 34720
rect -29120 34663 -29097 34697
rect -29063 34663 -29040 34697
rect -29120 34377 -29040 34663
rect -29120 34343 -29097 34377
rect -29063 34343 -29040 34377
rect -29120 34320 -29040 34343
rect -28960 34697 -28880 34720
rect -28960 34663 -28937 34697
rect -28903 34663 -28880 34697
rect -28960 34377 -28880 34663
rect -28960 34343 -28937 34377
rect -28903 34343 -28880 34377
rect -28960 34320 -28880 34343
rect -28800 34697 -28720 34720
rect -28800 34663 -28777 34697
rect -28743 34663 -28720 34697
rect -28800 34377 -28720 34663
rect -28800 34343 -28777 34377
rect -28743 34343 -28720 34377
rect -28800 34320 -28720 34343
rect -28640 34697 -28560 34720
rect -28640 34663 -28617 34697
rect -28583 34663 -28560 34697
rect -28640 34377 -28560 34663
rect -28640 34343 -28617 34377
rect -28583 34343 -28560 34377
rect -28640 34320 -28560 34343
rect -28480 34697 -28400 34720
rect -28480 34663 -28457 34697
rect -28423 34663 -28400 34697
rect -28480 34377 -28400 34663
rect -28480 34343 -28457 34377
rect -28423 34343 -28400 34377
rect -28480 34320 -28400 34343
rect -28320 34697 -28240 34720
rect -28320 34663 -28297 34697
rect -28263 34663 -28240 34697
rect -28320 34377 -28240 34663
rect -28320 34343 -28297 34377
rect -28263 34343 -28240 34377
rect -28320 34320 -28240 34343
rect -28160 34697 -28080 34720
rect -28160 34663 -28137 34697
rect -28103 34663 -28080 34697
rect -28160 34377 -28080 34663
rect -28160 34343 -28137 34377
rect -28103 34343 -28080 34377
rect -28160 34320 -28080 34343
rect -28000 34697 -27920 34720
rect -28000 34663 -27977 34697
rect -27943 34663 -27920 34697
rect -28000 34377 -27920 34663
rect -28000 34343 -27977 34377
rect -27943 34343 -27920 34377
rect -28000 34320 -27920 34343
rect -27840 34697 -27760 34720
rect -27840 34663 -27817 34697
rect -27783 34663 -27760 34697
rect -27840 34377 -27760 34663
rect -27840 34343 -27817 34377
rect -27783 34343 -27760 34377
rect -27840 34320 -27760 34343
rect -27680 34697 -27600 34720
rect -27680 34663 -27657 34697
rect -27623 34663 -27600 34697
rect -27680 34377 -27600 34663
rect -27680 34343 -27657 34377
rect -27623 34343 -27600 34377
rect -27680 34320 -27600 34343
rect -27520 34697 -27440 34720
rect -27520 34663 -27497 34697
rect -27463 34663 -27440 34697
rect -27520 34377 -27440 34663
rect -27520 34343 -27497 34377
rect -27463 34343 -27440 34377
rect -27520 34320 -27440 34343
rect -27360 34697 -27280 34720
rect -27360 34663 -27337 34697
rect -27303 34663 -27280 34697
rect -27360 34377 -27280 34663
rect -27360 34343 -27337 34377
rect -27303 34343 -27280 34377
rect -27360 34320 -27280 34343
rect -27200 34697 -27120 34720
rect -27200 34663 -27177 34697
rect -27143 34663 -27120 34697
rect -27200 34377 -27120 34663
rect -27200 34343 -27177 34377
rect -27143 34343 -27120 34377
rect -27200 34320 -27120 34343
rect -27040 34697 -26960 34720
rect -27040 34663 -27017 34697
rect -26983 34663 -26960 34697
rect -27040 34377 -26960 34663
rect -27040 34343 -27017 34377
rect -26983 34343 -26960 34377
rect -27040 34320 -26960 34343
rect -26880 34697 -26800 34720
rect -26880 34663 -26857 34697
rect -26823 34663 -26800 34697
rect -26880 34377 -26800 34663
rect -26880 34343 -26857 34377
rect -26823 34343 -26800 34377
rect -26880 34320 -26800 34343
rect -26720 34697 -26640 34720
rect -26720 34663 -26697 34697
rect -26663 34663 -26640 34697
rect -26720 34377 -26640 34663
rect -26720 34343 -26697 34377
rect -26663 34343 -26640 34377
rect -26720 34320 -26640 34343
rect -26560 34697 -26480 34720
rect -26560 34663 -26537 34697
rect -26503 34663 -26480 34697
rect -26560 34377 -26480 34663
rect -26560 34343 -26537 34377
rect -26503 34343 -26480 34377
rect -26560 34320 -26480 34343
rect -26400 34697 -26320 34720
rect -26400 34663 -26377 34697
rect -26343 34663 -26320 34697
rect -26400 34377 -26320 34663
rect -26400 34343 -26377 34377
rect -26343 34343 -26320 34377
rect -26400 34320 -26320 34343
rect -26240 34697 -26160 34720
rect -26240 34663 -26217 34697
rect -26183 34663 -26160 34697
rect -26240 34377 -26160 34663
rect -26240 34343 -26217 34377
rect -26183 34343 -26160 34377
rect -26240 34320 -26160 34343
rect -26080 34697 -26000 34720
rect -26080 34663 -26057 34697
rect -26023 34663 -26000 34697
rect -26080 34377 -26000 34663
rect -26080 34343 -26057 34377
rect -26023 34343 -26000 34377
rect -26080 34320 -26000 34343
rect -25920 34697 -25840 34720
rect -25920 34663 -25897 34697
rect -25863 34663 -25840 34697
rect -25920 34377 -25840 34663
rect -25920 34343 -25897 34377
rect -25863 34343 -25840 34377
rect -25920 34320 -25840 34343
rect -25760 34697 -25680 34720
rect -25760 34663 -25737 34697
rect -25703 34663 -25680 34697
rect -25760 34377 -25680 34663
rect -25760 34343 -25737 34377
rect -25703 34343 -25680 34377
rect -25760 34320 -25680 34343
rect -25600 34697 -25520 34720
rect -25600 34663 -25577 34697
rect -25543 34663 -25520 34697
rect -25600 34377 -25520 34663
rect -25600 34343 -25577 34377
rect -25543 34343 -25520 34377
rect -25600 34320 -25520 34343
rect -25440 34697 -25360 34720
rect -25440 34663 -25417 34697
rect -25383 34663 -25360 34697
rect -25440 34377 -25360 34663
rect -25440 34343 -25417 34377
rect -25383 34343 -25360 34377
rect -25440 34320 -25360 34343
rect -25280 34697 -25200 34720
rect -25280 34663 -25257 34697
rect -25223 34663 -25200 34697
rect -25280 34377 -25200 34663
rect -25280 34343 -25257 34377
rect -25223 34343 -25200 34377
rect -25280 34320 -25200 34343
rect -25120 34697 -25040 34720
rect -25120 34663 -25097 34697
rect -25063 34663 -25040 34697
rect -25120 34377 -25040 34663
rect -25120 34343 -25097 34377
rect -25063 34343 -25040 34377
rect -25120 34320 -25040 34343
rect -24960 34697 -24880 34720
rect -24960 34663 -24937 34697
rect -24903 34663 -24880 34697
rect -24960 34377 -24880 34663
rect -24960 34343 -24937 34377
rect -24903 34343 -24880 34377
rect -24960 34320 -24880 34343
rect -24800 34697 -24720 34720
rect -24800 34663 -24777 34697
rect -24743 34663 -24720 34697
rect -24800 34377 -24720 34663
rect -24800 34343 -24777 34377
rect -24743 34343 -24720 34377
rect -24800 34320 -24720 34343
rect -24640 34697 -24560 34720
rect -24640 34663 -24617 34697
rect -24583 34663 -24560 34697
rect -24640 34377 -24560 34663
rect -24640 34343 -24617 34377
rect -24583 34343 -24560 34377
rect -24640 34320 -24560 34343
rect -24480 34697 -24400 34720
rect -24480 34663 -24457 34697
rect -24423 34663 -24400 34697
rect -24480 34377 -24400 34663
rect -24480 34343 -24457 34377
rect -24423 34343 -24400 34377
rect -24480 34320 -24400 34343
rect -24320 34697 -24240 34720
rect -24320 34663 -24297 34697
rect -24263 34663 -24240 34697
rect -24320 34377 -24240 34663
rect -24320 34343 -24297 34377
rect -24263 34343 -24240 34377
rect -24320 34320 -24240 34343
rect -24160 34697 -24080 34720
rect -24160 34663 -24137 34697
rect -24103 34663 -24080 34697
rect -24160 34377 -24080 34663
rect -24160 34343 -24137 34377
rect -24103 34343 -24080 34377
rect -24160 34320 -24080 34343
rect -24000 34697 -23920 34720
rect -24000 34663 -23977 34697
rect -23943 34663 -23920 34697
rect -24000 34377 -23920 34663
rect -24000 34343 -23977 34377
rect -23943 34343 -23920 34377
rect -24000 34320 -23920 34343
rect -23840 34697 -23760 34720
rect -23840 34663 -23817 34697
rect -23783 34663 -23760 34697
rect -23840 34377 -23760 34663
rect -23840 34343 -23817 34377
rect -23783 34343 -23760 34377
rect -23840 34320 -23760 34343
rect -23680 34697 -23600 34720
rect -23680 34663 -23657 34697
rect -23623 34663 -23600 34697
rect -23680 34377 -23600 34663
rect -23680 34343 -23657 34377
rect -23623 34343 -23600 34377
rect -23680 34320 -23600 34343
rect -23520 34697 -23440 34720
rect -23520 34663 -23497 34697
rect -23463 34663 -23440 34697
rect -23520 34377 -23440 34663
rect -23520 34343 -23497 34377
rect -23463 34343 -23440 34377
rect -23520 34320 -23440 34343
rect -23360 34697 -23280 34720
rect -23360 34663 -23337 34697
rect -23303 34663 -23280 34697
rect -23360 34377 -23280 34663
rect -23360 34343 -23337 34377
rect -23303 34343 -23280 34377
rect -23360 34320 -23280 34343
rect -23200 34697 -23120 34720
rect -23200 34663 -23177 34697
rect -23143 34663 -23120 34697
rect -23200 34377 -23120 34663
rect -23200 34343 -23177 34377
rect -23143 34343 -23120 34377
rect -23200 34320 -23120 34343
rect -23040 34697 -22960 34720
rect -23040 34663 -23017 34697
rect -22983 34663 -22960 34697
rect -23040 34377 -22960 34663
rect -23040 34343 -23017 34377
rect -22983 34343 -22960 34377
rect -23040 34320 -22960 34343
rect -22880 34697 -22800 34720
rect -22880 34663 -22857 34697
rect -22823 34663 -22800 34697
rect -22880 34377 -22800 34663
rect -22880 34343 -22857 34377
rect -22823 34343 -22800 34377
rect -22880 34320 -22800 34343
rect -22720 34697 -22640 34720
rect -22720 34663 -22697 34697
rect -22663 34663 -22640 34697
rect -22720 34377 -22640 34663
rect -22720 34343 -22697 34377
rect -22663 34343 -22640 34377
rect -22720 34320 -22640 34343
rect -22560 34697 -22480 34720
rect -22560 34663 -22537 34697
rect -22503 34663 -22480 34697
rect -22560 34377 -22480 34663
rect -22560 34343 -22537 34377
rect -22503 34343 -22480 34377
rect -22560 34320 -22480 34343
rect -22400 34697 -22320 34720
rect -22400 34663 -22377 34697
rect -22343 34663 -22320 34697
rect -22400 34377 -22320 34663
rect -22400 34343 -22377 34377
rect -22343 34343 -22320 34377
rect -22400 34320 -22320 34343
rect -22240 34697 -22160 34720
rect -22240 34663 -22217 34697
rect -22183 34663 -22160 34697
rect -22240 34377 -22160 34663
rect -22240 34343 -22217 34377
rect -22183 34343 -22160 34377
rect -22240 34320 -22160 34343
rect -22080 34697 -22000 34720
rect -22080 34663 -22057 34697
rect -22023 34663 -22000 34697
rect -22080 34377 -22000 34663
rect -22080 34343 -22057 34377
rect -22023 34343 -22000 34377
rect -22080 34320 -22000 34343
rect -21920 34697 -21840 34720
rect -21920 34663 -21897 34697
rect -21863 34663 -21840 34697
rect -21920 34377 -21840 34663
rect -21920 34343 -21897 34377
rect -21863 34343 -21840 34377
rect -21920 34320 -21840 34343
rect -21760 34697 -21680 34720
rect -21760 34663 -21737 34697
rect -21703 34663 -21680 34697
rect -21760 34377 -21680 34663
rect -21760 34343 -21737 34377
rect -21703 34343 -21680 34377
rect -21760 34320 -21680 34343
rect -21600 34697 -21520 34720
rect -21600 34663 -21577 34697
rect -21543 34663 -21520 34697
rect -21600 34377 -21520 34663
rect -21600 34343 -21577 34377
rect -21543 34343 -21520 34377
rect -21600 34320 -21520 34343
rect -21440 34697 -21360 34720
rect -21440 34663 -21417 34697
rect -21383 34663 -21360 34697
rect -21440 34377 -21360 34663
rect -21440 34343 -21417 34377
rect -21383 34343 -21360 34377
rect -21440 34320 -21360 34343
rect -21280 34697 -21200 34720
rect -21280 34663 -21257 34697
rect -21223 34663 -21200 34697
rect -21280 34377 -21200 34663
rect -21280 34343 -21257 34377
rect -21223 34343 -21200 34377
rect -21280 34320 -21200 34343
rect -21120 34697 -21040 34720
rect -21120 34663 -21097 34697
rect -21063 34663 -21040 34697
rect -21120 34377 -21040 34663
rect -21120 34343 -21097 34377
rect -21063 34343 -21040 34377
rect -21120 34320 -21040 34343
rect -20960 34697 -20880 34720
rect -20960 34663 -20937 34697
rect -20903 34663 -20880 34697
rect -20960 34377 -20880 34663
rect -20960 34343 -20937 34377
rect -20903 34343 -20880 34377
rect -20960 34320 -20880 34343
rect -20800 34697 -20720 34720
rect -20800 34663 -20777 34697
rect -20743 34663 -20720 34697
rect -20800 34377 -20720 34663
rect -20800 34343 -20777 34377
rect -20743 34343 -20720 34377
rect -20800 34320 -20720 34343
rect -20640 34697 -20560 34720
rect -20640 34663 -20617 34697
rect -20583 34663 -20560 34697
rect -20640 34377 -20560 34663
rect -20640 34343 -20617 34377
rect -20583 34343 -20560 34377
rect -20640 34320 -20560 34343
rect -20480 34697 -20400 34720
rect -20480 34663 -20457 34697
rect -20423 34663 -20400 34697
rect -20480 34377 -20400 34663
rect -20480 34343 -20457 34377
rect -20423 34343 -20400 34377
rect -20480 34320 -20400 34343
rect -20320 34697 -20240 34720
rect -20320 34663 -20297 34697
rect -20263 34663 -20240 34697
rect -20320 34377 -20240 34663
rect -20320 34343 -20297 34377
rect -20263 34343 -20240 34377
rect -20320 34320 -20240 34343
rect -20160 34697 -20080 34720
rect -20160 34663 -20137 34697
rect -20103 34663 -20080 34697
rect -20160 34377 -20080 34663
rect -20160 34343 -20137 34377
rect -20103 34343 -20080 34377
rect -20160 34320 -20080 34343
rect -20000 34697 -19920 34720
rect -20000 34663 -19977 34697
rect -19943 34663 -19920 34697
rect -20000 34377 -19920 34663
rect -20000 34343 -19977 34377
rect -19943 34343 -19920 34377
rect -20000 34320 -19920 34343
rect -19840 34697 -19760 34720
rect -19840 34663 -19817 34697
rect -19783 34663 -19760 34697
rect -19840 34377 -19760 34663
rect -19840 34343 -19817 34377
rect -19783 34343 -19760 34377
rect -19840 34320 -19760 34343
rect -19680 34697 -19600 34720
rect -19680 34663 -19657 34697
rect -19623 34663 -19600 34697
rect -19680 34377 -19600 34663
rect -19680 34343 -19657 34377
rect -19623 34343 -19600 34377
rect -19680 34320 -19600 34343
rect -19520 34697 -19440 34720
rect -19520 34663 -19497 34697
rect -19463 34663 -19440 34697
rect -19520 34377 -19440 34663
rect -19520 34343 -19497 34377
rect -19463 34343 -19440 34377
rect -19520 34320 -19440 34343
rect -19360 34697 -19280 34720
rect -19360 34663 -19337 34697
rect -19303 34663 -19280 34697
rect -19360 34377 -19280 34663
rect -19360 34343 -19337 34377
rect -19303 34343 -19280 34377
rect -19360 34320 -19280 34343
rect -19200 34697 -19120 34720
rect -19200 34663 -19177 34697
rect -19143 34663 -19120 34697
rect -19200 34377 -19120 34663
rect -19200 34343 -19177 34377
rect -19143 34343 -19120 34377
rect -19200 34320 -19120 34343
rect -19040 34697 -18960 34720
rect -19040 34663 -19017 34697
rect -18983 34663 -18960 34697
rect -19040 34377 -18960 34663
rect -19040 34343 -19017 34377
rect -18983 34343 -18960 34377
rect -19040 34320 -18960 34343
rect -18880 34697 -18800 34720
rect -18880 34663 -18857 34697
rect -18823 34663 -18800 34697
rect -18880 34377 -18800 34663
rect -18880 34343 -18857 34377
rect -18823 34343 -18800 34377
rect -18880 34320 -18800 34343
rect -18720 34697 -18640 34720
rect -18720 34663 -18697 34697
rect -18663 34663 -18640 34697
rect -18720 34377 -18640 34663
rect -18720 34343 -18697 34377
rect -18663 34343 -18640 34377
rect -18720 34320 -18640 34343
rect -18560 34697 -18480 34720
rect -18560 34663 -18537 34697
rect -18503 34663 -18480 34697
rect -18560 34377 -18480 34663
rect -18560 34343 -18537 34377
rect -18503 34343 -18480 34377
rect -18560 34320 -18480 34343
rect -18400 34697 -18320 34720
rect -18400 34663 -18377 34697
rect -18343 34663 -18320 34697
rect -18400 34377 -18320 34663
rect -18400 34343 -18377 34377
rect -18343 34343 -18320 34377
rect -18400 34320 -18320 34343
rect -18240 34697 -18160 34720
rect -18240 34663 -18217 34697
rect -18183 34663 -18160 34697
rect -18240 34377 -18160 34663
rect -18240 34343 -18217 34377
rect -18183 34343 -18160 34377
rect -18240 34320 -18160 34343
rect -18080 34697 -18000 34720
rect -18080 34663 -18057 34697
rect -18023 34663 -18000 34697
rect -18080 34377 -18000 34663
rect -18080 34343 -18057 34377
rect -18023 34343 -18000 34377
rect -18080 34320 -18000 34343
rect -17920 34697 -17840 34720
rect -17920 34663 -17897 34697
rect -17863 34663 -17840 34697
rect -17920 34377 -17840 34663
rect -17920 34343 -17897 34377
rect -17863 34343 -17840 34377
rect -17920 34320 -17840 34343
rect -17760 34697 -17680 34720
rect -17760 34663 -17737 34697
rect -17703 34663 -17680 34697
rect -17760 34377 -17680 34663
rect -17760 34343 -17737 34377
rect -17703 34343 -17680 34377
rect -17760 34320 -17680 34343
rect -17600 34697 -17520 34720
rect -17600 34663 -17577 34697
rect -17543 34663 -17520 34697
rect -17600 34377 -17520 34663
rect -17600 34343 -17577 34377
rect -17543 34343 -17520 34377
rect -17600 34320 -17520 34343
rect -17440 34697 -17360 34720
rect -17440 34663 -17417 34697
rect -17383 34663 -17360 34697
rect -17440 34377 -17360 34663
rect -17440 34343 -17417 34377
rect -17383 34343 -17360 34377
rect -17440 34320 -17360 34343
rect -17280 34697 -17200 34720
rect -17280 34663 -17257 34697
rect -17223 34663 -17200 34697
rect -17280 34377 -17200 34663
rect -17280 34343 -17257 34377
rect -17223 34343 -17200 34377
rect -17280 34320 -17200 34343
rect -17120 34697 -17040 34720
rect -17120 34663 -17097 34697
rect -17063 34663 -17040 34697
rect -17120 34377 -17040 34663
rect -17120 34343 -17097 34377
rect -17063 34343 -17040 34377
rect -17120 34320 -17040 34343
rect -16960 34697 -16880 34720
rect -16960 34663 -16937 34697
rect -16903 34663 -16880 34697
rect -16960 34377 -16880 34663
rect -16960 34343 -16937 34377
rect -16903 34343 -16880 34377
rect -16960 34320 -16880 34343
rect -16800 34697 -16720 34720
rect -16800 34663 -16777 34697
rect -16743 34663 -16720 34697
rect -16800 34377 -16720 34663
rect -16800 34343 -16777 34377
rect -16743 34343 -16720 34377
rect -16800 34320 -16720 34343
rect -16640 34697 -16560 34720
rect -16640 34663 -16617 34697
rect -16583 34663 -16560 34697
rect -16640 34377 -16560 34663
rect -16640 34343 -16617 34377
rect -16583 34343 -16560 34377
rect -16640 34320 -16560 34343
rect -16480 34697 -16400 34720
rect -16480 34663 -16457 34697
rect -16423 34663 -16400 34697
rect -16480 34377 -16400 34663
rect -16480 34343 -16457 34377
rect -16423 34343 -16400 34377
rect -16480 34320 -16400 34343
rect -16320 34697 -16240 34720
rect -16320 34663 -16297 34697
rect -16263 34663 -16240 34697
rect -16320 34377 -16240 34663
rect -16320 34343 -16297 34377
rect -16263 34343 -16240 34377
rect -16320 34320 -16240 34343
rect -16160 34697 -16080 34720
rect -16160 34663 -16137 34697
rect -16103 34663 -16080 34697
rect -16160 34377 -16080 34663
rect -16160 34343 -16137 34377
rect -16103 34343 -16080 34377
rect -16160 34320 -16080 34343
rect -16000 34697 -15920 34720
rect -16000 34663 -15977 34697
rect -15943 34663 -15920 34697
rect -16000 34377 -15920 34663
rect -16000 34343 -15977 34377
rect -15943 34343 -15920 34377
rect -16000 34320 -15920 34343
rect -15840 34697 -15760 34720
rect -15840 34663 -15817 34697
rect -15783 34663 -15760 34697
rect -15840 34377 -15760 34663
rect -15840 34343 -15817 34377
rect -15783 34343 -15760 34377
rect -15840 34320 -15760 34343
rect -15680 34697 -15600 34720
rect -15680 34663 -15657 34697
rect -15623 34663 -15600 34697
rect -15680 34377 -15600 34663
rect -15680 34343 -15657 34377
rect -15623 34343 -15600 34377
rect -15680 34320 -15600 34343
rect -15520 34697 -15440 34720
rect -15520 34663 -15497 34697
rect -15463 34663 -15440 34697
rect -15520 34377 -15440 34663
rect -15520 34343 -15497 34377
rect -15463 34343 -15440 34377
rect -15520 34320 -15440 34343
rect -15360 34697 -15280 34720
rect -15360 34663 -15337 34697
rect -15303 34663 -15280 34697
rect -15360 34377 -15280 34663
rect -15360 34343 -15337 34377
rect -15303 34343 -15280 34377
rect -15360 34320 -15280 34343
rect -15200 34697 -15120 34720
rect -15200 34663 -15177 34697
rect -15143 34663 -15120 34697
rect -15200 34377 -15120 34663
rect -15200 34343 -15177 34377
rect -15143 34343 -15120 34377
rect -15200 34320 -15120 34343
rect -15040 34697 -14960 34720
rect -15040 34663 -15017 34697
rect -14983 34663 -14960 34697
rect -15040 34377 -14960 34663
rect -15040 34343 -15017 34377
rect -14983 34343 -14960 34377
rect -15040 34320 -14960 34343
rect -14880 34697 -14800 34720
rect -14880 34663 -14857 34697
rect -14823 34663 -14800 34697
rect -14880 34377 -14800 34663
rect -14880 34343 -14857 34377
rect -14823 34343 -14800 34377
rect -14880 34320 -14800 34343
rect -14720 34697 -14640 34720
rect -14720 34663 -14697 34697
rect -14663 34663 -14640 34697
rect -14720 34377 -14640 34663
rect -14720 34343 -14697 34377
rect -14663 34343 -14640 34377
rect -14720 34320 -14640 34343
rect -14560 34697 -14480 34720
rect -14560 34663 -14537 34697
rect -14503 34663 -14480 34697
rect -14560 34377 -14480 34663
rect -14560 34343 -14537 34377
rect -14503 34343 -14480 34377
rect -14560 34320 -14480 34343
rect -14400 34697 -14320 34720
rect -14400 34663 -14377 34697
rect -14343 34663 -14320 34697
rect -14400 34377 -14320 34663
rect -14400 34343 -14377 34377
rect -14343 34343 -14320 34377
rect -14400 34320 -14320 34343
rect -14240 34697 -14160 34720
rect -14240 34663 -14217 34697
rect -14183 34663 -14160 34697
rect -14240 34377 -14160 34663
rect -14240 34343 -14217 34377
rect -14183 34343 -14160 34377
rect -14240 34320 -14160 34343
rect -14080 34697 -14000 34720
rect -14080 34663 -14057 34697
rect -14023 34663 -14000 34697
rect -14080 34377 -14000 34663
rect -14080 34343 -14057 34377
rect -14023 34343 -14000 34377
rect -14080 34320 -14000 34343
rect -13920 34697 -13840 34720
rect -13920 34663 -13897 34697
rect -13863 34663 -13840 34697
rect -13920 34377 -13840 34663
rect -13920 34343 -13897 34377
rect -13863 34343 -13840 34377
rect -13920 34320 -13840 34343
rect -13760 34697 -13680 34720
rect -13760 34663 -13737 34697
rect -13703 34663 -13680 34697
rect -13760 34377 -13680 34663
rect -13760 34343 -13737 34377
rect -13703 34343 -13680 34377
rect -13760 34320 -13680 34343
rect -13600 34697 -13520 34720
rect -13600 34663 -13577 34697
rect -13543 34663 -13520 34697
rect -13600 34377 -13520 34663
rect -13600 34343 -13577 34377
rect -13543 34343 -13520 34377
rect -13600 34320 -13520 34343
rect -13440 34697 -13360 34720
rect -13440 34663 -13417 34697
rect -13383 34663 -13360 34697
rect -13440 34377 -13360 34663
rect -13440 34343 -13417 34377
rect -13383 34343 -13360 34377
rect -13440 34320 -13360 34343
rect -13280 34697 -13200 34720
rect -13280 34663 -13257 34697
rect -13223 34663 -13200 34697
rect -13280 34377 -13200 34663
rect -13280 34343 -13257 34377
rect -13223 34343 -13200 34377
rect -13280 34320 -13200 34343
rect -13120 34697 -13040 34720
rect -13120 34663 -13097 34697
rect -13063 34663 -13040 34697
rect -13120 34377 -13040 34663
rect -13120 34343 -13097 34377
rect -13063 34343 -13040 34377
rect -13120 34320 -13040 34343
rect -12960 34697 -12880 34720
rect -12960 34663 -12937 34697
rect -12903 34663 -12880 34697
rect -12960 34377 -12880 34663
rect -12960 34343 -12937 34377
rect -12903 34343 -12880 34377
rect -12960 34320 -12880 34343
rect -12800 34697 -12720 34720
rect -12800 34663 -12777 34697
rect -12743 34663 -12720 34697
rect -12800 34377 -12720 34663
rect -12800 34343 -12777 34377
rect -12743 34343 -12720 34377
rect -12800 34320 -12720 34343
rect -12640 34697 -12560 34720
rect -12640 34663 -12617 34697
rect -12583 34663 -12560 34697
rect -12640 34377 -12560 34663
rect -12640 34343 -12617 34377
rect -12583 34343 -12560 34377
rect -12640 34320 -12560 34343
rect -12480 34697 -12400 34720
rect -12480 34663 -12457 34697
rect -12423 34663 -12400 34697
rect -12480 34377 -12400 34663
rect -12480 34343 -12457 34377
rect -12423 34343 -12400 34377
rect -12480 34320 -12400 34343
rect -12320 34697 -12240 34720
rect -12320 34663 -12297 34697
rect -12263 34663 -12240 34697
rect -12320 34377 -12240 34663
rect -12320 34343 -12297 34377
rect -12263 34343 -12240 34377
rect -12320 34320 -12240 34343
rect -12160 34697 -12080 34720
rect -12160 34663 -12137 34697
rect -12103 34663 -12080 34697
rect -12160 34377 -12080 34663
rect -12160 34343 -12137 34377
rect -12103 34343 -12080 34377
rect -12160 34320 -12080 34343
rect -12000 34697 -11920 34720
rect -12000 34663 -11977 34697
rect -11943 34663 -11920 34697
rect -12000 34377 -11920 34663
rect -12000 34343 -11977 34377
rect -11943 34343 -11920 34377
rect -12000 34320 -11920 34343
rect -11840 34697 -11760 34720
rect -11840 34663 -11817 34697
rect -11783 34663 -11760 34697
rect -11840 34377 -11760 34663
rect -11840 34343 -11817 34377
rect -11783 34343 -11760 34377
rect -11840 34320 -11760 34343
rect -11680 34697 -11600 34720
rect -11680 34663 -11657 34697
rect -11623 34663 -11600 34697
rect -11680 34377 -11600 34663
rect -11680 34343 -11657 34377
rect -11623 34343 -11600 34377
rect -11680 34320 -11600 34343
rect -11520 34697 -11440 34720
rect -11520 34663 -11497 34697
rect -11463 34663 -11440 34697
rect -11520 34377 -11440 34663
rect -11520 34343 -11497 34377
rect -11463 34343 -11440 34377
rect -11520 34320 -11440 34343
rect -10880 34697 -10800 34720
rect -10880 34663 -10857 34697
rect -10823 34663 -10800 34697
rect -10880 34377 -10800 34663
rect -10880 34343 -10857 34377
rect -10823 34343 -10800 34377
rect -10880 34320 -10800 34343
rect -10560 34697 -10480 34720
rect -10560 34663 -10537 34697
rect -10503 34663 -10480 34697
rect -10560 34377 -10480 34663
rect -10560 34343 -10537 34377
rect -10503 34343 -10480 34377
rect -10560 34320 -10480 34343
rect -29920 32937 -29840 32960
rect -29920 32903 -29897 32937
rect -29863 32903 -29840 32937
rect -29920 32617 -29840 32903
rect -29920 32583 -29897 32617
rect -29863 32583 -29840 32617
rect -29920 32297 -29840 32583
rect -29920 32263 -29897 32297
rect -29863 32263 -29840 32297
rect -29920 31977 -29840 32263
rect -29920 31943 -29897 31977
rect -29863 31943 -29840 31977
rect -29920 31920 -29840 31943
rect -29760 32937 -29680 32960
rect -29760 32903 -29737 32937
rect -29703 32903 -29680 32937
rect -29760 32617 -29680 32903
rect -29760 32583 -29737 32617
rect -29703 32583 -29680 32617
rect -29760 32297 -29680 32583
rect -29760 32263 -29737 32297
rect -29703 32263 -29680 32297
rect -29760 31977 -29680 32263
rect -29760 31943 -29737 31977
rect -29703 31943 -29680 31977
rect -29760 31920 -29680 31943
rect -29600 32937 -29520 32960
rect -29600 32903 -29577 32937
rect -29543 32903 -29520 32937
rect -29600 32617 -29520 32903
rect -29600 32583 -29577 32617
rect -29543 32583 -29520 32617
rect -29600 32297 -29520 32583
rect -29600 32263 -29577 32297
rect -29543 32263 -29520 32297
rect -29600 31977 -29520 32263
rect -29600 31943 -29577 31977
rect -29543 31943 -29520 31977
rect -29600 31920 -29520 31943
rect -29440 32937 -29360 32960
rect -29440 32903 -29417 32937
rect -29383 32903 -29360 32937
rect -29440 32617 -29360 32903
rect -29440 32583 -29417 32617
rect -29383 32583 -29360 32617
rect -29440 32297 -29360 32583
rect -29440 32263 -29417 32297
rect -29383 32263 -29360 32297
rect -29440 31977 -29360 32263
rect -29440 31943 -29417 31977
rect -29383 31943 -29360 31977
rect -29440 31920 -29360 31943
rect -29280 32937 -29200 32960
rect -29280 32903 -29257 32937
rect -29223 32903 -29200 32937
rect -29280 32617 -29200 32903
rect -29280 32583 -29257 32617
rect -29223 32583 -29200 32617
rect -29280 32297 -29200 32583
rect -29280 32263 -29257 32297
rect -29223 32263 -29200 32297
rect -29280 31977 -29200 32263
rect -29280 31943 -29257 31977
rect -29223 31943 -29200 31977
rect -29280 31920 -29200 31943
rect -29120 32937 -29040 32960
rect -29120 32903 -29097 32937
rect -29063 32903 -29040 32937
rect -29120 32617 -29040 32903
rect -29120 32583 -29097 32617
rect -29063 32583 -29040 32617
rect -29120 32297 -29040 32583
rect -29120 32263 -29097 32297
rect -29063 32263 -29040 32297
rect -29120 31977 -29040 32263
rect -29120 31943 -29097 31977
rect -29063 31943 -29040 31977
rect -29120 31920 -29040 31943
rect -28960 32937 -28880 32960
rect -28960 32903 -28937 32937
rect -28903 32903 -28880 32937
rect -28960 32617 -28880 32903
rect -28960 32583 -28937 32617
rect -28903 32583 -28880 32617
rect -28960 32297 -28880 32583
rect -28960 32263 -28937 32297
rect -28903 32263 -28880 32297
rect -28960 31977 -28880 32263
rect -28960 31943 -28937 31977
rect -28903 31943 -28880 31977
rect -28960 31920 -28880 31943
rect -28800 32937 -28720 32960
rect -28800 32903 -28777 32937
rect -28743 32903 -28720 32937
rect -28800 32617 -28720 32903
rect -28800 32583 -28777 32617
rect -28743 32583 -28720 32617
rect -28800 32297 -28720 32583
rect -28800 32263 -28777 32297
rect -28743 32263 -28720 32297
rect -28800 31977 -28720 32263
rect -28800 31943 -28777 31977
rect -28743 31943 -28720 31977
rect -28800 31920 -28720 31943
rect -28640 32937 -28560 32960
rect -28640 32903 -28617 32937
rect -28583 32903 -28560 32937
rect -28640 32617 -28560 32903
rect -28640 32583 -28617 32617
rect -28583 32583 -28560 32617
rect -28640 32297 -28560 32583
rect -28640 32263 -28617 32297
rect -28583 32263 -28560 32297
rect -28640 31977 -28560 32263
rect -28640 31943 -28617 31977
rect -28583 31943 -28560 31977
rect -28640 31920 -28560 31943
rect -28480 32937 -28400 32960
rect -28480 32903 -28457 32937
rect -28423 32903 -28400 32937
rect -28480 32617 -28400 32903
rect -28480 32583 -28457 32617
rect -28423 32583 -28400 32617
rect -28480 32297 -28400 32583
rect -28480 32263 -28457 32297
rect -28423 32263 -28400 32297
rect -28480 31977 -28400 32263
rect -28480 31943 -28457 31977
rect -28423 31943 -28400 31977
rect -28480 31920 -28400 31943
rect -28320 32937 -28240 32960
rect -28320 32903 -28297 32937
rect -28263 32903 -28240 32937
rect -28320 32617 -28240 32903
rect -28320 32583 -28297 32617
rect -28263 32583 -28240 32617
rect -28320 32297 -28240 32583
rect -28320 32263 -28297 32297
rect -28263 32263 -28240 32297
rect -28320 31977 -28240 32263
rect -28320 31943 -28297 31977
rect -28263 31943 -28240 31977
rect -28320 31920 -28240 31943
rect -28160 32937 -28080 32960
rect -28160 32903 -28137 32937
rect -28103 32903 -28080 32937
rect -28160 32617 -28080 32903
rect -28160 32583 -28137 32617
rect -28103 32583 -28080 32617
rect -28160 32297 -28080 32583
rect -28160 32263 -28137 32297
rect -28103 32263 -28080 32297
rect -28160 31977 -28080 32263
rect -28160 31943 -28137 31977
rect -28103 31943 -28080 31977
rect -28160 31920 -28080 31943
rect -28000 32937 -27920 32960
rect -28000 32903 -27977 32937
rect -27943 32903 -27920 32937
rect -28000 32617 -27920 32903
rect -28000 32583 -27977 32617
rect -27943 32583 -27920 32617
rect -28000 32297 -27920 32583
rect -28000 32263 -27977 32297
rect -27943 32263 -27920 32297
rect -28000 31977 -27920 32263
rect -28000 31943 -27977 31977
rect -27943 31943 -27920 31977
rect -28000 31920 -27920 31943
rect -27840 32937 -27760 32960
rect -27840 32903 -27817 32937
rect -27783 32903 -27760 32937
rect -27840 32617 -27760 32903
rect -27840 32583 -27817 32617
rect -27783 32583 -27760 32617
rect -27840 32297 -27760 32583
rect -27840 32263 -27817 32297
rect -27783 32263 -27760 32297
rect -27840 31977 -27760 32263
rect -27840 31943 -27817 31977
rect -27783 31943 -27760 31977
rect -27840 31920 -27760 31943
rect -27680 32937 -27600 32960
rect -27680 32903 -27657 32937
rect -27623 32903 -27600 32937
rect -27680 32617 -27600 32903
rect -27680 32583 -27657 32617
rect -27623 32583 -27600 32617
rect -27680 32297 -27600 32583
rect -27680 32263 -27657 32297
rect -27623 32263 -27600 32297
rect -27680 31977 -27600 32263
rect -27680 31943 -27657 31977
rect -27623 31943 -27600 31977
rect -27680 31920 -27600 31943
rect -27520 32937 -27440 32960
rect -27520 32903 -27497 32937
rect -27463 32903 -27440 32937
rect -27520 32617 -27440 32903
rect -27520 32583 -27497 32617
rect -27463 32583 -27440 32617
rect -27520 32297 -27440 32583
rect -27520 32263 -27497 32297
rect -27463 32263 -27440 32297
rect -27520 31977 -27440 32263
rect -27520 31943 -27497 31977
rect -27463 31943 -27440 31977
rect -27520 31920 -27440 31943
rect -27360 32937 -27280 32960
rect -27360 32903 -27337 32937
rect -27303 32903 -27280 32937
rect -27360 32617 -27280 32903
rect -27360 32583 -27337 32617
rect -27303 32583 -27280 32617
rect -27360 32297 -27280 32583
rect -27360 32263 -27337 32297
rect -27303 32263 -27280 32297
rect -27360 31977 -27280 32263
rect -27360 31943 -27337 31977
rect -27303 31943 -27280 31977
rect -27360 31920 -27280 31943
rect -27200 32937 -27120 32960
rect -27200 32903 -27177 32937
rect -27143 32903 -27120 32937
rect -27200 32617 -27120 32903
rect -27200 32583 -27177 32617
rect -27143 32583 -27120 32617
rect -27200 32297 -27120 32583
rect -27200 32263 -27177 32297
rect -27143 32263 -27120 32297
rect -27200 31977 -27120 32263
rect -27200 31943 -27177 31977
rect -27143 31943 -27120 31977
rect -27200 31920 -27120 31943
rect -27040 32937 -26960 32960
rect -27040 32903 -27017 32937
rect -26983 32903 -26960 32937
rect -27040 32617 -26960 32903
rect -27040 32583 -27017 32617
rect -26983 32583 -26960 32617
rect -27040 32297 -26960 32583
rect -27040 32263 -27017 32297
rect -26983 32263 -26960 32297
rect -27040 31977 -26960 32263
rect -27040 31943 -27017 31977
rect -26983 31943 -26960 31977
rect -27040 31920 -26960 31943
rect -26880 32937 -26800 32960
rect -26880 32903 -26857 32937
rect -26823 32903 -26800 32937
rect -26880 32617 -26800 32903
rect -26880 32583 -26857 32617
rect -26823 32583 -26800 32617
rect -26880 32297 -26800 32583
rect -26880 32263 -26857 32297
rect -26823 32263 -26800 32297
rect -26880 31977 -26800 32263
rect -26880 31943 -26857 31977
rect -26823 31943 -26800 31977
rect -26880 31920 -26800 31943
rect -26720 32937 -26640 32960
rect -26720 32903 -26697 32937
rect -26663 32903 -26640 32937
rect -26720 32617 -26640 32903
rect -26720 32583 -26697 32617
rect -26663 32583 -26640 32617
rect -26720 32297 -26640 32583
rect -26720 32263 -26697 32297
rect -26663 32263 -26640 32297
rect -26720 31977 -26640 32263
rect -26720 31943 -26697 31977
rect -26663 31943 -26640 31977
rect -26720 31920 -26640 31943
rect -26560 32937 -26480 32960
rect -26560 32903 -26537 32937
rect -26503 32903 -26480 32937
rect -26560 32617 -26480 32903
rect -26560 32583 -26537 32617
rect -26503 32583 -26480 32617
rect -26560 32297 -26480 32583
rect -26560 32263 -26537 32297
rect -26503 32263 -26480 32297
rect -26560 31977 -26480 32263
rect -26560 31943 -26537 31977
rect -26503 31943 -26480 31977
rect -26560 31920 -26480 31943
rect -26400 32937 -26320 32960
rect -26400 32903 -26377 32937
rect -26343 32903 -26320 32937
rect -26400 32617 -26320 32903
rect -26400 32583 -26377 32617
rect -26343 32583 -26320 32617
rect -26400 32297 -26320 32583
rect -26400 32263 -26377 32297
rect -26343 32263 -26320 32297
rect -26400 31977 -26320 32263
rect -26400 31943 -26377 31977
rect -26343 31943 -26320 31977
rect -26400 31920 -26320 31943
rect -26240 32937 -26160 32960
rect -26240 32903 -26217 32937
rect -26183 32903 -26160 32937
rect -26240 32617 -26160 32903
rect -26240 32583 -26217 32617
rect -26183 32583 -26160 32617
rect -26240 32297 -26160 32583
rect -26240 32263 -26217 32297
rect -26183 32263 -26160 32297
rect -26240 31977 -26160 32263
rect -26240 31943 -26217 31977
rect -26183 31943 -26160 31977
rect -26240 31920 -26160 31943
rect -26080 32937 -26000 32960
rect -26080 32903 -26057 32937
rect -26023 32903 -26000 32937
rect -26080 32617 -26000 32903
rect -26080 32583 -26057 32617
rect -26023 32583 -26000 32617
rect -26080 32297 -26000 32583
rect -26080 32263 -26057 32297
rect -26023 32263 -26000 32297
rect -26080 31977 -26000 32263
rect -26080 31943 -26057 31977
rect -26023 31943 -26000 31977
rect -26080 31920 -26000 31943
rect -25920 32937 -25840 32960
rect -25920 32903 -25897 32937
rect -25863 32903 -25840 32937
rect -25920 32617 -25840 32903
rect -25920 32583 -25897 32617
rect -25863 32583 -25840 32617
rect -25920 32297 -25840 32583
rect -25920 32263 -25897 32297
rect -25863 32263 -25840 32297
rect -25920 31977 -25840 32263
rect -25920 31943 -25897 31977
rect -25863 31943 -25840 31977
rect -25920 31920 -25840 31943
rect -25760 32937 -25680 32960
rect -25760 32903 -25737 32937
rect -25703 32903 -25680 32937
rect -25760 32617 -25680 32903
rect -25760 32583 -25737 32617
rect -25703 32583 -25680 32617
rect -25760 32297 -25680 32583
rect -25760 32263 -25737 32297
rect -25703 32263 -25680 32297
rect -25760 31977 -25680 32263
rect -25760 31943 -25737 31977
rect -25703 31943 -25680 31977
rect -25760 31920 -25680 31943
rect -25600 32937 -25520 32960
rect -25600 32903 -25577 32937
rect -25543 32903 -25520 32937
rect -25600 32617 -25520 32903
rect -25600 32583 -25577 32617
rect -25543 32583 -25520 32617
rect -25600 32297 -25520 32583
rect -25600 32263 -25577 32297
rect -25543 32263 -25520 32297
rect -25600 31977 -25520 32263
rect -25600 31943 -25577 31977
rect -25543 31943 -25520 31977
rect -25600 31920 -25520 31943
rect -25440 32937 -25360 32960
rect -25440 32903 -25417 32937
rect -25383 32903 -25360 32937
rect -25440 32617 -25360 32903
rect -25440 32583 -25417 32617
rect -25383 32583 -25360 32617
rect -25440 32297 -25360 32583
rect -25440 32263 -25417 32297
rect -25383 32263 -25360 32297
rect -25440 31977 -25360 32263
rect -25440 31943 -25417 31977
rect -25383 31943 -25360 31977
rect -25440 31920 -25360 31943
rect -25280 32937 -25200 32960
rect -25280 32903 -25257 32937
rect -25223 32903 -25200 32937
rect -25280 32617 -25200 32903
rect -25280 32583 -25257 32617
rect -25223 32583 -25200 32617
rect -25280 32297 -25200 32583
rect -25280 32263 -25257 32297
rect -25223 32263 -25200 32297
rect -25280 31977 -25200 32263
rect -25280 31943 -25257 31977
rect -25223 31943 -25200 31977
rect -25280 31920 -25200 31943
rect -25120 32937 -25040 32960
rect -25120 32903 -25097 32937
rect -25063 32903 -25040 32937
rect -25120 32617 -25040 32903
rect -25120 32583 -25097 32617
rect -25063 32583 -25040 32617
rect -25120 32297 -25040 32583
rect -25120 32263 -25097 32297
rect -25063 32263 -25040 32297
rect -25120 31977 -25040 32263
rect -25120 31943 -25097 31977
rect -25063 31943 -25040 31977
rect -25120 31920 -25040 31943
rect -24960 32937 -24880 32960
rect -24960 32903 -24937 32937
rect -24903 32903 -24880 32937
rect -24960 32617 -24880 32903
rect -24960 32583 -24937 32617
rect -24903 32583 -24880 32617
rect -24960 32297 -24880 32583
rect -24960 32263 -24937 32297
rect -24903 32263 -24880 32297
rect -24960 31977 -24880 32263
rect -24960 31943 -24937 31977
rect -24903 31943 -24880 31977
rect -24960 31920 -24880 31943
rect -24800 32937 -24720 32960
rect -24800 32903 -24777 32937
rect -24743 32903 -24720 32937
rect -24800 32617 -24720 32903
rect -24800 32583 -24777 32617
rect -24743 32583 -24720 32617
rect -24800 32297 -24720 32583
rect -24800 32263 -24777 32297
rect -24743 32263 -24720 32297
rect -24800 31977 -24720 32263
rect -24800 31943 -24777 31977
rect -24743 31943 -24720 31977
rect -24800 31920 -24720 31943
rect -24640 32937 -24560 32960
rect -24640 32903 -24617 32937
rect -24583 32903 -24560 32937
rect -24640 32617 -24560 32903
rect -24640 32583 -24617 32617
rect -24583 32583 -24560 32617
rect -24640 32297 -24560 32583
rect -24640 32263 -24617 32297
rect -24583 32263 -24560 32297
rect -24640 31977 -24560 32263
rect -24640 31943 -24617 31977
rect -24583 31943 -24560 31977
rect -24640 31920 -24560 31943
rect -24480 32937 -24400 32960
rect -24480 32903 -24457 32937
rect -24423 32903 -24400 32937
rect -24480 32617 -24400 32903
rect -24480 32583 -24457 32617
rect -24423 32583 -24400 32617
rect -24480 32297 -24400 32583
rect -24480 32263 -24457 32297
rect -24423 32263 -24400 32297
rect -24480 31977 -24400 32263
rect -24480 31943 -24457 31977
rect -24423 31943 -24400 31977
rect -24480 31920 -24400 31943
rect -24320 32937 -24240 32960
rect -24320 32903 -24297 32937
rect -24263 32903 -24240 32937
rect -24320 32617 -24240 32903
rect -24320 32583 -24297 32617
rect -24263 32583 -24240 32617
rect -24320 32297 -24240 32583
rect -24320 32263 -24297 32297
rect -24263 32263 -24240 32297
rect -24320 31977 -24240 32263
rect -24320 31943 -24297 31977
rect -24263 31943 -24240 31977
rect -24320 31920 -24240 31943
rect -24160 32937 -24080 32960
rect -24160 32903 -24137 32937
rect -24103 32903 -24080 32937
rect -24160 32617 -24080 32903
rect -24160 32583 -24137 32617
rect -24103 32583 -24080 32617
rect -24160 32297 -24080 32583
rect -24160 32263 -24137 32297
rect -24103 32263 -24080 32297
rect -24160 31977 -24080 32263
rect -24160 31943 -24137 31977
rect -24103 31943 -24080 31977
rect -24160 31920 -24080 31943
rect -24000 32937 -23920 32960
rect -24000 32903 -23977 32937
rect -23943 32903 -23920 32937
rect -24000 32617 -23920 32903
rect -24000 32583 -23977 32617
rect -23943 32583 -23920 32617
rect -24000 32297 -23920 32583
rect -24000 32263 -23977 32297
rect -23943 32263 -23920 32297
rect -24000 31977 -23920 32263
rect -24000 31943 -23977 31977
rect -23943 31943 -23920 31977
rect -24000 31920 -23920 31943
rect -23840 32937 -23760 32960
rect -23840 32903 -23817 32937
rect -23783 32903 -23760 32937
rect -23840 32617 -23760 32903
rect -23840 32583 -23817 32617
rect -23783 32583 -23760 32617
rect -23840 32297 -23760 32583
rect -23840 32263 -23817 32297
rect -23783 32263 -23760 32297
rect -23840 31977 -23760 32263
rect -23840 31943 -23817 31977
rect -23783 31943 -23760 31977
rect -23840 31920 -23760 31943
rect -23680 32937 -23600 32960
rect -23680 32903 -23657 32937
rect -23623 32903 -23600 32937
rect -23680 32617 -23600 32903
rect -23680 32583 -23657 32617
rect -23623 32583 -23600 32617
rect -23680 32297 -23600 32583
rect -23680 32263 -23657 32297
rect -23623 32263 -23600 32297
rect -23680 31977 -23600 32263
rect -23680 31943 -23657 31977
rect -23623 31943 -23600 31977
rect -23680 31920 -23600 31943
rect -23520 32937 -23440 32960
rect -23520 32903 -23497 32937
rect -23463 32903 -23440 32937
rect -23520 32617 -23440 32903
rect -23520 32583 -23497 32617
rect -23463 32583 -23440 32617
rect -23520 32297 -23440 32583
rect -23520 32263 -23497 32297
rect -23463 32263 -23440 32297
rect -23520 31977 -23440 32263
rect -23520 31943 -23497 31977
rect -23463 31943 -23440 31977
rect -23520 31920 -23440 31943
rect -23360 32937 -23280 32960
rect -23360 32903 -23337 32937
rect -23303 32903 -23280 32937
rect -23360 32617 -23280 32903
rect -23360 32583 -23337 32617
rect -23303 32583 -23280 32617
rect -23360 32297 -23280 32583
rect -23360 32263 -23337 32297
rect -23303 32263 -23280 32297
rect -23360 31977 -23280 32263
rect -23360 31943 -23337 31977
rect -23303 31943 -23280 31977
rect -23360 31920 -23280 31943
rect -23200 32937 -23120 32960
rect -23200 32903 -23177 32937
rect -23143 32903 -23120 32937
rect -23200 32617 -23120 32903
rect -23200 32583 -23177 32617
rect -23143 32583 -23120 32617
rect -23200 32297 -23120 32583
rect -23200 32263 -23177 32297
rect -23143 32263 -23120 32297
rect -23200 31977 -23120 32263
rect -23200 31943 -23177 31977
rect -23143 31943 -23120 31977
rect -23200 31920 -23120 31943
rect -23040 32937 -22960 32960
rect -23040 32903 -23017 32937
rect -22983 32903 -22960 32937
rect -23040 32617 -22960 32903
rect -23040 32583 -23017 32617
rect -22983 32583 -22960 32617
rect -23040 32297 -22960 32583
rect -23040 32263 -23017 32297
rect -22983 32263 -22960 32297
rect -23040 31977 -22960 32263
rect -23040 31943 -23017 31977
rect -22983 31943 -22960 31977
rect -23040 31920 -22960 31943
rect -22880 32937 -22800 32960
rect -22880 32903 -22857 32937
rect -22823 32903 -22800 32937
rect -22880 32617 -22800 32903
rect -22880 32583 -22857 32617
rect -22823 32583 -22800 32617
rect -22880 32297 -22800 32583
rect -22880 32263 -22857 32297
rect -22823 32263 -22800 32297
rect -22880 31977 -22800 32263
rect -22880 31943 -22857 31977
rect -22823 31943 -22800 31977
rect -22880 31920 -22800 31943
rect -22720 32937 -22640 32960
rect -22720 32903 -22697 32937
rect -22663 32903 -22640 32937
rect -22720 32617 -22640 32903
rect -22720 32583 -22697 32617
rect -22663 32583 -22640 32617
rect -22720 32297 -22640 32583
rect -22720 32263 -22697 32297
rect -22663 32263 -22640 32297
rect -22720 31977 -22640 32263
rect -22720 31943 -22697 31977
rect -22663 31943 -22640 31977
rect -22720 31920 -22640 31943
rect -22560 32937 -22480 32960
rect -22560 32903 -22537 32937
rect -22503 32903 -22480 32937
rect -22560 32617 -22480 32903
rect -22560 32583 -22537 32617
rect -22503 32583 -22480 32617
rect -22560 32297 -22480 32583
rect -22560 32263 -22537 32297
rect -22503 32263 -22480 32297
rect -22560 31977 -22480 32263
rect -22560 31943 -22537 31977
rect -22503 31943 -22480 31977
rect -22560 31920 -22480 31943
rect -22400 32937 -22320 32960
rect -22400 32903 -22377 32937
rect -22343 32903 -22320 32937
rect -22400 32617 -22320 32903
rect -22400 32583 -22377 32617
rect -22343 32583 -22320 32617
rect -22400 32297 -22320 32583
rect -22400 32263 -22377 32297
rect -22343 32263 -22320 32297
rect -22400 31977 -22320 32263
rect -22400 31943 -22377 31977
rect -22343 31943 -22320 31977
rect -22400 31920 -22320 31943
rect -22240 32937 -22160 32960
rect -22240 32903 -22217 32937
rect -22183 32903 -22160 32937
rect -22240 32617 -22160 32903
rect -22240 32583 -22217 32617
rect -22183 32583 -22160 32617
rect -22240 32297 -22160 32583
rect -22240 32263 -22217 32297
rect -22183 32263 -22160 32297
rect -22240 31977 -22160 32263
rect -22240 31943 -22217 31977
rect -22183 31943 -22160 31977
rect -22240 31920 -22160 31943
rect -22080 32937 -22000 32960
rect -22080 32903 -22057 32937
rect -22023 32903 -22000 32937
rect -22080 32617 -22000 32903
rect -22080 32583 -22057 32617
rect -22023 32583 -22000 32617
rect -22080 32297 -22000 32583
rect -22080 32263 -22057 32297
rect -22023 32263 -22000 32297
rect -22080 31977 -22000 32263
rect -22080 31943 -22057 31977
rect -22023 31943 -22000 31977
rect -22080 31920 -22000 31943
rect -21920 32937 -21840 32960
rect -21920 32903 -21897 32937
rect -21863 32903 -21840 32937
rect -21920 32617 -21840 32903
rect -21920 32583 -21897 32617
rect -21863 32583 -21840 32617
rect -21920 32297 -21840 32583
rect -21920 32263 -21897 32297
rect -21863 32263 -21840 32297
rect -21920 31977 -21840 32263
rect -21920 31943 -21897 31977
rect -21863 31943 -21840 31977
rect -21920 31920 -21840 31943
rect -21760 32937 -21680 32960
rect -21760 32903 -21737 32937
rect -21703 32903 -21680 32937
rect -21760 32617 -21680 32903
rect -21760 32583 -21737 32617
rect -21703 32583 -21680 32617
rect -21760 32297 -21680 32583
rect -21760 32263 -21737 32297
rect -21703 32263 -21680 32297
rect -21760 31977 -21680 32263
rect -21760 31943 -21737 31977
rect -21703 31943 -21680 31977
rect -21760 31920 -21680 31943
rect -21600 32937 -21520 32960
rect -21600 32903 -21577 32937
rect -21543 32903 -21520 32937
rect -21600 32617 -21520 32903
rect -21600 32583 -21577 32617
rect -21543 32583 -21520 32617
rect -21600 32297 -21520 32583
rect -21600 32263 -21577 32297
rect -21543 32263 -21520 32297
rect -21600 31977 -21520 32263
rect -21600 31943 -21577 31977
rect -21543 31943 -21520 31977
rect -21600 31920 -21520 31943
rect -21440 32937 -21360 32960
rect -21440 32903 -21417 32937
rect -21383 32903 -21360 32937
rect -21440 32617 -21360 32903
rect -21440 32583 -21417 32617
rect -21383 32583 -21360 32617
rect -21440 32297 -21360 32583
rect -21440 32263 -21417 32297
rect -21383 32263 -21360 32297
rect -21440 31977 -21360 32263
rect -21440 31943 -21417 31977
rect -21383 31943 -21360 31977
rect -21440 31920 -21360 31943
rect -21280 32937 -21200 32960
rect -21280 32903 -21257 32937
rect -21223 32903 -21200 32937
rect -21280 32617 -21200 32903
rect -21280 32583 -21257 32617
rect -21223 32583 -21200 32617
rect -21280 32297 -21200 32583
rect -21280 32263 -21257 32297
rect -21223 32263 -21200 32297
rect -21280 31977 -21200 32263
rect -21280 31943 -21257 31977
rect -21223 31943 -21200 31977
rect -21280 31920 -21200 31943
rect -21120 32937 -21040 32960
rect -21120 32903 -21097 32937
rect -21063 32903 -21040 32937
rect -21120 32617 -21040 32903
rect -21120 32583 -21097 32617
rect -21063 32583 -21040 32617
rect -21120 32297 -21040 32583
rect -21120 32263 -21097 32297
rect -21063 32263 -21040 32297
rect -21120 31977 -21040 32263
rect -21120 31943 -21097 31977
rect -21063 31943 -21040 31977
rect -21120 31920 -21040 31943
rect -20960 32937 -20880 32960
rect -20960 32903 -20937 32937
rect -20903 32903 -20880 32937
rect -20960 32617 -20880 32903
rect -20960 32583 -20937 32617
rect -20903 32583 -20880 32617
rect -20960 32297 -20880 32583
rect -20960 32263 -20937 32297
rect -20903 32263 -20880 32297
rect -20960 31977 -20880 32263
rect -20960 31943 -20937 31977
rect -20903 31943 -20880 31977
rect -20960 31920 -20880 31943
rect -20800 32937 -20720 32960
rect -20800 32903 -20777 32937
rect -20743 32903 -20720 32937
rect -20800 32617 -20720 32903
rect -20800 32583 -20777 32617
rect -20743 32583 -20720 32617
rect -20800 32297 -20720 32583
rect -20800 32263 -20777 32297
rect -20743 32263 -20720 32297
rect -20800 31977 -20720 32263
rect -20800 31943 -20777 31977
rect -20743 31943 -20720 31977
rect -20800 31920 -20720 31943
rect -20640 32937 -20560 32960
rect -20640 32903 -20617 32937
rect -20583 32903 -20560 32937
rect -20640 32617 -20560 32903
rect -20640 32583 -20617 32617
rect -20583 32583 -20560 32617
rect -20640 32297 -20560 32583
rect -20640 32263 -20617 32297
rect -20583 32263 -20560 32297
rect -20640 31977 -20560 32263
rect -20640 31943 -20617 31977
rect -20583 31943 -20560 31977
rect -20640 31920 -20560 31943
rect -20480 32937 -20400 32960
rect -20480 32903 -20457 32937
rect -20423 32903 -20400 32937
rect -20480 32617 -20400 32903
rect -20480 32583 -20457 32617
rect -20423 32583 -20400 32617
rect -20480 32297 -20400 32583
rect -20480 32263 -20457 32297
rect -20423 32263 -20400 32297
rect -20480 31977 -20400 32263
rect -20480 31943 -20457 31977
rect -20423 31943 -20400 31977
rect -20480 31920 -20400 31943
rect -20320 32937 -20240 32960
rect -20320 32903 -20297 32937
rect -20263 32903 -20240 32937
rect -20320 32617 -20240 32903
rect -20320 32583 -20297 32617
rect -20263 32583 -20240 32617
rect -20320 32297 -20240 32583
rect -20320 32263 -20297 32297
rect -20263 32263 -20240 32297
rect -20320 31977 -20240 32263
rect -20320 31943 -20297 31977
rect -20263 31943 -20240 31977
rect -20320 31920 -20240 31943
rect -20160 32937 -20080 32960
rect -20160 32903 -20137 32937
rect -20103 32903 -20080 32937
rect -20160 32617 -20080 32903
rect -20160 32583 -20137 32617
rect -20103 32583 -20080 32617
rect -20160 32297 -20080 32583
rect -20160 32263 -20137 32297
rect -20103 32263 -20080 32297
rect -20160 31977 -20080 32263
rect -20160 31943 -20137 31977
rect -20103 31943 -20080 31977
rect -20160 31920 -20080 31943
rect -20000 32937 -19920 32960
rect -20000 32903 -19977 32937
rect -19943 32903 -19920 32937
rect -20000 32617 -19920 32903
rect -20000 32583 -19977 32617
rect -19943 32583 -19920 32617
rect -20000 32297 -19920 32583
rect -20000 32263 -19977 32297
rect -19943 32263 -19920 32297
rect -20000 31977 -19920 32263
rect -20000 31943 -19977 31977
rect -19943 31943 -19920 31977
rect -20000 31920 -19920 31943
rect -19840 32937 -19760 32960
rect -19840 32903 -19817 32937
rect -19783 32903 -19760 32937
rect -19840 32617 -19760 32903
rect -19840 32583 -19817 32617
rect -19783 32583 -19760 32617
rect -19840 32297 -19760 32583
rect -19840 32263 -19817 32297
rect -19783 32263 -19760 32297
rect -19840 31977 -19760 32263
rect -19840 31943 -19817 31977
rect -19783 31943 -19760 31977
rect -19840 31920 -19760 31943
rect -19680 32937 -19600 32960
rect -19680 32903 -19657 32937
rect -19623 32903 -19600 32937
rect -19680 32617 -19600 32903
rect -19680 32583 -19657 32617
rect -19623 32583 -19600 32617
rect -19680 32297 -19600 32583
rect -19680 32263 -19657 32297
rect -19623 32263 -19600 32297
rect -19680 31977 -19600 32263
rect -19680 31943 -19657 31977
rect -19623 31943 -19600 31977
rect -19680 31920 -19600 31943
rect -19520 32937 -19440 32960
rect -19520 32903 -19497 32937
rect -19463 32903 -19440 32937
rect -19520 32617 -19440 32903
rect -19520 32583 -19497 32617
rect -19463 32583 -19440 32617
rect -19520 32297 -19440 32583
rect -19520 32263 -19497 32297
rect -19463 32263 -19440 32297
rect -19520 31977 -19440 32263
rect -19520 31943 -19497 31977
rect -19463 31943 -19440 31977
rect -19520 31920 -19440 31943
rect -19360 32937 -19280 32960
rect -19360 32903 -19337 32937
rect -19303 32903 -19280 32937
rect -19360 32617 -19280 32903
rect -19360 32583 -19337 32617
rect -19303 32583 -19280 32617
rect -19360 32297 -19280 32583
rect -19360 32263 -19337 32297
rect -19303 32263 -19280 32297
rect -19360 31977 -19280 32263
rect -19360 31943 -19337 31977
rect -19303 31943 -19280 31977
rect -19360 31920 -19280 31943
rect -19200 32937 -19120 32960
rect -19200 32903 -19177 32937
rect -19143 32903 -19120 32937
rect -19200 32617 -19120 32903
rect -19200 32583 -19177 32617
rect -19143 32583 -19120 32617
rect -19200 32297 -19120 32583
rect -19200 32263 -19177 32297
rect -19143 32263 -19120 32297
rect -19200 31977 -19120 32263
rect -19200 31943 -19177 31977
rect -19143 31943 -19120 31977
rect -19200 31920 -19120 31943
rect -19040 32937 -18960 32960
rect -19040 32903 -19017 32937
rect -18983 32903 -18960 32937
rect -19040 32617 -18960 32903
rect -19040 32583 -19017 32617
rect -18983 32583 -18960 32617
rect -19040 32297 -18960 32583
rect -19040 32263 -19017 32297
rect -18983 32263 -18960 32297
rect -19040 31977 -18960 32263
rect -19040 31943 -19017 31977
rect -18983 31943 -18960 31977
rect -19040 31920 -18960 31943
rect -18880 32937 -18800 32960
rect -18880 32903 -18857 32937
rect -18823 32903 -18800 32937
rect -18880 32617 -18800 32903
rect -18880 32583 -18857 32617
rect -18823 32583 -18800 32617
rect -18880 32297 -18800 32583
rect -18880 32263 -18857 32297
rect -18823 32263 -18800 32297
rect -18880 31977 -18800 32263
rect -18880 31943 -18857 31977
rect -18823 31943 -18800 31977
rect -18880 31920 -18800 31943
rect -18720 32937 -18640 32960
rect -18720 32903 -18697 32937
rect -18663 32903 -18640 32937
rect -18720 32617 -18640 32903
rect -18720 32583 -18697 32617
rect -18663 32583 -18640 32617
rect -18720 32297 -18640 32583
rect -18720 32263 -18697 32297
rect -18663 32263 -18640 32297
rect -18720 31977 -18640 32263
rect -18720 31943 -18697 31977
rect -18663 31943 -18640 31977
rect -18720 31920 -18640 31943
rect -18560 32937 -18480 32960
rect -18560 32903 -18537 32937
rect -18503 32903 -18480 32937
rect -18560 32617 -18480 32903
rect -18560 32583 -18537 32617
rect -18503 32583 -18480 32617
rect -18560 32297 -18480 32583
rect -18560 32263 -18537 32297
rect -18503 32263 -18480 32297
rect -18560 31977 -18480 32263
rect -18560 31943 -18537 31977
rect -18503 31943 -18480 31977
rect -18560 31920 -18480 31943
rect -18400 32937 -18320 32960
rect -18400 32903 -18377 32937
rect -18343 32903 -18320 32937
rect -18400 32617 -18320 32903
rect -18400 32583 -18377 32617
rect -18343 32583 -18320 32617
rect -18400 32297 -18320 32583
rect -18400 32263 -18377 32297
rect -18343 32263 -18320 32297
rect -18400 31977 -18320 32263
rect -18400 31943 -18377 31977
rect -18343 31943 -18320 31977
rect -18400 31920 -18320 31943
rect -18240 32937 -18160 32960
rect -18240 32903 -18217 32937
rect -18183 32903 -18160 32937
rect -18240 32617 -18160 32903
rect -18240 32583 -18217 32617
rect -18183 32583 -18160 32617
rect -18240 32297 -18160 32583
rect -18240 32263 -18217 32297
rect -18183 32263 -18160 32297
rect -18240 31977 -18160 32263
rect -18240 31943 -18217 31977
rect -18183 31943 -18160 31977
rect -18240 31920 -18160 31943
rect -18080 32937 -18000 32960
rect -18080 32903 -18057 32937
rect -18023 32903 -18000 32937
rect -18080 32617 -18000 32903
rect -18080 32583 -18057 32617
rect -18023 32583 -18000 32617
rect -18080 32297 -18000 32583
rect -18080 32263 -18057 32297
rect -18023 32263 -18000 32297
rect -18080 31977 -18000 32263
rect -18080 31943 -18057 31977
rect -18023 31943 -18000 31977
rect -18080 31920 -18000 31943
rect -17920 32937 -17840 32960
rect -17920 32903 -17897 32937
rect -17863 32903 -17840 32937
rect -17920 32617 -17840 32903
rect -17920 32583 -17897 32617
rect -17863 32583 -17840 32617
rect -17920 32297 -17840 32583
rect -17920 32263 -17897 32297
rect -17863 32263 -17840 32297
rect -17920 31977 -17840 32263
rect -17920 31943 -17897 31977
rect -17863 31943 -17840 31977
rect -17920 31920 -17840 31943
rect -17760 32937 -17680 32960
rect -17760 32903 -17737 32937
rect -17703 32903 -17680 32937
rect -17760 32617 -17680 32903
rect -17760 32583 -17737 32617
rect -17703 32583 -17680 32617
rect -17760 32297 -17680 32583
rect -17760 32263 -17737 32297
rect -17703 32263 -17680 32297
rect -17760 31977 -17680 32263
rect -17760 31943 -17737 31977
rect -17703 31943 -17680 31977
rect -17760 31920 -17680 31943
rect -17600 32937 -17520 32960
rect -17600 32903 -17577 32937
rect -17543 32903 -17520 32937
rect -17600 32617 -17520 32903
rect -17600 32583 -17577 32617
rect -17543 32583 -17520 32617
rect -17600 32297 -17520 32583
rect -17600 32263 -17577 32297
rect -17543 32263 -17520 32297
rect -17600 31977 -17520 32263
rect -17600 31943 -17577 31977
rect -17543 31943 -17520 31977
rect -17600 31920 -17520 31943
rect -17440 32937 -17360 32960
rect -17440 32903 -17417 32937
rect -17383 32903 -17360 32937
rect -17440 32617 -17360 32903
rect -17440 32583 -17417 32617
rect -17383 32583 -17360 32617
rect -17440 32297 -17360 32583
rect -17440 32263 -17417 32297
rect -17383 32263 -17360 32297
rect -17440 31977 -17360 32263
rect -17440 31943 -17417 31977
rect -17383 31943 -17360 31977
rect -17440 31920 -17360 31943
rect -17280 32937 -17200 32960
rect -17280 32903 -17257 32937
rect -17223 32903 -17200 32937
rect -17280 32617 -17200 32903
rect -17280 32583 -17257 32617
rect -17223 32583 -17200 32617
rect -17280 32297 -17200 32583
rect -17280 32263 -17257 32297
rect -17223 32263 -17200 32297
rect -17280 31977 -17200 32263
rect -17280 31943 -17257 31977
rect -17223 31943 -17200 31977
rect -17280 31920 -17200 31943
rect -17120 32937 -17040 32960
rect -17120 32903 -17097 32937
rect -17063 32903 -17040 32937
rect -17120 32617 -17040 32903
rect -17120 32583 -17097 32617
rect -17063 32583 -17040 32617
rect -17120 32297 -17040 32583
rect -17120 32263 -17097 32297
rect -17063 32263 -17040 32297
rect -17120 31977 -17040 32263
rect -17120 31943 -17097 31977
rect -17063 31943 -17040 31977
rect -17120 31920 -17040 31943
rect -16960 32937 -16880 32960
rect -16960 32903 -16937 32937
rect -16903 32903 -16880 32937
rect -16960 32617 -16880 32903
rect -16960 32583 -16937 32617
rect -16903 32583 -16880 32617
rect -16960 32297 -16880 32583
rect -16960 32263 -16937 32297
rect -16903 32263 -16880 32297
rect -16960 31977 -16880 32263
rect -16960 31943 -16937 31977
rect -16903 31943 -16880 31977
rect -16960 31920 -16880 31943
rect -16800 32937 -16720 32960
rect -16800 32903 -16777 32937
rect -16743 32903 -16720 32937
rect -16800 32617 -16720 32903
rect -16800 32583 -16777 32617
rect -16743 32583 -16720 32617
rect -16800 32297 -16720 32583
rect -16800 32263 -16777 32297
rect -16743 32263 -16720 32297
rect -16800 31977 -16720 32263
rect -16800 31943 -16777 31977
rect -16743 31943 -16720 31977
rect -16800 31920 -16720 31943
rect -16640 32937 -16560 32960
rect -16640 32903 -16617 32937
rect -16583 32903 -16560 32937
rect -16640 32617 -16560 32903
rect -16640 32583 -16617 32617
rect -16583 32583 -16560 32617
rect -16640 32297 -16560 32583
rect -16640 32263 -16617 32297
rect -16583 32263 -16560 32297
rect -16640 31977 -16560 32263
rect -16640 31943 -16617 31977
rect -16583 31943 -16560 31977
rect -16640 31920 -16560 31943
rect -16480 32937 -16400 32960
rect -16480 32903 -16457 32937
rect -16423 32903 -16400 32937
rect -16480 32617 -16400 32903
rect -16480 32583 -16457 32617
rect -16423 32583 -16400 32617
rect -16480 32297 -16400 32583
rect -16480 32263 -16457 32297
rect -16423 32263 -16400 32297
rect -16480 31977 -16400 32263
rect -16480 31943 -16457 31977
rect -16423 31943 -16400 31977
rect -16480 31920 -16400 31943
rect -16320 32937 -16240 32960
rect -16320 32903 -16297 32937
rect -16263 32903 -16240 32937
rect -16320 32617 -16240 32903
rect -16320 32583 -16297 32617
rect -16263 32583 -16240 32617
rect -16320 32297 -16240 32583
rect -16320 32263 -16297 32297
rect -16263 32263 -16240 32297
rect -16320 31977 -16240 32263
rect -16320 31943 -16297 31977
rect -16263 31943 -16240 31977
rect -16320 31920 -16240 31943
rect -16160 32937 -16080 32960
rect -16160 32903 -16137 32937
rect -16103 32903 -16080 32937
rect -16160 32617 -16080 32903
rect -16160 32583 -16137 32617
rect -16103 32583 -16080 32617
rect -16160 32297 -16080 32583
rect -16160 32263 -16137 32297
rect -16103 32263 -16080 32297
rect -16160 31977 -16080 32263
rect -16160 31943 -16137 31977
rect -16103 31943 -16080 31977
rect -16160 31920 -16080 31943
rect -16000 32937 -15920 32960
rect -16000 32903 -15977 32937
rect -15943 32903 -15920 32937
rect -16000 32617 -15920 32903
rect -16000 32583 -15977 32617
rect -15943 32583 -15920 32617
rect -16000 32297 -15920 32583
rect -16000 32263 -15977 32297
rect -15943 32263 -15920 32297
rect -16000 31977 -15920 32263
rect -16000 31943 -15977 31977
rect -15943 31943 -15920 31977
rect -16000 31920 -15920 31943
rect -15840 32937 -15760 32960
rect -15840 32903 -15817 32937
rect -15783 32903 -15760 32937
rect -15840 32617 -15760 32903
rect -15840 32583 -15817 32617
rect -15783 32583 -15760 32617
rect -15840 32297 -15760 32583
rect -15840 32263 -15817 32297
rect -15783 32263 -15760 32297
rect -15840 31977 -15760 32263
rect -15840 31943 -15817 31977
rect -15783 31943 -15760 31977
rect -15840 31920 -15760 31943
rect -15680 32937 -15600 32960
rect -15680 32903 -15657 32937
rect -15623 32903 -15600 32937
rect -15680 32617 -15600 32903
rect -15680 32583 -15657 32617
rect -15623 32583 -15600 32617
rect -15680 32297 -15600 32583
rect -15680 32263 -15657 32297
rect -15623 32263 -15600 32297
rect -15680 31977 -15600 32263
rect -15680 31943 -15657 31977
rect -15623 31943 -15600 31977
rect -15680 31920 -15600 31943
rect -15520 32937 -15440 32960
rect -15520 32903 -15497 32937
rect -15463 32903 -15440 32937
rect -15520 32617 -15440 32903
rect -15520 32583 -15497 32617
rect -15463 32583 -15440 32617
rect -15520 32297 -15440 32583
rect -15520 32263 -15497 32297
rect -15463 32263 -15440 32297
rect -15520 31977 -15440 32263
rect -15520 31943 -15497 31977
rect -15463 31943 -15440 31977
rect -15520 31920 -15440 31943
rect -15360 32937 -15280 32960
rect -15360 32903 -15337 32937
rect -15303 32903 -15280 32937
rect -15360 32617 -15280 32903
rect -15360 32583 -15337 32617
rect -15303 32583 -15280 32617
rect -15360 32297 -15280 32583
rect -15360 32263 -15337 32297
rect -15303 32263 -15280 32297
rect -15360 31977 -15280 32263
rect -15360 31943 -15337 31977
rect -15303 31943 -15280 31977
rect -15360 31920 -15280 31943
rect -15200 32937 -15120 32960
rect -15200 32903 -15177 32937
rect -15143 32903 -15120 32937
rect -15200 32617 -15120 32903
rect -15200 32583 -15177 32617
rect -15143 32583 -15120 32617
rect -15200 32297 -15120 32583
rect -15200 32263 -15177 32297
rect -15143 32263 -15120 32297
rect -15200 31977 -15120 32263
rect -15200 31943 -15177 31977
rect -15143 31943 -15120 31977
rect -15200 31920 -15120 31943
rect -15040 32937 -14960 32960
rect -15040 32903 -15017 32937
rect -14983 32903 -14960 32937
rect -15040 32617 -14960 32903
rect -15040 32583 -15017 32617
rect -14983 32583 -14960 32617
rect -15040 32297 -14960 32583
rect -15040 32263 -15017 32297
rect -14983 32263 -14960 32297
rect -15040 31977 -14960 32263
rect -15040 31943 -15017 31977
rect -14983 31943 -14960 31977
rect -15040 31920 -14960 31943
rect -14880 32937 -14800 32960
rect -14880 32903 -14857 32937
rect -14823 32903 -14800 32937
rect -14880 32617 -14800 32903
rect -14880 32583 -14857 32617
rect -14823 32583 -14800 32617
rect -14880 32297 -14800 32583
rect -14880 32263 -14857 32297
rect -14823 32263 -14800 32297
rect -14880 31977 -14800 32263
rect -14880 31943 -14857 31977
rect -14823 31943 -14800 31977
rect -14880 31920 -14800 31943
rect -14720 32937 -14640 32960
rect -14720 32903 -14697 32937
rect -14663 32903 -14640 32937
rect -14720 32617 -14640 32903
rect -14720 32583 -14697 32617
rect -14663 32583 -14640 32617
rect -14720 32297 -14640 32583
rect -14720 32263 -14697 32297
rect -14663 32263 -14640 32297
rect -14720 31977 -14640 32263
rect -14720 31943 -14697 31977
rect -14663 31943 -14640 31977
rect -14720 31920 -14640 31943
rect -14560 32937 -14480 32960
rect -14560 32903 -14537 32937
rect -14503 32903 -14480 32937
rect -14560 32617 -14480 32903
rect -14560 32583 -14537 32617
rect -14503 32583 -14480 32617
rect -14560 32297 -14480 32583
rect -14560 32263 -14537 32297
rect -14503 32263 -14480 32297
rect -14560 31977 -14480 32263
rect -14560 31943 -14537 31977
rect -14503 31943 -14480 31977
rect -14560 31920 -14480 31943
rect -14400 32937 -14320 32960
rect -14400 32903 -14377 32937
rect -14343 32903 -14320 32937
rect -14400 32617 -14320 32903
rect -14400 32583 -14377 32617
rect -14343 32583 -14320 32617
rect -14400 32297 -14320 32583
rect -14400 32263 -14377 32297
rect -14343 32263 -14320 32297
rect -14400 31977 -14320 32263
rect -14400 31943 -14377 31977
rect -14343 31943 -14320 31977
rect -14400 31920 -14320 31943
rect -14240 32937 -14160 32960
rect -14240 32903 -14217 32937
rect -14183 32903 -14160 32937
rect -14240 32617 -14160 32903
rect -14240 32583 -14217 32617
rect -14183 32583 -14160 32617
rect -14240 32297 -14160 32583
rect -14240 32263 -14217 32297
rect -14183 32263 -14160 32297
rect -14240 31977 -14160 32263
rect -14240 31943 -14217 31977
rect -14183 31943 -14160 31977
rect -14240 31920 -14160 31943
rect -14080 32937 -14000 32960
rect -14080 32903 -14057 32937
rect -14023 32903 -14000 32937
rect -14080 32617 -14000 32903
rect -14080 32583 -14057 32617
rect -14023 32583 -14000 32617
rect -14080 32297 -14000 32583
rect -14080 32263 -14057 32297
rect -14023 32263 -14000 32297
rect -14080 31977 -14000 32263
rect -14080 31943 -14057 31977
rect -14023 31943 -14000 31977
rect -14080 31920 -14000 31943
rect -13920 32937 -13840 32960
rect -13920 32903 -13897 32937
rect -13863 32903 -13840 32937
rect -13920 32617 -13840 32903
rect -13920 32583 -13897 32617
rect -13863 32583 -13840 32617
rect -13920 32297 -13840 32583
rect -13920 32263 -13897 32297
rect -13863 32263 -13840 32297
rect -13920 31977 -13840 32263
rect -13920 31943 -13897 31977
rect -13863 31943 -13840 31977
rect -13920 31920 -13840 31943
rect -13760 32937 -13680 32960
rect -13760 32903 -13737 32937
rect -13703 32903 -13680 32937
rect -13760 32617 -13680 32903
rect -13760 32583 -13737 32617
rect -13703 32583 -13680 32617
rect -13760 32297 -13680 32583
rect -13760 32263 -13737 32297
rect -13703 32263 -13680 32297
rect -13760 31977 -13680 32263
rect -13760 31943 -13737 31977
rect -13703 31943 -13680 31977
rect -13760 31920 -13680 31943
rect -13600 32937 -13520 32960
rect -13600 32903 -13577 32937
rect -13543 32903 -13520 32937
rect -13600 32617 -13520 32903
rect -13600 32583 -13577 32617
rect -13543 32583 -13520 32617
rect -13600 32297 -13520 32583
rect -13600 32263 -13577 32297
rect -13543 32263 -13520 32297
rect -13600 31977 -13520 32263
rect -13600 31943 -13577 31977
rect -13543 31943 -13520 31977
rect -13600 31920 -13520 31943
rect -13440 32937 -13360 32960
rect -13440 32903 -13417 32937
rect -13383 32903 -13360 32937
rect -13440 32617 -13360 32903
rect -13440 32583 -13417 32617
rect -13383 32583 -13360 32617
rect -13440 32297 -13360 32583
rect -13440 32263 -13417 32297
rect -13383 32263 -13360 32297
rect -13440 31977 -13360 32263
rect -13440 31943 -13417 31977
rect -13383 31943 -13360 31977
rect -13440 31920 -13360 31943
rect -13280 32937 -13200 32960
rect -13280 32903 -13257 32937
rect -13223 32903 -13200 32937
rect -13280 32617 -13200 32903
rect -13280 32583 -13257 32617
rect -13223 32583 -13200 32617
rect -13280 32297 -13200 32583
rect -13280 32263 -13257 32297
rect -13223 32263 -13200 32297
rect -13280 31977 -13200 32263
rect -13280 31943 -13257 31977
rect -13223 31943 -13200 31977
rect -13280 31920 -13200 31943
rect -13120 32937 -13040 32960
rect -13120 32903 -13097 32937
rect -13063 32903 -13040 32937
rect -13120 32617 -13040 32903
rect -13120 32583 -13097 32617
rect -13063 32583 -13040 32617
rect -13120 32297 -13040 32583
rect -13120 32263 -13097 32297
rect -13063 32263 -13040 32297
rect -13120 31977 -13040 32263
rect -13120 31943 -13097 31977
rect -13063 31943 -13040 31977
rect -13120 31920 -13040 31943
rect -12960 32937 -12880 32960
rect -12960 32903 -12937 32937
rect -12903 32903 -12880 32937
rect -12960 32617 -12880 32903
rect -12960 32583 -12937 32617
rect -12903 32583 -12880 32617
rect -12960 32297 -12880 32583
rect -12960 32263 -12937 32297
rect -12903 32263 -12880 32297
rect -12960 31977 -12880 32263
rect -12960 31943 -12937 31977
rect -12903 31943 -12880 31977
rect -12960 31920 -12880 31943
rect -12800 32937 -12720 32960
rect -12800 32903 -12777 32937
rect -12743 32903 -12720 32937
rect -12800 32617 -12720 32903
rect -12800 32583 -12777 32617
rect -12743 32583 -12720 32617
rect -12800 32297 -12720 32583
rect -12800 32263 -12777 32297
rect -12743 32263 -12720 32297
rect -12800 31977 -12720 32263
rect -12800 31943 -12777 31977
rect -12743 31943 -12720 31977
rect -12800 31920 -12720 31943
rect -12640 32937 -12560 32960
rect -12640 32903 -12617 32937
rect -12583 32903 -12560 32937
rect -12640 32617 -12560 32903
rect -12640 32583 -12617 32617
rect -12583 32583 -12560 32617
rect -12640 32297 -12560 32583
rect -12640 32263 -12617 32297
rect -12583 32263 -12560 32297
rect -12640 31977 -12560 32263
rect -12640 31943 -12617 31977
rect -12583 31943 -12560 31977
rect -12640 31920 -12560 31943
rect -12480 32937 -12400 32960
rect -12480 32903 -12457 32937
rect -12423 32903 -12400 32937
rect -12480 32617 -12400 32903
rect -12480 32583 -12457 32617
rect -12423 32583 -12400 32617
rect -12480 32297 -12400 32583
rect -12480 32263 -12457 32297
rect -12423 32263 -12400 32297
rect -12480 31977 -12400 32263
rect -12480 31943 -12457 31977
rect -12423 31943 -12400 31977
rect -12480 31920 -12400 31943
rect -12320 32937 -12240 32960
rect -12320 32903 -12297 32937
rect -12263 32903 -12240 32937
rect -12320 32617 -12240 32903
rect -12320 32583 -12297 32617
rect -12263 32583 -12240 32617
rect -12320 32297 -12240 32583
rect -12320 32263 -12297 32297
rect -12263 32263 -12240 32297
rect -12320 31977 -12240 32263
rect -12320 31943 -12297 31977
rect -12263 31943 -12240 31977
rect -12320 31920 -12240 31943
rect -12160 32937 -12080 32960
rect -12160 32903 -12137 32937
rect -12103 32903 -12080 32937
rect -12160 32617 -12080 32903
rect -12160 32583 -12137 32617
rect -12103 32583 -12080 32617
rect -12160 32297 -12080 32583
rect -12160 32263 -12137 32297
rect -12103 32263 -12080 32297
rect -12160 31977 -12080 32263
rect -12160 31943 -12137 31977
rect -12103 31943 -12080 31977
rect -12160 31920 -12080 31943
rect -12000 32937 -11920 32960
rect -12000 32903 -11977 32937
rect -11943 32903 -11920 32937
rect -12000 32617 -11920 32903
rect -12000 32583 -11977 32617
rect -11943 32583 -11920 32617
rect -12000 32297 -11920 32583
rect -12000 32263 -11977 32297
rect -11943 32263 -11920 32297
rect -12000 31977 -11920 32263
rect -12000 31943 -11977 31977
rect -11943 31943 -11920 31977
rect -12000 31920 -11920 31943
rect -11840 32937 -11760 32960
rect -11840 32903 -11817 32937
rect -11783 32903 -11760 32937
rect -11840 32617 -11760 32903
rect -11840 32583 -11817 32617
rect -11783 32583 -11760 32617
rect -11840 32297 -11760 32583
rect -11840 32263 -11817 32297
rect -11783 32263 -11760 32297
rect -11840 31977 -11760 32263
rect -11840 31943 -11817 31977
rect -11783 31943 -11760 31977
rect -11840 31920 -11760 31943
rect -11680 32937 -11600 32960
rect -11680 32903 -11657 32937
rect -11623 32903 -11600 32937
rect -11680 32617 -11600 32903
rect -11680 32583 -11657 32617
rect -11623 32583 -11600 32617
rect -11680 32297 -11600 32583
rect -11680 32263 -11657 32297
rect -11623 32263 -11600 32297
rect -11680 31977 -11600 32263
rect -11680 31943 -11657 31977
rect -11623 31943 -11600 31977
rect -11680 31920 -11600 31943
rect -11520 32937 -11440 32960
rect -11520 32903 -11497 32937
rect -11463 32903 -11440 32937
rect -11520 32617 -11440 32903
rect -11520 32583 -11497 32617
rect -11463 32583 -11440 32617
rect -11520 32297 -11440 32583
rect -11200 32937 -11120 32960
rect -11200 32903 -11177 32937
rect -11143 32903 -11120 32937
rect -11200 32617 -11120 32903
rect -11200 32583 -11177 32617
rect -11143 32583 -11120 32617
rect -11520 32263 -11497 32297
rect -11463 32263 -11440 32297
rect -11520 31977 -11440 32263
rect -11520 31943 -11497 31977
rect -11463 31943 -11440 31977
rect -11520 31920 -11440 31943
rect -11360 32297 -11280 32320
rect -11360 32263 -11337 32297
rect -11303 32263 -11280 32297
rect -11360 31977 -11280 32263
rect -11360 31943 -11337 31977
rect -11303 31943 -11280 31977
rect -11360 31920 -11280 31943
rect -11200 32297 -11120 32583
rect -11200 32263 -11177 32297
rect -11143 32263 -11120 32297
rect -11200 31977 -11120 32263
rect -11200 31943 -11177 31977
rect -11143 31943 -11120 31977
rect -11200 31920 -11120 31943
rect -10880 32937 -10800 32960
rect -10880 32903 -10857 32937
rect -10823 32903 -10800 32937
rect -10880 32617 -10800 32903
rect -10880 32583 -10857 32617
rect -10823 32583 -10800 32617
rect -10880 32297 -10800 32583
rect -10880 32263 -10857 32297
rect -10823 32263 -10800 32297
rect -10880 31977 -10800 32263
rect -10880 31943 -10857 31977
rect -10823 31943 -10800 31977
rect -10880 31920 -10800 31943
rect -10720 32937 -10640 32960
rect -10720 32903 -10697 32937
rect -10663 32903 -10640 32937
rect -10720 32617 -10640 32903
rect -10720 32583 -10697 32617
rect -10663 32583 -10640 32617
rect -10720 32297 -10640 32583
rect -10720 32263 -10697 32297
rect -10663 32263 -10640 32297
rect -10720 31977 -10640 32263
rect -10720 31943 -10697 31977
rect -10663 31943 -10640 31977
rect -10720 31920 -10640 31943
rect -10560 32937 -10480 32960
rect -10560 32903 -10537 32937
rect -10503 32903 -10480 32937
rect -10560 32617 -10480 32903
rect -10560 32583 -10537 32617
rect -10503 32583 -10480 32617
rect -10560 32297 -10480 32583
rect -10560 32263 -10537 32297
rect -10503 32263 -10480 32297
rect -10560 31977 -10480 32263
rect -10560 31943 -10537 31977
rect -10503 31943 -10480 31977
rect -10560 31920 -10480 31943
rect -10400 32937 -10320 32960
rect -10400 32903 -10377 32937
rect -10343 32903 -10320 32937
rect -10400 32617 -10320 32903
rect -10400 32583 -10377 32617
rect -10343 32583 -10320 32617
rect -10400 32297 -10320 32583
rect -10400 32263 -10377 32297
rect -10343 32263 -10320 32297
rect -10400 31977 -10320 32263
rect -10400 31943 -10377 31977
rect -10343 31943 -10320 31977
rect -10400 31920 -10320 31943
rect -10240 32937 -10160 32960
rect -10240 32903 -10217 32937
rect -10183 32903 -10160 32937
rect -10240 32617 -10160 32903
rect -10240 32583 -10217 32617
rect -10183 32583 -10160 32617
rect -10240 32297 -10160 32583
rect -10240 32263 -10217 32297
rect -10183 32263 -10160 32297
rect -10240 31977 -10160 32263
rect -10240 31943 -10217 31977
rect -10183 31943 -10160 31977
rect -10240 31920 -10160 31943
rect -10080 32937 -10000 32960
rect -10080 32903 -10057 32937
rect -10023 32903 -10000 32937
rect -10080 32617 -10000 32903
rect -10080 32583 -10057 32617
rect -10023 32583 -10000 32617
rect -10080 32297 -10000 32583
rect -10080 32263 -10057 32297
rect -10023 32263 -10000 32297
rect -10080 31977 -10000 32263
rect -10080 31943 -10057 31977
rect -10023 31943 -10000 31977
rect -10080 31920 -10000 31943
rect -9920 32937 -9840 32960
rect -9920 32903 -9897 32937
rect -9863 32903 -9840 32937
rect -9920 32617 -9840 32903
rect -9920 32583 -9897 32617
rect -9863 32583 -9840 32617
rect -9920 32297 -9840 32583
rect -9920 32263 -9897 32297
rect -9863 32263 -9840 32297
rect -9920 31977 -9840 32263
rect -9920 31943 -9897 31977
rect -9863 31943 -9840 31977
rect -9920 31920 -9840 31943
rect -9760 32937 -9680 32960
rect -9760 32903 -9737 32937
rect -9703 32903 -9680 32937
rect -9760 32617 -9680 32903
rect -9760 32583 -9737 32617
rect -9703 32583 -9680 32617
rect -9760 32297 -9680 32583
rect -9760 32263 -9737 32297
rect -9703 32263 -9680 32297
rect -9760 31977 -9680 32263
rect -9760 31943 -9737 31977
rect -9703 31943 -9680 31977
rect -9760 31920 -9680 31943
rect -9600 32937 -9520 32960
rect -9600 32903 -9577 32937
rect -9543 32903 -9520 32937
rect -9600 32617 -9520 32903
rect -9600 32583 -9577 32617
rect -9543 32583 -9520 32617
rect -9600 32297 -9520 32583
rect -9600 32263 -9577 32297
rect -9543 32263 -9520 32297
rect -9600 31977 -9520 32263
rect -9600 31943 -9577 31977
rect -9543 31943 -9520 31977
rect -9600 31920 -9520 31943
rect -9440 32937 -9360 32960
rect -9440 32903 -9417 32937
rect -9383 32903 -9360 32937
rect -9440 32617 -9360 32903
rect -9440 32583 -9417 32617
rect -9383 32583 -9360 32617
rect -9440 32297 -9360 32583
rect -9440 32263 -9417 32297
rect -9383 32263 -9360 32297
rect -9440 31977 -9360 32263
rect -9440 31943 -9417 31977
rect -9383 31943 -9360 31977
rect -9440 31920 -9360 31943
rect -9280 32937 -9200 32960
rect -9280 32903 -9257 32937
rect -9223 32903 -9200 32937
rect -9280 32617 -9200 32903
rect -9280 32583 -9257 32617
rect -9223 32583 -9200 32617
rect -9280 32297 -9200 32583
rect -9280 32263 -9257 32297
rect -9223 32263 -9200 32297
rect -9280 31977 -9200 32263
rect -9280 31943 -9257 31977
rect -9223 31943 -9200 31977
rect -9280 31920 -9200 31943
rect -9120 32937 -9040 32960
rect -9120 32903 -9097 32937
rect -9063 32903 -9040 32937
rect -9120 32617 -9040 32903
rect -9120 32583 -9097 32617
rect -9063 32583 -9040 32617
rect -9120 32297 -9040 32583
rect -9120 32263 -9097 32297
rect -9063 32263 -9040 32297
rect -9120 31977 -9040 32263
rect -9120 31943 -9097 31977
rect -9063 31943 -9040 31977
rect -9120 31920 -9040 31943
rect -8960 32937 -8880 32960
rect -8960 32903 -8937 32937
rect -8903 32903 -8880 32937
rect -8960 32617 -8880 32903
rect -8960 32583 -8937 32617
rect -8903 32583 -8880 32617
rect -8960 32297 -8880 32583
rect -8960 32263 -8937 32297
rect -8903 32263 -8880 32297
rect -8960 31977 -8880 32263
rect -8960 31943 -8937 31977
rect -8903 31943 -8880 31977
rect -8960 31920 -8880 31943
rect -8800 32937 -8720 32960
rect -8800 32903 -8777 32937
rect -8743 32903 -8720 32937
rect -8800 32617 -8720 32903
rect -8800 32583 -8777 32617
rect -8743 32583 -8720 32617
rect -8800 32297 -8720 32583
rect -8800 32263 -8777 32297
rect -8743 32263 -8720 32297
rect -8800 31977 -8720 32263
rect -8800 31943 -8777 31977
rect -8743 31943 -8720 31977
rect -8800 31920 -8720 31943
rect -8640 32937 -8560 32960
rect -8640 32903 -8617 32937
rect -8583 32903 -8560 32937
rect -8640 32617 -8560 32903
rect -8640 32583 -8617 32617
rect -8583 32583 -8560 32617
rect -8640 32297 -8560 32583
rect -8640 32263 -8617 32297
rect -8583 32263 -8560 32297
rect -8640 31977 -8560 32263
rect -8640 31943 -8617 31977
rect -8583 31943 -8560 31977
rect -8640 31920 -8560 31943
rect -8480 32937 -8400 32960
rect -8480 32903 -8457 32937
rect -8423 32903 -8400 32937
rect -8480 32617 -8400 32903
rect -8480 32583 -8457 32617
rect -8423 32583 -8400 32617
rect -8480 32297 -8400 32583
rect -8480 32263 -8457 32297
rect -8423 32263 -8400 32297
rect -8480 31977 -8400 32263
rect -8480 31943 -8457 31977
rect -8423 31943 -8400 31977
rect -8480 31920 -8400 31943
rect -8320 32937 -8240 32960
rect -8320 32903 -8297 32937
rect -8263 32903 -8240 32937
rect -8320 32617 -8240 32903
rect -8320 32583 -8297 32617
rect -8263 32583 -8240 32617
rect -8320 32297 -8240 32583
rect -8320 32263 -8297 32297
rect -8263 32263 -8240 32297
rect -8320 31977 -8240 32263
rect -8320 31943 -8297 31977
rect -8263 31943 -8240 31977
rect -8320 31920 -8240 31943
rect -8160 32937 -8080 32960
rect -8160 32903 -8137 32937
rect -8103 32903 -8080 32937
rect -8160 32617 -8080 32903
rect -8160 32583 -8137 32617
rect -8103 32583 -8080 32617
rect -8160 32297 -8080 32583
rect -8160 32263 -8137 32297
rect -8103 32263 -8080 32297
rect -8160 31977 -8080 32263
rect -8160 31943 -8137 31977
rect -8103 31943 -8080 31977
rect -8160 31920 -8080 31943
rect -8000 32937 -7920 32960
rect -8000 32903 -7977 32937
rect -7943 32903 -7920 32937
rect -8000 32617 -7920 32903
rect -8000 32583 -7977 32617
rect -7943 32583 -7920 32617
rect -8000 32297 -7920 32583
rect -8000 32263 -7977 32297
rect -7943 32263 -7920 32297
rect -8000 31977 -7920 32263
rect -8000 31943 -7977 31977
rect -7943 31943 -7920 31977
rect -8000 31920 -7920 31943
rect -7840 32937 -7760 32960
rect -7840 32903 -7817 32937
rect -7783 32903 -7760 32937
rect -7840 32617 -7760 32903
rect -7840 32583 -7817 32617
rect -7783 32583 -7760 32617
rect -7840 32297 -7760 32583
rect -7840 32263 -7817 32297
rect -7783 32263 -7760 32297
rect -7840 31977 -7760 32263
rect -7840 31943 -7817 31977
rect -7783 31943 -7760 31977
rect -7840 31920 -7760 31943
rect -7680 32937 -7600 32960
rect -7680 32903 -7657 32937
rect -7623 32903 -7600 32937
rect -7680 32617 -7600 32903
rect -7680 32583 -7657 32617
rect -7623 32583 -7600 32617
rect -7680 32297 -7600 32583
rect -7680 32263 -7657 32297
rect -7623 32263 -7600 32297
rect -7680 31977 -7600 32263
rect -7680 31943 -7657 31977
rect -7623 31943 -7600 31977
rect -7680 31920 -7600 31943
rect -7520 32937 -7440 32960
rect -7520 32903 -7497 32937
rect -7463 32903 -7440 32937
rect -7520 32617 -7440 32903
rect -7520 32583 -7497 32617
rect -7463 32583 -7440 32617
rect -7520 32297 -7440 32583
rect -7520 32263 -7497 32297
rect -7463 32263 -7440 32297
rect -7520 31977 -7440 32263
rect -7520 31943 -7497 31977
rect -7463 31943 -7440 31977
rect -7520 31920 -7440 31943
rect -7360 32937 -7280 32960
rect -7360 32903 -7337 32937
rect -7303 32903 -7280 32937
rect -7360 32617 -7280 32903
rect -7360 32583 -7337 32617
rect -7303 32583 -7280 32617
rect -7360 32297 -7280 32583
rect -7360 32263 -7337 32297
rect -7303 32263 -7280 32297
rect -7360 31977 -7280 32263
rect -7360 31943 -7337 31977
rect -7303 31943 -7280 31977
rect -7360 31920 -7280 31943
rect -7200 32937 -7120 32960
rect -7200 32903 -7177 32937
rect -7143 32903 -7120 32937
rect -7200 32617 -7120 32903
rect -7200 32583 -7177 32617
rect -7143 32583 -7120 32617
rect -7200 32297 -7120 32583
rect -7200 32263 -7177 32297
rect -7143 32263 -7120 32297
rect -7200 31977 -7120 32263
rect -7200 31943 -7177 31977
rect -7143 31943 -7120 31977
rect -7200 31920 -7120 31943
rect -7040 32937 -6960 32960
rect -7040 32903 -7017 32937
rect -6983 32903 -6960 32937
rect -7040 32617 -6960 32903
rect -7040 32583 -7017 32617
rect -6983 32583 -6960 32617
rect -7040 32297 -6960 32583
rect -7040 32263 -7017 32297
rect -6983 32263 -6960 32297
rect -7040 31977 -6960 32263
rect -7040 31943 -7017 31977
rect -6983 31943 -6960 31977
rect -7040 31920 -6960 31943
rect -6880 32937 -6800 32960
rect -6880 32903 -6857 32937
rect -6823 32903 -6800 32937
rect -6880 32617 -6800 32903
rect -6880 32583 -6857 32617
rect -6823 32583 -6800 32617
rect -6880 32297 -6800 32583
rect -6880 32263 -6857 32297
rect -6823 32263 -6800 32297
rect -6880 31977 -6800 32263
rect -6880 31943 -6857 31977
rect -6823 31943 -6800 31977
rect -6880 31920 -6800 31943
rect -6720 32937 -6640 32960
rect -6720 32903 -6697 32937
rect -6663 32903 -6640 32937
rect -6720 32617 -6640 32903
rect -6720 32583 -6697 32617
rect -6663 32583 -6640 32617
rect -6720 32297 -6640 32583
rect -6720 32263 -6697 32297
rect -6663 32263 -6640 32297
rect -6720 31977 -6640 32263
rect -6720 31943 -6697 31977
rect -6663 31943 -6640 31977
rect -6720 31920 -6640 31943
rect -6560 32937 -6480 32960
rect -6560 32903 -6537 32937
rect -6503 32903 -6480 32937
rect -6560 32617 -6480 32903
rect -6560 32583 -6537 32617
rect -6503 32583 -6480 32617
rect -6560 32297 -6480 32583
rect -6560 32263 -6537 32297
rect -6503 32263 -6480 32297
rect -6560 31977 -6480 32263
rect -6560 31943 -6537 31977
rect -6503 31943 -6480 31977
rect -6560 31920 -6480 31943
rect -6400 32937 -6320 32960
rect -6400 32903 -6377 32937
rect -6343 32903 -6320 32937
rect -6400 32617 -6320 32903
rect -6400 32583 -6377 32617
rect -6343 32583 -6320 32617
rect -6400 32297 -6320 32583
rect -6400 32263 -6377 32297
rect -6343 32263 -6320 32297
rect -6400 31977 -6320 32263
rect -6400 31943 -6377 31977
rect -6343 31943 -6320 31977
rect -6400 31920 -6320 31943
rect -6240 32937 -6160 32960
rect -6240 32903 -6217 32937
rect -6183 32903 -6160 32937
rect -6240 32617 -6160 32903
rect -6240 32583 -6217 32617
rect -6183 32583 -6160 32617
rect -6240 32297 -6160 32583
rect -6240 32263 -6217 32297
rect -6183 32263 -6160 32297
rect -6240 31977 -6160 32263
rect -6240 31943 -6217 31977
rect -6183 31943 -6160 31977
rect -6240 31920 -6160 31943
rect -6080 32937 -6000 32960
rect -6080 32903 -6057 32937
rect -6023 32903 -6000 32937
rect -6080 32617 -6000 32903
rect -6080 32583 -6057 32617
rect -6023 32583 -6000 32617
rect -6080 32297 -6000 32583
rect -6080 32263 -6057 32297
rect -6023 32263 -6000 32297
rect -6080 31977 -6000 32263
rect -6080 31943 -6057 31977
rect -6023 31943 -6000 31977
rect -6080 31920 -6000 31943
rect -5920 32937 -5840 32960
rect -5920 32903 -5897 32937
rect -5863 32903 -5840 32937
rect -5920 32617 -5840 32903
rect -5920 32583 -5897 32617
rect -5863 32583 -5840 32617
rect -5920 32297 -5840 32583
rect -5920 32263 -5897 32297
rect -5863 32263 -5840 32297
rect -5920 31977 -5840 32263
rect -5920 31943 -5897 31977
rect -5863 31943 -5840 31977
rect -5920 31920 -5840 31943
rect -5760 32937 -5680 32960
rect -5760 32903 -5737 32937
rect -5703 32903 -5680 32937
rect -5760 32617 -5680 32903
rect -5760 32583 -5737 32617
rect -5703 32583 -5680 32617
rect -5760 32297 -5680 32583
rect -5760 32263 -5737 32297
rect -5703 32263 -5680 32297
rect -5760 31977 -5680 32263
rect -5760 31943 -5737 31977
rect -5703 31943 -5680 31977
rect -5760 31920 -5680 31943
rect -5600 32937 -5520 32960
rect -5600 32903 -5577 32937
rect -5543 32903 -5520 32937
rect -5600 32617 -5520 32903
rect -5600 32583 -5577 32617
rect -5543 32583 -5520 32617
rect -5600 32297 -5520 32583
rect -5600 32263 -5577 32297
rect -5543 32263 -5520 32297
rect -5600 31977 -5520 32263
rect -5600 31943 -5577 31977
rect -5543 31943 -5520 31977
rect -5600 31920 -5520 31943
rect -5440 32937 -5360 32960
rect -5440 32903 -5417 32937
rect -5383 32903 -5360 32937
rect -5440 32617 -5360 32903
rect -5440 32583 -5417 32617
rect -5383 32583 -5360 32617
rect -5440 32297 -5360 32583
rect -5440 32263 -5417 32297
rect -5383 32263 -5360 32297
rect -5440 31977 -5360 32263
rect -5440 31943 -5417 31977
rect -5383 31943 -5360 31977
rect -5440 31920 -5360 31943
rect -5280 32937 -5200 32960
rect -5280 32903 -5257 32937
rect -5223 32903 -5200 32937
rect -5280 32617 -5200 32903
rect -5280 32583 -5257 32617
rect -5223 32583 -5200 32617
rect -5280 32297 -5200 32583
rect -5280 32263 -5257 32297
rect -5223 32263 -5200 32297
rect -5280 31977 -5200 32263
rect -5280 31943 -5257 31977
rect -5223 31943 -5200 31977
rect -5280 31920 -5200 31943
rect -5120 32937 -5040 32960
rect -5120 32903 -5097 32937
rect -5063 32903 -5040 32937
rect -5120 32617 -5040 32903
rect -5120 32583 -5097 32617
rect -5063 32583 -5040 32617
rect -5120 32297 -5040 32583
rect -5120 32263 -5097 32297
rect -5063 32263 -5040 32297
rect -5120 31977 -5040 32263
rect -5120 31943 -5097 31977
rect -5063 31943 -5040 31977
rect -5120 31920 -5040 31943
rect -4960 32937 -4880 32960
rect -4960 32903 -4937 32937
rect -4903 32903 -4880 32937
rect -4960 32617 -4880 32903
rect -4960 32583 -4937 32617
rect -4903 32583 -4880 32617
rect -4960 32297 -4880 32583
rect -4960 32263 -4937 32297
rect -4903 32263 -4880 32297
rect -4960 31977 -4880 32263
rect -4960 31943 -4937 31977
rect -4903 31943 -4880 31977
rect -4960 31920 -4880 31943
rect -4800 32937 -4720 32960
rect -4800 32903 -4777 32937
rect -4743 32903 -4720 32937
rect -4800 32617 -4720 32903
rect -4800 32583 -4777 32617
rect -4743 32583 -4720 32617
rect -4800 32297 -4720 32583
rect -4800 32263 -4777 32297
rect -4743 32263 -4720 32297
rect -4800 31977 -4720 32263
rect -4800 31943 -4777 31977
rect -4743 31943 -4720 31977
rect -4800 31920 -4720 31943
rect -4640 32937 -4560 32960
rect -4640 32903 -4617 32937
rect -4583 32903 -4560 32937
rect -4640 32617 -4560 32903
rect -4640 32583 -4617 32617
rect -4583 32583 -4560 32617
rect -4640 32297 -4560 32583
rect -4640 32263 -4617 32297
rect -4583 32263 -4560 32297
rect -4640 31977 -4560 32263
rect -4640 31943 -4617 31977
rect -4583 31943 -4560 31977
rect -4640 31920 -4560 31943
rect -4480 32937 -4400 32960
rect -4480 32903 -4457 32937
rect -4423 32903 -4400 32937
rect -4480 32617 -4400 32903
rect -4480 32583 -4457 32617
rect -4423 32583 -4400 32617
rect -4480 32297 -4400 32583
rect -4480 32263 -4457 32297
rect -4423 32263 -4400 32297
rect -4480 31977 -4400 32263
rect -4480 31943 -4457 31977
rect -4423 31943 -4400 31977
rect -4480 31920 -4400 31943
rect -4320 32937 -4240 32960
rect -4320 32903 -4297 32937
rect -4263 32903 -4240 32937
rect -4320 32617 -4240 32903
rect -4320 32583 -4297 32617
rect -4263 32583 -4240 32617
rect -4320 32297 -4240 32583
rect -4320 32263 -4297 32297
rect -4263 32263 -4240 32297
rect -4320 31977 -4240 32263
rect -4320 31943 -4297 31977
rect -4263 31943 -4240 31977
rect -4320 31920 -4240 31943
rect -4160 32937 -4080 32960
rect -4160 32903 -4137 32937
rect -4103 32903 -4080 32937
rect -4160 32617 -4080 32903
rect -4160 32583 -4137 32617
rect -4103 32583 -4080 32617
rect -4160 32297 -4080 32583
rect -4160 32263 -4137 32297
rect -4103 32263 -4080 32297
rect -4160 31977 -4080 32263
rect -4160 31943 -4137 31977
rect -4103 31943 -4080 31977
rect -4160 31920 -4080 31943
rect -4000 32937 -3920 32960
rect -4000 32903 -3977 32937
rect -3943 32903 -3920 32937
rect -4000 32617 -3920 32903
rect -4000 32583 -3977 32617
rect -3943 32583 -3920 32617
rect -4000 32297 -3920 32583
rect -4000 32263 -3977 32297
rect -3943 32263 -3920 32297
rect -4000 31977 -3920 32263
rect -4000 31943 -3977 31977
rect -3943 31943 -3920 31977
rect -4000 31920 -3920 31943
rect -3840 31840 -3760 34880
rect -3680 32937 -3600 32960
rect -3680 32903 -3657 32937
rect -3623 32903 -3600 32937
rect -3680 32617 -3600 32903
rect -3680 32583 -3657 32617
rect -3623 32583 -3600 32617
rect -3680 32297 -3600 32583
rect -3680 32263 -3657 32297
rect -3623 32263 -3600 32297
rect -3680 31977 -3600 32263
rect -3680 31943 -3657 31977
rect -3623 31943 -3600 31977
rect -3680 31920 -3600 31943
rect -3520 32937 -3440 32960
rect -3520 32903 -3497 32937
rect -3463 32903 -3440 32937
rect -3520 32617 -3440 32903
rect -3520 32583 -3497 32617
rect -3463 32583 -3440 32617
rect -3520 32297 -3440 32583
rect -3520 32263 -3497 32297
rect -3463 32263 -3440 32297
rect -3520 31977 -3440 32263
rect -3520 31943 -3497 31977
rect -3463 31943 -3440 31977
rect -3520 31920 -3440 31943
rect -3360 32937 -3280 32960
rect -3360 32903 -3337 32937
rect -3303 32903 -3280 32937
rect -3360 32617 -3280 32903
rect -3360 32583 -3337 32617
rect -3303 32583 -3280 32617
rect -3360 32297 -3280 32583
rect -3360 32263 -3337 32297
rect -3303 32263 -3280 32297
rect -3360 31977 -3280 32263
rect -3360 31943 -3337 31977
rect -3303 31943 -3280 31977
rect -3360 31920 -3280 31943
rect -3200 32937 -3120 32960
rect -3200 32903 -3177 32937
rect -3143 32903 -3120 32937
rect -3200 32617 -3120 32903
rect -3200 32583 -3177 32617
rect -3143 32583 -3120 32617
rect -3200 32297 -3120 32583
rect -3200 32263 -3177 32297
rect -3143 32263 -3120 32297
rect -3200 31977 -3120 32263
rect -3200 31943 -3177 31977
rect -3143 31943 -3120 31977
rect -3200 31920 -3120 31943
rect -3040 32937 -2960 32960
rect -3040 32903 -3017 32937
rect -2983 32903 -2960 32937
rect -3040 32617 -2960 32903
rect -3040 32583 -3017 32617
rect -2983 32583 -2960 32617
rect -3040 32297 -2960 32583
rect -3040 32263 -3017 32297
rect -2983 32263 -2960 32297
rect -3040 31977 -2960 32263
rect -3040 31943 -3017 31977
rect -2983 31943 -2960 31977
rect -3040 31920 -2960 31943
rect -2880 32937 -2800 32960
rect -2880 32903 -2857 32937
rect -2823 32903 -2800 32937
rect -2880 32617 -2800 32903
rect -2880 32583 -2857 32617
rect -2823 32583 -2800 32617
rect -2880 32297 -2800 32583
rect -2880 32263 -2857 32297
rect -2823 32263 -2800 32297
rect -2880 31977 -2800 32263
rect -2880 31943 -2857 31977
rect -2823 31943 -2800 31977
rect -2880 31920 -2800 31943
rect -2720 32937 -2640 32960
rect -2720 32903 -2697 32937
rect -2663 32903 -2640 32937
rect -2720 32617 -2640 32903
rect -2720 32583 -2697 32617
rect -2663 32583 -2640 32617
rect -2720 32297 -2640 32583
rect -2720 32263 -2697 32297
rect -2663 32263 -2640 32297
rect -2720 31977 -2640 32263
rect -2720 31943 -2697 31977
rect -2663 31943 -2640 31977
rect -2720 31920 -2640 31943
rect -2400 32937 -2320 32960
rect -2400 32903 -2377 32937
rect -2343 32903 -2320 32937
rect -2400 32617 -2320 32903
rect -2400 32583 -2377 32617
rect -2343 32583 -2320 32617
rect -2400 32297 -2320 32583
rect -2400 32263 -2377 32297
rect -2343 32263 -2320 32297
rect -2400 31977 -2320 32263
rect -2400 31943 -2377 31977
rect -2343 31943 -2320 31977
rect -2400 31920 -2320 31943
rect -2080 32937 -2000 32960
rect -2080 32903 -2057 32937
rect -2023 32903 -2000 32937
rect -2080 32617 -2000 32903
rect -2080 32583 -2057 32617
rect -2023 32583 -2000 32617
rect -2080 32297 -2000 32583
rect -2080 32263 -2057 32297
rect -2023 32263 -2000 32297
rect -2080 31977 -2000 32263
rect -2080 31943 -2057 31977
rect -2023 31943 -2000 31977
rect -2080 31920 -2000 31943
rect -1760 32937 -1680 32960
rect -1760 32903 -1737 32937
rect -1703 32903 -1680 32937
rect -1760 32617 -1680 32903
rect -1760 32583 -1737 32617
rect -1703 32583 -1680 32617
rect -1760 32297 -1680 32583
rect -1760 32263 -1737 32297
rect -1703 32263 -1680 32297
rect -1760 31977 -1680 32263
rect -1760 31943 -1737 31977
rect -1703 31943 -1680 31977
rect -1760 31920 -1680 31943
rect -1440 32937 -1360 32960
rect -1440 32903 -1417 32937
rect -1383 32903 -1360 32937
rect -1440 32617 -1360 32903
rect -1440 32583 -1417 32617
rect -1383 32583 -1360 32617
rect -1440 32297 -1360 32583
rect -1440 32263 -1417 32297
rect -1383 32263 -1360 32297
rect -1440 31977 -1360 32263
rect -1440 31943 -1417 31977
rect -1383 31943 -1360 31977
rect -1440 31920 -1360 31943
rect -1120 32937 -1040 32960
rect -1120 32903 -1097 32937
rect -1063 32903 -1040 32937
rect -1120 32617 -1040 32903
rect -1120 32583 -1097 32617
rect -1063 32583 -1040 32617
rect -1120 32297 -1040 32583
rect -1120 32263 -1097 32297
rect -1063 32263 -1040 32297
rect -1120 31977 -1040 32263
rect -1120 31943 -1097 31977
rect -1063 31943 -1040 31977
rect -1120 31920 -1040 31943
<< viali >>
rect -29897 42823 -29863 42857
rect -29897 42503 -29863 42537
rect -29897 42183 -29863 42217
rect -29897 41863 -29863 41897
rect -29737 42823 -29703 42857
rect -29737 42503 -29703 42537
rect -29737 42183 -29703 42217
rect -29737 41863 -29703 41897
rect -29577 42823 -29543 42857
rect -29577 42503 -29543 42537
rect -29577 42183 -29543 42217
rect -29577 41863 -29543 41897
rect -29417 42823 -29383 42857
rect -29417 42503 -29383 42537
rect -29417 42183 -29383 42217
rect -29417 41863 -29383 41897
rect -29257 42823 -29223 42857
rect -29257 42503 -29223 42537
rect -29257 42183 -29223 42217
rect -29257 41863 -29223 41897
rect -29097 42823 -29063 42857
rect -29097 42503 -29063 42537
rect -29097 42183 -29063 42217
rect -29097 41863 -29063 41897
rect -28937 42823 -28903 42857
rect -28937 42503 -28903 42537
rect -28937 42183 -28903 42217
rect -28937 41863 -28903 41897
rect -28777 42823 -28743 42857
rect -28777 42503 -28743 42537
rect -28777 42183 -28743 42217
rect -28777 41863 -28743 41897
rect -28617 42823 -28583 42857
rect -28617 42503 -28583 42537
rect -28617 42183 -28583 42217
rect -28617 41863 -28583 41897
rect -28457 42823 -28423 42857
rect -28457 42503 -28423 42537
rect -28457 42183 -28423 42217
rect -28457 41863 -28423 41897
rect -28297 42823 -28263 42857
rect -28297 42503 -28263 42537
rect -28297 42183 -28263 42217
rect -28297 41863 -28263 41897
rect -28137 42823 -28103 42857
rect -28137 42503 -28103 42537
rect -28137 42183 -28103 42217
rect -28137 41863 -28103 41897
rect -27977 42823 -27943 42857
rect -27977 42503 -27943 42537
rect -27977 42183 -27943 42217
rect -27977 41863 -27943 41897
rect -27817 42823 -27783 42857
rect -27817 42503 -27783 42537
rect -27817 42183 -27783 42217
rect -27817 41863 -27783 41897
rect -27657 42823 -27623 42857
rect -27657 42503 -27623 42537
rect -27657 42183 -27623 42217
rect -27657 41863 -27623 41897
rect -27497 42823 -27463 42857
rect -27497 42503 -27463 42537
rect -27497 42183 -27463 42217
rect -27497 41863 -27463 41897
rect -27337 42823 -27303 42857
rect -27337 42503 -27303 42537
rect -27337 42183 -27303 42217
rect -27337 41863 -27303 41897
rect -27177 42823 -27143 42857
rect -27177 42503 -27143 42537
rect -27177 42183 -27143 42217
rect -27177 41863 -27143 41897
rect -27017 42823 -26983 42857
rect -27017 42503 -26983 42537
rect -27017 42183 -26983 42217
rect -27017 41863 -26983 41897
rect -26857 42823 -26823 42857
rect -26857 42503 -26823 42537
rect -26857 42183 -26823 42217
rect -26857 41863 -26823 41897
rect -26697 42823 -26663 42857
rect -26697 42503 -26663 42537
rect -26697 42183 -26663 42217
rect -26697 41863 -26663 41897
rect -26537 42823 -26503 42857
rect -26537 42503 -26503 42537
rect -26537 42183 -26503 42217
rect -26537 41863 -26503 41897
rect -26377 42823 -26343 42857
rect -26377 42503 -26343 42537
rect -26377 42183 -26343 42217
rect -26377 41863 -26343 41897
rect -26217 42823 -26183 42857
rect -26217 42503 -26183 42537
rect -26217 42183 -26183 42217
rect -26217 41863 -26183 41897
rect -26057 42823 -26023 42857
rect -26057 42503 -26023 42537
rect -26057 42183 -26023 42217
rect -26057 41863 -26023 41897
rect -25897 42823 -25863 42857
rect -25897 42503 -25863 42537
rect -25897 42183 -25863 42217
rect -25897 41863 -25863 41897
rect -25737 42823 -25703 42857
rect -25737 42503 -25703 42537
rect -25737 42183 -25703 42217
rect -25737 41863 -25703 41897
rect -25577 42823 -25543 42857
rect -25577 42503 -25543 42537
rect -25577 42183 -25543 42217
rect -25577 41863 -25543 41897
rect -25417 42823 -25383 42857
rect -25417 42503 -25383 42537
rect -25417 42183 -25383 42217
rect -25417 41863 -25383 41897
rect -25257 42823 -25223 42857
rect -25257 42503 -25223 42537
rect -25257 42183 -25223 42217
rect -25257 41863 -25223 41897
rect -25097 42823 -25063 42857
rect -25097 42503 -25063 42537
rect -25097 42183 -25063 42217
rect -25097 41863 -25063 41897
rect -24937 42823 -24903 42857
rect -24937 42503 -24903 42537
rect -24937 42183 -24903 42217
rect -24937 41863 -24903 41897
rect -24777 42823 -24743 42857
rect -24777 42503 -24743 42537
rect -24777 42183 -24743 42217
rect -24777 41863 -24743 41897
rect -24617 42823 -24583 42857
rect -24617 42503 -24583 42537
rect -24617 42183 -24583 42217
rect -24617 41863 -24583 41897
rect -24457 42823 -24423 42857
rect -24457 42503 -24423 42537
rect -24457 42183 -24423 42217
rect -24457 41863 -24423 41897
rect -24297 42823 -24263 42857
rect -24297 42503 -24263 42537
rect -24297 42183 -24263 42217
rect -24297 41863 -24263 41897
rect -24137 42823 -24103 42857
rect -24137 42503 -24103 42537
rect -24137 42183 -24103 42217
rect -24137 41863 -24103 41897
rect -23977 42823 -23943 42857
rect -23977 42503 -23943 42537
rect -23977 42183 -23943 42217
rect -23977 41863 -23943 41897
rect -23817 42823 -23783 42857
rect -23817 42503 -23783 42537
rect -23817 42183 -23783 42217
rect -23817 41863 -23783 41897
rect -23657 42823 -23623 42857
rect -23657 42503 -23623 42537
rect -23657 42183 -23623 42217
rect -23657 41863 -23623 41897
rect -23497 42823 -23463 42857
rect -23497 42503 -23463 42537
rect -23497 42183 -23463 42217
rect -23497 41863 -23463 41897
rect -23337 42823 -23303 42857
rect -23337 42503 -23303 42537
rect -23337 42183 -23303 42217
rect -23337 41863 -23303 41897
rect -23177 42823 -23143 42857
rect -23177 42503 -23143 42537
rect -23177 42183 -23143 42217
rect -23177 41863 -23143 41897
rect -23017 42823 -22983 42857
rect -23017 42503 -22983 42537
rect -23017 42183 -22983 42217
rect -23017 41863 -22983 41897
rect -22857 42823 -22823 42857
rect -22857 42503 -22823 42537
rect -22857 42183 -22823 42217
rect -22857 41863 -22823 41897
rect -22697 42823 -22663 42857
rect -22697 42503 -22663 42537
rect -22697 42183 -22663 42217
rect -22697 41863 -22663 41897
rect -22537 42823 -22503 42857
rect -22537 42503 -22503 42537
rect -22537 42183 -22503 42217
rect -22537 41863 -22503 41897
rect -22377 42823 -22343 42857
rect -22377 42503 -22343 42537
rect -22377 42183 -22343 42217
rect -22377 41863 -22343 41897
rect -22217 42823 -22183 42857
rect -22217 42503 -22183 42537
rect -22217 42183 -22183 42217
rect -22217 41863 -22183 41897
rect -22057 42823 -22023 42857
rect -22057 42503 -22023 42537
rect -22057 42183 -22023 42217
rect -22057 41863 -22023 41897
rect -21897 42823 -21863 42857
rect -21897 42503 -21863 42537
rect -21897 42183 -21863 42217
rect -21897 41863 -21863 41897
rect -21737 42823 -21703 42857
rect -21737 42503 -21703 42537
rect -21737 42183 -21703 42217
rect -21737 41863 -21703 41897
rect -21577 42823 -21543 42857
rect -21577 42503 -21543 42537
rect -21577 42183 -21543 42217
rect -21577 41863 -21543 41897
rect -21417 42823 -21383 42857
rect -21417 42503 -21383 42537
rect -21417 42183 -21383 42217
rect -21417 41863 -21383 41897
rect -21257 42823 -21223 42857
rect -21257 42503 -21223 42537
rect -21257 42183 -21223 42217
rect -21257 41863 -21223 41897
rect -21097 42823 -21063 42857
rect -21097 42503 -21063 42537
rect -21097 42183 -21063 42217
rect -21097 41863 -21063 41897
rect -20937 42823 -20903 42857
rect -20937 42503 -20903 42537
rect -20937 42183 -20903 42217
rect -20937 41863 -20903 41897
rect -20777 42823 -20743 42857
rect -20777 42503 -20743 42537
rect -20777 42183 -20743 42217
rect -20777 41863 -20743 41897
rect -20617 42823 -20583 42857
rect -20617 42503 -20583 42537
rect -20617 42183 -20583 42217
rect -20617 41863 -20583 41897
rect -20457 42823 -20423 42857
rect -20457 42503 -20423 42537
rect -20457 42183 -20423 42217
rect -20457 41863 -20423 41897
rect -20297 42823 -20263 42857
rect -20297 42503 -20263 42537
rect -20297 42183 -20263 42217
rect -20297 41863 -20263 41897
rect -20137 42823 -20103 42857
rect -20137 42503 -20103 42537
rect -20137 42183 -20103 42217
rect -20137 41863 -20103 41897
rect -19977 42823 -19943 42857
rect -19977 42503 -19943 42537
rect -19977 42183 -19943 42217
rect -19977 41863 -19943 41897
rect -19817 42823 -19783 42857
rect -19817 42503 -19783 42537
rect -19817 42183 -19783 42217
rect -19817 41863 -19783 41897
rect -19657 42823 -19623 42857
rect -19657 42503 -19623 42537
rect -19657 42183 -19623 42217
rect -19657 41863 -19623 41897
rect -19497 42823 -19463 42857
rect -19497 42503 -19463 42537
rect -19497 42183 -19463 42217
rect -19497 41863 -19463 41897
rect -19337 42823 -19303 42857
rect -19337 42503 -19303 42537
rect -19337 42183 -19303 42217
rect -19337 41863 -19303 41897
rect -19177 42823 -19143 42857
rect -19177 42503 -19143 42537
rect -19177 42183 -19143 42217
rect -19177 41863 -19143 41897
rect -19017 42823 -18983 42857
rect -19017 42503 -18983 42537
rect -19017 42183 -18983 42217
rect -19017 41863 -18983 41897
rect -18857 42823 -18823 42857
rect -18857 42503 -18823 42537
rect -18857 42183 -18823 42217
rect -18857 41863 -18823 41897
rect -18697 42823 -18663 42857
rect -18697 42503 -18663 42537
rect -18697 42183 -18663 42217
rect -18697 41863 -18663 41897
rect -18537 42823 -18503 42857
rect -18537 42503 -18503 42537
rect -18537 42183 -18503 42217
rect -18537 41863 -18503 41897
rect -18377 42823 -18343 42857
rect -18377 42503 -18343 42537
rect -18377 42183 -18343 42217
rect -18377 41863 -18343 41897
rect -18217 42823 -18183 42857
rect -18217 42503 -18183 42537
rect -18217 42183 -18183 42217
rect -18217 41863 -18183 41897
rect -18057 42823 -18023 42857
rect -18057 42503 -18023 42537
rect -18057 42183 -18023 42217
rect -18057 41863 -18023 41897
rect -17897 42823 -17863 42857
rect -17897 42503 -17863 42537
rect -17897 42183 -17863 42217
rect -17897 41863 -17863 41897
rect -17737 42823 -17703 42857
rect -17737 42503 -17703 42537
rect -17737 42183 -17703 42217
rect -17737 41863 -17703 41897
rect -17577 42823 -17543 42857
rect -17577 42503 -17543 42537
rect -17577 42183 -17543 42217
rect -17577 41863 -17543 41897
rect -17417 42823 -17383 42857
rect -17417 42503 -17383 42537
rect -17417 42183 -17383 42217
rect -17417 41863 -17383 41897
rect -17257 42823 -17223 42857
rect -17257 42503 -17223 42537
rect -17257 42183 -17223 42217
rect -17257 41863 -17223 41897
rect -17097 42823 -17063 42857
rect -17097 42503 -17063 42537
rect -17097 42183 -17063 42217
rect -17097 41863 -17063 41897
rect -16937 42823 -16903 42857
rect -16937 42503 -16903 42537
rect -16937 42183 -16903 42217
rect -16937 41863 -16903 41897
rect -16777 42823 -16743 42857
rect -16777 42503 -16743 42537
rect -16777 42183 -16743 42217
rect -16777 41863 -16743 41897
rect -16617 42823 -16583 42857
rect -16617 42503 -16583 42537
rect -16617 42183 -16583 42217
rect -16617 41863 -16583 41897
rect -16457 42823 -16423 42857
rect -16457 42503 -16423 42537
rect -16457 42183 -16423 42217
rect -16457 41863 -16423 41897
rect -16297 42823 -16263 42857
rect -16297 42503 -16263 42537
rect -16297 42183 -16263 42217
rect -16297 41863 -16263 41897
rect -16137 42823 -16103 42857
rect -16137 42503 -16103 42537
rect -16137 42183 -16103 42217
rect -16137 41863 -16103 41897
rect -15977 42823 -15943 42857
rect -15977 42503 -15943 42537
rect -15977 42183 -15943 42217
rect -15977 41863 -15943 41897
rect -15817 42823 -15783 42857
rect -15817 42503 -15783 42537
rect -15817 42183 -15783 42217
rect -15817 41863 -15783 41897
rect -15657 42823 -15623 42857
rect -15657 42503 -15623 42537
rect -15657 42183 -15623 42217
rect -15657 41863 -15623 41897
rect -15497 42823 -15463 42857
rect -15497 42503 -15463 42537
rect -15497 42183 -15463 42217
rect -15497 41863 -15463 41897
rect -15337 42823 -15303 42857
rect -15337 42503 -15303 42537
rect -15337 42183 -15303 42217
rect -15337 41863 -15303 41897
rect -15177 42823 -15143 42857
rect -15177 42503 -15143 42537
rect -15177 42183 -15143 42217
rect -15177 41863 -15143 41897
rect -15017 42823 -14983 42857
rect -15017 42503 -14983 42537
rect -15017 42183 -14983 42217
rect -15017 41863 -14983 41897
rect -14857 42823 -14823 42857
rect -14857 42503 -14823 42537
rect -14857 42183 -14823 42217
rect -14857 41863 -14823 41897
rect -14697 42823 -14663 42857
rect -14697 42503 -14663 42537
rect -14697 42183 -14663 42217
rect -14697 41863 -14663 41897
rect -14537 42823 -14503 42857
rect -14537 42503 -14503 42537
rect -14537 42183 -14503 42217
rect -14537 41863 -14503 41897
rect -14377 42823 -14343 42857
rect -14377 42503 -14343 42537
rect -14377 42183 -14343 42217
rect -14377 41863 -14343 41897
rect -14217 42823 -14183 42857
rect -14217 42503 -14183 42537
rect -14217 42183 -14183 42217
rect -14217 41863 -14183 41897
rect -14057 42823 -14023 42857
rect -14057 42503 -14023 42537
rect -14057 42183 -14023 42217
rect -14057 41863 -14023 41897
rect -13897 42823 -13863 42857
rect -13897 42503 -13863 42537
rect -13897 42183 -13863 42217
rect -13897 41863 -13863 41897
rect -13737 42823 -13703 42857
rect -13737 42503 -13703 42537
rect -13737 42183 -13703 42217
rect -13737 41863 -13703 41897
rect -13577 42823 -13543 42857
rect -13577 42503 -13543 42537
rect -13577 42183 -13543 42217
rect -13577 41863 -13543 41897
rect -13417 42823 -13383 42857
rect -13417 42503 -13383 42537
rect -13417 42183 -13383 42217
rect -13417 41863 -13383 41897
rect -13257 42823 -13223 42857
rect -13257 42503 -13223 42537
rect -13257 42183 -13223 42217
rect -13257 41863 -13223 41897
rect -13097 42823 -13063 42857
rect -13097 42503 -13063 42537
rect -13097 42183 -13063 42217
rect -13097 41863 -13063 41897
rect -12937 42823 -12903 42857
rect -12937 42503 -12903 42537
rect -12937 42183 -12903 42217
rect -12937 41863 -12903 41897
rect -12777 42823 -12743 42857
rect -12777 42503 -12743 42537
rect -12777 42183 -12743 42217
rect -12777 41863 -12743 41897
rect -12617 42823 -12583 42857
rect -12617 42503 -12583 42537
rect -12617 42183 -12583 42217
rect -12617 41863 -12583 41897
rect -12457 42823 -12423 42857
rect -12457 42503 -12423 42537
rect -12457 42183 -12423 42217
rect -12457 41863 -12423 41897
rect -12297 42823 -12263 42857
rect -12297 42503 -12263 42537
rect -12297 42183 -12263 42217
rect -12297 41863 -12263 41897
rect -11337 42823 -11303 42857
rect -11337 42503 -11303 42537
rect -11337 42183 -11303 42217
rect -11337 41863 -11303 41897
rect -11177 42823 -11143 42857
rect -11177 42503 -11143 42537
rect -11177 42183 -11143 42217
rect -11177 41863 -11143 41897
rect -11017 42823 -10983 42857
rect -11017 42503 -10983 42537
rect -11017 42183 -10983 42217
rect -11017 41863 -10983 41897
rect -10857 42823 -10823 42857
rect -10857 42503 -10823 42537
rect -10857 42183 -10823 42217
rect -10857 41863 -10823 41897
rect -10697 42823 -10663 42857
rect -10697 42503 -10663 42537
rect -10697 42183 -10663 42217
rect -10697 41863 -10663 41897
rect -10537 42823 -10503 42857
rect -10537 42503 -10503 42537
rect -10537 42183 -10503 42217
rect -10537 41863 -10503 41897
rect -10377 42823 -10343 42857
rect -10377 42503 -10343 42537
rect -10377 42183 -10343 42217
rect -10377 41863 -10343 41897
rect -10217 42823 -10183 42857
rect -10217 42503 -10183 42537
rect -10217 42183 -10183 42217
rect -10217 41863 -10183 41897
rect -10057 42823 -10023 42857
rect -10057 42503 -10023 42537
rect -10057 42183 -10023 42217
rect -10057 41863 -10023 41897
rect -9897 42823 -9863 42857
rect -9897 42503 -9863 42537
rect -9897 42183 -9863 42217
rect -9897 41863 -9863 41897
rect -9737 42823 -9703 42857
rect -9737 42503 -9703 42537
rect -9737 42183 -9703 42217
rect -9737 41863 -9703 41897
rect -9577 42823 -9543 42857
rect -9577 42503 -9543 42537
rect -9577 42183 -9543 42217
rect -9577 41863 -9543 41897
rect -9417 42823 -9383 42857
rect -9417 42503 -9383 42537
rect -9417 42183 -9383 42217
rect -9417 41863 -9383 41897
rect -9257 42823 -9223 42857
rect -9257 42503 -9223 42537
rect -9257 42183 -9223 42217
rect -9257 41863 -9223 41897
rect -9097 42823 -9063 42857
rect -9097 42503 -9063 42537
rect -9097 42183 -9063 42217
rect -9097 41863 -9063 41897
rect -8937 42823 -8903 42857
rect -8937 42503 -8903 42537
rect -8937 42183 -8903 42217
rect -8937 41863 -8903 41897
rect -8777 42823 -8743 42857
rect -8777 42503 -8743 42537
rect -8777 42183 -8743 42217
rect -8777 41863 -8743 41897
rect -8617 42823 -8583 42857
rect -8617 42503 -8583 42537
rect -8617 42183 -8583 42217
rect -8617 41863 -8583 41897
rect -8457 42823 -8423 42857
rect -8457 42503 -8423 42537
rect -8457 42183 -8423 42217
rect -8457 41863 -8423 41897
rect -8297 42823 -8263 42857
rect -8297 42503 -8263 42537
rect -8297 42183 -8263 42217
rect -8297 41863 -8263 41897
rect -8137 42823 -8103 42857
rect -8137 42503 -8103 42537
rect -8137 42183 -8103 42217
rect -8137 41863 -8103 41897
rect -7977 42823 -7943 42857
rect -7977 42503 -7943 42537
rect -7977 42183 -7943 42217
rect -7977 41863 -7943 41897
rect -7817 42823 -7783 42857
rect -7817 42503 -7783 42537
rect -7817 42183 -7783 42217
rect -7817 41863 -7783 41897
rect -7657 42823 -7623 42857
rect -7657 42503 -7623 42537
rect -7657 42183 -7623 42217
rect -7657 41863 -7623 41897
rect -7497 42823 -7463 42857
rect -7497 42503 -7463 42537
rect -7497 42183 -7463 42217
rect -7497 41863 -7463 41897
rect -7337 42823 -7303 42857
rect -7337 42503 -7303 42537
rect -7337 42183 -7303 42217
rect -7337 41863 -7303 41897
rect -7177 42823 -7143 42857
rect -7177 42503 -7143 42537
rect -7177 42183 -7143 42217
rect -7177 41863 -7143 41897
rect -7017 42823 -6983 42857
rect -7017 42503 -6983 42537
rect -7017 42183 -6983 42217
rect -7017 41863 -6983 41897
rect -6857 42823 -6823 42857
rect -6857 42503 -6823 42537
rect -6857 42183 -6823 42217
rect -6857 41863 -6823 41897
rect -6697 42823 -6663 42857
rect -6697 42503 -6663 42537
rect -6697 42183 -6663 42217
rect -6697 41863 -6663 41897
rect -6537 42823 -6503 42857
rect -6537 42503 -6503 42537
rect -6537 42183 -6503 42217
rect -6537 41863 -6503 41897
rect -6377 42823 -6343 42857
rect -6377 42503 -6343 42537
rect -6377 42183 -6343 42217
rect -6377 41863 -6343 41897
rect -6217 42823 -6183 42857
rect -6217 42503 -6183 42537
rect -6217 42183 -6183 42217
rect -6217 41863 -6183 41897
rect -6057 42823 -6023 42857
rect -6057 42503 -6023 42537
rect -6057 42183 -6023 42217
rect -6057 41863 -6023 41897
rect -5897 42823 -5863 42857
rect -5897 42503 -5863 42537
rect -5897 42183 -5863 42217
rect -5897 41863 -5863 41897
rect -5737 42823 -5703 42857
rect -5737 42503 -5703 42537
rect -5737 42183 -5703 42217
rect -5737 41863 -5703 41897
rect -5577 42823 -5543 42857
rect -5577 42503 -5543 42537
rect -5577 42183 -5543 42217
rect -5577 41863 -5543 41897
rect -5417 42823 -5383 42857
rect -5417 42503 -5383 42537
rect -5417 42183 -5383 42217
rect -5417 41863 -5383 41897
rect -5257 42823 -5223 42857
rect -5257 42503 -5223 42537
rect -5257 42183 -5223 42217
rect -5257 41863 -5223 41897
rect -5097 42823 -5063 42857
rect -5097 42503 -5063 42537
rect -5097 42183 -5063 42217
rect -5097 41863 -5063 41897
rect -4937 42823 -4903 42857
rect -4937 42503 -4903 42537
rect -4937 42183 -4903 42217
rect -4937 41863 -4903 41897
rect -4777 42823 -4743 42857
rect -4777 42503 -4743 42537
rect -4777 42183 -4743 42217
rect -4777 41863 -4743 41897
rect -4617 42823 -4583 42857
rect -4617 42503 -4583 42537
rect -4617 42183 -4583 42217
rect -4617 41863 -4583 41897
rect -4457 42823 -4423 42857
rect -4457 42503 -4423 42537
rect -4457 42183 -4423 42217
rect -4457 41863 -4423 41897
rect -4297 42823 -4263 42857
rect -4297 42503 -4263 42537
rect -4297 42183 -4263 42217
rect -4297 41863 -4263 41897
rect -4137 42823 -4103 42857
rect -4137 42503 -4103 42537
rect -4137 42183 -4103 42217
rect -4137 41863 -4103 41897
rect -3977 42823 -3943 42857
rect -3977 42503 -3943 42537
rect -3977 42183 -3943 42217
rect -3977 41863 -3943 41897
rect -33097 41303 -33063 41337
rect -33097 40983 -33063 41017
rect -32937 41303 -32903 41337
rect -32937 40983 -32903 41017
rect -32777 41303 -32743 41337
rect -32777 40983 -32743 41017
rect -32617 41303 -32583 41337
rect -32617 40983 -32583 41017
rect -32457 41303 -32423 41337
rect -32457 40983 -32423 41017
rect -32297 41303 -32263 41337
rect -32297 40983 -32263 41017
rect -32137 41303 -32103 41337
rect -32137 40983 -32103 41017
rect -31977 41303 -31943 41337
rect -31977 40983 -31943 41017
rect -31817 41303 -31783 41337
rect -31817 40983 -31783 41017
rect -31657 41303 -31623 41337
rect -31657 40983 -31623 41017
rect -31497 41303 -31463 41337
rect -31497 40983 -31463 41017
rect -31337 41303 -31303 41337
rect -31337 40983 -31303 41017
rect -31177 41303 -31143 41337
rect -31177 40983 -31143 41017
rect -29897 41303 -29863 41337
rect -29897 40983 -29863 41017
rect -29737 41303 -29703 41337
rect -29737 40983 -29703 41017
rect -29577 41303 -29543 41337
rect -29577 40983 -29543 41017
rect -29417 41303 -29383 41337
rect -29417 40983 -29383 41017
rect -29257 41303 -29223 41337
rect -29257 40983 -29223 41017
rect -29097 41303 -29063 41337
rect -29097 40983 -29063 41017
rect -28937 41303 -28903 41337
rect -28937 40983 -28903 41017
rect -28777 41303 -28743 41337
rect -28777 40983 -28743 41017
rect -28617 41303 -28583 41337
rect -28617 40983 -28583 41017
rect -28457 41303 -28423 41337
rect -28457 40983 -28423 41017
rect -28297 41303 -28263 41337
rect -28297 40983 -28263 41017
rect -28137 41303 -28103 41337
rect -28137 40983 -28103 41017
rect -27977 41303 -27943 41337
rect -27977 40983 -27943 41017
rect -27817 41303 -27783 41337
rect -27817 40983 -27783 41017
rect -27657 41303 -27623 41337
rect -27657 40983 -27623 41017
rect -27497 41303 -27463 41337
rect -27497 40983 -27463 41017
rect -27337 41303 -27303 41337
rect -27337 40983 -27303 41017
rect -27177 41303 -27143 41337
rect -27177 40983 -27143 41017
rect -27017 41303 -26983 41337
rect -27017 40983 -26983 41017
rect -26857 41303 -26823 41337
rect -26857 40983 -26823 41017
rect -26697 41303 -26663 41337
rect -26697 40983 -26663 41017
rect -26537 41303 -26503 41337
rect -26537 40983 -26503 41017
rect -26377 41303 -26343 41337
rect -26377 40983 -26343 41017
rect -26217 41303 -26183 41337
rect -26217 40983 -26183 41017
rect -26057 41303 -26023 41337
rect -26057 40983 -26023 41017
rect -25897 41303 -25863 41337
rect -25897 40983 -25863 41017
rect -25737 41303 -25703 41337
rect -25737 40983 -25703 41017
rect -25577 41303 -25543 41337
rect -25577 40983 -25543 41017
rect -25417 41303 -25383 41337
rect -25417 40983 -25383 41017
rect -25257 41303 -25223 41337
rect -25257 40983 -25223 41017
rect -25097 41303 -25063 41337
rect -25097 40983 -25063 41017
rect -24937 41303 -24903 41337
rect -24937 40983 -24903 41017
rect -24777 41303 -24743 41337
rect -24777 40983 -24743 41017
rect -24617 41303 -24583 41337
rect -24617 40983 -24583 41017
rect -24457 41303 -24423 41337
rect -24457 40983 -24423 41017
rect -24297 41303 -24263 41337
rect -24297 40983 -24263 41017
rect -24137 41303 -24103 41337
rect -24137 40983 -24103 41017
rect -23977 41303 -23943 41337
rect -23977 40983 -23943 41017
rect -23817 41303 -23783 41337
rect -23817 40983 -23783 41017
rect -23657 41303 -23623 41337
rect -23657 40983 -23623 41017
rect -23497 41303 -23463 41337
rect -23497 40983 -23463 41017
rect -23337 41303 -23303 41337
rect -23337 40983 -23303 41017
rect -23177 41303 -23143 41337
rect -23177 40983 -23143 41017
rect -23017 41303 -22983 41337
rect -23017 40983 -22983 41017
rect -22857 41303 -22823 41337
rect -22857 40983 -22823 41017
rect -22697 41303 -22663 41337
rect -22697 40983 -22663 41017
rect -22537 41303 -22503 41337
rect -22537 40983 -22503 41017
rect -22377 41303 -22343 41337
rect -22377 40983 -22343 41017
rect -22217 41303 -22183 41337
rect -22217 40983 -22183 41017
rect -22057 41303 -22023 41337
rect -22057 40983 -22023 41017
rect -21897 41303 -21863 41337
rect -21897 40983 -21863 41017
rect -21737 41303 -21703 41337
rect -21737 40983 -21703 41017
rect -21577 41303 -21543 41337
rect -21577 40983 -21543 41017
rect -21417 41303 -21383 41337
rect -21417 40983 -21383 41017
rect -21257 41303 -21223 41337
rect -21257 40983 -21223 41017
rect -21097 41303 -21063 41337
rect -21097 40983 -21063 41017
rect -20937 41303 -20903 41337
rect -20937 40983 -20903 41017
rect -20777 41303 -20743 41337
rect -20777 40983 -20743 41017
rect -20617 41303 -20583 41337
rect -20617 40983 -20583 41017
rect -20457 41303 -20423 41337
rect -20457 40983 -20423 41017
rect -20297 41303 -20263 41337
rect -20297 40983 -20263 41017
rect -20137 41303 -20103 41337
rect -20137 40983 -20103 41017
rect -19977 41303 -19943 41337
rect -19977 40983 -19943 41017
rect -19817 41303 -19783 41337
rect -19817 40983 -19783 41017
rect -19657 41303 -19623 41337
rect -19657 40983 -19623 41017
rect -19497 41303 -19463 41337
rect -19497 40983 -19463 41017
rect -19337 41303 -19303 41337
rect -19337 40983 -19303 41017
rect -19177 41303 -19143 41337
rect -19177 40983 -19143 41017
rect -19017 41303 -18983 41337
rect -19017 40983 -18983 41017
rect -18857 41303 -18823 41337
rect -18857 40983 -18823 41017
rect -18697 41303 -18663 41337
rect -18697 40983 -18663 41017
rect -18537 41303 -18503 41337
rect -18537 40983 -18503 41017
rect -18377 41303 -18343 41337
rect -18377 40983 -18343 41017
rect -18217 41303 -18183 41337
rect -18217 40983 -18183 41017
rect -18057 41303 -18023 41337
rect -18057 40983 -18023 41017
rect -17897 41303 -17863 41337
rect -17897 40983 -17863 41017
rect -17737 41303 -17703 41337
rect -17737 40983 -17703 41017
rect -17577 41303 -17543 41337
rect -17577 40983 -17543 41017
rect -17417 41303 -17383 41337
rect -17417 40983 -17383 41017
rect -17257 41303 -17223 41337
rect -17257 40983 -17223 41017
rect -17097 41303 -17063 41337
rect -17097 40983 -17063 41017
rect -16937 41303 -16903 41337
rect -16937 40983 -16903 41017
rect -16777 41303 -16743 41337
rect -16777 40983 -16743 41017
rect -16617 41303 -16583 41337
rect -16617 40983 -16583 41017
rect -16457 41303 -16423 41337
rect -16457 40983 -16423 41017
rect -16297 41303 -16263 41337
rect -16297 40983 -16263 41017
rect -16137 41303 -16103 41337
rect -16137 40983 -16103 41017
rect -15977 41303 -15943 41337
rect -15977 40983 -15943 41017
rect -15817 41303 -15783 41337
rect -15817 40983 -15783 41017
rect -15657 41303 -15623 41337
rect -15657 40983 -15623 41017
rect -15497 41303 -15463 41337
rect -15497 40983 -15463 41017
rect -15337 41303 -15303 41337
rect -15337 40983 -15303 41017
rect -15177 41303 -15143 41337
rect -15177 40983 -15143 41017
rect -15017 41303 -14983 41337
rect -15017 40983 -14983 41017
rect -14857 41303 -14823 41337
rect -14857 40983 -14823 41017
rect -14697 41303 -14663 41337
rect -14697 40983 -14663 41017
rect -14537 41303 -14503 41337
rect -14537 40983 -14503 41017
rect -14377 41303 -14343 41337
rect -14377 40983 -14343 41017
rect -14217 41303 -14183 41337
rect -14217 40983 -14183 41017
rect -14057 41303 -14023 41337
rect -14057 40983 -14023 41017
rect -13897 41303 -13863 41337
rect -13897 40983 -13863 41017
rect -13737 41303 -13703 41337
rect -13737 40983 -13703 41017
rect -13577 41303 -13543 41337
rect -13577 40983 -13543 41017
rect -13417 41303 -13383 41337
rect -13417 40983 -13383 41017
rect -13257 41303 -13223 41337
rect -13257 40983 -13223 41017
rect -13097 41303 -13063 41337
rect -13097 40983 -13063 41017
rect -12937 41303 -12903 41337
rect -12937 40983 -12903 41017
rect -12777 41303 -12743 41337
rect -12777 40983 -12743 41017
rect -12617 41303 -12583 41337
rect -12617 40983 -12583 41017
rect -12457 41303 -12423 41337
rect -12457 40983 -12423 41017
rect -12297 41303 -12263 41337
rect -12297 40983 -12263 41017
rect -11337 41303 -11303 41337
rect -11337 40983 -11303 41017
rect -11177 41303 -11143 41337
rect -11177 40983 -11143 41017
rect -11017 41303 -10983 41337
rect -11017 40983 -10983 41017
rect -10857 41303 -10823 41337
rect -10857 40983 -10823 41017
rect -10697 41303 -10663 41337
rect -10697 40983 -10663 41017
rect -10537 41303 -10503 41337
rect -10537 40983 -10503 41017
rect -10377 41303 -10343 41337
rect -10377 40983 -10343 41017
rect -10217 41303 -10183 41337
rect -10217 40983 -10183 41017
rect -10057 41303 -10023 41337
rect -10057 40983 -10023 41017
rect -9897 41303 -9863 41337
rect -9897 40983 -9863 41017
rect -9737 41303 -9703 41337
rect -9737 40983 -9703 41017
rect -9577 41303 -9543 41337
rect -9577 40983 -9543 41017
rect -9417 41303 -9383 41337
rect -9417 40983 -9383 41017
rect -9257 41303 -9223 41337
rect -9257 40983 -9223 41017
rect -9097 41303 -9063 41337
rect -9097 40983 -9063 41017
rect -8937 41303 -8903 41337
rect -8937 40983 -8903 41017
rect -8777 41303 -8743 41337
rect -8777 40983 -8743 41017
rect -8617 41303 -8583 41337
rect -8617 40983 -8583 41017
rect -8457 41303 -8423 41337
rect -8457 40983 -8423 41017
rect -8297 41303 -8263 41337
rect -8297 40983 -8263 41017
rect -8137 41303 -8103 41337
rect -8137 40983 -8103 41017
rect -7977 41303 -7943 41337
rect -7977 40983 -7943 41017
rect -7817 41303 -7783 41337
rect -7817 40983 -7783 41017
rect -7657 41303 -7623 41337
rect -7657 40983 -7623 41017
rect -7497 41303 -7463 41337
rect -7497 40983 -7463 41017
rect -7337 41303 -7303 41337
rect -7337 40983 -7303 41017
rect -7177 41303 -7143 41337
rect -7177 40983 -7143 41017
rect -7017 41303 -6983 41337
rect -7017 40983 -6983 41017
rect -6857 41303 -6823 41337
rect -6857 40983 -6823 41017
rect -6697 41303 -6663 41337
rect -6697 40983 -6663 41017
rect -6537 41303 -6503 41337
rect -6537 40983 -6503 41017
rect -6377 41303 -6343 41337
rect -6377 40983 -6343 41017
rect -6217 41303 -6183 41337
rect -6217 40983 -6183 41017
rect -6057 41303 -6023 41337
rect -6057 40983 -6023 41017
rect -5897 41303 -5863 41337
rect -5897 40983 -5863 41017
rect -5737 41303 -5703 41337
rect -5737 40983 -5703 41017
rect -5577 41303 -5543 41337
rect -5577 40983 -5543 41017
rect -5417 41303 -5383 41337
rect -5417 40983 -5383 41017
rect -5257 41303 -5223 41337
rect -5257 40983 -5223 41017
rect -5097 41303 -5063 41337
rect -5097 40983 -5063 41017
rect -4937 41303 -4903 41337
rect -4937 40983 -4903 41017
rect -4777 41303 -4743 41337
rect -4777 40983 -4743 41017
rect -4617 41303 -4583 41337
rect -4617 40983 -4583 41017
rect -4457 41303 -4423 41337
rect -4457 40983 -4423 41017
rect -4297 41303 -4263 41337
rect -4297 40983 -4263 41017
rect -4137 41303 -4103 41337
rect -4137 40983 -4103 41017
rect -3977 41303 -3943 41337
rect -3977 40983 -3943 41017
rect -3657 42823 -3623 42857
rect -3657 42503 -3623 42537
rect -3657 42183 -3623 42217
rect -3657 41863 -3623 41897
rect -3497 42823 -3463 42857
rect -3497 42503 -3463 42537
rect -3497 42183 -3463 42217
rect -3497 41863 -3463 41897
rect -3337 42823 -3303 42857
rect -3337 42503 -3303 42537
rect -3337 42183 -3303 42217
rect -3337 41863 -3303 41897
rect -3017 42823 -2983 42857
rect -3017 42503 -2983 42537
rect -3017 42183 -2983 42217
rect -3017 41863 -2983 41897
rect -2697 42823 -2663 42857
rect -2697 42503 -2663 42537
rect -2697 42183 -2663 42217
rect -2697 41863 -2663 41897
rect -2537 42823 -2503 42857
rect -2537 42503 -2503 42537
rect -2537 42183 -2503 42217
rect -2537 41863 -2503 41897
rect -2377 42823 -2343 42857
rect -2377 42503 -2343 42537
rect -2377 42183 -2343 42217
rect -2377 41863 -2343 41897
rect -2217 42823 -2183 42857
rect -2217 42503 -2183 42537
rect -2217 42183 -2183 42217
rect -2217 41863 -2183 41897
rect -2057 42823 -2023 42857
rect -2057 42503 -2023 42537
rect -2057 42183 -2023 42217
rect -2057 41863 -2023 41897
rect -1737 42823 -1703 42857
rect -1737 42503 -1703 42537
rect -1737 42183 -1703 42217
rect -1737 41863 -1703 41897
rect -1417 42823 -1383 42857
rect -1417 42503 -1383 42537
rect -1417 42183 -1383 42217
rect -1417 41863 -1383 41897
rect -1097 42823 -1063 42857
rect -1097 42503 -1063 42537
rect -1097 42183 -1063 42217
rect -1097 41863 -1063 41897
rect -3817 41303 -3783 41337
rect -3817 40983 -3783 41017
rect -10537 40663 -10503 40697
rect -10537 40343 -10503 40377
rect -10217 40663 -10183 40697
rect -10217 40343 -10183 40377
rect -10057 40663 -10023 40697
rect -10057 40343 -10023 40377
rect -9897 40663 -9863 40697
rect -9897 40343 -9863 40377
rect -9737 40663 -9703 40697
rect -9737 40343 -9703 40377
rect -9577 40663 -9543 40697
rect -9577 40343 -9543 40377
rect -9417 40663 -9383 40697
rect -9417 40343 -9383 40377
rect -9257 40663 -9223 40697
rect -9257 40343 -9223 40377
rect -9097 40663 -9063 40697
rect -9097 40343 -9063 40377
rect -8937 40663 -8903 40697
rect -8937 40343 -8903 40377
rect -8777 40663 -8743 40697
rect -8777 40343 -8743 40377
rect -8617 40663 -8583 40697
rect -8617 40343 -8583 40377
rect -8457 40663 -8423 40697
rect -8457 40343 -8423 40377
rect -8297 40663 -8263 40697
rect -8297 40343 -8263 40377
rect -8137 40663 -8103 40697
rect -8137 40343 -8103 40377
rect -7977 40663 -7943 40697
rect -7977 40343 -7943 40377
rect -7817 40663 -7783 40697
rect -7817 40343 -7783 40377
rect -7657 40663 -7623 40697
rect -7657 40343 -7623 40377
rect -7497 40663 -7463 40697
rect -7497 40343 -7463 40377
rect -7337 40663 -7303 40697
rect -7337 40343 -7303 40377
rect -7177 40663 -7143 40697
rect -7177 40343 -7143 40377
rect -7017 40663 -6983 40697
rect -7017 40343 -6983 40377
rect -6857 40663 -6823 40697
rect -6857 40343 -6823 40377
rect -6697 40663 -6663 40697
rect -6697 40343 -6663 40377
rect -6537 40663 -6503 40697
rect -6537 40343 -6503 40377
rect -6377 40663 -6343 40697
rect -6377 40343 -6343 40377
rect -6217 40663 -6183 40697
rect -6217 40343 -6183 40377
rect -6057 40663 -6023 40697
rect -6057 40343 -6023 40377
rect -5897 40663 -5863 40697
rect -5897 40343 -5863 40377
rect -5737 40663 -5703 40697
rect -5737 40343 -5703 40377
rect -5577 40663 -5543 40697
rect -5577 40343 -5543 40377
rect -5417 40663 -5383 40697
rect -5417 40343 -5383 40377
rect -5257 40663 -5223 40697
rect -5257 40343 -5223 40377
rect -5097 40663 -5063 40697
rect -5097 40343 -5063 40377
rect -4937 40663 -4903 40697
rect -4937 40343 -4903 40377
rect -4777 40663 -4743 40697
rect -4777 40343 -4743 40377
rect -4617 40663 -4583 40697
rect -4617 40343 -4583 40377
rect -4457 40663 -4423 40697
rect -4457 40343 -4423 40377
rect -4297 40663 -4263 40697
rect -4297 40343 -4263 40377
rect -4137 40663 -4103 40697
rect -4137 40343 -4103 40377
rect -3977 40663 -3943 40697
rect -3977 40343 -3943 40377
rect -3657 41303 -3623 41337
rect -3657 40983 -3623 41017
rect -3497 41303 -3463 41337
rect -3497 40983 -3463 41017
rect 41063 41303 41097 41337
rect 41063 40983 41097 41017
rect 41223 41303 41257 41337
rect 41223 40983 41257 41017
rect 41383 41303 41417 41337
rect 41383 40983 41417 41017
rect 41543 41303 41577 41337
rect 41543 40983 41577 41017
rect 41703 41303 41737 41337
rect 41703 40983 41737 41017
rect 41863 41303 41897 41337
rect 41863 40983 41897 41017
rect 42023 41303 42057 41337
rect 42023 40983 42057 41017
rect 42183 41303 42217 41337
rect 42183 40983 42217 41017
rect 42343 41303 42377 41337
rect 42343 40983 42377 41017
rect 42503 41303 42537 41337
rect 42503 40983 42537 41017
rect 42663 41303 42697 41337
rect 42663 40983 42697 41017
rect 42823 41303 42857 41337
rect 42823 40983 42857 41017
rect 42983 41303 43017 41337
rect 42983 40983 43017 41017
rect 43143 41303 43177 41337
rect 43143 40983 43177 41017
rect -3657 40663 -3623 40697
rect -3657 40343 -3623 40377
rect -3497 40663 -3463 40697
rect -3497 40343 -3463 40377
rect 41063 40023 41097 40057
rect 41063 39703 41097 39737
rect 41223 40023 41257 40057
rect 41223 39703 41257 39737
rect 41383 40023 41417 40057
rect 41383 39703 41417 39737
rect 41543 40023 41577 40057
rect 41543 39703 41577 39737
rect 41703 40023 41737 40057
rect 41703 39703 41737 39737
rect 41863 40023 41897 40057
rect 41863 39703 41897 39737
rect 42023 40023 42057 40057
rect 42023 39703 42057 39737
rect 42183 40023 42217 40057
rect 42183 39703 42217 39737
rect 42343 40023 42377 40057
rect 42343 39703 42377 39737
rect 42503 40023 42537 40057
rect 42503 39703 42537 39737
rect 42663 40023 42697 40057
rect 42663 39703 42697 39737
rect 42823 40023 42857 40057
rect 42823 39703 42857 39737
rect 42983 40023 43017 40057
rect 42983 39703 43017 39737
rect 43143 40023 43177 40057
rect 43143 39703 43177 39737
rect -33097 37703 -33063 37737
rect -33097 37383 -33063 37417
rect -33097 37063 -33063 37097
rect -32937 37703 -32903 37737
rect -32937 37383 -32903 37417
rect -32937 37063 -32903 37097
rect -32777 37703 -32743 37737
rect -32777 37383 -32743 37417
rect -32777 37063 -32743 37097
rect -32617 37703 -32583 37737
rect -32617 37383 -32583 37417
rect -32617 37063 -32583 37097
rect -32457 37703 -32423 37737
rect -32457 37383 -32423 37417
rect -32457 37063 -32423 37097
rect -32297 37703 -32263 37737
rect -32297 37383 -32263 37417
rect -32297 37063 -32263 37097
rect -32137 37703 -32103 37737
rect -32137 37383 -32103 37417
rect -32137 37063 -32103 37097
rect -31977 37703 -31943 37737
rect -31977 37383 -31943 37417
rect -31977 37063 -31943 37097
rect -31817 37703 -31783 37737
rect -31817 37383 -31783 37417
rect -31817 37063 -31783 37097
rect -31657 37703 -31623 37737
rect -31657 37383 -31623 37417
rect -31657 37063 -31623 37097
rect -31497 37703 -31463 37737
rect -31497 37383 -31463 37417
rect -31497 37063 -31463 37097
rect -31337 37703 -31303 37737
rect -31337 37383 -31303 37417
rect -31337 37063 -31303 37097
rect -31177 37703 -31143 37737
rect -31177 37383 -31143 37417
rect -31177 37063 -31143 37097
rect 41063 36023 41097 36057
rect 41063 35703 41097 35737
rect 41223 36023 41257 36057
rect 41223 35703 41257 35737
rect 41383 36023 41417 36057
rect 41383 35703 41417 35737
rect 41543 36023 41577 36057
rect 41543 35703 41577 35737
rect 41703 36023 41737 36057
rect 41703 35703 41737 35737
rect 41863 36023 41897 36057
rect 41863 35703 41897 35737
rect 42023 36023 42057 36057
rect 42023 35703 42057 35737
rect 42183 36023 42217 36057
rect 42183 35703 42217 35737
rect 42343 36023 42377 36057
rect 42343 35703 42377 35737
rect 42503 36023 42537 36057
rect 42503 35703 42537 35737
rect 42663 36023 42697 36057
rect 42663 35703 42697 35737
rect 42823 36023 42857 36057
rect 42823 35703 42857 35737
rect 42983 36023 43017 36057
rect 42983 35703 43017 35737
rect 43143 36023 43177 36057
rect 43143 35703 43177 35737
rect -33097 34663 -33063 34697
rect -33097 34343 -33063 34377
rect -32937 34663 -32903 34697
rect -32937 34343 -32903 34377
rect -32777 34663 -32743 34697
rect -32777 34343 -32743 34377
rect -32617 34663 -32583 34697
rect -32617 34343 -32583 34377
rect -32457 34663 -32423 34697
rect -32457 34343 -32423 34377
rect -32297 34663 -32263 34697
rect -32297 34343 -32263 34377
rect -32137 34663 -32103 34697
rect -32137 34343 -32103 34377
rect -31977 34663 -31943 34697
rect -31977 34343 -31943 34377
rect -31817 34663 -31783 34697
rect -31817 34343 -31783 34377
rect -31657 34663 -31623 34697
rect -31657 34343 -31623 34377
rect -31497 34663 -31463 34697
rect -31497 34343 -31463 34377
rect -31337 34663 -31303 34697
rect -31337 34343 -31303 34377
rect -31177 34663 -31143 34697
rect -31177 34343 -31143 34377
rect -29897 34663 -29863 34697
rect -29897 34343 -29863 34377
rect -29737 34663 -29703 34697
rect -29737 34343 -29703 34377
rect -29577 34663 -29543 34697
rect -29577 34343 -29543 34377
rect -29417 34663 -29383 34697
rect -29417 34343 -29383 34377
rect -29257 34663 -29223 34697
rect -29257 34343 -29223 34377
rect -29097 34663 -29063 34697
rect -29097 34343 -29063 34377
rect -28937 34663 -28903 34697
rect -28937 34343 -28903 34377
rect -28777 34663 -28743 34697
rect -28777 34343 -28743 34377
rect -28617 34663 -28583 34697
rect -28617 34343 -28583 34377
rect -28457 34663 -28423 34697
rect -28457 34343 -28423 34377
rect -28297 34663 -28263 34697
rect -28297 34343 -28263 34377
rect -28137 34663 -28103 34697
rect -28137 34343 -28103 34377
rect -27977 34663 -27943 34697
rect -27977 34343 -27943 34377
rect -27817 34663 -27783 34697
rect -27817 34343 -27783 34377
rect -27657 34663 -27623 34697
rect -27657 34343 -27623 34377
rect -27497 34663 -27463 34697
rect -27497 34343 -27463 34377
rect -27337 34663 -27303 34697
rect -27337 34343 -27303 34377
rect -27177 34663 -27143 34697
rect -27177 34343 -27143 34377
rect -27017 34663 -26983 34697
rect -27017 34343 -26983 34377
rect -26857 34663 -26823 34697
rect -26857 34343 -26823 34377
rect -26697 34663 -26663 34697
rect -26697 34343 -26663 34377
rect -26537 34663 -26503 34697
rect -26537 34343 -26503 34377
rect -26377 34663 -26343 34697
rect -26377 34343 -26343 34377
rect -26217 34663 -26183 34697
rect -26217 34343 -26183 34377
rect -26057 34663 -26023 34697
rect -26057 34343 -26023 34377
rect -25897 34663 -25863 34697
rect -25897 34343 -25863 34377
rect -25737 34663 -25703 34697
rect -25737 34343 -25703 34377
rect -25577 34663 -25543 34697
rect -25577 34343 -25543 34377
rect -25417 34663 -25383 34697
rect -25417 34343 -25383 34377
rect -25257 34663 -25223 34697
rect -25257 34343 -25223 34377
rect -25097 34663 -25063 34697
rect -25097 34343 -25063 34377
rect -24937 34663 -24903 34697
rect -24937 34343 -24903 34377
rect -24777 34663 -24743 34697
rect -24777 34343 -24743 34377
rect -24617 34663 -24583 34697
rect -24617 34343 -24583 34377
rect -24457 34663 -24423 34697
rect -24457 34343 -24423 34377
rect -24297 34663 -24263 34697
rect -24297 34343 -24263 34377
rect -24137 34663 -24103 34697
rect -24137 34343 -24103 34377
rect -23977 34663 -23943 34697
rect -23977 34343 -23943 34377
rect -23817 34663 -23783 34697
rect -23817 34343 -23783 34377
rect -23657 34663 -23623 34697
rect -23657 34343 -23623 34377
rect -23497 34663 -23463 34697
rect -23497 34343 -23463 34377
rect -23337 34663 -23303 34697
rect -23337 34343 -23303 34377
rect -23177 34663 -23143 34697
rect -23177 34343 -23143 34377
rect -23017 34663 -22983 34697
rect -23017 34343 -22983 34377
rect -22857 34663 -22823 34697
rect -22857 34343 -22823 34377
rect -22697 34663 -22663 34697
rect -22697 34343 -22663 34377
rect -22537 34663 -22503 34697
rect -22537 34343 -22503 34377
rect -22377 34663 -22343 34697
rect -22377 34343 -22343 34377
rect -22217 34663 -22183 34697
rect -22217 34343 -22183 34377
rect -22057 34663 -22023 34697
rect -22057 34343 -22023 34377
rect -21897 34663 -21863 34697
rect -21897 34343 -21863 34377
rect -21737 34663 -21703 34697
rect -21737 34343 -21703 34377
rect -21577 34663 -21543 34697
rect -21577 34343 -21543 34377
rect -21417 34663 -21383 34697
rect -21417 34343 -21383 34377
rect -21257 34663 -21223 34697
rect -21257 34343 -21223 34377
rect -21097 34663 -21063 34697
rect -21097 34343 -21063 34377
rect -20937 34663 -20903 34697
rect -20937 34343 -20903 34377
rect -20777 34663 -20743 34697
rect -20777 34343 -20743 34377
rect -20617 34663 -20583 34697
rect -20617 34343 -20583 34377
rect -20457 34663 -20423 34697
rect -20457 34343 -20423 34377
rect -20297 34663 -20263 34697
rect -20297 34343 -20263 34377
rect -20137 34663 -20103 34697
rect -20137 34343 -20103 34377
rect -19977 34663 -19943 34697
rect -19977 34343 -19943 34377
rect -19817 34663 -19783 34697
rect -19817 34343 -19783 34377
rect -19657 34663 -19623 34697
rect -19657 34343 -19623 34377
rect -19497 34663 -19463 34697
rect -19497 34343 -19463 34377
rect -19337 34663 -19303 34697
rect -19337 34343 -19303 34377
rect -19177 34663 -19143 34697
rect -19177 34343 -19143 34377
rect -19017 34663 -18983 34697
rect -19017 34343 -18983 34377
rect -18857 34663 -18823 34697
rect -18857 34343 -18823 34377
rect -18697 34663 -18663 34697
rect -18697 34343 -18663 34377
rect -18537 34663 -18503 34697
rect -18537 34343 -18503 34377
rect -18377 34663 -18343 34697
rect -18377 34343 -18343 34377
rect -18217 34663 -18183 34697
rect -18217 34343 -18183 34377
rect -18057 34663 -18023 34697
rect -18057 34343 -18023 34377
rect -17897 34663 -17863 34697
rect -17897 34343 -17863 34377
rect -17737 34663 -17703 34697
rect -17737 34343 -17703 34377
rect -17577 34663 -17543 34697
rect -17577 34343 -17543 34377
rect -17417 34663 -17383 34697
rect -17417 34343 -17383 34377
rect -17257 34663 -17223 34697
rect -17257 34343 -17223 34377
rect -17097 34663 -17063 34697
rect -17097 34343 -17063 34377
rect -16937 34663 -16903 34697
rect -16937 34343 -16903 34377
rect -16777 34663 -16743 34697
rect -16777 34343 -16743 34377
rect -16617 34663 -16583 34697
rect -16617 34343 -16583 34377
rect -16457 34663 -16423 34697
rect -16457 34343 -16423 34377
rect -16297 34663 -16263 34697
rect -16297 34343 -16263 34377
rect -16137 34663 -16103 34697
rect -16137 34343 -16103 34377
rect -15977 34663 -15943 34697
rect -15977 34343 -15943 34377
rect -15817 34663 -15783 34697
rect -15817 34343 -15783 34377
rect -15657 34663 -15623 34697
rect -15657 34343 -15623 34377
rect -15497 34663 -15463 34697
rect -15497 34343 -15463 34377
rect -15337 34663 -15303 34697
rect -15337 34343 -15303 34377
rect -15177 34663 -15143 34697
rect -15177 34343 -15143 34377
rect -15017 34663 -14983 34697
rect -15017 34343 -14983 34377
rect -14857 34663 -14823 34697
rect -14857 34343 -14823 34377
rect -14697 34663 -14663 34697
rect -14697 34343 -14663 34377
rect -14537 34663 -14503 34697
rect -14537 34343 -14503 34377
rect -14377 34663 -14343 34697
rect -14377 34343 -14343 34377
rect -14217 34663 -14183 34697
rect -14217 34343 -14183 34377
rect -14057 34663 -14023 34697
rect -14057 34343 -14023 34377
rect -13897 34663 -13863 34697
rect -13897 34343 -13863 34377
rect -13737 34663 -13703 34697
rect -13737 34343 -13703 34377
rect -13577 34663 -13543 34697
rect -13577 34343 -13543 34377
rect -13417 34663 -13383 34697
rect -13417 34343 -13383 34377
rect -13257 34663 -13223 34697
rect -13257 34343 -13223 34377
rect -13097 34663 -13063 34697
rect -13097 34343 -13063 34377
rect -12937 34663 -12903 34697
rect -12937 34343 -12903 34377
rect -12777 34663 -12743 34697
rect -12777 34343 -12743 34377
rect -12617 34663 -12583 34697
rect -12617 34343 -12583 34377
rect -12457 34663 -12423 34697
rect -12457 34343 -12423 34377
rect -12297 34663 -12263 34697
rect -12297 34343 -12263 34377
rect -12137 34663 -12103 34697
rect -12137 34343 -12103 34377
rect -11977 34663 -11943 34697
rect -11977 34343 -11943 34377
rect -11817 34663 -11783 34697
rect -11817 34343 -11783 34377
rect -11657 34663 -11623 34697
rect -11657 34343 -11623 34377
rect -11497 34663 -11463 34697
rect -11497 34343 -11463 34377
rect -10857 34663 -10823 34697
rect -10857 34343 -10823 34377
rect -10537 34663 -10503 34697
rect -10537 34343 -10503 34377
rect -29897 32903 -29863 32937
rect -29897 32583 -29863 32617
rect -29897 32263 -29863 32297
rect -29897 31943 -29863 31977
rect -29737 32903 -29703 32937
rect -29737 32583 -29703 32617
rect -29737 32263 -29703 32297
rect -29737 31943 -29703 31977
rect -29577 32903 -29543 32937
rect -29577 32583 -29543 32617
rect -29577 32263 -29543 32297
rect -29577 31943 -29543 31977
rect -29417 32903 -29383 32937
rect -29417 32583 -29383 32617
rect -29417 32263 -29383 32297
rect -29417 31943 -29383 31977
rect -29257 32903 -29223 32937
rect -29257 32583 -29223 32617
rect -29257 32263 -29223 32297
rect -29257 31943 -29223 31977
rect -29097 32903 -29063 32937
rect -29097 32583 -29063 32617
rect -29097 32263 -29063 32297
rect -29097 31943 -29063 31977
rect -28937 32903 -28903 32937
rect -28937 32583 -28903 32617
rect -28937 32263 -28903 32297
rect -28937 31943 -28903 31977
rect -28777 32903 -28743 32937
rect -28777 32583 -28743 32617
rect -28777 32263 -28743 32297
rect -28777 31943 -28743 31977
rect -28617 32903 -28583 32937
rect -28617 32583 -28583 32617
rect -28617 32263 -28583 32297
rect -28617 31943 -28583 31977
rect -28457 32903 -28423 32937
rect -28457 32583 -28423 32617
rect -28457 32263 -28423 32297
rect -28457 31943 -28423 31977
rect -28297 32903 -28263 32937
rect -28297 32583 -28263 32617
rect -28297 32263 -28263 32297
rect -28297 31943 -28263 31977
rect -28137 32903 -28103 32937
rect -28137 32583 -28103 32617
rect -28137 32263 -28103 32297
rect -28137 31943 -28103 31977
rect -27977 32903 -27943 32937
rect -27977 32583 -27943 32617
rect -27977 32263 -27943 32297
rect -27977 31943 -27943 31977
rect -27817 32903 -27783 32937
rect -27817 32583 -27783 32617
rect -27817 32263 -27783 32297
rect -27817 31943 -27783 31977
rect -27657 32903 -27623 32937
rect -27657 32583 -27623 32617
rect -27657 32263 -27623 32297
rect -27657 31943 -27623 31977
rect -27497 32903 -27463 32937
rect -27497 32583 -27463 32617
rect -27497 32263 -27463 32297
rect -27497 31943 -27463 31977
rect -27337 32903 -27303 32937
rect -27337 32583 -27303 32617
rect -27337 32263 -27303 32297
rect -27337 31943 -27303 31977
rect -27177 32903 -27143 32937
rect -27177 32583 -27143 32617
rect -27177 32263 -27143 32297
rect -27177 31943 -27143 31977
rect -27017 32903 -26983 32937
rect -27017 32583 -26983 32617
rect -27017 32263 -26983 32297
rect -27017 31943 -26983 31977
rect -26857 32903 -26823 32937
rect -26857 32583 -26823 32617
rect -26857 32263 -26823 32297
rect -26857 31943 -26823 31977
rect -26697 32903 -26663 32937
rect -26697 32583 -26663 32617
rect -26697 32263 -26663 32297
rect -26697 31943 -26663 31977
rect -26537 32903 -26503 32937
rect -26537 32583 -26503 32617
rect -26537 32263 -26503 32297
rect -26537 31943 -26503 31977
rect -26377 32903 -26343 32937
rect -26377 32583 -26343 32617
rect -26377 32263 -26343 32297
rect -26377 31943 -26343 31977
rect -26217 32903 -26183 32937
rect -26217 32583 -26183 32617
rect -26217 32263 -26183 32297
rect -26217 31943 -26183 31977
rect -26057 32903 -26023 32937
rect -26057 32583 -26023 32617
rect -26057 32263 -26023 32297
rect -26057 31943 -26023 31977
rect -25897 32903 -25863 32937
rect -25897 32583 -25863 32617
rect -25897 32263 -25863 32297
rect -25897 31943 -25863 31977
rect -25737 32903 -25703 32937
rect -25737 32583 -25703 32617
rect -25737 32263 -25703 32297
rect -25737 31943 -25703 31977
rect -25577 32903 -25543 32937
rect -25577 32583 -25543 32617
rect -25577 32263 -25543 32297
rect -25577 31943 -25543 31977
rect -25417 32903 -25383 32937
rect -25417 32583 -25383 32617
rect -25417 32263 -25383 32297
rect -25417 31943 -25383 31977
rect -25257 32903 -25223 32937
rect -25257 32583 -25223 32617
rect -25257 32263 -25223 32297
rect -25257 31943 -25223 31977
rect -25097 32903 -25063 32937
rect -25097 32583 -25063 32617
rect -25097 32263 -25063 32297
rect -25097 31943 -25063 31977
rect -24937 32903 -24903 32937
rect -24937 32583 -24903 32617
rect -24937 32263 -24903 32297
rect -24937 31943 -24903 31977
rect -24777 32903 -24743 32937
rect -24777 32583 -24743 32617
rect -24777 32263 -24743 32297
rect -24777 31943 -24743 31977
rect -24617 32903 -24583 32937
rect -24617 32583 -24583 32617
rect -24617 32263 -24583 32297
rect -24617 31943 -24583 31977
rect -24457 32903 -24423 32937
rect -24457 32583 -24423 32617
rect -24457 32263 -24423 32297
rect -24457 31943 -24423 31977
rect -24297 32903 -24263 32937
rect -24297 32583 -24263 32617
rect -24297 32263 -24263 32297
rect -24297 31943 -24263 31977
rect -24137 32903 -24103 32937
rect -24137 32583 -24103 32617
rect -24137 32263 -24103 32297
rect -24137 31943 -24103 31977
rect -23977 32903 -23943 32937
rect -23977 32583 -23943 32617
rect -23977 32263 -23943 32297
rect -23977 31943 -23943 31977
rect -23817 32903 -23783 32937
rect -23817 32583 -23783 32617
rect -23817 32263 -23783 32297
rect -23817 31943 -23783 31977
rect -23657 32903 -23623 32937
rect -23657 32583 -23623 32617
rect -23657 32263 -23623 32297
rect -23657 31943 -23623 31977
rect -23497 32903 -23463 32937
rect -23497 32583 -23463 32617
rect -23497 32263 -23463 32297
rect -23497 31943 -23463 31977
rect -23337 32903 -23303 32937
rect -23337 32583 -23303 32617
rect -23337 32263 -23303 32297
rect -23337 31943 -23303 31977
rect -23177 32903 -23143 32937
rect -23177 32583 -23143 32617
rect -23177 32263 -23143 32297
rect -23177 31943 -23143 31977
rect -23017 32903 -22983 32937
rect -23017 32583 -22983 32617
rect -23017 32263 -22983 32297
rect -23017 31943 -22983 31977
rect -22857 32903 -22823 32937
rect -22857 32583 -22823 32617
rect -22857 32263 -22823 32297
rect -22857 31943 -22823 31977
rect -22697 32903 -22663 32937
rect -22697 32583 -22663 32617
rect -22697 32263 -22663 32297
rect -22697 31943 -22663 31977
rect -22537 32903 -22503 32937
rect -22537 32583 -22503 32617
rect -22537 32263 -22503 32297
rect -22537 31943 -22503 31977
rect -22377 32903 -22343 32937
rect -22377 32583 -22343 32617
rect -22377 32263 -22343 32297
rect -22377 31943 -22343 31977
rect -22217 32903 -22183 32937
rect -22217 32583 -22183 32617
rect -22217 32263 -22183 32297
rect -22217 31943 -22183 31977
rect -22057 32903 -22023 32937
rect -22057 32583 -22023 32617
rect -22057 32263 -22023 32297
rect -22057 31943 -22023 31977
rect -21897 32903 -21863 32937
rect -21897 32583 -21863 32617
rect -21897 32263 -21863 32297
rect -21897 31943 -21863 31977
rect -21737 32903 -21703 32937
rect -21737 32583 -21703 32617
rect -21737 32263 -21703 32297
rect -21737 31943 -21703 31977
rect -21577 32903 -21543 32937
rect -21577 32583 -21543 32617
rect -21577 32263 -21543 32297
rect -21577 31943 -21543 31977
rect -21417 32903 -21383 32937
rect -21417 32583 -21383 32617
rect -21417 32263 -21383 32297
rect -21417 31943 -21383 31977
rect -21257 32903 -21223 32937
rect -21257 32583 -21223 32617
rect -21257 32263 -21223 32297
rect -21257 31943 -21223 31977
rect -21097 32903 -21063 32937
rect -21097 32583 -21063 32617
rect -21097 32263 -21063 32297
rect -21097 31943 -21063 31977
rect -20937 32903 -20903 32937
rect -20937 32583 -20903 32617
rect -20937 32263 -20903 32297
rect -20937 31943 -20903 31977
rect -20777 32903 -20743 32937
rect -20777 32583 -20743 32617
rect -20777 32263 -20743 32297
rect -20777 31943 -20743 31977
rect -20617 32903 -20583 32937
rect -20617 32583 -20583 32617
rect -20617 32263 -20583 32297
rect -20617 31943 -20583 31977
rect -20457 32903 -20423 32937
rect -20457 32583 -20423 32617
rect -20457 32263 -20423 32297
rect -20457 31943 -20423 31977
rect -20297 32903 -20263 32937
rect -20297 32583 -20263 32617
rect -20297 32263 -20263 32297
rect -20297 31943 -20263 31977
rect -20137 32903 -20103 32937
rect -20137 32583 -20103 32617
rect -20137 32263 -20103 32297
rect -20137 31943 -20103 31977
rect -19977 32903 -19943 32937
rect -19977 32583 -19943 32617
rect -19977 32263 -19943 32297
rect -19977 31943 -19943 31977
rect -19817 32903 -19783 32937
rect -19817 32583 -19783 32617
rect -19817 32263 -19783 32297
rect -19817 31943 -19783 31977
rect -19657 32903 -19623 32937
rect -19657 32583 -19623 32617
rect -19657 32263 -19623 32297
rect -19657 31943 -19623 31977
rect -19497 32903 -19463 32937
rect -19497 32583 -19463 32617
rect -19497 32263 -19463 32297
rect -19497 31943 -19463 31977
rect -19337 32903 -19303 32937
rect -19337 32583 -19303 32617
rect -19337 32263 -19303 32297
rect -19337 31943 -19303 31977
rect -19177 32903 -19143 32937
rect -19177 32583 -19143 32617
rect -19177 32263 -19143 32297
rect -19177 31943 -19143 31977
rect -19017 32903 -18983 32937
rect -19017 32583 -18983 32617
rect -19017 32263 -18983 32297
rect -19017 31943 -18983 31977
rect -18857 32903 -18823 32937
rect -18857 32583 -18823 32617
rect -18857 32263 -18823 32297
rect -18857 31943 -18823 31977
rect -18697 32903 -18663 32937
rect -18697 32583 -18663 32617
rect -18697 32263 -18663 32297
rect -18697 31943 -18663 31977
rect -18537 32903 -18503 32937
rect -18537 32583 -18503 32617
rect -18537 32263 -18503 32297
rect -18537 31943 -18503 31977
rect -18377 32903 -18343 32937
rect -18377 32583 -18343 32617
rect -18377 32263 -18343 32297
rect -18377 31943 -18343 31977
rect -18217 32903 -18183 32937
rect -18217 32583 -18183 32617
rect -18217 32263 -18183 32297
rect -18217 31943 -18183 31977
rect -18057 32903 -18023 32937
rect -18057 32583 -18023 32617
rect -18057 32263 -18023 32297
rect -18057 31943 -18023 31977
rect -17897 32903 -17863 32937
rect -17897 32583 -17863 32617
rect -17897 32263 -17863 32297
rect -17897 31943 -17863 31977
rect -17737 32903 -17703 32937
rect -17737 32583 -17703 32617
rect -17737 32263 -17703 32297
rect -17737 31943 -17703 31977
rect -17577 32903 -17543 32937
rect -17577 32583 -17543 32617
rect -17577 32263 -17543 32297
rect -17577 31943 -17543 31977
rect -17417 32903 -17383 32937
rect -17417 32583 -17383 32617
rect -17417 32263 -17383 32297
rect -17417 31943 -17383 31977
rect -17257 32903 -17223 32937
rect -17257 32583 -17223 32617
rect -17257 32263 -17223 32297
rect -17257 31943 -17223 31977
rect -17097 32903 -17063 32937
rect -17097 32583 -17063 32617
rect -17097 32263 -17063 32297
rect -17097 31943 -17063 31977
rect -16937 32903 -16903 32937
rect -16937 32583 -16903 32617
rect -16937 32263 -16903 32297
rect -16937 31943 -16903 31977
rect -16777 32903 -16743 32937
rect -16777 32583 -16743 32617
rect -16777 32263 -16743 32297
rect -16777 31943 -16743 31977
rect -16617 32903 -16583 32937
rect -16617 32583 -16583 32617
rect -16617 32263 -16583 32297
rect -16617 31943 -16583 31977
rect -16457 32903 -16423 32937
rect -16457 32583 -16423 32617
rect -16457 32263 -16423 32297
rect -16457 31943 -16423 31977
rect -16297 32903 -16263 32937
rect -16297 32583 -16263 32617
rect -16297 32263 -16263 32297
rect -16297 31943 -16263 31977
rect -16137 32903 -16103 32937
rect -16137 32583 -16103 32617
rect -16137 32263 -16103 32297
rect -16137 31943 -16103 31977
rect -15977 32903 -15943 32937
rect -15977 32583 -15943 32617
rect -15977 32263 -15943 32297
rect -15977 31943 -15943 31977
rect -15817 32903 -15783 32937
rect -15817 32583 -15783 32617
rect -15817 32263 -15783 32297
rect -15817 31943 -15783 31977
rect -15657 32903 -15623 32937
rect -15657 32583 -15623 32617
rect -15657 32263 -15623 32297
rect -15657 31943 -15623 31977
rect -15497 32903 -15463 32937
rect -15497 32583 -15463 32617
rect -15497 32263 -15463 32297
rect -15497 31943 -15463 31977
rect -15337 32903 -15303 32937
rect -15337 32583 -15303 32617
rect -15337 32263 -15303 32297
rect -15337 31943 -15303 31977
rect -15177 32903 -15143 32937
rect -15177 32583 -15143 32617
rect -15177 32263 -15143 32297
rect -15177 31943 -15143 31977
rect -15017 32903 -14983 32937
rect -15017 32583 -14983 32617
rect -15017 32263 -14983 32297
rect -15017 31943 -14983 31977
rect -14857 32903 -14823 32937
rect -14857 32583 -14823 32617
rect -14857 32263 -14823 32297
rect -14857 31943 -14823 31977
rect -14697 32903 -14663 32937
rect -14697 32583 -14663 32617
rect -14697 32263 -14663 32297
rect -14697 31943 -14663 31977
rect -14537 32903 -14503 32937
rect -14537 32583 -14503 32617
rect -14537 32263 -14503 32297
rect -14537 31943 -14503 31977
rect -14377 32903 -14343 32937
rect -14377 32583 -14343 32617
rect -14377 32263 -14343 32297
rect -14377 31943 -14343 31977
rect -14217 32903 -14183 32937
rect -14217 32583 -14183 32617
rect -14217 32263 -14183 32297
rect -14217 31943 -14183 31977
rect -14057 32903 -14023 32937
rect -14057 32583 -14023 32617
rect -14057 32263 -14023 32297
rect -14057 31943 -14023 31977
rect -13897 32903 -13863 32937
rect -13897 32583 -13863 32617
rect -13897 32263 -13863 32297
rect -13897 31943 -13863 31977
rect -13737 32903 -13703 32937
rect -13737 32583 -13703 32617
rect -13737 32263 -13703 32297
rect -13737 31943 -13703 31977
rect -13577 32903 -13543 32937
rect -13577 32583 -13543 32617
rect -13577 32263 -13543 32297
rect -13577 31943 -13543 31977
rect -13417 32903 -13383 32937
rect -13417 32583 -13383 32617
rect -13417 32263 -13383 32297
rect -13417 31943 -13383 31977
rect -13257 32903 -13223 32937
rect -13257 32583 -13223 32617
rect -13257 32263 -13223 32297
rect -13257 31943 -13223 31977
rect -13097 32903 -13063 32937
rect -13097 32583 -13063 32617
rect -13097 32263 -13063 32297
rect -13097 31943 -13063 31977
rect -12937 32903 -12903 32937
rect -12937 32583 -12903 32617
rect -12937 32263 -12903 32297
rect -12937 31943 -12903 31977
rect -12777 32903 -12743 32937
rect -12777 32583 -12743 32617
rect -12777 32263 -12743 32297
rect -12777 31943 -12743 31977
rect -12617 32903 -12583 32937
rect -12617 32583 -12583 32617
rect -12617 32263 -12583 32297
rect -12617 31943 -12583 31977
rect -12457 32903 -12423 32937
rect -12457 32583 -12423 32617
rect -12457 32263 -12423 32297
rect -12457 31943 -12423 31977
rect -12297 32903 -12263 32937
rect -12297 32583 -12263 32617
rect -12297 32263 -12263 32297
rect -12297 31943 -12263 31977
rect -12137 32903 -12103 32937
rect -12137 32583 -12103 32617
rect -12137 32263 -12103 32297
rect -12137 31943 -12103 31977
rect -11977 32903 -11943 32937
rect -11977 32583 -11943 32617
rect -11977 32263 -11943 32297
rect -11977 31943 -11943 31977
rect -11817 32903 -11783 32937
rect -11817 32583 -11783 32617
rect -11817 32263 -11783 32297
rect -11817 31943 -11783 31977
rect -11657 32903 -11623 32937
rect -11657 32583 -11623 32617
rect -11657 32263 -11623 32297
rect -11657 31943 -11623 31977
rect -11497 32903 -11463 32937
rect -11497 32583 -11463 32617
rect -11177 32903 -11143 32937
rect -11177 32583 -11143 32617
rect -11497 32263 -11463 32297
rect -11497 31943 -11463 31977
rect -11337 32263 -11303 32297
rect -11337 31943 -11303 31977
rect -11177 32263 -11143 32297
rect -11177 31943 -11143 31977
rect -10857 32903 -10823 32937
rect -10857 32583 -10823 32617
rect -10857 32263 -10823 32297
rect -10857 31943 -10823 31977
rect -10697 32903 -10663 32937
rect -10697 32583 -10663 32617
rect -10697 32263 -10663 32297
rect -10697 31943 -10663 31977
rect -10537 32903 -10503 32937
rect -10537 32583 -10503 32617
rect -10537 32263 -10503 32297
rect -10537 31943 -10503 31977
rect -10377 32903 -10343 32937
rect -10377 32583 -10343 32617
rect -10377 32263 -10343 32297
rect -10377 31943 -10343 31977
rect -10217 32903 -10183 32937
rect -10217 32583 -10183 32617
rect -10217 32263 -10183 32297
rect -10217 31943 -10183 31977
rect -10057 32903 -10023 32937
rect -10057 32583 -10023 32617
rect -10057 32263 -10023 32297
rect -10057 31943 -10023 31977
rect -9897 32903 -9863 32937
rect -9897 32583 -9863 32617
rect -9897 32263 -9863 32297
rect -9897 31943 -9863 31977
rect -9737 32903 -9703 32937
rect -9737 32583 -9703 32617
rect -9737 32263 -9703 32297
rect -9737 31943 -9703 31977
rect -9577 32903 -9543 32937
rect -9577 32583 -9543 32617
rect -9577 32263 -9543 32297
rect -9577 31943 -9543 31977
rect -9417 32903 -9383 32937
rect -9417 32583 -9383 32617
rect -9417 32263 -9383 32297
rect -9417 31943 -9383 31977
rect -9257 32903 -9223 32937
rect -9257 32583 -9223 32617
rect -9257 32263 -9223 32297
rect -9257 31943 -9223 31977
rect -9097 32903 -9063 32937
rect -9097 32583 -9063 32617
rect -9097 32263 -9063 32297
rect -9097 31943 -9063 31977
rect -8937 32903 -8903 32937
rect -8937 32583 -8903 32617
rect -8937 32263 -8903 32297
rect -8937 31943 -8903 31977
rect -8777 32903 -8743 32937
rect -8777 32583 -8743 32617
rect -8777 32263 -8743 32297
rect -8777 31943 -8743 31977
rect -8617 32903 -8583 32937
rect -8617 32583 -8583 32617
rect -8617 32263 -8583 32297
rect -8617 31943 -8583 31977
rect -8457 32903 -8423 32937
rect -8457 32583 -8423 32617
rect -8457 32263 -8423 32297
rect -8457 31943 -8423 31977
rect -8297 32903 -8263 32937
rect -8297 32583 -8263 32617
rect -8297 32263 -8263 32297
rect -8297 31943 -8263 31977
rect -8137 32903 -8103 32937
rect -8137 32583 -8103 32617
rect -8137 32263 -8103 32297
rect -8137 31943 -8103 31977
rect -7977 32903 -7943 32937
rect -7977 32583 -7943 32617
rect -7977 32263 -7943 32297
rect -7977 31943 -7943 31977
rect -7817 32903 -7783 32937
rect -7817 32583 -7783 32617
rect -7817 32263 -7783 32297
rect -7817 31943 -7783 31977
rect -7657 32903 -7623 32937
rect -7657 32583 -7623 32617
rect -7657 32263 -7623 32297
rect -7657 31943 -7623 31977
rect -7497 32903 -7463 32937
rect -7497 32583 -7463 32617
rect -7497 32263 -7463 32297
rect -7497 31943 -7463 31977
rect -7337 32903 -7303 32937
rect -7337 32583 -7303 32617
rect -7337 32263 -7303 32297
rect -7337 31943 -7303 31977
rect -7177 32903 -7143 32937
rect -7177 32583 -7143 32617
rect -7177 32263 -7143 32297
rect -7177 31943 -7143 31977
rect -7017 32903 -6983 32937
rect -7017 32583 -6983 32617
rect -7017 32263 -6983 32297
rect -7017 31943 -6983 31977
rect -6857 32903 -6823 32937
rect -6857 32583 -6823 32617
rect -6857 32263 -6823 32297
rect -6857 31943 -6823 31977
rect -6697 32903 -6663 32937
rect -6697 32583 -6663 32617
rect -6697 32263 -6663 32297
rect -6697 31943 -6663 31977
rect -6537 32903 -6503 32937
rect -6537 32583 -6503 32617
rect -6537 32263 -6503 32297
rect -6537 31943 -6503 31977
rect -6377 32903 -6343 32937
rect -6377 32583 -6343 32617
rect -6377 32263 -6343 32297
rect -6377 31943 -6343 31977
rect -6217 32903 -6183 32937
rect -6217 32583 -6183 32617
rect -6217 32263 -6183 32297
rect -6217 31943 -6183 31977
rect -6057 32903 -6023 32937
rect -6057 32583 -6023 32617
rect -6057 32263 -6023 32297
rect -6057 31943 -6023 31977
rect -5897 32903 -5863 32937
rect -5897 32583 -5863 32617
rect -5897 32263 -5863 32297
rect -5897 31943 -5863 31977
rect -5737 32903 -5703 32937
rect -5737 32583 -5703 32617
rect -5737 32263 -5703 32297
rect -5737 31943 -5703 31977
rect -5577 32903 -5543 32937
rect -5577 32583 -5543 32617
rect -5577 32263 -5543 32297
rect -5577 31943 -5543 31977
rect -5417 32903 -5383 32937
rect -5417 32583 -5383 32617
rect -5417 32263 -5383 32297
rect -5417 31943 -5383 31977
rect -5257 32903 -5223 32937
rect -5257 32583 -5223 32617
rect -5257 32263 -5223 32297
rect -5257 31943 -5223 31977
rect -5097 32903 -5063 32937
rect -5097 32583 -5063 32617
rect -5097 32263 -5063 32297
rect -5097 31943 -5063 31977
rect -4937 32903 -4903 32937
rect -4937 32583 -4903 32617
rect -4937 32263 -4903 32297
rect -4937 31943 -4903 31977
rect -4777 32903 -4743 32937
rect -4777 32583 -4743 32617
rect -4777 32263 -4743 32297
rect -4777 31943 -4743 31977
rect -4617 32903 -4583 32937
rect -4617 32583 -4583 32617
rect -4617 32263 -4583 32297
rect -4617 31943 -4583 31977
rect -4457 32903 -4423 32937
rect -4457 32583 -4423 32617
rect -4457 32263 -4423 32297
rect -4457 31943 -4423 31977
rect -4297 32903 -4263 32937
rect -4297 32583 -4263 32617
rect -4297 32263 -4263 32297
rect -4297 31943 -4263 31977
rect -4137 32903 -4103 32937
rect -4137 32583 -4103 32617
rect -4137 32263 -4103 32297
rect -4137 31943 -4103 31977
rect -3977 32903 -3943 32937
rect -3977 32583 -3943 32617
rect -3977 32263 -3943 32297
rect -3977 31943 -3943 31977
rect -3657 32903 -3623 32937
rect -3657 32583 -3623 32617
rect -3657 32263 -3623 32297
rect -3657 31943 -3623 31977
rect -3497 32903 -3463 32937
rect -3497 32583 -3463 32617
rect -3497 32263 -3463 32297
rect -3497 31943 -3463 31977
rect -3337 32903 -3303 32937
rect -3337 32583 -3303 32617
rect -3337 32263 -3303 32297
rect -3337 31943 -3303 31977
rect -3177 32903 -3143 32937
rect -3177 32583 -3143 32617
rect -3177 32263 -3143 32297
rect -3177 31943 -3143 31977
rect -3017 32903 -2983 32937
rect -3017 32583 -2983 32617
rect -3017 32263 -2983 32297
rect -3017 31943 -2983 31977
rect -2857 32903 -2823 32937
rect -2857 32583 -2823 32617
rect -2857 32263 -2823 32297
rect -2857 31943 -2823 31977
rect -2697 32903 -2663 32937
rect -2697 32583 -2663 32617
rect -2697 32263 -2663 32297
rect -2697 31943 -2663 31977
rect -2377 32903 -2343 32937
rect -2377 32583 -2343 32617
rect -2377 32263 -2343 32297
rect -2377 31943 -2343 31977
rect -2057 32903 -2023 32937
rect -2057 32583 -2023 32617
rect -2057 32263 -2023 32297
rect -2057 31943 -2023 31977
rect -1737 32903 -1703 32937
rect -1737 32583 -1703 32617
rect -1737 32263 -1703 32297
rect -1737 31943 -1703 31977
rect -1417 32903 -1383 32937
rect -1417 32583 -1383 32617
rect -1417 32263 -1383 32297
rect -1417 31943 -1383 31977
rect -1097 32903 -1063 32937
rect -1097 32583 -1063 32617
rect -1097 32263 -1063 32297
rect -1097 31943 -1063 31977
<< metal1 >>
rect -29920 42866 -29840 42880
rect -29920 42814 -29906 42866
rect -29854 42814 -29840 42866
rect -29920 42800 -29840 42814
rect -29760 42866 -29680 42880
rect -29760 42814 -29746 42866
rect -29694 42814 -29680 42866
rect -29760 42800 -29680 42814
rect -29600 42866 -29520 42880
rect -29600 42814 -29586 42866
rect -29534 42814 -29520 42866
rect -29600 42800 -29520 42814
rect -29440 42866 -29360 42880
rect -29440 42814 -29426 42866
rect -29374 42814 -29360 42866
rect -29440 42800 -29360 42814
rect -29280 42866 -29200 42880
rect -29280 42814 -29266 42866
rect -29214 42814 -29200 42866
rect -29280 42800 -29200 42814
rect -29120 42866 -29040 42880
rect -29120 42814 -29106 42866
rect -29054 42814 -29040 42866
rect -29120 42800 -29040 42814
rect -28960 42866 -28880 42880
rect -28960 42814 -28946 42866
rect -28894 42814 -28880 42866
rect -28960 42800 -28880 42814
rect -28800 42866 -28720 42880
rect -28800 42814 -28786 42866
rect -28734 42814 -28720 42866
rect -28800 42800 -28720 42814
rect -28640 42866 -28560 42880
rect -28640 42814 -28626 42866
rect -28574 42814 -28560 42866
rect -28640 42800 -28560 42814
rect -28480 42866 -28400 42880
rect -28480 42814 -28466 42866
rect -28414 42814 -28400 42866
rect -28480 42800 -28400 42814
rect -28320 42866 -28240 42880
rect -28320 42814 -28306 42866
rect -28254 42814 -28240 42866
rect -28320 42800 -28240 42814
rect -28160 42866 -28080 42880
rect -28160 42814 -28146 42866
rect -28094 42814 -28080 42866
rect -28160 42800 -28080 42814
rect -28000 42866 -27920 42880
rect -28000 42814 -27986 42866
rect -27934 42814 -27920 42866
rect -28000 42800 -27920 42814
rect -27840 42866 -27760 42880
rect -27840 42814 -27826 42866
rect -27774 42814 -27760 42866
rect -27840 42800 -27760 42814
rect -27680 42866 -27600 42880
rect -27680 42814 -27666 42866
rect -27614 42814 -27600 42866
rect -27680 42800 -27600 42814
rect -27520 42866 -27440 42880
rect -27520 42814 -27506 42866
rect -27454 42814 -27440 42866
rect -27520 42800 -27440 42814
rect -27360 42866 -27280 42880
rect -27360 42814 -27346 42866
rect -27294 42814 -27280 42866
rect -27360 42800 -27280 42814
rect -27200 42866 -27120 42880
rect -27200 42814 -27186 42866
rect -27134 42814 -27120 42866
rect -27200 42800 -27120 42814
rect -27040 42866 -26960 42880
rect -27040 42814 -27026 42866
rect -26974 42814 -26960 42866
rect -27040 42800 -26960 42814
rect -26880 42866 -26800 42880
rect -26880 42814 -26866 42866
rect -26814 42814 -26800 42866
rect -26880 42800 -26800 42814
rect -26720 42866 -26640 42880
rect -26720 42814 -26706 42866
rect -26654 42814 -26640 42866
rect -26720 42800 -26640 42814
rect -26560 42866 -26480 42880
rect -26560 42814 -26546 42866
rect -26494 42814 -26480 42866
rect -26560 42800 -26480 42814
rect -26400 42866 -26320 42880
rect -26400 42814 -26386 42866
rect -26334 42814 -26320 42866
rect -26400 42800 -26320 42814
rect -26240 42866 -26160 42880
rect -26240 42814 -26226 42866
rect -26174 42814 -26160 42866
rect -26240 42800 -26160 42814
rect -26080 42866 -26000 42880
rect -26080 42814 -26066 42866
rect -26014 42814 -26000 42866
rect -26080 42800 -26000 42814
rect -25920 42866 -25840 42880
rect -25920 42814 -25906 42866
rect -25854 42814 -25840 42866
rect -25920 42800 -25840 42814
rect -25760 42866 -25680 42880
rect -25760 42814 -25746 42866
rect -25694 42814 -25680 42866
rect -25760 42800 -25680 42814
rect -25600 42866 -25520 42880
rect -25600 42814 -25586 42866
rect -25534 42814 -25520 42866
rect -25600 42800 -25520 42814
rect -25440 42866 -25360 42880
rect -25440 42814 -25426 42866
rect -25374 42814 -25360 42866
rect -25440 42800 -25360 42814
rect -25280 42866 -25200 42880
rect -25280 42814 -25266 42866
rect -25214 42814 -25200 42866
rect -25280 42800 -25200 42814
rect -25120 42866 -25040 42880
rect -25120 42814 -25106 42866
rect -25054 42814 -25040 42866
rect -25120 42800 -25040 42814
rect -24960 42866 -24880 42880
rect -24960 42814 -24946 42866
rect -24894 42814 -24880 42866
rect -24960 42800 -24880 42814
rect -24800 42866 -24720 42880
rect -24800 42814 -24786 42866
rect -24734 42814 -24720 42866
rect -24800 42800 -24720 42814
rect -24640 42866 -24560 42880
rect -24640 42814 -24626 42866
rect -24574 42814 -24560 42866
rect -24640 42800 -24560 42814
rect -24480 42866 -24400 42880
rect -24480 42814 -24466 42866
rect -24414 42814 -24400 42866
rect -24480 42800 -24400 42814
rect -24320 42866 -24240 42880
rect -24320 42814 -24306 42866
rect -24254 42814 -24240 42866
rect -24320 42800 -24240 42814
rect -24160 42866 -24080 42880
rect -24160 42814 -24146 42866
rect -24094 42814 -24080 42866
rect -24160 42800 -24080 42814
rect -24000 42866 -23920 42880
rect -24000 42814 -23986 42866
rect -23934 42814 -23920 42866
rect -24000 42800 -23920 42814
rect -23840 42866 -23760 42880
rect -23840 42814 -23826 42866
rect -23774 42814 -23760 42866
rect -23840 42800 -23760 42814
rect -23680 42866 -23600 42880
rect -23680 42814 -23666 42866
rect -23614 42814 -23600 42866
rect -23680 42800 -23600 42814
rect -23520 42866 -23440 42880
rect -23520 42814 -23506 42866
rect -23454 42814 -23440 42866
rect -23520 42800 -23440 42814
rect -23360 42866 -23280 42880
rect -23360 42814 -23346 42866
rect -23294 42814 -23280 42866
rect -23360 42800 -23280 42814
rect -23200 42866 -23120 42880
rect -23200 42814 -23186 42866
rect -23134 42814 -23120 42866
rect -23200 42800 -23120 42814
rect -23040 42866 -22960 42880
rect -23040 42814 -23026 42866
rect -22974 42814 -22960 42866
rect -23040 42800 -22960 42814
rect -22880 42866 -22800 42880
rect -22880 42814 -22866 42866
rect -22814 42814 -22800 42866
rect -22880 42800 -22800 42814
rect -22720 42866 -22640 42880
rect -22720 42814 -22706 42866
rect -22654 42814 -22640 42866
rect -22720 42800 -22640 42814
rect -22560 42866 -22480 42880
rect -22560 42814 -22546 42866
rect -22494 42814 -22480 42866
rect -22560 42800 -22480 42814
rect -22400 42866 -22320 42880
rect -22400 42814 -22386 42866
rect -22334 42814 -22320 42866
rect -22400 42800 -22320 42814
rect -22240 42866 -22160 42880
rect -22240 42814 -22226 42866
rect -22174 42814 -22160 42866
rect -22240 42800 -22160 42814
rect -22080 42866 -22000 42880
rect -22080 42814 -22066 42866
rect -22014 42814 -22000 42866
rect -22080 42800 -22000 42814
rect -21920 42866 -21840 42880
rect -21920 42814 -21906 42866
rect -21854 42814 -21840 42866
rect -21920 42800 -21840 42814
rect -21760 42866 -21680 42880
rect -21760 42814 -21746 42866
rect -21694 42814 -21680 42866
rect -21760 42800 -21680 42814
rect -21600 42866 -21520 42880
rect -21600 42814 -21586 42866
rect -21534 42814 -21520 42866
rect -21600 42800 -21520 42814
rect -21440 42866 -21360 42880
rect -21440 42814 -21426 42866
rect -21374 42814 -21360 42866
rect -21440 42800 -21360 42814
rect -21280 42866 -21200 42880
rect -21280 42814 -21266 42866
rect -21214 42814 -21200 42866
rect -21280 42800 -21200 42814
rect -21120 42866 -21040 42880
rect -21120 42814 -21106 42866
rect -21054 42814 -21040 42866
rect -21120 42800 -21040 42814
rect -20960 42866 -20880 42880
rect -20960 42814 -20946 42866
rect -20894 42814 -20880 42866
rect -20960 42800 -20880 42814
rect -20800 42866 -20720 42880
rect -20800 42814 -20786 42866
rect -20734 42814 -20720 42866
rect -20800 42800 -20720 42814
rect -20640 42866 -20560 42880
rect -20640 42814 -20626 42866
rect -20574 42814 -20560 42866
rect -20640 42800 -20560 42814
rect -20480 42866 -20400 42880
rect -20480 42814 -20466 42866
rect -20414 42814 -20400 42866
rect -20480 42800 -20400 42814
rect -20320 42866 -20240 42880
rect -20320 42814 -20306 42866
rect -20254 42814 -20240 42866
rect -20320 42800 -20240 42814
rect -20160 42866 -20080 42880
rect -20160 42814 -20146 42866
rect -20094 42814 -20080 42866
rect -20160 42800 -20080 42814
rect -20000 42866 -19920 42880
rect -20000 42814 -19986 42866
rect -19934 42814 -19920 42866
rect -20000 42800 -19920 42814
rect -19840 42866 -19760 42880
rect -19840 42814 -19826 42866
rect -19774 42814 -19760 42866
rect -19840 42800 -19760 42814
rect -19680 42866 -19600 42880
rect -19680 42814 -19666 42866
rect -19614 42814 -19600 42866
rect -19680 42800 -19600 42814
rect -19520 42866 -19440 42880
rect -19520 42814 -19506 42866
rect -19454 42814 -19440 42866
rect -19520 42800 -19440 42814
rect -19360 42866 -19280 42880
rect -19360 42814 -19346 42866
rect -19294 42814 -19280 42866
rect -19360 42800 -19280 42814
rect -19200 42866 -19120 42880
rect -19200 42814 -19186 42866
rect -19134 42814 -19120 42866
rect -19200 42800 -19120 42814
rect -19040 42866 -18960 42880
rect -19040 42814 -19026 42866
rect -18974 42814 -18960 42866
rect -19040 42800 -18960 42814
rect -18880 42866 -18800 42880
rect -18880 42814 -18866 42866
rect -18814 42814 -18800 42866
rect -18880 42800 -18800 42814
rect -18720 42866 -18640 42880
rect -18720 42814 -18706 42866
rect -18654 42814 -18640 42866
rect -18720 42800 -18640 42814
rect -18560 42866 -18480 42880
rect -18560 42814 -18546 42866
rect -18494 42814 -18480 42866
rect -18560 42800 -18480 42814
rect -18400 42866 -18320 42880
rect -18400 42814 -18386 42866
rect -18334 42814 -18320 42866
rect -18400 42800 -18320 42814
rect -18240 42866 -18160 42880
rect -18240 42814 -18226 42866
rect -18174 42814 -18160 42866
rect -18240 42800 -18160 42814
rect -18080 42866 -18000 42880
rect -18080 42814 -18066 42866
rect -18014 42814 -18000 42866
rect -18080 42800 -18000 42814
rect -17920 42866 -17840 42880
rect -17920 42814 -17906 42866
rect -17854 42814 -17840 42866
rect -17920 42800 -17840 42814
rect -17760 42866 -17680 42880
rect -17760 42814 -17746 42866
rect -17694 42814 -17680 42866
rect -17760 42800 -17680 42814
rect -17600 42866 -17520 42880
rect -17600 42814 -17586 42866
rect -17534 42814 -17520 42866
rect -17600 42800 -17520 42814
rect -17440 42866 -17360 42880
rect -17440 42814 -17426 42866
rect -17374 42814 -17360 42866
rect -17440 42800 -17360 42814
rect -17280 42866 -17200 42880
rect -17280 42814 -17266 42866
rect -17214 42814 -17200 42866
rect -17280 42800 -17200 42814
rect -17120 42866 -17040 42880
rect -17120 42814 -17106 42866
rect -17054 42814 -17040 42866
rect -17120 42800 -17040 42814
rect -16960 42866 -16880 42880
rect -16960 42814 -16946 42866
rect -16894 42814 -16880 42866
rect -16960 42800 -16880 42814
rect -16800 42866 -16720 42880
rect -16800 42814 -16786 42866
rect -16734 42814 -16720 42866
rect -16800 42800 -16720 42814
rect -16640 42866 -16560 42880
rect -16640 42814 -16626 42866
rect -16574 42814 -16560 42866
rect -16640 42800 -16560 42814
rect -16480 42866 -16400 42880
rect -16480 42814 -16466 42866
rect -16414 42814 -16400 42866
rect -16480 42800 -16400 42814
rect -16320 42866 -16240 42880
rect -16320 42814 -16306 42866
rect -16254 42814 -16240 42866
rect -16320 42800 -16240 42814
rect -16160 42866 -16080 42880
rect -16160 42814 -16146 42866
rect -16094 42814 -16080 42866
rect -16160 42800 -16080 42814
rect -16000 42866 -15920 42880
rect -16000 42814 -15986 42866
rect -15934 42814 -15920 42866
rect -16000 42800 -15920 42814
rect -15840 42866 -15760 42880
rect -15840 42814 -15826 42866
rect -15774 42814 -15760 42866
rect -15840 42800 -15760 42814
rect -15680 42866 -15600 42880
rect -15680 42814 -15666 42866
rect -15614 42814 -15600 42866
rect -15680 42800 -15600 42814
rect -15520 42866 -15440 42880
rect -15520 42814 -15506 42866
rect -15454 42814 -15440 42866
rect -15520 42800 -15440 42814
rect -15360 42866 -15280 42880
rect -15360 42814 -15346 42866
rect -15294 42814 -15280 42866
rect -15360 42800 -15280 42814
rect -15200 42866 -15120 42880
rect -15200 42814 -15186 42866
rect -15134 42814 -15120 42866
rect -15200 42800 -15120 42814
rect -15040 42866 -14960 42880
rect -15040 42814 -15026 42866
rect -14974 42814 -14960 42866
rect -15040 42800 -14960 42814
rect -14880 42866 -14800 42880
rect -14880 42814 -14866 42866
rect -14814 42814 -14800 42866
rect -14880 42800 -14800 42814
rect -14720 42866 -14640 42880
rect -14720 42814 -14706 42866
rect -14654 42814 -14640 42866
rect -14720 42800 -14640 42814
rect -14560 42866 -14480 42880
rect -14560 42814 -14546 42866
rect -14494 42814 -14480 42866
rect -14560 42800 -14480 42814
rect -14400 42866 -14320 42880
rect -14400 42814 -14386 42866
rect -14334 42814 -14320 42866
rect -14400 42800 -14320 42814
rect -14240 42866 -14160 42880
rect -14240 42814 -14226 42866
rect -14174 42814 -14160 42866
rect -14240 42800 -14160 42814
rect -14080 42866 -14000 42880
rect -14080 42814 -14066 42866
rect -14014 42814 -14000 42866
rect -14080 42800 -14000 42814
rect -13920 42866 -13840 42880
rect -13920 42814 -13906 42866
rect -13854 42814 -13840 42866
rect -13920 42800 -13840 42814
rect -13760 42866 -13680 42880
rect -13760 42814 -13746 42866
rect -13694 42814 -13680 42866
rect -13760 42800 -13680 42814
rect -13600 42866 -13520 42880
rect -13600 42814 -13586 42866
rect -13534 42814 -13520 42866
rect -13600 42800 -13520 42814
rect -13440 42866 -13360 42880
rect -13440 42814 -13426 42866
rect -13374 42814 -13360 42866
rect -13440 42800 -13360 42814
rect -13280 42866 -13200 42880
rect -13280 42814 -13266 42866
rect -13214 42814 -13200 42866
rect -13280 42800 -13200 42814
rect -13120 42866 -13040 42880
rect -13120 42814 -13106 42866
rect -13054 42814 -13040 42866
rect -13120 42800 -13040 42814
rect -12960 42866 -12880 42880
rect -12960 42814 -12946 42866
rect -12894 42814 -12880 42866
rect -12960 42800 -12880 42814
rect -12800 42866 -12720 42880
rect -12800 42814 -12786 42866
rect -12734 42814 -12720 42866
rect -12800 42800 -12720 42814
rect -12640 42866 -12560 42880
rect -12640 42814 -12626 42866
rect -12574 42814 -12560 42866
rect -12640 42800 -12560 42814
rect -12480 42866 -12400 42880
rect -12480 42814 -12466 42866
rect -12414 42814 -12400 42866
rect -12480 42800 -12400 42814
rect -12320 42866 -12240 42880
rect -12320 42814 -12306 42866
rect -12254 42814 -12240 42866
rect -12320 42800 -12240 42814
rect -11360 42866 -11280 42880
rect -11360 42814 -11346 42866
rect -11294 42814 -11280 42866
rect -11360 42800 -11280 42814
rect -11200 42866 -11120 42880
rect -11200 42814 -11186 42866
rect -11134 42814 -11120 42866
rect -11200 42800 -11120 42814
rect -11040 42866 -10960 42880
rect -11040 42814 -11026 42866
rect -10974 42814 -10960 42866
rect -11040 42800 -10960 42814
rect -10880 42866 -10800 42880
rect -10880 42814 -10866 42866
rect -10814 42814 -10800 42866
rect -10880 42800 -10800 42814
rect -10720 42866 -10640 42880
rect -10720 42814 -10706 42866
rect -10654 42814 -10640 42866
rect -10720 42800 -10640 42814
rect -10560 42866 -10480 42880
rect -10560 42814 -10546 42866
rect -10494 42814 -10480 42866
rect -10560 42800 -10480 42814
rect -10400 42866 -10320 42880
rect -10400 42814 -10386 42866
rect -10334 42814 -10320 42866
rect -10400 42800 -10320 42814
rect -10240 42866 -10160 42880
rect -10240 42814 -10226 42866
rect -10174 42814 -10160 42866
rect -10240 42800 -10160 42814
rect -10080 42866 -10000 42880
rect -10080 42814 -10066 42866
rect -10014 42814 -10000 42866
rect -10080 42800 -10000 42814
rect -9920 42866 -9840 42880
rect -9920 42814 -9906 42866
rect -9854 42814 -9840 42866
rect -9920 42800 -9840 42814
rect -9760 42866 -9680 42880
rect -9760 42814 -9746 42866
rect -9694 42814 -9680 42866
rect -9760 42800 -9680 42814
rect -9600 42866 -9520 42880
rect -9600 42814 -9586 42866
rect -9534 42814 -9520 42866
rect -9600 42800 -9520 42814
rect -9440 42866 -9360 42880
rect -9440 42814 -9426 42866
rect -9374 42814 -9360 42866
rect -9440 42800 -9360 42814
rect -9280 42866 -9200 42880
rect -9280 42814 -9266 42866
rect -9214 42814 -9200 42866
rect -9280 42800 -9200 42814
rect -9120 42866 -9040 42880
rect -9120 42814 -9106 42866
rect -9054 42814 -9040 42866
rect -9120 42800 -9040 42814
rect -8960 42866 -8880 42880
rect -8960 42814 -8946 42866
rect -8894 42814 -8880 42866
rect -8960 42800 -8880 42814
rect -8800 42866 -8720 42880
rect -8800 42814 -8786 42866
rect -8734 42814 -8720 42866
rect -8800 42800 -8720 42814
rect -8640 42866 -8560 42880
rect -8640 42814 -8626 42866
rect -8574 42814 -8560 42866
rect -8640 42800 -8560 42814
rect -8480 42866 -8400 42880
rect -8480 42814 -8466 42866
rect -8414 42814 -8400 42866
rect -8480 42800 -8400 42814
rect -8320 42866 -8240 42880
rect -8320 42814 -8306 42866
rect -8254 42814 -8240 42866
rect -8320 42800 -8240 42814
rect -8160 42866 -8080 42880
rect -8160 42814 -8146 42866
rect -8094 42814 -8080 42866
rect -8160 42800 -8080 42814
rect -8000 42866 -7920 42880
rect -8000 42814 -7986 42866
rect -7934 42814 -7920 42866
rect -8000 42800 -7920 42814
rect -7840 42866 -7760 42880
rect -7840 42814 -7826 42866
rect -7774 42814 -7760 42866
rect -7840 42800 -7760 42814
rect -7680 42866 -7600 42880
rect -7680 42814 -7666 42866
rect -7614 42814 -7600 42866
rect -7680 42800 -7600 42814
rect -7520 42866 -7440 42880
rect -7520 42814 -7506 42866
rect -7454 42814 -7440 42866
rect -7520 42800 -7440 42814
rect -7360 42866 -7280 42880
rect -7360 42814 -7346 42866
rect -7294 42814 -7280 42866
rect -7360 42800 -7280 42814
rect -7200 42866 -7120 42880
rect -7200 42814 -7186 42866
rect -7134 42814 -7120 42866
rect -7200 42800 -7120 42814
rect -7040 42866 -6960 42880
rect -7040 42814 -7026 42866
rect -6974 42814 -6960 42866
rect -7040 42800 -6960 42814
rect -6880 42866 -6800 42880
rect -6880 42814 -6866 42866
rect -6814 42814 -6800 42866
rect -6880 42800 -6800 42814
rect -6720 42866 -6640 42880
rect -6720 42814 -6706 42866
rect -6654 42814 -6640 42866
rect -6720 42800 -6640 42814
rect -6560 42866 -6480 42880
rect -6560 42814 -6546 42866
rect -6494 42814 -6480 42866
rect -6560 42800 -6480 42814
rect -6400 42866 -6320 42880
rect -6400 42814 -6386 42866
rect -6334 42814 -6320 42866
rect -6400 42800 -6320 42814
rect -6240 42866 -6160 42880
rect -6240 42814 -6226 42866
rect -6174 42814 -6160 42866
rect -6240 42800 -6160 42814
rect -6080 42866 -6000 42880
rect -6080 42814 -6066 42866
rect -6014 42814 -6000 42866
rect -6080 42800 -6000 42814
rect -5920 42866 -5840 42880
rect -5920 42814 -5906 42866
rect -5854 42814 -5840 42866
rect -5920 42800 -5840 42814
rect -5760 42866 -5680 42880
rect -5760 42814 -5746 42866
rect -5694 42814 -5680 42866
rect -5760 42800 -5680 42814
rect -5600 42866 -5520 42880
rect -5600 42814 -5586 42866
rect -5534 42814 -5520 42866
rect -5600 42800 -5520 42814
rect -5440 42866 -5360 42880
rect -5440 42814 -5426 42866
rect -5374 42814 -5360 42866
rect -5440 42800 -5360 42814
rect -5280 42866 -5200 42880
rect -5280 42814 -5266 42866
rect -5214 42814 -5200 42866
rect -5280 42800 -5200 42814
rect -5120 42866 -5040 42880
rect -5120 42814 -5106 42866
rect -5054 42814 -5040 42866
rect -5120 42800 -5040 42814
rect -4960 42866 -4880 42880
rect -4960 42814 -4946 42866
rect -4894 42814 -4880 42866
rect -4960 42800 -4880 42814
rect -4800 42866 -4720 42880
rect -4800 42814 -4786 42866
rect -4734 42814 -4720 42866
rect -4800 42800 -4720 42814
rect -4640 42866 -4560 42880
rect -4640 42814 -4626 42866
rect -4574 42814 -4560 42866
rect -4640 42800 -4560 42814
rect -4480 42866 -4400 42880
rect -4480 42814 -4466 42866
rect -4414 42814 -4400 42866
rect -4480 42800 -4400 42814
rect -4320 42866 -4240 42880
rect -4320 42814 -4306 42866
rect -4254 42814 -4240 42866
rect -4320 42800 -4240 42814
rect -4160 42866 -4080 42880
rect -4160 42814 -4146 42866
rect -4094 42814 -4080 42866
rect -4160 42800 -4080 42814
rect -4000 42866 -3920 42880
rect -4000 42814 -3986 42866
rect -3934 42814 -3920 42866
rect -4000 42800 -3920 42814
rect -3680 42866 -3600 42880
rect -3680 42814 -3666 42866
rect -3614 42814 -3600 42866
rect -3680 42800 -3600 42814
rect -3520 42866 -3440 42880
rect -3520 42814 -3506 42866
rect -3454 42814 -3440 42866
rect -3520 42800 -3440 42814
rect -3360 42866 -3280 42880
rect -3360 42814 -3346 42866
rect -3294 42814 -3280 42866
rect -3360 42800 -3280 42814
rect -3040 42866 -2960 42880
rect -3040 42814 -3026 42866
rect -2974 42814 -2960 42866
rect -3040 42800 -2960 42814
rect -2720 42866 -2640 42880
rect -2720 42814 -2706 42866
rect -2654 42814 -2640 42866
rect -2720 42800 -2640 42814
rect -2560 42866 -2480 42880
rect -2560 42814 -2546 42866
rect -2494 42814 -2480 42866
rect -2560 42800 -2480 42814
rect -2400 42866 -2320 42880
rect -2400 42814 -2386 42866
rect -2334 42814 -2320 42866
rect -2400 42800 -2320 42814
rect -2240 42866 -2160 42880
rect -2240 42814 -2226 42866
rect -2174 42814 -2160 42866
rect -2240 42800 -2160 42814
rect -2080 42866 -2000 42880
rect -2080 42814 -2066 42866
rect -2014 42814 -2000 42866
rect -2080 42800 -2000 42814
rect -1760 42866 -1680 42880
rect -1760 42814 -1746 42866
rect -1694 42814 -1680 42866
rect -1760 42800 -1680 42814
rect -1440 42866 -1360 42880
rect -1440 42814 -1426 42866
rect -1374 42814 -1360 42866
rect -1440 42800 -1360 42814
rect -1120 42866 -1040 42880
rect -1120 42814 -1106 42866
rect -1054 42814 -1040 42866
rect -1120 42800 -1040 42814
rect -29920 42546 -29840 42560
rect -29920 42494 -29906 42546
rect -29854 42494 -29840 42546
rect -29920 42480 -29840 42494
rect -29760 42546 -29680 42560
rect -29760 42494 -29746 42546
rect -29694 42494 -29680 42546
rect -29760 42480 -29680 42494
rect -29600 42546 -29520 42560
rect -29600 42494 -29586 42546
rect -29534 42494 -29520 42546
rect -29600 42480 -29520 42494
rect -29440 42546 -29360 42560
rect -29440 42494 -29426 42546
rect -29374 42494 -29360 42546
rect -29440 42480 -29360 42494
rect -29280 42546 -29200 42560
rect -29280 42494 -29266 42546
rect -29214 42494 -29200 42546
rect -29280 42480 -29200 42494
rect -29120 42546 -29040 42560
rect -29120 42494 -29106 42546
rect -29054 42494 -29040 42546
rect -29120 42480 -29040 42494
rect -28960 42546 -28880 42560
rect -28960 42494 -28946 42546
rect -28894 42494 -28880 42546
rect -28960 42480 -28880 42494
rect -28800 42546 -28720 42560
rect -28800 42494 -28786 42546
rect -28734 42494 -28720 42546
rect -28800 42480 -28720 42494
rect -28640 42546 -28560 42560
rect -28640 42494 -28626 42546
rect -28574 42494 -28560 42546
rect -28640 42480 -28560 42494
rect -28480 42546 -28400 42560
rect -28480 42494 -28466 42546
rect -28414 42494 -28400 42546
rect -28480 42480 -28400 42494
rect -28320 42546 -28240 42560
rect -28320 42494 -28306 42546
rect -28254 42494 -28240 42546
rect -28320 42480 -28240 42494
rect -28160 42546 -28080 42560
rect -28160 42494 -28146 42546
rect -28094 42494 -28080 42546
rect -28160 42480 -28080 42494
rect -28000 42546 -27920 42560
rect -28000 42494 -27986 42546
rect -27934 42494 -27920 42546
rect -28000 42480 -27920 42494
rect -27840 42546 -27760 42560
rect -27840 42494 -27826 42546
rect -27774 42494 -27760 42546
rect -27840 42480 -27760 42494
rect -27680 42546 -27600 42560
rect -27680 42494 -27666 42546
rect -27614 42494 -27600 42546
rect -27680 42480 -27600 42494
rect -27520 42546 -27440 42560
rect -27520 42494 -27506 42546
rect -27454 42494 -27440 42546
rect -27520 42480 -27440 42494
rect -27360 42546 -27280 42560
rect -27360 42494 -27346 42546
rect -27294 42494 -27280 42546
rect -27360 42480 -27280 42494
rect -27200 42546 -27120 42560
rect -27200 42494 -27186 42546
rect -27134 42494 -27120 42546
rect -27200 42480 -27120 42494
rect -27040 42546 -26960 42560
rect -27040 42494 -27026 42546
rect -26974 42494 -26960 42546
rect -27040 42480 -26960 42494
rect -26880 42546 -26800 42560
rect -26880 42494 -26866 42546
rect -26814 42494 -26800 42546
rect -26880 42480 -26800 42494
rect -26720 42546 -26640 42560
rect -26720 42494 -26706 42546
rect -26654 42494 -26640 42546
rect -26720 42480 -26640 42494
rect -26560 42546 -26480 42560
rect -26560 42494 -26546 42546
rect -26494 42494 -26480 42546
rect -26560 42480 -26480 42494
rect -26400 42546 -26320 42560
rect -26400 42494 -26386 42546
rect -26334 42494 -26320 42546
rect -26400 42480 -26320 42494
rect -26240 42546 -26160 42560
rect -26240 42494 -26226 42546
rect -26174 42494 -26160 42546
rect -26240 42480 -26160 42494
rect -26080 42546 -26000 42560
rect -26080 42494 -26066 42546
rect -26014 42494 -26000 42546
rect -26080 42480 -26000 42494
rect -25920 42546 -25840 42560
rect -25920 42494 -25906 42546
rect -25854 42494 -25840 42546
rect -25920 42480 -25840 42494
rect -25760 42546 -25680 42560
rect -25760 42494 -25746 42546
rect -25694 42494 -25680 42546
rect -25760 42480 -25680 42494
rect -25600 42546 -25520 42560
rect -25600 42494 -25586 42546
rect -25534 42494 -25520 42546
rect -25600 42480 -25520 42494
rect -25440 42546 -25360 42560
rect -25440 42494 -25426 42546
rect -25374 42494 -25360 42546
rect -25440 42480 -25360 42494
rect -25280 42546 -25200 42560
rect -25280 42494 -25266 42546
rect -25214 42494 -25200 42546
rect -25280 42480 -25200 42494
rect -25120 42546 -25040 42560
rect -25120 42494 -25106 42546
rect -25054 42494 -25040 42546
rect -25120 42480 -25040 42494
rect -24960 42546 -24880 42560
rect -24960 42494 -24946 42546
rect -24894 42494 -24880 42546
rect -24960 42480 -24880 42494
rect -24800 42546 -24720 42560
rect -24800 42494 -24786 42546
rect -24734 42494 -24720 42546
rect -24800 42480 -24720 42494
rect -24640 42546 -24560 42560
rect -24640 42494 -24626 42546
rect -24574 42494 -24560 42546
rect -24640 42480 -24560 42494
rect -24480 42546 -24400 42560
rect -24480 42494 -24466 42546
rect -24414 42494 -24400 42546
rect -24480 42480 -24400 42494
rect -24320 42546 -24240 42560
rect -24320 42494 -24306 42546
rect -24254 42494 -24240 42546
rect -24320 42480 -24240 42494
rect -24160 42546 -24080 42560
rect -24160 42494 -24146 42546
rect -24094 42494 -24080 42546
rect -24160 42480 -24080 42494
rect -24000 42546 -23920 42560
rect -24000 42494 -23986 42546
rect -23934 42494 -23920 42546
rect -24000 42480 -23920 42494
rect -23840 42546 -23760 42560
rect -23840 42494 -23826 42546
rect -23774 42494 -23760 42546
rect -23840 42480 -23760 42494
rect -23680 42546 -23600 42560
rect -23680 42494 -23666 42546
rect -23614 42494 -23600 42546
rect -23680 42480 -23600 42494
rect -23520 42546 -23440 42560
rect -23520 42494 -23506 42546
rect -23454 42494 -23440 42546
rect -23520 42480 -23440 42494
rect -23360 42546 -23280 42560
rect -23360 42494 -23346 42546
rect -23294 42494 -23280 42546
rect -23360 42480 -23280 42494
rect -23200 42546 -23120 42560
rect -23200 42494 -23186 42546
rect -23134 42494 -23120 42546
rect -23200 42480 -23120 42494
rect -23040 42546 -22960 42560
rect -23040 42494 -23026 42546
rect -22974 42494 -22960 42546
rect -23040 42480 -22960 42494
rect -22880 42546 -22800 42560
rect -22880 42494 -22866 42546
rect -22814 42494 -22800 42546
rect -22880 42480 -22800 42494
rect -22720 42546 -22640 42560
rect -22720 42494 -22706 42546
rect -22654 42494 -22640 42546
rect -22720 42480 -22640 42494
rect -22560 42546 -22480 42560
rect -22560 42494 -22546 42546
rect -22494 42494 -22480 42546
rect -22560 42480 -22480 42494
rect -22400 42546 -22320 42560
rect -22400 42494 -22386 42546
rect -22334 42494 -22320 42546
rect -22400 42480 -22320 42494
rect -22240 42546 -22160 42560
rect -22240 42494 -22226 42546
rect -22174 42494 -22160 42546
rect -22240 42480 -22160 42494
rect -22080 42546 -22000 42560
rect -22080 42494 -22066 42546
rect -22014 42494 -22000 42546
rect -22080 42480 -22000 42494
rect -21920 42546 -21840 42560
rect -21920 42494 -21906 42546
rect -21854 42494 -21840 42546
rect -21920 42480 -21840 42494
rect -21760 42546 -21680 42560
rect -21760 42494 -21746 42546
rect -21694 42494 -21680 42546
rect -21760 42480 -21680 42494
rect -21600 42546 -21520 42560
rect -21600 42494 -21586 42546
rect -21534 42494 -21520 42546
rect -21600 42480 -21520 42494
rect -21440 42546 -21360 42560
rect -21440 42494 -21426 42546
rect -21374 42494 -21360 42546
rect -21440 42480 -21360 42494
rect -21280 42546 -21200 42560
rect -21280 42494 -21266 42546
rect -21214 42494 -21200 42546
rect -21280 42480 -21200 42494
rect -21120 42546 -21040 42560
rect -21120 42494 -21106 42546
rect -21054 42494 -21040 42546
rect -21120 42480 -21040 42494
rect -20960 42546 -20880 42560
rect -20960 42494 -20946 42546
rect -20894 42494 -20880 42546
rect -20960 42480 -20880 42494
rect -20800 42546 -20720 42560
rect -20800 42494 -20786 42546
rect -20734 42494 -20720 42546
rect -20800 42480 -20720 42494
rect -20640 42546 -20560 42560
rect -20640 42494 -20626 42546
rect -20574 42494 -20560 42546
rect -20640 42480 -20560 42494
rect -20480 42546 -20400 42560
rect -20480 42494 -20466 42546
rect -20414 42494 -20400 42546
rect -20480 42480 -20400 42494
rect -20320 42546 -20240 42560
rect -20320 42494 -20306 42546
rect -20254 42494 -20240 42546
rect -20320 42480 -20240 42494
rect -20160 42546 -20080 42560
rect -20160 42494 -20146 42546
rect -20094 42494 -20080 42546
rect -20160 42480 -20080 42494
rect -20000 42546 -19920 42560
rect -20000 42494 -19986 42546
rect -19934 42494 -19920 42546
rect -20000 42480 -19920 42494
rect -19840 42546 -19760 42560
rect -19840 42494 -19826 42546
rect -19774 42494 -19760 42546
rect -19840 42480 -19760 42494
rect -19680 42546 -19600 42560
rect -19680 42494 -19666 42546
rect -19614 42494 -19600 42546
rect -19680 42480 -19600 42494
rect -19520 42546 -19440 42560
rect -19520 42494 -19506 42546
rect -19454 42494 -19440 42546
rect -19520 42480 -19440 42494
rect -19360 42546 -19280 42560
rect -19360 42494 -19346 42546
rect -19294 42494 -19280 42546
rect -19360 42480 -19280 42494
rect -19200 42546 -19120 42560
rect -19200 42494 -19186 42546
rect -19134 42494 -19120 42546
rect -19200 42480 -19120 42494
rect -19040 42546 -18960 42560
rect -19040 42494 -19026 42546
rect -18974 42494 -18960 42546
rect -19040 42480 -18960 42494
rect -18880 42546 -18800 42560
rect -18880 42494 -18866 42546
rect -18814 42494 -18800 42546
rect -18880 42480 -18800 42494
rect -18720 42546 -18640 42560
rect -18720 42494 -18706 42546
rect -18654 42494 -18640 42546
rect -18720 42480 -18640 42494
rect -18560 42546 -18480 42560
rect -18560 42494 -18546 42546
rect -18494 42494 -18480 42546
rect -18560 42480 -18480 42494
rect -18400 42546 -18320 42560
rect -18400 42494 -18386 42546
rect -18334 42494 -18320 42546
rect -18400 42480 -18320 42494
rect -18240 42546 -18160 42560
rect -18240 42494 -18226 42546
rect -18174 42494 -18160 42546
rect -18240 42480 -18160 42494
rect -18080 42546 -18000 42560
rect -18080 42494 -18066 42546
rect -18014 42494 -18000 42546
rect -18080 42480 -18000 42494
rect -17920 42546 -17840 42560
rect -17920 42494 -17906 42546
rect -17854 42494 -17840 42546
rect -17920 42480 -17840 42494
rect -17760 42546 -17680 42560
rect -17760 42494 -17746 42546
rect -17694 42494 -17680 42546
rect -17760 42480 -17680 42494
rect -17600 42546 -17520 42560
rect -17600 42494 -17586 42546
rect -17534 42494 -17520 42546
rect -17600 42480 -17520 42494
rect -17440 42546 -17360 42560
rect -17440 42494 -17426 42546
rect -17374 42494 -17360 42546
rect -17440 42480 -17360 42494
rect -17280 42546 -17200 42560
rect -17280 42494 -17266 42546
rect -17214 42494 -17200 42546
rect -17280 42480 -17200 42494
rect -17120 42546 -17040 42560
rect -17120 42494 -17106 42546
rect -17054 42494 -17040 42546
rect -17120 42480 -17040 42494
rect -16960 42546 -16880 42560
rect -16960 42494 -16946 42546
rect -16894 42494 -16880 42546
rect -16960 42480 -16880 42494
rect -16800 42546 -16720 42560
rect -16800 42494 -16786 42546
rect -16734 42494 -16720 42546
rect -16800 42480 -16720 42494
rect -16640 42546 -16560 42560
rect -16640 42494 -16626 42546
rect -16574 42494 -16560 42546
rect -16640 42480 -16560 42494
rect -16480 42546 -16400 42560
rect -16480 42494 -16466 42546
rect -16414 42494 -16400 42546
rect -16480 42480 -16400 42494
rect -16320 42546 -16240 42560
rect -16320 42494 -16306 42546
rect -16254 42494 -16240 42546
rect -16320 42480 -16240 42494
rect -16160 42546 -16080 42560
rect -16160 42494 -16146 42546
rect -16094 42494 -16080 42546
rect -16160 42480 -16080 42494
rect -16000 42546 -15920 42560
rect -16000 42494 -15986 42546
rect -15934 42494 -15920 42546
rect -16000 42480 -15920 42494
rect -15840 42546 -15760 42560
rect -15840 42494 -15826 42546
rect -15774 42494 -15760 42546
rect -15840 42480 -15760 42494
rect -15680 42546 -15600 42560
rect -15680 42494 -15666 42546
rect -15614 42494 -15600 42546
rect -15680 42480 -15600 42494
rect -15520 42546 -15440 42560
rect -15520 42494 -15506 42546
rect -15454 42494 -15440 42546
rect -15520 42480 -15440 42494
rect -15360 42546 -15280 42560
rect -15360 42494 -15346 42546
rect -15294 42494 -15280 42546
rect -15360 42480 -15280 42494
rect -15200 42546 -15120 42560
rect -15200 42494 -15186 42546
rect -15134 42494 -15120 42546
rect -15200 42480 -15120 42494
rect -15040 42546 -14960 42560
rect -15040 42494 -15026 42546
rect -14974 42494 -14960 42546
rect -15040 42480 -14960 42494
rect -14880 42546 -14800 42560
rect -14880 42494 -14866 42546
rect -14814 42494 -14800 42546
rect -14880 42480 -14800 42494
rect -14720 42546 -14640 42560
rect -14720 42494 -14706 42546
rect -14654 42494 -14640 42546
rect -14720 42480 -14640 42494
rect -14560 42546 -14480 42560
rect -14560 42494 -14546 42546
rect -14494 42494 -14480 42546
rect -14560 42480 -14480 42494
rect -14400 42546 -14320 42560
rect -14400 42494 -14386 42546
rect -14334 42494 -14320 42546
rect -14400 42480 -14320 42494
rect -14240 42546 -14160 42560
rect -14240 42494 -14226 42546
rect -14174 42494 -14160 42546
rect -14240 42480 -14160 42494
rect -14080 42546 -14000 42560
rect -14080 42494 -14066 42546
rect -14014 42494 -14000 42546
rect -14080 42480 -14000 42494
rect -13920 42546 -13840 42560
rect -13920 42494 -13906 42546
rect -13854 42494 -13840 42546
rect -13920 42480 -13840 42494
rect -13760 42546 -13680 42560
rect -13760 42494 -13746 42546
rect -13694 42494 -13680 42546
rect -13760 42480 -13680 42494
rect -13600 42546 -13520 42560
rect -13600 42494 -13586 42546
rect -13534 42494 -13520 42546
rect -13600 42480 -13520 42494
rect -13440 42546 -13360 42560
rect -13440 42494 -13426 42546
rect -13374 42494 -13360 42546
rect -13440 42480 -13360 42494
rect -13280 42546 -13200 42560
rect -13280 42494 -13266 42546
rect -13214 42494 -13200 42546
rect -13280 42480 -13200 42494
rect -13120 42546 -13040 42560
rect -13120 42494 -13106 42546
rect -13054 42494 -13040 42546
rect -13120 42480 -13040 42494
rect -12960 42546 -12880 42560
rect -12960 42494 -12946 42546
rect -12894 42494 -12880 42546
rect -12960 42480 -12880 42494
rect -12800 42546 -12720 42560
rect -12800 42494 -12786 42546
rect -12734 42494 -12720 42546
rect -12800 42480 -12720 42494
rect -12640 42546 -12560 42560
rect -12640 42494 -12626 42546
rect -12574 42494 -12560 42546
rect -12640 42480 -12560 42494
rect -12480 42546 -12400 42560
rect -12480 42494 -12466 42546
rect -12414 42494 -12400 42546
rect -12480 42480 -12400 42494
rect -12320 42546 -12240 42560
rect -12320 42494 -12306 42546
rect -12254 42494 -12240 42546
rect -12320 42480 -12240 42494
rect -11360 42546 -11280 42560
rect -11360 42494 -11346 42546
rect -11294 42494 -11280 42546
rect -11360 42480 -11280 42494
rect -11200 42546 -11120 42560
rect -11200 42494 -11186 42546
rect -11134 42494 -11120 42546
rect -11200 42480 -11120 42494
rect -11040 42546 -10960 42560
rect -11040 42494 -11026 42546
rect -10974 42494 -10960 42546
rect -11040 42480 -10960 42494
rect -10880 42546 -10800 42560
rect -10880 42494 -10866 42546
rect -10814 42494 -10800 42546
rect -10880 42480 -10800 42494
rect -10720 42546 -10640 42560
rect -10720 42494 -10706 42546
rect -10654 42494 -10640 42546
rect -10720 42480 -10640 42494
rect -10560 42546 -10480 42560
rect -10560 42494 -10546 42546
rect -10494 42494 -10480 42546
rect -10560 42480 -10480 42494
rect -10400 42546 -10320 42560
rect -10400 42494 -10386 42546
rect -10334 42494 -10320 42546
rect -10400 42480 -10320 42494
rect -10240 42546 -10160 42560
rect -10240 42494 -10226 42546
rect -10174 42494 -10160 42546
rect -10240 42480 -10160 42494
rect -10080 42546 -10000 42560
rect -10080 42494 -10066 42546
rect -10014 42494 -10000 42546
rect -10080 42480 -10000 42494
rect -9920 42546 -9840 42560
rect -9920 42494 -9906 42546
rect -9854 42494 -9840 42546
rect -9920 42480 -9840 42494
rect -9760 42546 -9680 42560
rect -9760 42494 -9746 42546
rect -9694 42494 -9680 42546
rect -9760 42480 -9680 42494
rect -9600 42546 -9520 42560
rect -9600 42494 -9586 42546
rect -9534 42494 -9520 42546
rect -9600 42480 -9520 42494
rect -9440 42546 -9360 42560
rect -9440 42494 -9426 42546
rect -9374 42494 -9360 42546
rect -9440 42480 -9360 42494
rect -9280 42546 -9200 42560
rect -9280 42494 -9266 42546
rect -9214 42494 -9200 42546
rect -9280 42480 -9200 42494
rect -9120 42546 -9040 42560
rect -9120 42494 -9106 42546
rect -9054 42494 -9040 42546
rect -9120 42480 -9040 42494
rect -8960 42546 -8880 42560
rect -8960 42494 -8946 42546
rect -8894 42494 -8880 42546
rect -8960 42480 -8880 42494
rect -8800 42546 -8720 42560
rect -8800 42494 -8786 42546
rect -8734 42494 -8720 42546
rect -8800 42480 -8720 42494
rect -8640 42546 -8560 42560
rect -8640 42494 -8626 42546
rect -8574 42494 -8560 42546
rect -8640 42480 -8560 42494
rect -8480 42546 -8400 42560
rect -8480 42494 -8466 42546
rect -8414 42494 -8400 42546
rect -8480 42480 -8400 42494
rect -8320 42546 -8240 42560
rect -8320 42494 -8306 42546
rect -8254 42494 -8240 42546
rect -8320 42480 -8240 42494
rect -8160 42546 -8080 42560
rect -8160 42494 -8146 42546
rect -8094 42494 -8080 42546
rect -8160 42480 -8080 42494
rect -8000 42546 -7920 42560
rect -8000 42494 -7986 42546
rect -7934 42494 -7920 42546
rect -8000 42480 -7920 42494
rect -7840 42546 -7760 42560
rect -7840 42494 -7826 42546
rect -7774 42494 -7760 42546
rect -7840 42480 -7760 42494
rect -7680 42546 -7600 42560
rect -7680 42494 -7666 42546
rect -7614 42494 -7600 42546
rect -7680 42480 -7600 42494
rect -7520 42546 -7440 42560
rect -7520 42494 -7506 42546
rect -7454 42494 -7440 42546
rect -7520 42480 -7440 42494
rect -7360 42546 -7280 42560
rect -7360 42494 -7346 42546
rect -7294 42494 -7280 42546
rect -7360 42480 -7280 42494
rect -7200 42546 -7120 42560
rect -7200 42494 -7186 42546
rect -7134 42494 -7120 42546
rect -7200 42480 -7120 42494
rect -7040 42546 -6960 42560
rect -7040 42494 -7026 42546
rect -6974 42494 -6960 42546
rect -7040 42480 -6960 42494
rect -6880 42546 -6800 42560
rect -6880 42494 -6866 42546
rect -6814 42494 -6800 42546
rect -6880 42480 -6800 42494
rect -6720 42546 -6640 42560
rect -6720 42494 -6706 42546
rect -6654 42494 -6640 42546
rect -6720 42480 -6640 42494
rect -6560 42546 -6480 42560
rect -6560 42494 -6546 42546
rect -6494 42494 -6480 42546
rect -6560 42480 -6480 42494
rect -6400 42546 -6320 42560
rect -6400 42494 -6386 42546
rect -6334 42494 -6320 42546
rect -6400 42480 -6320 42494
rect -6240 42546 -6160 42560
rect -6240 42494 -6226 42546
rect -6174 42494 -6160 42546
rect -6240 42480 -6160 42494
rect -6080 42546 -6000 42560
rect -6080 42494 -6066 42546
rect -6014 42494 -6000 42546
rect -6080 42480 -6000 42494
rect -5920 42546 -5840 42560
rect -5920 42494 -5906 42546
rect -5854 42494 -5840 42546
rect -5920 42480 -5840 42494
rect -5760 42546 -5680 42560
rect -5760 42494 -5746 42546
rect -5694 42494 -5680 42546
rect -5760 42480 -5680 42494
rect -5600 42546 -5520 42560
rect -5600 42494 -5586 42546
rect -5534 42494 -5520 42546
rect -5600 42480 -5520 42494
rect -5440 42546 -5360 42560
rect -5440 42494 -5426 42546
rect -5374 42494 -5360 42546
rect -5440 42480 -5360 42494
rect -5280 42546 -5200 42560
rect -5280 42494 -5266 42546
rect -5214 42494 -5200 42546
rect -5280 42480 -5200 42494
rect -5120 42546 -5040 42560
rect -5120 42494 -5106 42546
rect -5054 42494 -5040 42546
rect -5120 42480 -5040 42494
rect -4960 42546 -4880 42560
rect -4960 42494 -4946 42546
rect -4894 42494 -4880 42546
rect -4960 42480 -4880 42494
rect -4800 42546 -4720 42560
rect -4800 42494 -4786 42546
rect -4734 42494 -4720 42546
rect -4800 42480 -4720 42494
rect -4640 42546 -4560 42560
rect -4640 42494 -4626 42546
rect -4574 42494 -4560 42546
rect -4640 42480 -4560 42494
rect -4480 42546 -4400 42560
rect -4480 42494 -4466 42546
rect -4414 42494 -4400 42546
rect -4480 42480 -4400 42494
rect -4320 42546 -4240 42560
rect -4320 42494 -4306 42546
rect -4254 42494 -4240 42546
rect -4320 42480 -4240 42494
rect -4160 42546 -4080 42560
rect -4160 42494 -4146 42546
rect -4094 42494 -4080 42546
rect -4160 42480 -4080 42494
rect -4000 42546 -3920 42560
rect -4000 42494 -3986 42546
rect -3934 42494 -3920 42546
rect -4000 42480 -3920 42494
rect -3680 42546 -3600 42560
rect -3680 42494 -3666 42546
rect -3614 42494 -3600 42546
rect -3680 42480 -3600 42494
rect -3520 42546 -3440 42560
rect -3520 42494 -3506 42546
rect -3454 42494 -3440 42546
rect -3520 42480 -3440 42494
rect -3360 42546 -3280 42560
rect -3360 42494 -3346 42546
rect -3294 42494 -3280 42546
rect -3360 42480 -3280 42494
rect -3040 42546 -2960 42560
rect -3040 42494 -3026 42546
rect -2974 42494 -2960 42546
rect -3040 42480 -2960 42494
rect -2720 42546 -2640 42560
rect -2720 42494 -2706 42546
rect -2654 42494 -2640 42546
rect -2720 42480 -2640 42494
rect -2560 42546 -2480 42560
rect -2560 42494 -2546 42546
rect -2494 42494 -2480 42546
rect -2560 42480 -2480 42494
rect -2400 42546 -2320 42560
rect -2400 42494 -2386 42546
rect -2334 42494 -2320 42546
rect -2400 42480 -2320 42494
rect -2240 42546 -2160 42560
rect -2240 42494 -2226 42546
rect -2174 42494 -2160 42546
rect -2240 42480 -2160 42494
rect -2080 42546 -2000 42560
rect -2080 42494 -2066 42546
rect -2014 42494 -2000 42546
rect -2080 42480 -2000 42494
rect -1760 42546 -1680 42560
rect -1760 42494 -1746 42546
rect -1694 42494 -1680 42546
rect -1760 42480 -1680 42494
rect -1440 42546 -1360 42560
rect -1440 42494 -1426 42546
rect -1374 42494 -1360 42546
rect -1440 42480 -1360 42494
rect -1120 42546 -1040 42560
rect -1120 42494 -1106 42546
rect -1054 42494 -1040 42546
rect -1120 42480 -1040 42494
rect -29920 42226 -29840 42240
rect -29920 42174 -29906 42226
rect -29854 42174 -29840 42226
rect -29920 42160 -29840 42174
rect -29760 42226 -29680 42240
rect -29760 42174 -29746 42226
rect -29694 42174 -29680 42226
rect -29760 42160 -29680 42174
rect -29600 42226 -29520 42240
rect -29600 42174 -29586 42226
rect -29534 42174 -29520 42226
rect -29600 42160 -29520 42174
rect -29440 42226 -29360 42240
rect -29440 42174 -29426 42226
rect -29374 42174 -29360 42226
rect -29440 42160 -29360 42174
rect -29280 42226 -29200 42240
rect -29280 42174 -29266 42226
rect -29214 42174 -29200 42226
rect -29280 42160 -29200 42174
rect -29120 42226 -29040 42240
rect -29120 42174 -29106 42226
rect -29054 42174 -29040 42226
rect -29120 42160 -29040 42174
rect -28960 42226 -28880 42240
rect -28960 42174 -28946 42226
rect -28894 42174 -28880 42226
rect -28960 42160 -28880 42174
rect -28800 42226 -28720 42240
rect -28800 42174 -28786 42226
rect -28734 42174 -28720 42226
rect -28800 42160 -28720 42174
rect -28640 42226 -28560 42240
rect -28640 42174 -28626 42226
rect -28574 42174 -28560 42226
rect -28640 42160 -28560 42174
rect -28480 42226 -28400 42240
rect -28480 42174 -28466 42226
rect -28414 42174 -28400 42226
rect -28480 42160 -28400 42174
rect -28320 42226 -28240 42240
rect -28320 42174 -28306 42226
rect -28254 42174 -28240 42226
rect -28320 42160 -28240 42174
rect -28160 42226 -28080 42240
rect -28160 42174 -28146 42226
rect -28094 42174 -28080 42226
rect -28160 42160 -28080 42174
rect -28000 42226 -27920 42240
rect -28000 42174 -27986 42226
rect -27934 42174 -27920 42226
rect -28000 42160 -27920 42174
rect -27840 42226 -27760 42240
rect -27840 42174 -27826 42226
rect -27774 42174 -27760 42226
rect -27840 42160 -27760 42174
rect -27680 42226 -27600 42240
rect -27680 42174 -27666 42226
rect -27614 42174 -27600 42226
rect -27680 42160 -27600 42174
rect -27520 42226 -27440 42240
rect -27520 42174 -27506 42226
rect -27454 42174 -27440 42226
rect -27520 42160 -27440 42174
rect -27360 42226 -27280 42240
rect -27360 42174 -27346 42226
rect -27294 42174 -27280 42226
rect -27360 42160 -27280 42174
rect -27200 42226 -27120 42240
rect -27200 42174 -27186 42226
rect -27134 42174 -27120 42226
rect -27200 42160 -27120 42174
rect -27040 42226 -26960 42240
rect -27040 42174 -27026 42226
rect -26974 42174 -26960 42226
rect -27040 42160 -26960 42174
rect -26880 42226 -26800 42240
rect -26880 42174 -26866 42226
rect -26814 42174 -26800 42226
rect -26880 42160 -26800 42174
rect -26720 42226 -26640 42240
rect -26720 42174 -26706 42226
rect -26654 42174 -26640 42226
rect -26720 42160 -26640 42174
rect -26560 42226 -26480 42240
rect -26560 42174 -26546 42226
rect -26494 42174 -26480 42226
rect -26560 42160 -26480 42174
rect -26400 42226 -26320 42240
rect -26400 42174 -26386 42226
rect -26334 42174 -26320 42226
rect -26400 42160 -26320 42174
rect -26240 42226 -26160 42240
rect -26240 42174 -26226 42226
rect -26174 42174 -26160 42226
rect -26240 42160 -26160 42174
rect -26080 42226 -26000 42240
rect -26080 42174 -26066 42226
rect -26014 42174 -26000 42226
rect -26080 42160 -26000 42174
rect -25920 42226 -25840 42240
rect -25920 42174 -25906 42226
rect -25854 42174 -25840 42226
rect -25920 42160 -25840 42174
rect -25760 42226 -25680 42240
rect -25760 42174 -25746 42226
rect -25694 42174 -25680 42226
rect -25760 42160 -25680 42174
rect -25600 42226 -25520 42240
rect -25600 42174 -25586 42226
rect -25534 42174 -25520 42226
rect -25600 42160 -25520 42174
rect -25440 42226 -25360 42240
rect -25440 42174 -25426 42226
rect -25374 42174 -25360 42226
rect -25440 42160 -25360 42174
rect -25280 42226 -25200 42240
rect -25280 42174 -25266 42226
rect -25214 42174 -25200 42226
rect -25280 42160 -25200 42174
rect -25120 42226 -25040 42240
rect -25120 42174 -25106 42226
rect -25054 42174 -25040 42226
rect -25120 42160 -25040 42174
rect -24960 42226 -24880 42240
rect -24960 42174 -24946 42226
rect -24894 42174 -24880 42226
rect -24960 42160 -24880 42174
rect -24800 42226 -24720 42240
rect -24800 42174 -24786 42226
rect -24734 42174 -24720 42226
rect -24800 42160 -24720 42174
rect -24640 42226 -24560 42240
rect -24640 42174 -24626 42226
rect -24574 42174 -24560 42226
rect -24640 42160 -24560 42174
rect -24480 42226 -24400 42240
rect -24480 42174 -24466 42226
rect -24414 42174 -24400 42226
rect -24480 42160 -24400 42174
rect -24320 42226 -24240 42240
rect -24320 42174 -24306 42226
rect -24254 42174 -24240 42226
rect -24320 42160 -24240 42174
rect -24160 42226 -24080 42240
rect -24160 42174 -24146 42226
rect -24094 42174 -24080 42226
rect -24160 42160 -24080 42174
rect -24000 42226 -23920 42240
rect -24000 42174 -23986 42226
rect -23934 42174 -23920 42226
rect -24000 42160 -23920 42174
rect -23840 42226 -23760 42240
rect -23840 42174 -23826 42226
rect -23774 42174 -23760 42226
rect -23840 42160 -23760 42174
rect -23680 42226 -23600 42240
rect -23680 42174 -23666 42226
rect -23614 42174 -23600 42226
rect -23680 42160 -23600 42174
rect -23520 42226 -23440 42240
rect -23520 42174 -23506 42226
rect -23454 42174 -23440 42226
rect -23520 42160 -23440 42174
rect -23360 42226 -23280 42240
rect -23360 42174 -23346 42226
rect -23294 42174 -23280 42226
rect -23360 42160 -23280 42174
rect -23200 42226 -23120 42240
rect -23200 42174 -23186 42226
rect -23134 42174 -23120 42226
rect -23200 42160 -23120 42174
rect -23040 42226 -22960 42240
rect -23040 42174 -23026 42226
rect -22974 42174 -22960 42226
rect -23040 42160 -22960 42174
rect -22880 42226 -22800 42240
rect -22880 42174 -22866 42226
rect -22814 42174 -22800 42226
rect -22880 42160 -22800 42174
rect -22720 42226 -22640 42240
rect -22720 42174 -22706 42226
rect -22654 42174 -22640 42226
rect -22720 42160 -22640 42174
rect -22560 42226 -22480 42240
rect -22560 42174 -22546 42226
rect -22494 42174 -22480 42226
rect -22560 42160 -22480 42174
rect -22400 42226 -22320 42240
rect -22400 42174 -22386 42226
rect -22334 42174 -22320 42226
rect -22400 42160 -22320 42174
rect -22240 42226 -22160 42240
rect -22240 42174 -22226 42226
rect -22174 42174 -22160 42226
rect -22240 42160 -22160 42174
rect -22080 42226 -22000 42240
rect -22080 42174 -22066 42226
rect -22014 42174 -22000 42226
rect -22080 42160 -22000 42174
rect -21920 42226 -21840 42240
rect -21920 42174 -21906 42226
rect -21854 42174 -21840 42226
rect -21920 42160 -21840 42174
rect -21760 42226 -21680 42240
rect -21760 42174 -21746 42226
rect -21694 42174 -21680 42226
rect -21760 42160 -21680 42174
rect -21600 42226 -21520 42240
rect -21600 42174 -21586 42226
rect -21534 42174 -21520 42226
rect -21600 42160 -21520 42174
rect -21440 42226 -21360 42240
rect -21440 42174 -21426 42226
rect -21374 42174 -21360 42226
rect -21440 42160 -21360 42174
rect -21280 42226 -21200 42240
rect -21280 42174 -21266 42226
rect -21214 42174 -21200 42226
rect -21280 42160 -21200 42174
rect -21120 42226 -21040 42240
rect -21120 42174 -21106 42226
rect -21054 42174 -21040 42226
rect -21120 42160 -21040 42174
rect -20960 42226 -20880 42240
rect -20960 42174 -20946 42226
rect -20894 42174 -20880 42226
rect -20960 42160 -20880 42174
rect -20800 42226 -20720 42240
rect -20800 42174 -20786 42226
rect -20734 42174 -20720 42226
rect -20800 42160 -20720 42174
rect -20640 42226 -20560 42240
rect -20640 42174 -20626 42226
rect -20574 42174 -20560 42226
rect -20640 42160 -20560 42174
rect -20480 42226 -20400 42240
rect -20480 42174 -20466 42226
rect -20414 42174 -20400 42226
rect -20480 42160 -20400 42174
rect -20320 42226 -20240 42240
rect -20320 42174 -20306 42226
rect -20254 42174 -20240 42226
rect -20320 42160 -20240 42174
rect -20160 42226 -20080 42240
rect -20160 42174 -20146 42226
rect -20094 42174 -20080 42226
rect -20160 42160 -20080 42174
rect -20000 42226 -19920 42240
rect -20000 42174 -19986 42226
rect -19934 42174 -19920 42226
rect -20000 42160 -19920 42174
rect -19840 42226 -19760 42240
rect -19840 42174 -19826 42226
rect -19774 42174 -19760 42226
rect -19840 42160 -19760 42174
rect -19680 42226 -19600 42240
rect -19680 42174 -19666 42226
rect -19614 42174 -19600 42226
rect -19680 42160 -19600 42174
rect -19520 42226 -19440 42240
rect -19520 42174 -19506 42226
rect -19454 42174 -19440 42226
rect -19520 42160 -19440 42174
rect -19360 42226 -19280 42240
rect -19360 42174 -19346 42226
rect -19294 42174 -19280 42226
rect -19360 42160 -19280 42174
rect -19200 42226 -19120 42240
rect -19200 42174 -19186 42226
rect -19134 42174 -19120 42226
rect -19200 42160 -19120 42174
rect -19040 42226 -18960 42240
rect -19040 42174 -19026 42226
rect -18974 42174 -18960 42226
rect -19040 42160 -18960 42174
rect -18880 42226 -18800 42240
rect -18880 42174 -18866 42226
rect -18814 42174 -18800 42226
rect -18880 42160 -18800 42174
rect -18720 42226 -18640 42240
rect -18720 42174 -18706 42226
rect -18654 42174 -18640 42226
rect -18720 42160 -18640 42174
rect -18560 42226 -18480 42240
rect -18560 42174 -18546 42226
rect -18494 42174 -18480 42226
rect -18560 42160 -18480 42174
rect -18400 42226 -18320 42240
rect -18400 42174 -18386 42226
rect -18334 42174 -18320 42226
rect -18400 42160 -18320 42174
rect -18240 42226 -18160 42240
rect -18240 42174 -18226 42226
rect -18174 42174 -18160 42226
rect -18240 42160 -18160 42174
rect -18080 42226 -18000 42240
rect -18080 42174 -18066 42226
rect -18014 42174 -18000 42226
rect -18080 42160 -18000 42174
rect -17920 42226 -17840 42240
rect -17920 42174 -17906 42226
rect -17854 42174 -17840 42226
rect -17920 42160 -17840 42174
rect -17760 42226 -17680 42240
rect -17760 42174 -17746 42226
rect -17694 42174 -17680 42226
rect -17760 42160 -17680 42174
rect -17600 42226 -17520 42240
rect -17600 42174 -17586 42226
rect -17534 42174 -17520 42226
rect -17600 42160 -17520 42174
rect -17440 42226 -17360 42240
rect -17440 42174 -17426 42226
rect -17374 42174 -17360 42226
rect -17440 42160 -17360 42174
rect -17280 42226 -17200 42240
rect -17280 42174 -17266 42226
rect -17214 42174 -17200 42226
rect -17280 42160 -17200 42174
rect -17120 42226 -17040 42240
rect -17120 42174 -17106 42226
rect -17054 42174 -17040 42226
rect -17120 42160 -17040 42174
rect -16960 42226 -16880 42240
rect -16960 42174 -16946 42226
rect -16894 42174 -16880 42226
rect -16960 42160 -16880 42174
rect -16800 42226 -16720 42240
rect -16800 42174 -16786 42226
rect -16734 42174 -16720 42226
rect -16800 42160 -16720 42174
rect -16640 42226 -16560 42240
rect -16640 42174 -16626 42226
rect -16574 42174 -16560 42226
rect -16640 42160 -16560 42174
rect -16480 42226 -16400 42240
rect -16480 42174 -16466 42226
rect -16414 42174 -16400 42226
rect -16480 42160 -16400 42174
rect -16320 42226 -16240 42240
rect -16320 42174 -16306 42226
rect -16254 42174 -16240 42226
rect -16320 42160 -16240 42174
rect -16160 42226 -16080 42240
rect -16160 42174 -16146 42226
rect -16094 42174 -16080 42226
rect -16160 42160 -16080 42174
rect -16000 42226 -15920 42240
rect -16000 42174 -15986 42226
rect -15934 42174 -15920 42226
rect -16000 42160 -15920 42174
rect -15840 42226 -15760 42240
rect -15840 42174 -15826 42226
rect -15774 42174 -15760 42226
rect -15840 42160 -15760 42174
rect -15680 42226 -15600 42240
rect -15680 42174 -15666 42226
rect -15614 42174 -15600 42226
rect -15680 42160 -15600 42174
rect -15520 42226 -15440 42240
rect -15520 42174 -15506 42226
rect -15454 42174 -15440 42226
rect -15520 42160 -15440 42174
rect -15360 42226 -15280 42240
rect -15360 42174 -15346 42226
rect -15294 42174 -15280 42226
rect -15360 42160 -15280 42174
rect -15200 42226 -15120 42240
rect -15200 42174 -15186 42226
rect -15134 42174 -15120 42226
rect -15200 42160 -15120 42174
rect -15040 42226 -14960 42240
rect -15040 42174 -15026 42226
rect -14974 42174 -14960 42226
rect -15040 42160 -14960 42174
rect -14880 42226 -14800 42240
rect -14880 42174 -14866 42226
rect -14814 42174 -14800 42226
rect -14880 42160 -14800 42174
rect -14720 42226 -14640 42240
rect -14720 42174 -14706 42226
rect -14654 42174 -14640 42226
rect -14720 42160 -14640 42174
rect -14560 42226 -14480 42240
rect -14560 42174 -14546 42226
rect -14494 42174 -14480 42226
rect -14560 42160 -14480 42174
rect -14400 42226 -14320 42240
rect -14400 42174 -14386 42226
rect -14334 42174 -14320 42226
rect -14400 42160 -14320 42174
rect -14240 42226 -14160 42240
rect -14240 42174 -14226 42226
rect -14174 42174 -14160 42226
rect -14240 42160 -14160 42174
rect -14080 42226 -14000 42240
rect -14080 42174 -14066 42226
rect -14014 42174 -14000 42226
rect -14080 42160 -14000 42174
rect -13920 42226 -13840 42240
rect -13920 42174 -13906 42226
rect -13854 42174 -13840 42226
rect -13920 42160 -13840 42174
rect -13760 42226 -13680 42240
rect -13760 42174 -13746 42226
rect -13694 42174 -13680 42226
rect -13760 42160 -13680 42174
rect -13600 42226 -13520 42240
rect -13600 42174 -13586 42226
rect -13534 42174 -13520 42226
rect -13600 42160 -13520 42174
rect -13440 42226 -13360 42240
rect -13440 42174 -13426 42226
rect -13374 42174 -13360 42226
rect -13440 42160 -13360 42174
rect -13280 42226 -13200 42240
rect -13280 42174 -13266 42226
rect -13214 42174 -13200 42226
rect -13280 42160 -13200 42174
rect -13120 42226 -13040 42240
rect -13120 42174 -13106 42226
rect -13054 42174 -13040 42226
rect -13120 42160 -13040 42174
rect -12960 42226 -12880 42240
rect -12960 42174 -12946 42226
rect -12894 42174 -12880 42226
rect -12960 42160 -12880 42174
rect -12800 42226 -12720 42240
rect -12800 42174 -12786 42226
rect -12734 42174 -12720 42226
rect -12800 42160 -12720 42174
rect -12640 42226 -12560 42240
rect -12640 42174 -12626 42226
rect -12574 42174 -12560 42226
rect -12640 42160 -12560 42174
rect -12480 42226 -12400 42240
rect -12480 42174 -12466 42226
rect -12414 42174 -12400 42226
rect -12480 42160 -12400 42174
rect -12320 42226 -12240 42240
rect -12320 42174 -12306 42226
rect -12254 42174 -12240 42226
rect -12320 42160 -12240 42174
rect -11360 42226 -11280 42240
rect -11360 42174 -11346 42226
rect -11294 42174 -11280 42226
rect -11360 42160 -11280 42174
rect -11200 42226 -11120 42240
rect -11200 42174 -11186 42226
rect -11134 42174 -11120 42226
rect -11200 42160 -11120 42174
rect -11040 42226 -10960 42240
rect -11040 42174 -11026 42226
rect -10974 42174 -10960 42226
rect -11040 42160 -10960 42174
rect -10880 42226 -10800 42240
rect -10880 42174 -10866 42226
rect -10814 42174 -10800 42226
rect -10880 42160 -10800 42174
rect -10720 42226 -10640 42240
rect -10720 42174 -10706 42226
rect -10654 42174 -10640 42226
rect -10720 42160 -10640 42174
rect -10560 42226 -10480 42240
rect -10560 42174 -10546 42226
rect -10494 42174 -10480 42226
rect -10560 42160 -10480 42174
rect -10400 42226 -10320 42240
rect -10400 42174 -10386 42226
rect -10334 42174 -10320 42226
rect -10400 42160 -10320 42174
rect -10240 42226 -10160 42240
rect -10240 42174 -10226 42226
rect -10174 42174 -10160 42226
rect -10240 42160 -10160 42174
rect -10080 42226 -10000 42240
rect -10080 42174 -10066 42226
rect -10014 42174 -10000 42226
rect -10080 42160 -10000 42174
rect -9920 42226 -9840 42240
rect -9920 42174 -9906 42226
rect -9854 42174 -9840 42226
rect -9920 42160 -9840 42174
rect -9760 42226 -9680 42240
rect -9760 42174 -9746 42226
rect -9694 42174 -9680 42226
rect -9760 42160 -9680 42174
rect -9600 42226 -9520 42240
rect -9600 42174 -9586 42226
rect -9534 42174 -9520 42226
rect -9600 42160 -9520 42174
rect -9440 42226 -9360 42240
rect -9440 42174 -9426 42226
rect -9374 42174 -9360 42226
rect -9440 42160 -9360 42174
rect -9280 42226 -9200 42240
rect -9280 42174 -9266 42226
rect -9214 42174 -9200 42226
rect -9280 42160 -9200 42174
rect -9120 42226 -9040 42240
rect -9120 42174 -9106 42226
rect -9054 42174 -9040 42226
rect -9120 42160 -9040 42174
rect -8960 42226 -8880 42240
rect -8960 42174 -8946 42226
rect -8894 42174 -8880 42226
rect -8960 42160 -8880 42174
rect -8800 42226 -8720 42240
rect -8800 42174 -8786 42226
rect -8734 42174 -8720 42226
rect -8800 42160 -8720 42174
rect -8640 42226 -8560 42240
rect -8640 42174 -8626 42226
rect -8574 42174 -8560 42226
rect -8640 42160 -8560 42174
rect -8480 42226 -8400 42240
rect -8480 42174 -8466 42226
rect -8414 42174 -8400 42226
rect -8480 42160 -8400 42174
rect -8320 42226 -8240 42240
rect -8320 42174 -8306 42226
rect -8254 42174 -8240 42226
rect -8320 42160 -8240 42174
rect -8160 42226 -8080 42240
rect -8160 42174 -8146 42226
rect -8094 42174 -8080 42226
rect -8160 42160 -8080 42174
rect -8000 42226 -7920 42240
rect -8000 42174 -7986 42226
rect -7934 42174 -7920 42226
rect -8000 42160 -7920 42174
rect -7840 42226 -7760 42240
rect -7840 42174 -7826 42226
rect -7774 42174 -7760 42226
rect -7840 42160 -7760 42174
rect -7680 42226 -7600 42240
rect -7680 42174 -7666 42226
rect -7614 42174 -7600 42226
rect -7680 42160 -7600 42174
rect -7520 42226 -7440 42240
rect -7520 42174 -7506 42226
rect -7454 42174 -7440 42226
rect -7520 42160 -7440 42174
rect -7360 42226 -7280 42240
rect -7360 42174 -7346 42226
rect -7294 42174 -7280 42226
rect -7360 42160 -7280 42174
rect -7200 42226 -7120 42240
rect -7200 42174 -7186 42226
rect -7134 42174 -7120 42226
rect -7200 42160 -7120 42174
rect -7040 42226 -6960 42240
rect -7040 42174 -7026 42226
rect -6974 42174 -6960 42226
rect -7040 42160 -6960 42174
rect -6880 42226 -6800 42240
rect -6880 42174 -6866 42226
rect -6814 42174 -6800 42226
rect -6880 42160 -6800 42174
rect -6720 42226 -6640 42240
rect -6720 42174 -6706 42226
rect -6654 42174 -6640 42226
rect -6720 42160 -6640 42174
rect -6560 42226 -6480 42240
rect -6560 42174 -6546 42226
rect -6494 42174 -6480 42226
rect -6560 42160 -6480 42174
rect -6400 42226 -6320 42240
rect -6400 42174 -6386 42226
rect -6334 42174 -6320 42226
rect -6400 42160 -6320 42174
rect -6240 42226 -6160 42240
rect -6240 42174 -6226 42226
rect -6174 42174 -6160 42226
rect -6240 42160 -6160 42174
rect -6080 42226 -6000 42240
rect -6080 42174 -6066 42226
rect -6014 42174 -6000 42226
rect -6080 42160 -6000 42174
rect -5920 42226 -5840 42240
rect -5920 42174 -5906 42226
rect -5854 42174 -5840 42226
rect -5920 42160 -5840 42174
rect -5760 42226 -5680 42240
rect -5760 42174 -5746 42226
rect -5694 42174 -5680 42226
rect -5760 42160 -5680 42174
rect -5600 42226 -5520 42240
rect -5600 42174 -5586 42226
rect -5534 42174 -5520 42226
rect -5600 42160 -5520 42174
rect -5440 42226 -5360 42240
rect -5440 42174 -5426 42226
rect -5374 42174 -5360 42226
rect -5440 42160 -5360 42174
rect -5280 42226 -5200 42240
rect -5280 42174 -5266 42226
rect -5214 42174 -5200 42226
rect -5280 42160 -5200 42174
rect -5120 42226 -5040 42240
rect -5120 42174 -5106 42226
rect -5054 42174 -5040 42226
rect -5120 42160 -5040 42174
rect -4960 42226 -4880 42240
rect -4960 42174 -4946 42226
rect -4894 42174 -4880 42226
rect -4960 42160 -4880 42174
rect -4800 42226 -4720 42240
rect -4800 42174 -4786 42226
rect -4734 42174 -4720 42226
rect -4800 42160 -4720 42174
rect -4640 42226 -4560 42240
rect -4640 42174 -4626 42226
rect -4574 42174 -4560 42226
rect -4640 42160 -4560 42174
rect -4480 42226 -4400 42240
rect -4480 42174 -4466 42226
rect -4414 42174 -4400 42226
rect -4480 42160 -4400 42174
rect -4320 42226 -4240 42240
rect -4320 42174 -4306 42226
rect -4254 42174 -4240 42226
rect -4320 42160 -4240 42174
rect -4160 42226 -4080 42240
rect -4160 42174 -4146 42226
rect -4094 42174 -4080 42226
rect -4160 42160 -4080 42174
rect -4000 42226 -3920 42240
rect -4000 42174 -3986 42226
rect -3934 42174 -3920 42226
rect -4000 42160 -3920 42174
rect -3680 42226 -3600 42240
rect -3680 42174 -3666 42226
rect -3614 42174 -3600 42226
rect -3680 42160 -3600 42174
rect -3520 42226 -3440 42240
rect -3520 42174 -3506 42226
rect -3454 42174 -3440 42226
rect -3520 42160 -3440 42174
rect -3360 42226 -3280 42240
rect -3360 42174 -3346 42226
rect -3294 42174 -3280 42226
rect -3360 42160 -3280 42174
rect -3040 42226 -2960 42240
rect -3040 42174 -3026 42226
rect -2974 42174 -2960 42226
rect -3040 42160 -2960 42174
rect -2720 42226 -2640 42240
rect -2720 42174 -2706 42226
rect -2654 42174 -2640 42226
rect -2720 42160 -2640 42174
rect -2560 42226 -2480 42240
rect -2560 42174 -2546 42226
rect -2494 42174 -2480 42226
rect -2560 42160 -2480 42174
rect -2400 42226 -2320 42240
rect -2400 42174 -2386 42226
rect -2334 42174 -2320 42226
rect -2400 42160 -2320 42174
rect -2240 42226 -2160 42240
rect -2240 42174 -2226 42226
rect -2174 42174 -2160 42226
rect -2240 42160 -2160 42174
rect -2080 42226 -2000 42240
rect -2080 42174 -2066 42226
rect -2014 42174 -2000 42226
rect -2080 42160 -2000 42174
rect -1760 42226 -1680 42240
rect -1760 42174 -1746 42226
rect -1694 42174 -1680 42226
rect -1760 42160 -1680 42174
rect -1440 42226 -1360 42240
rect -1440 42174 -1426 42226
rect -1374 42174 -1360 42226
rect -1440 42160 -1360 42174
rect -1120 42226 -1040 42240
rect -1120 42174 -1106 42226
rect -1054 42174 -1040 42226
rect -1120 42160 -1040 42174
rect -29920 41906 -29840 41920
rect -29920 41854 -29906 41906
rect -29854 41854 -29840 41906
rect -29920 41840 -29840 41854
rect -29760 41906 -29680 41920
rect -29760 41854 -29746 41906
rect -29694 41854 -29680 41906
rect -29760 41840 -29680 41854
rect -29600 41906 -29520 41920
rect -29600 41854 -29586 41906
rect -29534 41854 -29520 41906
rect -29600 41840 -29520 41854
rect -29440 41906 -29360 41920
rect -29440 41854 -29426 41906
rect -29374 41854 -29360 41906
rect -29440 41840 -29360 41854
rect -29280 41906 -29200 41920
rect -29280 41854 -29266 41906
rect -29214 41854 -29200 41906
rect -29280 41840 -29200 41854
rect -29120 41906 -29040 41920
rect -29120 41854 -29106 41906
rect -29054 41854 -29040 41906
rect -29120 41840 -29040 41854
rect -28960 41906 -28880 41920
rect -28960 41854 -28946 41906
rect -28894 41854 -28880 41906
rect -28960 41840 -28880 41854
rect -28800 41906 -28720 41920
rect -28800 41854 -28786 41906
rect -28734 41854 -28720 41906
rect -28800 41840 -28720 41854
rect -28640 41906 -28560 41920
rect -28640 41854 -28626 41906
rect -28574 41854 -28560 41906
rect -28640 41840 -28560 41854
rect -28480 41906 -28400 41920
rect -28480 41854 -28466 41906
rect -28414 41854 -28400 41906
rect -28480 41840 -28400 41854
rect -28320 41906 -28240 41920
rect -28320 41854 -28306 41906
rect -28254 41854 -28240 41906
rect -28320 41840 -28240 41854
rect -28160 41906 -28080 41920
rect -28160 41854 -28146 41906
rect -28094 41854 -28080 41906
rect -28160 41840 -28080 41854
rect -28000 41906 -27920 41920
rect -28000 41854 -27986 41906
rect -27934 41854 -27920 41906
rect -28000 41840 -27920 41854
rect -27840 41906 -27760 41920
rect -27840 41854 -27826 41906
rect -27774 41854 -27760 41906
rect -27840 41840 -27760 41854
rect -27680 41906 -27600 41920
rect -27680 41854 -27666 41906
rect -27614 41854 -27600 41906
rect -27680 41840 -27600 41854
rect -27520 41906 -27440 41920
rect -27520 41854 -27506 41906
rect -27454 41854 -27440 41906
rect -27520 41840 -27440 41854
rect -27360 41906 -27280 41920
rect -27360 41854 -27346 41906
rect -27294 41854 -27280 41906
rect -27360 41840 -27280 41854
rect -27200 41906 -27120 41920
rect -27200 41854 -27186 41906
rect -27134 41854 -27120 41906
rect -27200 41840 -27120 41854
rect -27040 41906 -26960 41920
rect -27040 41854 -27026 41906
rect -26974 41854 -26960 41906
rect -27040 41840 -26960 41854
rect -26880 41906 -26800 41920
rect -26880 41854 -26866 41906
rect -26814 41854 -26800 41906
rect -26880 41840 -26800 41854
rect -26720 41906 -26640 41920
rect -26720 41854 -26706 41906
rect -26654 41854 -26640 41906
rect -26720 41840 -26640 41854
rect -26560 41906 -26480 41920
rect -26560 41854 -26546 41906
rect -26494 41854 -26480 41906
rect -26560 41840 -26480 41854
rect -26400 41906 -26320 41920
rect -26400 41854 -26386 41906
rect -26334 41854 -26320 41906
rect -26400 41840 -26320 41854
rect -26240 41906 -26160 41920
rect -26240 41854 -26226 41906
rect -26174 41854 -26160 41906
rect -26240 41840 -26160 41854
rect -26080 41906 -26000 41920
rect -26080 41854 -26066 41906
rect -26014 41854 -26000 41906
rect -26080 41840 -26000 41854
rect -25920 41906 -25840 41920
rect -25920 41854 -25906 41906
rect -25854 41854 -25840 41906
rect -25920 41840 -25840 41854
rect -25760 41906 -25680 41920
rect -25760 41854 -25746 41906
rect -25694 41854 -25680 41906
rect -25760 41840 -25680 41854
rect -25600 41906 -25520 41920
rect -25600 41854 -25586 41906
rect -25534 41854 -25520 41906
rect -25600 41840 -25520 41854
rect -25440 41906 -25360 41920
rect -25440 41854 -25426 41906
rect -25374 41854 -25360 41906
rect -25440 41840 -25360 41854
rect -25280 41906 -25200 41920
rect -25280 41854 -25266 41906
rect -25214 41854 -25200 41906
rect -25280 41840 -25200 41854
rect -25120 41906 -25040 41920
rect -25120 41854 -25106 41906
rect -25054 41854 -25040 41906
rect -25120 41840 -25040 41854
rect -24960 41906 -24880 41920
rect -24960 41854 -24946 41906
rect -24894 41854 -24880 41906
rect -24960 41840 -24880 41854
rect -24800 41906 -24720 41920
rect -24800 41854 -24786 41906
rect -24734 41854 -24720 41906
rect -24800 41840 -24720 41854
rect -24640 41906 -24560 41920
rect -24640 41854 -24626 41906
rect -24574 41854 -24560 41906
rect -24640 41840 -24560 41854
rect -24480 41906 -24400 41920
rect -24480 41854 -24466 41906
rect -24414 41854 -24400 41906
rect -24480 41840 -24400 41854
rect -24320 41906 -24240 41920
rect -24320 41854 -24306 41906
rect -24254 41854 -24240 41906
rect -24320 41840 -24240 41854
rect -24160 41906 -24080 41920
rect -24160 41854 -24146 41906
rect -24094 41854 -24080 41906
rect -24160 41840 -24080 41854
rect -24000 41906 -23920 41920
rect -24000 41854 -23986 41906
rect -23934 41854 -23920 41906
rect -24000 41840 -23920 41854
rect -23840 41906 -23760 41920
rect -23840 41854 -23826 41906
rect -23774 41854 -23760 41906
rect -23840 41840 -23760 41854
rect -23680 41906 -23600 41920
rect -23680 41854 -23666 41906
rect -23614 41854 -23600 41906
rect -23680 41840 -23600 41854
rect -23520 41906 -23440 41920
rect -23520 41854 -23506 41906
rect -23454 41854 -23440 41906
rect -23520 41840 -23440 41854
rect -23360 41906 -23280 41920
rect -23360 41854 -23346 41906
rect -23294 41854 -23280 41906
rect -23360 41840 -23280 41854
rect -23200 41906 -23120 41920
rect -23200 41854 -23186 41906
rect -23134 41854 -23120 41906
rect -23200 41840 -23120 41854
rect -23040 41906 -22960 41920
rect -23040 41854 -23026 41906
rect -22974 41854 -22960 41906
rect -23040 41840 -22960 41854
rect -22880 41906 -22800 41920
rect -22880 41854 -22866 41906
rect -22814 41854 -22800 41906
rect -22880 41840 -22800 41854
rect -22720 41906 -22640 41920
rect -22720 41854 -22706 41906
rect -22654 41854 -22640 41906
rect -22720 41840 -22640 41854
rect -22560 41906 -22480 41920
rect -22560 41854 -22546 41906
rect -22494 41854 -22480 41906
rect -22560 41840 -22480 41854
rect -22400 41906 -22320 41920
rect -22400 41854 -22386 41906
rect -22334 41854 -22320 41906
rect -22400 41840 -22320 41854
rect -22240 41906 -22160 41920
rect -22240 41854 -22226 41906
rect -22174 41854 -22160 41906
rect -22240 41840 -22160 41854
rect -22080 41906 -22000 41920
rect -22080 41854 -22066 41906
rect -22014 41854 -22000 41906
rect -22080 41840 -22000 41854
rect -21920 41906 -21840 41920
rect -21920 41854 -21906 41906
rect -21854 41854 -21840 41906
rect -21920 41840 -21840 41854
rect -21760 41906 -21680 41920
rect -21760 41854 -21746 41906
rect -21694 41854 -21680 41906
rect -21760 41840 -21680 41854
rect -21600 41906 -21520 41920
rect -21600 41854 -21586 41906
rect -21534 41854 -21520 41906
rect -21600 41840 -21520 41854
rect -21440 41906 -21360 41920
rect -21440 41854 -21426 41906
rect -21374 41854 -21360 41906
rect -21440 41840 -21360 41854
rect -21280 41906 -21200 41920
rect -21280 41854 -21266 41906
rect -21214 41854 -21200 41906
rect -21280 41840 -21200 41854
rect -21120 41906 -21040 41920
rect -21120 41854 -21106 41906
rect -21054 41854 -21040 41906
rect -21120 41840 -21040 41854
rect -20960 41906 -20880 41920
rect -20960 41854 -20946 41906
rect -20894 41854 -20880 41906
rect -20960 41840 -20880 41854
rect -20800 41906 -20720 41920
rect -20800 41854 -20786 41906
rect -20734 41854 -20720 41906
rect -20800 41840 -20720 41854
rect -20640 41906 -20560 41920
rect -20640 41854 -20626 41906
rect -20574 41854 -20560 41906
rect -20640 41840 -20560 41854
rect -20480 41906 -20400 41920
rect -20480 41854 -20466 41906
rect -20414 41854 -20400 41906
rect -20480 41840 -20400 41854
rect -20320 41906 -20240 41920
rect -20320 41854 -20306 41906
rect -20254 41854 -20240 41906
rect -20320 41840 -20240 41854
rect -20160 41906 -20080 41920
rect -20160 41854 -20146 41906
rect -20094 41854 -20080 41906
rect -20160 41840 -20080 41854
rect -20000 41906 -19920 41920
rect -20000 41854 -19986 41906
rect -19934 41854 -19920 41906
rect -20000 41840 -19920 41854
rect -19840 41906 -19760 41920
rect -19840 41854 -19826 41906
rect -19774 41854 -19760 41906
rect -19840 41840 -19760 41854
rect -19680 41906 -19600 41920
rect -19680 41854 -19666 41906
rect -19614 41854 -19600 41906
rect -19680 41840 -19600 41854
rect -19520 41906 -19440 41920
rect -19520 41854 -19506 41906
rect -19454 41854 -19440 41906
rect -19520 41840 -19440 41854
rect -19360 41906 -19280 41920
rect -19360 41854 -19346 41906
rect -19294 41854 -19280 41906
rect -19360 41840 -19280 41854
rect -19200 41906 -19120 41920
rect -19200 41854 -19186 41906
rect -19134 41854 -19120 41906
rect -19200 41840 -19120 41854
rect -19040 41906 -18960 41920
rect -19040 41854 -19026 41906
rect -18974 41854 -18960 41906
rect -19040 41840 -18960 41854
rect -18880 41906 -18800 41920
rect -18880 41854 -18866 41906
rect -18814 41854 -18800 41906
rect -18880 41840 -18800 41854
rect -18720 41906 -18640 41920
rect -18720 41854 -18706 41906
rect -18654 41854 -18640 41906
rect -18720 41840 -18640 41854
rect -18560 41906 -18480 41920
rect -18560 41854 -18546 41906
rect -18494 41854 -18480 41906
rect -18560 41840 -18480 41854
rect -18400 41906 -18320 41920
rect -18400 41854 -18386 41906
rect -18334 41854 -18320 41906
rect -18400 41840 -18320 41854
rect -18240 41906 -18160 41920
rect -18240 41854 -18226 41906
rect -18174 41854 -18160 41906
rect -18240 41840 -18160 41854
rect -18080 41906 -18000 41920
rect -18080 41854 -18066 41906
rect -18014 41854 -18000 41906
rect -18080 41840 -18000 41854
rect -17920 41906 -17840 41920
rect -17920 41854 -17906 41906
rect -17854 41854 -17840 41906
rect -17920 41840 -17840 41854
rect -17760 41906 -17680 41920
rect -17760 41854 -17746 41906
rect -17694 41854 -17680 41906
rect -17760 41840 -17680 41854
rect -17600 41906 -17520 41920
rect -17600 41854 -17586 41906
rect -17534 41854 -17520 41906
rect -17600 41840 -17520 41854
rect -17440 41906 -17360 41920
rect -17440 41854 -17426 41906
rect -17374 41854 -17360 41906
rect -17440 41840 -17360 41854
rect -17280 41906 -17200 41920
rect -17280 41854 -17266 41906
rect -17214 41854 -17200 41906
rect -17280 41840 -17200 41854
rect -17120 41906 -17040 41920
rect -17120 41854 -17106 41906
rect -17054 41854 -17040 41906
rect -17120 41840 -17040 41854
rect -16960 41906 -16880 41920
rect -16960 41854 -16946 41906
rect -16894 41854 -16880 41906
rect -16960 41840 -16880 41854
rect -16800 41906 -16720 41920
rect -16800 41854 -16786 41906
rect -16734 41854 -16720 41906
rect -16800 41840 -16720 41854
rect -16640 41906 -16560 41920
rect -16640 41854 -16626 41906
rect -16574 41854 -16560 41906
rect -16640 41840 -16560 41854
rect -16480 41906 -16400 41920
rect -16480 41854 -16466 41906
rect -16414 41854 -16400 41906
rect -16480 41840 -16400 41854
rect -16320 41906 -16240 41920
rect -16320 41854 -16306 41906
rect -16254 41854 -16240 41906
rect -16320 41840 -16240 41854
rect -16160 41906 -16080 41920
rect -16160 41854 -16146 41906
rect -16094 41854 -16080 41906
rect -16160 41840 -16080 41854
rect -16000 41906 -15920 41920
rect -16000 41854 -15986 41906
rect -15934 41854 -15920 41906
rect -16000 41840 -15920 41854
rect -15840 41906 -15760 41920
rect -15840 41854 -15826 41906
rect -15774 41854 -15760 41906
rect -15840 41840 -15760 41854
rect -15680 41906 -15600 41920
rect -15680 41854 -15666 41906
rect -15614 41854 -15600 41906
rect -15680 41840 -15600 41854
rect -15520 41906 -15440 41920
rect -15520 41854 -15506 41906
rect -15454 41854 -15440 41906
rect -15520 41840 -15440 41854
rect -15360 41906 -15280 41920
rect -15360 41854 -15346 41906
rect -15294 41854 -15280 41906
rect -15360 41840 -15280 41854
rect -15200 41906 -15120 41920
rect -15200 41854 -15186 41906
rect -15134 41854 -15120 41906
rect -15200 41840 -15120 41854
rect -15040 41906 -14960 41920
rect -15040 41854 -15026 41906
rect -14974 41854 -14960 41906
rect -15040 41840 -14960 41854
rect -14880 41906 -14800 41920
rect -14880 41854 -14866 41906
rect -14814 41854 -14800 41906
rect -14880 41840 -14800 41854
rect -14720 41906 -14640 41920
rect -14720 41854 -14706 41906
rect -14654 41854 -14640 41906
rect -14720 41840 -14640 41854
rect -14560 41906 -14480 41920
rect -14560 41854 -14546 41906
rect -14494 41854 -14480 41906
rect -14560 41840 -14480 41854
rect -14400 41906 -14320 41920
rect -14400 41854 -14386 41906
rect -14334 41854 -14320 41906
rect -14400 41840 -14320 41854
rect -14240 41906 -14160 41920
rect -14240 41854 -14226 41906
rect -14174 41854 -14160 41906
rect -14240 41840 -14160 41854
rect -14080 41906 -14000 41920
rect -14080 41854 -14066 41906
rect -14014 41854 -14000 41906
rect -14080 41840 -14000 41854
rect -13920 41906 -13840 41920
rect -13920 41854 -13906 41906
rect -13854 41854 -13840 41906
rect -13920 41840 -13840 41854
rect -13760 41906 -13680 41920
rect -13760 41854 -13746 41906
rect -13694 41854 -13680 41906
rect -13760 41840 -13680 41854
rect -13600 41906 -13520 41920
rect -13600 41854 -13586 41906
rect -13534 41854 -13520 41906
rect -13600 41840 -13520 41854
rect -13440 41906 -13360 41920
rect -13440 41854 -13426 41906
rect -13374 41854 -13360 41906
rect -13440 41840 -13360 41854
rect -13280 41906 -13200 41920
rect -13280 41854 -13266 41906
rect -13214 41854 -13200 41906
rect -13280 41840 -13200 41854
rect -13120 41906 -13040 41920
rect -13120 41854 -13106 41906
rect -13054 41854 -13040 41906
rect -13120 41840 -13040 41854
rect -12960 41906 -12880 41920
rect -12960 41854 -12946 41906
rect -12894 41854 -12880 41906
rect -12960 41840 -12880 41854
rect -12800 41906 -12720 41920
rect -12800 41854 -12786 41906
rect -12734 41854 -12720 41906
rect -12800 41840 -12720 41854
rect -12640 41906 -12560 41920
rect -12640 41854 -12626 41906
rect -12574 41854 -12560 41906
rect -12640 41840 -12560 41854
rect -12480 41906 -12400 41920
rect -12480 41854 -12466 41906
rect -12414 41854 -12400 41906
rect -12480 41840 -12400 41854
rect -12320 41906 -12240 41920
rect -12320 41854 -12306 41906
rect -12254 41854 -12240 41906
rect -12320 41840 -12240 41854
rect -11360 41906 -11280 41920
rect -11360 41854 -11346 41906
rect -11294 41854 -11280 41906
rect -11360 41840 -11280 41854
rect -11200 41906 -11120 41920
rect -11200 41854 -11186 41906
rect -11134 41854 -11120 41906
rect -11200 41840 -11120 41854
rect -11040 41906 -10960 41920
rect -11040 41854 -11026 41906
rect -10974 41854 -10960 41906
rect -11040 41840 -10960 41854
rect -10880 41906 -10800 41920
rect -10880 41854 -10866 41906
rect -10814 41854 -10800 41906
rect -10880 41840 -10800 41854
rect -10720 41906 -10640 41920
rect -10720 41854 -10706 41906
rect -10654 41854 -10640 41906
rect -10720 41840 -10640 41854
rect -10560 41906 -10480 41920
rect -10560 41854 -10546 41906
rect -10494 41854 -10480 41906
rect -10560 41840 -10480 41854
rect -10400 41906 -10320 41920
rect -10400 41854 -10386 41906
rect -10334 41854 -10320 41906
rect -10400 41840 -10320 41854
rect -10240 41906 -10160 41920
rect -10240 41854 -10226 41906
rect -10174 41854 -10160 41906
rect -10240 41840 -10160 41854
rect -10080 41906 -10000 41920
rect -10080 41854 -10066 41906
rect -10014 41854 -10000 41906
rect -10080 41840 -10000 41854
rect -9920 41906 -9840 41920
rect -9920 41854 -9906 41906
rect -9854 41854 -9840 41906
rect -9920 41840 -9840 41854
rect -9760 41906 -9680 41920
rect -9760 41854 -9746 41906
rect -9694 41854 -9680 41906
rect -9760 41840 -9680 41854
rect -9600 41906 -9520 41920
rect -9600 41854 -9586 41906
rect -9534 41854 -9520 41906
rect -9600 41840 -9520 41854
rect -9440 41906 -9360 41920
rect -9440 41854 -9426 41906
rect -9374 41854 -9360 41906
rect -9440 41840 -9360 41854
rect -9280 41906 -9200 41920
rect -9280 41854 -9266 41906
rect -9214 41854 -9200 41906
rect -9280 41840 -9200 41854
rect -9120 41906 -9040 41920
rect -9120 41854 -9106 41906
rect -9054 41854 -9040 41906
rect -9120 41840 -9040 41854
rect -8960 41906 -8880 41920
rect -8960 41854 -8946 41906
rect -8894 41854 -8880 41906
rect -8960 41840 -8880 41854
rect -8800 41906 -8720 41920
rect -8800 41854 -8786 41906
rect -8734 41854 -8720 41906
rect -8800 41840 -8720 41854
rect -8640 41906 -8560 41920
rect -8640 41854 -8626 41906
rect -8574 41854 -8560 41906
rect -8640 41840 -8560 41854
rect -8480 41906 -8400 41920
rect -8480 41854 -8466 41906
rect -8414 41854 -8400 41906
rect -8480 41840 -8400 41854
rect -8320 41906 -8240 41920
rect -8320 41854 -8306 41906
rect -8254 41854 -8240 41906
rect -8320 41840 -8240 41854
rect -8160 41906 -8080 41920
rect -8160 41854 -8146 41906
rect -8094 41854 -8080 41906
rect -8160 41840 -8080 41854
rect -8000 41906 -7920 41920
rect -8000 41854 -7986 41906
rect -7934 41854 -7920 41906
rect -8000 41840 -7920 41854
rect -7840 41906 -7760 41920
rect -7840 41854 -7826 41906
rect -7774 41854 -7760 41906
rect -7840 41840 -7760 41854
rect -7680 41906 -7600 41920
rect -7680 41854 -7666 41906
rect -7614 41854 -7600 41906
rect -7680 41840 -7600 41854
rect -7520 41906 -7440 41920
rect -7520 41854 -7506 41906
rect -7454 41854 -7440 41906
rect -7520 41840 -7440 41854
rect -7360 41906 -7280 41920
rect -7360 41854 -7346 41906
rect -7294 41854 -7280 41906
rect -7360 41840 -7280 41854
rect -7200 41906 -7120 41920
rect -7200 41854 -7186 41906
rect -7134 41854 -7120 41906
rect -7200 41840 -7120 41854
rect -7040 41906 -6960 41920
rect -7040 41854 -7026 41906
rect -6974 41854 -6960 41906
rect -7040 41840 -6960 41854
rect -6880 41906 -6800 41920
rect -6880 41854 -6866 41906
rect -6814 41854 -6800 41906
rect -6880 41840 -6800 41854
rect -6720 41906 -6640 41920
rect -6720 41854 -6706 41906
rect -6654 41854 -6640 41906
rect -6720 41840 -6640 41854
rect -6560 41906 -6480 41920
rect -6560 41854 -6546 41906
rect -6494 41854 -6480 41906
rect -6560 41840 -6480 41854
rect -6400 41906 -6320 41920
rect -6400 41854 -6386 41906
rect -6334 41854 -6320 41906
rect -6400 41840 -6320 41854
rect -6240 41906 -6160 41920
rect -6240 41854 -6226 41906
rect -6174 41854 -6160 41906
rect -6240 41840 -6160 41854
rect -6080 41906 -6000 41920
rect -6080 41854 -6066 41906
rect -6014 41854 -6000 41906
rect -6080 41840 -6000 41854
rect -5920 41906 -5840 41920
rect -5920 41854 -5906 41906
rect -5854 41854 -5840 41906
rect -5920 41840 -5840 41854
rect -5760 41906 -5680 41920
rect -5760 41854 -5746 41906
rect -5694 41854 -5680 41906
rect -5760 41840 -5680 41854
rect -5600 41906 -5520 41920
rect -5600 41854 -5586 41906
rect -5534 41854 -5520 41906
rect -5600 41840 -5520 41854
rect -5440 41906 -5360 41920
rect -5440 41854 -5426 41906
rect -5374 41854 -5360 41906
rect -5440 41840 -5360 41854
rect -5280 41906 -5200 41920
rect -5280 41854 -5266 41906
rect -5214 41854 -5200 41906
rect -5280 41840 -5200 41854
rect -5120 41906 -5040 41920
rect -5120 41854 -5106 41906
rect -5054 41854 -5040 41906
rect -5120 41840 -5040 41854
rect -4960 41906 -4880 41920
rect -4960 41854 -4946 41906
rect -4894 41854 -4880 41906
rect -4960 41840 -4880 41854
rect -4800 41906 -4720 41920
rect -4800 41854 -4786 41906
rect -4734 41854 -4720 41906
rect -4800 41840 -4720 41854
rect -4640 41906 -4560 41920
rect -4640 41854 -4626 41906
rect -4574 41854 -4560 41906
rect -4640 41840 -4560 41854
rect -4480 41906 -4400 41920
rect -4480 41854 -4466 41906
rect -4414 41854 -4400 41906
rect -4480 41840 -4400 41854
rect -4320 41906 -4240 41920
rect -4320 41854 -4306 41906
rect -4254 41854 -4240 41906
rect -4320 41840 -4240 41854
rect -4160 41906 -4080 41920
rect -4160 41854 -4146 41906
rect -4094 41854 -4080 41906
rect -4160 41840 -4080 41854
rect -4000 41906 -3920 41920
rect -4000 41854 -3986 41906
rect -3934 41854 -3920 41906
rect -4000 41840 -3920 41854
rect -3680 41906 -3600 41920
rect -3680 41854 -3666 41906
rect -3614 41854 -3600 41906
rect -3680 41840 -3600 41854
rect -3520 41906 -3440 41920
rect -3520 41854 -3506 41906
rect -3454 41854 -3440 41906
rect -3520 41840 -3440 41854
rect -3360 41906 -3280 41920
rect -3360 41854 -3346 41906
rect -3294 41854 -3280 41906
rect -3360 41840 -3280 41854
rect -3040 41906 -2960 41920
rect -3040 41854 -3026 41906
rect -2974 41854 -2960 41906
rect -3040 41840 -2960 41854
rect -2720 41906 -2640 41920
rect -2720 41854 -2706 41906
rect -2654 41854 -2640 41906
rect -2720 41840 -2640 41854
rect -2560 41906 -2480 41920
rect -2560 41854 -2546 41906
rect -2494 41854 -2480 41906
rect -2560 41840 -2480 41854
rect -2400 41906 -2320 41920
rect -2400 41854 -2386 41906
rect -2334 41854 -2320 41906
rect -2400 41840 -2320 41854
rect -2240 41906 -2160 41920
rect -2240 41854 -2226 41906
rect -2174 41854 -2160 41906
rect -2240 41840 -2160 41854
rect -2080 41906 -2000 41920
rect -2080 41854 -2066 41906
rect -2014 41854 -2000 41906
rect -2080 41840 -2000 41854
rect -1760 41906 -1680 41920
rect -1760 41854 -1746 41906
rect -1694 41854 -1680 41906
rect -1760 41840 -1680 41854
rect -1440 41906 -1360 41920
rect -1440 41854 -1426 41906
rect -1374 41854 -1360 41906
rect -1440 41840 -1360 41854
rect -1120 41906 -1040 41920
rect -1120 41854 -1106 41906
rect -1054 41854 -1040 41906
rect -1120 41840 -1040 41854
rect -33120 41346 -33040 41360
rect -33120 41294 -33106 41346
rect -33054 41294 -33040 41346
rect -33120 41280 -33040 41294
rect -32960 41346 -32880 41360
rect -32960 41294 -32946 41346
rect -32894 41294 -32880 41346
rect -32960 41280 -32880 41294
rect -32800 41346 -32720 41360
rect -32800 41294 -32786 41346
rect -32734 41294 -32720 41346
rect -32800 41280 -32720 41294
rect -32640 41346 -32560 41360
rect -32640 41294 -32626 41346
rect -32574 41294 -32560 41346
rect -32640 41280 -32560 41294
rect -32480 41346 -32400 41360
rect -32480 41294 -32466 41346
rect -32414 41294 -32400 41346
rect -32480 41280 -32400 41294
rect -32320 41346 -32240 41360
rect -32320 41294 -32306 41346
rect -32254 41294 -32240 41346
rect -32320 41280 -32240 41294
rect -32160 41346 -32080 41360
rect -32160 41294 -32146 41346
rect -32094 41294 -32080 41346
rect -32160 41280 -32080 41294
rect -32000 41346 -31920 41360
rect -32000 41294 -31986 41346
rect -31934 41294 -31920 41346
rect -32000 41280 -31920 41294
rect -31840 41346 -31760 41360
rect -31840 41294 -31826 41346
rect -31774 41294 -31760 41346
rect -31840 41280 -31760 41294
rect -31680 41346 -31600 41360
rect -31680 41294 -31666 41346
rect -31614 41294 -31600 41346
rect -31680 41280 -31600 41294
rect -31520 41346 -31440 41360
rect -31520 41294 -31506 41346
rect -31454 41294 -31440 41346
rect -31520 41280 -31440 41294
rect -31360 41346 -31280 41360
rect -31360 41294 -31346 41346
rect -31294 41294 -31280 41346
rect -31360 41280 -31280 41294
rect -31200 41346 -31120 41360
rect -31200 41294 -31186 41346
rect -31134 41294 -31120 41346
rect -31200 41280 -31120 41294
rect -29920 41346 -29840 41360
rect -29920 41294 -29906 41346
rect -29854 41294 -29840 41346
rect -29920 41280 -29840 41294
rect -29760 41346 -29680 41360
rect -29760 41294 -29746 41346
rect -29694 41294 -29680 41346
rect -29760 41280 -29680 41294
rect -29600 41346 -29520 41360
rect -29600 41294 -29586 41346
rect -29534 41294 -29520 41346
rect -29600 41280 -29520 41294
rect -29440 41346 -29360 41360
rect -29440 41294 -29426 41346
rect -29374 41294 -29360 41346
rect -29440 41280 -29360 41294
rect -29280 41346 -29200 41360
rect -29280 41294 -29266 41346
rect -29214 41294 -29200 41346
rect -29280 41280 -29200 41294
rect -29120 41346 -29040 41360
rect -29120 41294 -29106 41346
rect -29054 41294 -29040 41346
rect -29120 41280 -29040 41294
rect -28960 41346 -28880 41360
rect -28960 41294 -28946 41346
rect -28894 41294 -28880 41346
rect -28960 41280 -28880 41294
rect -28800 41346 -28720 41360
rect -28800 41294 -28786 41346
rect -28734 41294 -28720 41346
rect -28800 41280 -28720 41294
rect -28640 41346 -28560 41360
rect -28640 41294 -28626 41346
rect -28574 41294 -28560 41346
rect -28640 41280 -28560 41294
rect -28480 41346 -28400 41360
rect -28480 41294 -28466 41346
rect -28414 41294 -28400 41346
rect -28480 41280 -28400 41294
rect -28320 41346 -28240 41360
rect -28320 41294 -28306 41346
rect -28254 41294 -28240 41346
rect -28320 41280 -28240 41294
rect -28160 41346 -28080 41360
rect -28160 41294 -28146 41346
rect -28094 41294 -28080 41346
rect -28160 41280 -28080 41294
rect -28000 41346 -27920 41360
rect -28000 41294 -27986 41346
rect -27934 41294 -27920 41346
rect -28000 41280 -27920 41294
rect -27840 41346 -27760 41360
rect -27840 41294 -27826 41346
rect -27774 41294 -27760 41346
rect -27840 41280 -27760 41294
rect -27680 41346 -27600 41360
rect -27680 41294 -27666 41346
rect -27614 41294 -27600 41346
rect -27680 41280 -27600 41294
rect -27520 41346 -27440 41360
rect -27520 41294 -27506 41346
rect -27454 41294 -27440 41346
rect -27520 41280 -27440 41294
rect -27360 41346 -27280 41360
rect -27360 41294 -27346 41346
rect -27294 41294 -27280 41346
rect -27360 41280 -27280 41294
rect -27200 41346 -27120 41360
rect -27200 41294 -27186 41346
rect -27134 41294 -27120 41346
rect -27200 41280 -27120 41294
rect -27040 41346 -26960 41360
rect -27040 41294 -27026 41346
rect -26974 41294 -26960 41346
rect -27040 41280 -26960 41294
rect -26880 41346 -26800 41360
rect -26880 41294 -26866 41346
rect -26814 41294 -26800 41346
rect -26880 41280 -26800 41294
rect -26720 41346 -26640 41360
rect -26720 41294 -26706 41346
rect -26654 41294 -26640 41346
rect -26720 41280 -26640 41294
rect -26560 41346 -26480 41360
rect -26560 41294 -26546 41346
rect -26494 41294 -26480 41346
rect -26560 41280 -26480 41294
rect -26400 41346 -26320 41360
rect -26400 41294 -26386 41346
rect -26334 41294 -26320 41346
rect -26400 41280 -26320 41294
rect -26240 41346 -26160 41360
rect -26240 41294 -26226 41346
rect -26174 41294 -26160 41346
rect -26240 41280 -26160 41294
rect -26080 41346 -26000 41360
rect -26080 41294 -26066 41346
rect -26014 41294 -26000 41346
rect -26080 41280 -26000 41294
rect -25920 41346 -25840 41360
rect -25920 41294 -25906 41346
rect -25854 41294 -25840 41346
rect -25920 41280 -25840 41294
rect -25760 41346 -25680 41360
rect -25760 41294 -25746 41346
rect -25694 41294 -25680 41346
rect -25760 41280 -25680 41294
rect -25600 41346 -25520 41360
rect -25600 41294 -25586 41346
rect -25534 41294 -25520 41346
rect -25600 41280 -25520 41294
rect -25440 41346 -25360 41360
rect -25440 41294 -25426 41346
rect -25374 41294 -25360 41346
rect -25440 41280 -25360 41294
rect -25280 41346 -25200 41360
rect -25280 41294 -25266 41346
rect -25214 41294 -25200 41346
rect -25280 41280 -25200 41294
rect -25120 41346 -25040 41360
rect -25120 41294 -25106 41346
rect -25054 41294 -25040 41346
rect -25120 41280 -25040 41294
rect -24960 41346 -24880 41360
rect -24960 41294 -24946 41346
rect -24894 41294 -24880 41346
rect -24960 41280 -24880 41294
rect -24800 41346 -24720 41360
rect -24800 41294 -24786 41346
rect -24734 41294 -24720 41346
rect -24800 41280 -24720 41294
rect -24640 41346 -24560 41360
rect -24640 41294 -24626 41346
rect -24574 41294 -24560 41346
rect -24640 41280 -24560 41294
rect -24480 41346 -24400 41360
rect -24480 41294 -24466 41346
rect -24414 41294 -24400 41346
rect -24480 41280 -24400 41294
rect -24320 41346 -24240 41360
rect -24320 41294 -24306 41346
rect -24254 41294 -24240 41346
rect -24320 41280 -24240 41294
rect -24160 41346 -24080 41360
rect -24160 41294 -24146 41346
rect -24094 41294 -24080 41346
rect -24160 41280 -24080 41294
rect -24000 41346 -23920 41360
rect -24000 41294 -23986 41346
rect -23934 41294 -23920 41346
rect -24000 41280 -23920 41294
rect -23840 41346 -23760 41360
rect -23840 41294 -23826 41346
rect -23774 41294 -23760 41346
rect -23840 41280 -23760 41294
rect -23680 41346 -23600 41360
rect -23680 41294 -23666 41346
rect -23614 41294 -23600 41346
rect -23680 41280 -23600 41294
rect -23520 41346 -23440 41360
rect -23520 41294 -23506 41346
rect -23454 41294 -23440 41346
rect -23520 41280 -23440 41294
rect -23360 41346 -23280 41360
rect -23360 41294 -23346 41346
rect -23294 41294 -23280 41346
rect -23360 41280 -23280 41294
rect -23200 41346 -23120 41360
rect -23200 41294 -23186 41346
rect -23134 41294 -23120 41346
rect -23200 41280 -23120 41294
rect -23040 41346 -22960 41360
rect -23040 41294 -23026 41346
rect -22974 41294 -22960 41346
rect -23040 41280 -22960 41294
rect -22880 41346 -22800 41360
rect -22880 41294 -22866 41346
rect -22814 41294 -22800 41346
rect -22880 41280 -22800 41294
rect -22720 41346 -22640 41360
rect -22720 41294 -22706 41346
rect -22654 41294 -22640 41346
rect -22720 41280 -22640 41294
rect -22560 41346 -22480 41360
rect -22560 41294 -22546 41346
rect -22494 41294 -22480 41346
rect -22560 41280 -22480 41294
rect -22400 41346 -22320 41360
rect -22400 41294 -22386 41346
rect -22334 41294 -22320 41346
rect -22400 41280 -22320 41294
rect -22240 41346 -22160 41360
rect -22240 41294 -22226 41346
rect -22174 41294 -22160 41346
rect -22240 41280 -22160 41294
rect -22080 41346 -22000 41360
rect -22080 41294 -22066 41346
rect -22014 41294 -22000 41346
rect -22080 41280 -22000 41294
rect -21920 41346 -21840 41360
rect -21920 41294 -21906 41346
rect -21854 41294 -21840 41346
rect -21920 41280 -21840 41294
rect -21760 41346 -21680 41360
rect -21760 41294 -21746 41346
rect -21694 41294 -21680 41346
rect -21760 41280 -21680 41294
rect -21600 41346 -21520 41360
rect -21600 41294 -21586 41346
rect -21534 41294 -21520 41346
rect -21600 41280 -21520 41294
rect -21440 41346 -21360 41360
rect -21440 41294 -21426 41346
rect -21374 41294 -21360 41346
rect -21440 41280 -21360 41294
rect -21280 41346 -21200 41360
rect -21280 41294 -21266 41346
rect -21214 41294 -21200 41346
rect -21280 41280 -21200 41294
rect -21120 41346 -21040 41360
rect -21120 41294 -21106 41346
rect -21054 41294 -21040 41346
rect -21120 41280 -21040 41294
rect -20960 41346 -20880 41360
rect -20960 41294 -20946 41346
rect -20894 41294 -20880 41346
rect -20960 41280 -20880 41294
rect -20800 41346 -20720 41360
rect -20800 41294 -20786 41346
rect -20734 41294 -20720 41346
rect -20800 41280 -20720 41294
rect -20640 41346 -20560 41360
rect -20640 41294 -20626 41346
rect -20574 41294 -20560 41346
rect -20640 41280 -20560 41294
rect -20480 41346 -20400 41360
rect -20480 41294 -20466 41346
rect -20414 41294 -20400 41346
rect -20480 41280 -20400 41294
rect -20320 41346 -20240 41360
rect -20320 41294 -20306 41346
rect -20254 41294 -20240 41346
rect -20320 41280 -20240 41294
rect -20160 41346 -20080 41360
rect -20160 41294 -20146 41346
rect -20094 41294 -20080 41346
rect -20160 41280 -20080 41294
rect -20000 41346 -19920 41360
rect -20000 41294 -19986 41346
rect -19934 41294 -19920 41346
rect -20000 41280 -19920 41294
rect -19840 41346 -19760 41360
rect -19840 41294 -19826 41346
rect -19774 41294 -19760 41346
rect -19840 41280 -19760 41294
rect -19680 41346 -19600 41360
rect -19680 41294 -19666 41346
rect -19614 41294 -19600 41346
rect -19680 41280 -19600 41294
rect -19520 41346 -19440 41360
rect -19520 41294 -19506 41346
rect -19454 41294 -19440 41346
rect -19520 41280 -19440 41294
rect -19360 41346 -19280 41360
rect -19360 41294 -19346 41346
rect -19294 41294 -19280 41346
rect -19360 41280 -19280 41294
rect -19200 41346 -19120 41360
rect -19200 41294 -19186 41346
rect -19134 41294 -19120 41346
rect -19200 41280 -19120 41294
rect -19040 41346 -18960 41360
rect -19040 41294 -19026 41346
rect -18974 41294 -18960 41346
rect -19040 41280 -18960 41294
rect -18880 41346 -18800 41360
rect -18880 41294 -18866 41346
rect -18814 41294 -18800 41346
rect -18880 41280 -18800 41294
rect -18720 41346 -18640 41360
rect -18720 41294 -18706 41346
rect -18654 41294 -18640 41346
rect -18720 41280 -18640 41294
rect -18560 41346 -18480 41360
rect -18560 41294 -18546 41346
rect -18494 41294 -18480 41346
rect -18560 41280 -18480 41294
rect -18400 41346 -18320 41360
rect -18400 41294 -18386 41346
rect -18334 41294 -18320 41346
rect -18400 41280 -18320 41294
rect -18240 41346 -18160 41360
rect -18240 41294 -18226 41346
rect -18174 41294 -18160 41346
rect -18240 41280 -18160 41294
rect -18080 41346 -18000 41360
rect -18080 41294 -18066 41346
rect -18014 41294 -18000 41346
rect -18080 41280 -18000 41294
rect -17920 41346 -17840 41360
rect -17920 41294 -17906 41346
rect -17854 41294 -17840 41346
rect -17920 41280 -17840 41294
rect -17760 41346 -17680 41360
rect -17760 41294 -17746 41346
rect -17694 41294 -17680 41346
rect -17760 41280 -17680 41294
rect -17600 41346 -17520 41360
rect -17600 41294 -17586 41346
rect -17534 41294 -17520 41346
rect -17600 41280 -17520 41294
rect -17440 41346 -17360 41360
rect -17440 41294 -17426 41346
rect -17374 41294 -17360 41346
rect -17440 41280 -17360 41294
rect -17280 41346 -17200 41360
rect -17280 41294 -17266 41346
rect -17214 41294 -17200 41346
rect -17280 41280 -17200 41294
rect -17120 41346 -17040 41360
rect -17120 41294 -17106 41346
rect -17054 41294 -17040 41346
rect -17120 41280 -17040 41294
rect -16960 41346 -16880 41360
rect -16960 41294 -16946 41346
rect -16894 41294 -16880 41346
rect -16960 41280 -16880 41294
rect -16800 41346 -16720 41360
rect -16800 41294 -16786 41346
rect -16734 41294 -16720 41346
rect -16800 41280 -16720 41294
rect -16640 41346 -16560 41360
rect -16640 41294 -16626 41346
rect -16574 41294 -16560 41346
rect -16640 41280 -16560 41294
rect -16480 41346 -16400 41360
rect -16480 41294 -16466 41346
rect -16414 41294 -16400 41346
rect -16480 41280 -16400 41294
rect -16320 41346 -16240 41360
rect -16320 41294 -16306 41346
rect -16254 41294 -16240 41346
rect -16320 41280 -16240 41294
rect -16160 41346 -16080 41360
rect -16160 41294 -16146 41346
rect -16094 41294 -16080 41346
rect -16160 41280 -16080 41294
rect -16000 41346 -15920 41360
rect -16000 41294 -15986 41346
rect -15934 41294 -15920 41346
rect -16000 41280 -15920 41294
rect -15840 41346 -15760 41360
rect -15840 41294 -15826 41346
rect -15774 41294 -15760 41346
rect -15840 41280 -15760 41294
rect -15680 41346 -15600 41360
rect -15680 41294 -15666 41346
rect -15614 41294 -15600 41346
rect -15680 41280 -15600 41294
rect -15520 41346 -15440 41360
rect -15520 41294 -15506 41346
rect -15454 41294 -15440 41346
rect -15520 41280 -15440 41294
rect -15360 41346 -15280 41360
rect -15360 41294 -15346 41346
rect -15294 41294 -15280 41346
rect -15360 41280 -15280 41294
rect -15200 41346 -15120 41360
rect -15200 41294 -15186 41346
rect -15134 41294 -15120 41346
rect -15200 41280 -15120 41294
rect -15040 41346 -14960 41360
rect -15040 41294 -15026 41346
rect -14974 41294 -14960 41346
rect -15040 41280 -14960 41294
rect -14880 41346 -14800 41360
rect -14880 41294 -14866 41346
rect -14814 41294 -14800 41346
rect -14880 41280 -14800 41294
rect -14720 41346 -14640 41360
rect -14720 41294 -14706 41346
rect -14654 41294 -14640 41346
rect -14720 41280 -14640 41294
rect -14560 41346 -14480 41360
rect -14560 41294 -14546 41346
rect -14494 41294 -14480 41346
rect -14560 41280 -14480 41294
rect -14400 41346 -14320 41360
rect -14400 41294 -14386 41346
rect -14334 41294 -14320 41346
rect -14400 41280 -14320 41294
rect -14240 41346 -14160 41360
rect -14240 41294 -14226 41346
rect -14174 41294 -14160 41346
rect -14240 41280 -14160 41294
rect -14080 41346 -14000 41360
rect -14080 41294 -14066 41346
rect -14014 41294 -14000 41346
rect -14080 41280 -14000 41294
rect -13920 41346 -13840 41360
rect -13920 41294 -13906 41346
rect -13854 41294 -13840 41346
rect -13920 41280 -13840 41294
rect -13760 41346 -13680 41360
rect -13760 41294 -13746 41346
rect -13694 41294 -13680 41346
rect -13760 41280 -13680 41294
rect -13600 41346 -13520 41360
rect -13600 41294 -13586 41346
rect -13534 41294 -13520 41346
rect -13600 41280 -13520 41294
rect -13440 41346 -13360 41360
rect -13440 41294 -13426 41346
rect -13374 41294 -13360 41346
rect -13440 41280 -13360 41294
rect -13280 41346 -13200 41360
rect -13280 41294 -13266 41346
rect -13214 41294 -13200 41346
rect -13280 41280 -13200 41294
rect -13120 41346 -13040 41360
rect -13120 41294 -13106 41346
rect -13054 41294 -13040 41346
rect -13120 41280 -13040 41294
rect -12960 41346 -12880 41360
rect -12960 41294 -12946 41346
rect -12894 41294 -12880 41346
rect -12960 41280 -12880 41294
rect -12800 41346 -12720 41360
rect -12800 41294 -12786 41346
rect -12734 41294 -12720 41346
rect -12800 41280 -12720 41294
rect -12640 41346 -12560 41360
rect -12640 41294 -12626 41346
rect -12574 41294 -12560 41346
rect -12640 41280 -12560 41294
rect -12480 41346 -12400 41360
rect -12480 41294 -12466 41346
rect -12414 41294 -12400 41346
rect -12480 41280 -12400 41294
rect -12320 41346 -12240 41360
rect -12320 41294 -12306 41346
rect -12254 41294 -12240 41346
rect -12320 41280 -12240 41294
rect -11360 41346 -11280 41360
rect -11360 41294 -11346 41346
rect -11294 41294 -11280 41346
rect -11360 41280 -11280 41294
rect -11200 41346 -11120 41360
rect -11200 41294 -11186 41346
rect -11134 41294 -11120 41346
rect -11200 41280 -11120 41294
rect -11040 41346 -10960 41360
rect -11040 41294 -11026 41346
rect -10974 41294 -10960 41346
rect -11040 41280 -10960 41294
rect -10880 41346 -10800 41360
rect -10880 41294 -10866 41346
rect -10814 41294 -10800 41346
rect -10880 41280 -10800 41294
rect -10720 41346 -10640 41360
rect -10720 41294 -10706 41346
rect -10654 41294 -10640 41346
rect -10720 41280 -10640 41294
rect -10560 41346 -10480 41360
rect -10560 41294 -10546 41346
rect -10494 41294 -10480 41346
rect -10560 41280 -10480 41294
rect -10400 41346 -10320 41360
rect -10400 41294 -10386 41346
rect -10334 41294 -10320 41346
rect -10400 41280 -10320 41294
rect -10240 41346 -10160 41360
rect -10240 41294 -10226 41346
rect -10174 41294 -10160 41346
rect -10240 41280 -10160 41294
rect -10080 41346 -10000 41360
rect -10080 41294 -10066 41346
rect -10014 41294 -10000 41346
rect -10080 41280 -10000 41294
rect -9920 41346 -9840 41360
rect -9920 41294 -9906 41346
rect -9854 41294 -9840 41346
rect -9920 41280 -9840 41294
rect -9760 41346 -9680 41360
rect -9760 41294 -9746 41346
rect -9694 41294 -9680 41346
rect -9760 41280 -9680 41294
rect -9600 41346 -9520 41360
rect -9600 41294 -9586 41346
rect -9534 41294 -9520 41346
rect -9600 41280 -9520 41294
rect -9440 41346 -9360 41360
rect -9440 41294 -9426 41346
rect -9374 41294 -9360 41346
rect -9440 41280 -9360 41294
rect -9280 41346 -9200 41360
rect -9280 41294 -9266 41346
rect -9214 41294 -9200 41346
rect -9280 41280 -9200 41294
rect -9120 41346 -9040 41360
rect -9120 41294 -9106 41346
rect -9054 41294 -9040 41346
rect -9120 41280 -9040 41294
rect -8960 41346 -8880 41360
rect -8960 41294 -8946 41346
rect -8894 41294 -8880 41346
rect -8960 41280 -8880 41294
rect -8800 41346 -8720 41360
rect -8800 41294 -8786 41346
rect -8734 41294 -8720 41346
rect -8800 41280 -8720 41294
rect -8640 41346 -8560 41360
rect -8640 41294 -8626 41346
rect -8574 41294 -8560 41346
rect -8640 41280 -8560 41294
rect -8480 41346 -8400 41360
rect -8480 41294 -8466 41346
rect -8414 41294 -8400 41346
rect -8480 41280 -8400 41294
rect -8320 41346 -8240 41360
rect -8320 41294 -8306 41346
rect -8254 41294 -8240 41346
rect -8320 41280 -8240 41294
rect -8160 41346 -8080 41360
rect -8160 41294 -8146 41346
rect -8094 41294 -8080 41346
rect -8160 41280 -8080 41294
rect -8000 41346 -7920 41360
rect -8000 41294 -7986 41346
rect -7934 41294 -7920 41346
rect -8000 41280 -7920 41294
rect -7840 41346 -7760 41360
rect -7840 41294 -7826 41346
rect -7774 41294 -7760 41346
rect -7840 41280 -7760 41294
rect -7680 41346 -7600 41360
rect -7680 41294 -7666 41346
rect -7614 41294 -7600 41346
rect -7680 41280 -7600 41294
rect -7520 41346 -7440 41360
rect -7520 41294 -7506 41346
rect -7454 41294 -7440 41346
rect -7520 41280 -7440 41294
rect -7360 41346 -7280 41360
rect -7360 41294 -7346 41346
rect -7294 41294 -7280 41346
rect -7360 41280 -7280 41294
rect -7200 41346 -7120 41360
rect -7200 41294 -7186 41346
rect -7134 41294 -7120 41346
rect -7200 41280 -7120 41294
rect -7040 41346 -6960 41360
rect -7040 41294 -7026 41346
rect -6974 41294 -6960 41346
rect -7040 41280 -6960 41294
rect -6880 41346 -6800 41360
rect -6880 41294 -6866 41346
rect -6814 41294 -6800 41346
rect -6880 41280 -6800 41294
rect -6720 41346 -6640 41360
rect -6720 41294 -6706 41346
rect -6654 41294 -6640 41346
rect -6720 41280 -6640 41294
rect -6560 41346 -6480 41360
rect -6560 41294 -6546 41346
rect -6494 41294 -6480 41346
rect -6560 41280 -6480 41294
rect -6400 41346 -6320 41360
rect -6400 41294 -6386 41346
rect -6334 41294 -6320 41346
rect -6400 41280 -6320 41294
rect -6240 41346 -6160 41360
rect -6240 41294 -6226 41346
rect -6174 41294 -6160 41346
rect -6240 41280 -6160 41294
rect -6080 41346 -6000 41360
rect -6080 41294 -6066 41346
rect -6014 41294 -6000 41346
rect -6080 41280 -6000 41294
rect -5920 41346 -5840 41360
rect -5920 41294 -5906 41346
rect -5854 41294 -5840 41346
rect -5920 41280 -5840 41294
rect -5760 41346 -5680 41360
rect -5760 41294 -5746 41346
rect -5694 41294 -5680 41346
rect -5760 41280 -5680 41294
rect -5600 41346 -5520 41360
rect -5600 41294 -5586 41346
rect -5534 41294 -5520 41346
rect -5600 41280 -5520 41294
rect -5440 41346 -5360 41360
rect -5440 41294 -5426 41346
rect -5374 41294 -5360 41346
rect -5440 41280 -5360 41294
rect -5280 41346 -5200 41360
rect -5280 41294 -5266 41346
rect -5214 41294 -5200 41346
rect -5280 41280 -5200 41294
rect -5120 41346 -5040 41360
rect -5120 41294 -5106 41346
rect -5054 41294 -5040 41346
rect -5120 41280 -5040 41294
rect -4960 41346 -4880 41360
rect -4960 41294 -4946 41346
rect -4894 41294 -4880 41346
rect -4960 41280 -4880 41294
rect -4800 41346 -4720 41360
rect -4800 41294 -4786 41346
rect -4734 41294 -4720 41346
rect -4800 41280 -4720 41294
rect -4640 41346 -4560 41360
rect -4640 41294 -4626 41346
rect -4574 41294 -4560 41346
rect -4640 41280 -4560 41294
rect -4480 41346 -4400 41360
rect -4480 41294 -4466 41346
rect -4414 41294 -4400 41346
rect -4480 41280 -4400 41294
rect -4320 41346 -4240 41360
rect -4320 41294 -4306 41346
rect -4254 41294 -4240 41346
rect -4320 41280 -4240 41294
rect -4160 41346 -4080 41360
rect -4160 41294 -4146 41346
rect -4094 41294 -4080 41346
rect -4160 41280 -4080 41294
rect -4000 41346 -3920 41360
rect -4000 41294 -3986 41346
rect -3934 41294 -3920 41346
rect -4000 41280 -3920 41294
rect -3840 41337 -3760 41360
rect -3840 41303 -3817 41337
rect -3783 41303 -3760 41337
rect -3840 41280 -3760 41303
rect -3680 41346 -3600 41360
rect -3680 41294 -3666 41346
rect -3614 41294 -3600 41346
rect -3680 41280 -3600 41294
rect -3520 41346 -3440 41360
rect -3520 41294 -3506 41346
rect -3454 41294 -3440 41346
rect -3520 41280 -3440 41294
rect 41040 41346 41120 41360
rect 41040 41294 41054 41346
rect 41106 41294 41120 41346
rect 41040 41280 41120 41294
rect 41200 41346 41280 41360
rect 41200 41294 41214 41346
rect 41266 41294 41280 41346
rect 41200 41280 41280 41294
rect 41360 41346 41440 41360
rect 41360 41294 41374 41346
rect 41426 41294 41440 41346
rect 41360 41280 41440 41294
rect 41520 41346 41600 41360
rect 41520 41294 41534 41346
rect 41586 41294 41600 41346
rect 41520 41280 41600 41294
rect 41680 41346 41760 41360
rect 41680 41294 41694 41346
rect 41746 41294 41760 41346
rect 41680 41280 41760 41294
rect 41840 41346 41920 41360
rect 41840 41294 41854 41346
rect 41906 41294 41920 41346
rect 41840 41280 41920 41294
rect 42000 41346 42080 41360
rect 42000 41294 42014 41346
rect 42066 41294 42080 41346
rect 42000 41280 42080 41294
rect 42160 41346 42240 41360
rect 42160 41294 42174 41346
rect 42226 41294 42240 41346
rect 42160 41280 42240 41294
rect 42320 41346 42400 41360
rect 42320 41294 42334 41346
rect 42386 41294 42400 41346
rect 42320 41280 42400 41294
rect 42480 41346 42560 41360
rect 42480 41294 42494 41346
rect 42546 41294 42560 41346
rect 42480 41280 42560 41294
rect 42640 41346 42720 41360
rect 42640 41294 42654 41346
rect 42706 41294 42720 41346
rect 42640 41280 42720 41294
rect 42800 41346 42880 41360
rect 42800 41294 42814 41346
rect 42866 41294 42880 41346
rect 42800 41280 42880 41294
rect 42960 41346 43040 41360
rect 42960 41294 42974 41346
rect 43026 41294 43040 41346
rect 42960 41280 43040 41294
rect 43120 41346 43200 41360
rect 43120 41294 43134 41346
rect 43186 41294 43200 41346
rect 43120 41280 43200 41294
rect -33120 41026 -33040 41040
rect -33120 40974 -33106 41026
rect -33054 40974 -33040 41026
rect -33120 40960 -33040 40974
rect -32960 41026 -32880 41040
rect -32960 40974 -32946 41026
rect -32894 40974 -32880 41026
rect -32960 40960 -32880 40974
rect -32800 41026 -32720 41040
rect -32800 40974 -32786 41026
rect -32734 40974 -32720 41026
rect -32800 40960 -32720 40974
rect -32640 41026 -32560 41040
rect -32640 40974 -32626 41026
rect -32574 40974 -32560 41026
rect -32640 40960 -32560 40974
rect -32480 41026 -32400 41040
rect -32480 40974 -32466 41026
rect -32414 40974 -32400 41026
rect -32480 40960 -32400 40974
rect -32320 41026 -32240 41040
rect -32320 40974 -32306 41026
rect -32254 40974 -32240 41026
rect -32320 40960 -32240 40974
rect -32160 41026 -32080 41040
rect -32160 40974 -32146 41026
rect -32094 40974 -32080 41026
rect -32160 40960 -32080 40974
rect -32000 41026 -31920 41040
rect -32000 40974 -31986 41026
rect -31934 40974 -31920 41026
rect -32000 40960 -31920 40974
rect -31840 41026 -31760 41040
rect -31840 40974 -31826 41026
rect -31774 40974 -31760 41026
rect -31840 40960 -31760 40974
rect -31680 41026 -31600 41040
rect -31680 40974 -31666 41026
rect -31614 40974 -31600 41026
rect -31680 40960 -31600 40974
rect -31520 41026 -31440 41040
rect -31520 40974 -31506 41026
rect -31454 40974 -31440 41026
rect -31520 40960 -31440 40974
rect -31360 41026 -31280 41040
rect -31360 40974 -31346 41026
rect -31294 40974 -31280 41026
rect -31360 40960 -31280 40974
rect -31200 41026 -31120 41040
rect -31200 40974 -31186 41026
rect -31134 40974 -31120 41026
rect -31200 40960 -31120 40974
rect -29920 41026 -29840 41040
rect -29920 40974 -29906 41026
rect -29854 40974 -29840 41026
rect -29920 40960 -29840 40974
rect -29760 41026 -29680 41040
rect -29760 40974 -29746 41026
rect -29694 40974 -29680 41026
rect -29760 40960 -29680 40974
rect -29600 41026 -29520 41040
rect -29600 40974 -29586 41026
rect -29534 40974 -29520 41026
rect -29600 40960 -29520 40974
rect -29440 41026 -29360 41040
rect -29440 40974 -29426 41026
rect -29374 40974 -29360 41026
rect -29440 40960 -29360 40974
rect -29280 41026 -29200 41040
rect -29280 40974 -29266 41026
rect -29214 40974 -29200 41026
rect -29280 40960 -29200 40974
rect -29120 41026 -29040 41040
rect -29120 40974 -29106 41026
rect -29054 40974 -29040 41026
rect -29120 40960 -29040 40974
rect -28960 41026 -28880 41040
rect -28960 40974 -28946 41026
rect -28894 40974 -28880 41026
rect -28960 40960 -28880 40974
rect -28800 41026 -28720 41040
rect -28800 40974 -28786 41026
rect -28734 40974 -28720 41026
rect -28800 40960 -28720 40974
rect -28640 41026 -28560 41040
rect -28640 40974 -28626 41026
rect -28574 40974 -28560 41026
rect -28640 40960 -28560 40974
rect -28480 41026 -28400 41040
rect -28480 40974 -28466 41026
rect -28414 40974 -28400 41026
rect -28480 40960 -28400 40974
rect -28320 41026 -28240 41040
rect -28320 40974 -28306 41026
rect -28254 40974 -28240 41026
rect -28320 40960 -28240 40974
rect -28160 41026 -28080 41040
rect -28160 40974 -28146 41026
rect -28094 40974 -28080 41026
rect -28160 40960 -28080 40974
rect -28000 41026 -27920 41040
rect -28000 40974 -27986 41026
rect -27934 40974 -27920 41026
rect -28000 40960 -27920 40974
rect -27840 41026 -27760 41040
rect -27840 40974 -27826 41026
rect -27774 40974 -27760 41026
rect -27840 40960 -27760 40974
rect -27680 41026 -27600 41040
rect -27680 40974 -27666 41026
rect -27614 40974 -27600 41026
rect -27680 40960 -27600 40974
rect -27520 41026 -27440 41040
rect -27520 40974 -27506 41026
rect -27454 40974 -27440 41026
rect -27520 40960 -27440 40974
rect -27360 41026 -27280 41040
rect -27360 40974 -27346 41026
rect -27294 40974 -27280 41026
rect -27360 40960 -27280 40974
rect -27200 41026 -27120 41040
rect -27200 40974 -27186 41026
rect -27134 40974 -27120 41026
rect -27200 40960 -27120 40974
rect -27040 41026 -26960 41040
rect -27040 40974 -27026 41026
rect -26974 40974 -26960 41026
rect -27040 40960 -26960 40974
rect -26880 41026 -26800 41040
rect -26880 40974 -26866 41026
rect -26814 40974 -26800 41026
rect -26880 40960 -26800 40974
rect -26720 41026 -26640 41040
rect -26720 40974 -26706 41026
rect -26654 40974 -26640 41026
rect -26720 40960 -26640 40974
rect -26560 41026 -26480 41040
rect -26560 40974 -26546 41026
rect -26494 40974 -26480 41026
rect -26560 40960 -26480 40974
rect -26400 41026 -26320 41040
rect -26400 40974 -26386 41026
rect -26334 40974 -26320 41026
rect -26400 40960 -26320 40974
rect -26240 41026 -26160 41040
rect -26240 40974 -26226 41026
rect -26174 40974 -26160 41026
rect -26240 40960 -26160 40974
rect -26080 41026 -26000 41040
rect -26080 40974 -26066 41026
rect -26014 40974 -26000 41026
rect -26080 40960 -26000 40974
rect -25920 41026 -25840 41040
rect -25920 40974 -25906 41026
rect -25854 40974 -25840 41026
rect -25920 40960 -25840 40974
rect -25760 41026 -25680 41040
rect -25760 40974 -25746 41026
rect -25694 40974 -25680 41026
rect -25760 40960 -25680 40974
rect -25600 41026 -25520 41040
rect -25600 40974 -25586 41026
rect -25534 40974 -25520 41026
rect -25600 40960 -25520 40974
rect -25440 41026 -25360 41040
rect -25440 40974 -25426 41026
rect -25374 40974 -25360 41026
rect -25440 40960 -25360 40974
rect -25280 41026 -25200 41040
rect -25280 40974 -25266 41026
rect -25214 40974 -25200 41026
rect -25280 40960 -25200 40974
rect -25120 41026 -25040 41040
rect -25120 40974 -25106 41026
rect -25054 40974 -25040 41026
rect -25120 40960 -25040 40974
rect -24960 41026 -24880 41040
rect -24960 40974 -24946 41026
rect -24894 40974 -24880 41026
rect -24960 40960 -24880 40974
rect -24800 41026 -24720 41040
rect -24800 40974 -24786 41026
rect -24734 40974 -24720 41026
rect -24800 40960 -24720 40974
rect -24640 41026 -24560 41040
rect -24640 40974 -24626 41026
rect -24574 40974 -24560 41026
rect -24640 40960 -24560 40974
rect -24480 41026 -24400 41040
rect -24480 40974 -24466 41026
rect -24414 40974 -24400 41026
rect -24480 40960 -24400 40974
rect -24320 41026 -24240 41040
rect -24320 40974 -24306 41026
rect -24254 40974 -24240 41026
rect -24320 40960 -24240 40974
rect -24160 41026 -24080 41040
rect -24160 40974 -24146 41026
rect -24094 40974 -24080 41026
rect -24160 40960 -24080 40974
rect -24000 41026 -23920 41040
rect -24000 40974 -23986 41026
rect -23934 40974 -23920 41026
rect -24000 40960 -23920 40974
rect -23840 41026 -23760 41040
rect -23840 40974 -23826 41026
rect -23774 40974 -23760 41026
rect -23840 40960 -23760 40974
rect -23680 41026 -23600 41040
rect -23680 40974 -23666 41026
rect -23614 40974 -23600 41026
rect -23680 40960 -23600 40974
rect -23520 41026 -23440 41040
rect -23520 40974 -23506 41026
rect -23454 40974 -23440 41026
rect -23520 40960 -23440 40974
rect -23360 41026 -23280 41040
rect -23360 40974 -23346 41026
rect -23294 40974 -23280 41026
rect -23360 40960 -23280 40974
rect -23200 41026 -23120 41040
rect -23200 40974 -23186 41026
rect -23134 40974 -23120 41026
rect -23200 40960 -23120 40974
rect -23040 41026 -22960 41040
rect -23040 40974 -23026 41026
rect -22974 40974 -22960 41026
rect -23040 40960 -22960 40974
rect -22880 41026 -22800 41040
rect -22880 40974 -22866 41026
rect -22814 40974 -22800 41026
rect -22880 40960 -22800 40974
rect -22720 41026 -22640 41040
rect -22720 40974 -22706 41026
rect -22654 40974 -22640 41026
rect -22720 40960 -22640 40974
rect -22560 41026 -22480 41040
rect -22560 40974 -22546 41026
rect -22494 40974 -22480 41026
rect -22560 40960 -22480 40974
rect -22400 41026 -22320 41040
rect -22400 40974 -22386 41026
rect -22334 40974 -22320 41026
rect -22400 40960 -22320 40974
rect -22240 41026 -22160 41040
rect -22240 40974 -22226 41026
rect -22174 40974 -22160 41026
rect -22240 40960 -22160 40974
rect -22080 41026 -22000 41040
rect -22080 40974 -22066 41026
rect -22014 40974 -22000 41026
rect -22080 40960 -22000 40974
rect -21920 41026 -21840 41040
rect -21920 40974 -21906 41026
rect -21854 40974 -21840 41026
rect -21920 40960 -21840 40974
rect -21760 41026 -21680 41040
rect -21760 40974 -21746 41026
rect -21694 40974 -21680 41026
rect -21760 40960 -21680 40974
rect -21600 41026 -21520 41040
rect -21600 40974 -21586 41026
rect -21534 40974 -21520 41026
rect -21600 40960 -21520 40974
rect -21440 41026 -21360 41040
rect -21440 40974 -21426 41026
rect -21374 40974 -21360 41026
rect -21440 40960 -21360 40974
rect -21280 41026 -21200 41040
rect -21280 40974 -21266 41026
rect -21214 40974 -21200 41026
rect -21280 40960 -21200 40974
rect -21120 41026 -21040 41040
rect -21120 40974 -21106 41026
rect -21054 40974 -21040 41026
rect -21120 40960 -21040 40974
rect -20960 41026 -20880 41040
rect -20960 40974 -20946 41026
rect -20894 40974 -20880 41026
rect -20960 40960 -20880 40974
rect -20800 41026 -20720 41040
rect -20800 40974 -20786 41026
rect -20734 40974 -20720 41026
rect -20800 40960 -20720 40974
rect -20640 41026 -20560 41040
rect -20640 40974 -20626 41026
rect -20574 40974 -20560 41026
rect -20640 40960 -20560 40974
rect -20480 41026 -20400 41040
rect -20480 40974 -20466 41026
rect -20414 40974 -20400 41026
rect -20480 40960 -20400 40974
rect -20320 41026 -20240 41040
rect -20320 40974 -20306 41026
rect -20254 40974 -20240 41026
rect -20320 40960 -20240 40974
rect -20160 41026 -20080 41040
rect -20160 40974 -20146 41026
rect -20094 40974 -20080 41026
rect -20160 40960 -20080 40974
rect -20000 41026 -19920 41040
rect -20000 40974 -19986 41026
rect -19934 40974 -19920 41026
rect -20000 40960 -19920 40974
rect -19840 41026 -19760 41040
rect -19840 40974 -19826 41026
rect -19774 40974 -19760 41026
rect -19840 40960 -19760 40974
rect -19680 41026 -19600 41040
rect -19680 40974 -19666 41026
rect -19614 40974 -19600 41026
rect -19680 40960 -19600 40974
rect -19520 41026 -19440 41040
rect -19520 40974 -19506 41026
rect -19454 40974 -19440 41026
rect -19520 40960 -19440 40974
rect -19360 41026 -19280 41040
rect -19360 40974 -19346 41026
rect -19294 40974 -19280 41026
rect -19360 40960 -19280 40974
rect -19200 41026 -19120 41040
rect -19200 40974 -19186 41026
rect -19134 40974 -19120 41026
rect -19200 40960 -19120 40974
rect -19040 41026 -18960 41040
rect -19040 40974 -19026 41026
rect -18974 40974 -18960 41026
rect -19040 40960 -18960 40974
rect -18880 41026 -18800 41040
rect -18880 40974 -18866 41026
rect -18814 40974 -18800 41026
rect -18880 40960 -18800 40974
rect -18720 41026 -18640 41040
rect -18720 40974 -18706 41026
rect -18654 40974 -18640 41026
rect -18720 40960 -18640 40974
rect -18560 41026 -18480 41040
rect -18560 40974 -18546 41026
rect -18494 40974 -18480 41026
rect -18560 40960 -18480 40974
rect -18400 41026 -18320 41040
rect -18400 40974 -18386 41026
rect -18334 40974 -18320 41026
rect -18400 40960 -18320 40974
rect -18240 41026 -18160 41040
rect -18240 40974 -18226 41026
rect -18174 40974 -18160 41026
rect -18240 40960 -18160 40974
rect -18080 41026 -18000 41040
rect -18080 40974 -18066 41026
rect -18014 40974 -18000 41026
rect -18080 40960 -18000 40974
rect -17920 41026 -17840 41040
rect -17920 40974 -17906 41026
rect -17854 40974 -17840 41026
rect -17920 40960 -17840 40974
rect -17760 41026 -17680 41040
rect -17760 40974 -17746 41026
rect -17694 40974 -17680 41026
rect -17760 40960 -17680 40974
rect -17600 41026 -17520 41040
rect -17600 40974 -17586 41026
rect -17534 40974 -17520 41026
rect -17600 40960 -17520 40974
rect -17440 41026 -17360 41040
rect -17440 40974 -17426 41026
rect -17374 40974 -17360 41026
rect -17440 40960 -17360 40974
rect -17280 41026 -17200 41040
rect -17280 40974 -17266 41026
rect -17214 40974 -17200 41026
rect -17280 40960 -17200 40974
rect -17120 41026 -17040 41040
rect -17120 40974 -17106 41026
rect -17054 40974 -17040 41026
rect -17120 40960 -17040 40974
rect -16960 41026 -16880 41040
rect -16960 40974 -16946 41026
rect -16894 40974 -16880 41026
rect -16960 40960 -16880 40974
rect -16800 41026 -16720 41040
rect -16800 40974 -16786 41026
rect -16734 40974 -16720 41026
rect -16800 40960 -16720 40974
rect -16640 41026 -16560 41040
rect -16640 40974 -16626 41026
rect -16574 40974 -16560 41026
rect -16640 40960 -16560 40974
rect -16480 41026 -16400 41040
rect -16480 40974 -16466 41026
rect -16414 40974 -16400 41026
rect -16480 40960 -16400 40974
rect -16320 41026 -16240 41040
rect -16320 40974 -16306 41026
rect -16254 40974 -16240 41026
rect -16320 40960 -16240 40974
rect -16160 41026 -16080 41040
rect -16160 40974 -16146 41026
rect -16094 40974 -16080 41026
rect -16160 40960 -16080 40974
rect -16000 41026 -15920 41040
rect -16000 40974 -15986 41026
rect -15934 40974 -15920 41026
rect -16000 40960 -15920 40974
rect -15840 41026 -15760 41040
rect -15840 40974 -15826 41026
rect -15774 40974 -15760 41026
rect -15840 40960 -15760 40974
rect -15680 41026 -15600 41040
rect -15680 40974 -15666 41026
rect -15614 40974 -15600 41026
rect -15680 40960 -15600 40974
rect -15520 41026 -15440 41040
rect -15520 40974 -15506 41026
rect -15454 40974 -15440 41026
rect -15520 40960 -15440 40974
rect -15360 41026 -15280 41040
rect -15360 40974 -15346 41026
rect -15294 40974 -15280 41026
rect -15360 40960 -15280 40974
rect -15200 41026 -15120 41040
rect -15200 40974 -15186 41026
rect -15134 40974 -15120 41026
rect -15200 40960 -15120 40974
rect -15040 41026 -14960 41040
rect -15040 40974 -15026 41026
rect -14974 40974 -14960 41026
rect -15040 40960 -14960 40974
rect -14880 41026 -14800 41040
rect -14880 40974 -14866 41026
rect -14814 40974 -14800 41026
rect -14880 40960 -14800 40974
rect -14720 41026 -14640 41040
rect -14720 40974 -14706 41026
rect -14654 40974 -14640 41026
rect -14720 40960 -14640 40974
rect -14560 41026 -14480 41040
rect -14560 40974 -14546 41026
rect -14494 40974 -14480 41026
rect -14560 40960 -14480 40974
rect -14400 41026 -14320 41040
rect -14400 40974 -14386 41026
rect -14334 40974 -14320 41026
rect -14400 40960 -14320 40974
rect -14240 41026 -14160 41040
rect -14240 40974 -14226 41026
rect -14174 40974 -14160 41026
rect -14240 40960 -14160 40974
rect -14080 41026 -14000 41040
rect -14080 40974 -14066 41026
rect -14014 40974 -14000 41026
rect -14080 40960 -14000 40974
rect -13920 41026 -13840 41040
rect -13920 40974 -13906 41026
rect -13854 40974 -13840 41026
rect -13920 40960 -13840 40974
rect -13760 41026 -13680 41040
rect -13760 40974 -13746 41026
rect -13694 40974 -13680 41026
rect -13760 40960 -13680 40974
rect -13600 41026 -13520 41040
rect -13600 40974 -13586 41026
rect -13534 40974 -13520 41026
rect -13600 40960 -13520 40974
rect -13440 41026 -13360 41040
rect -13440 40974 -13426 41026
rect -13374 40974 -13360 41026
rect -13440 40960 -13360 40974
rect -13280 41026 -13200 41040
rect -13280 40974 -13266 41026
rect -13214 40974 -13200 41026
rect -13280 40960 -13200 40974
rect -13120 41026 -13040 41040
rect -13120 40974 -13106 41026
rect -13054 40974 -13040 41026
rect -13120 40960 -13040 40974
rect -12960 41026 -12880 41040
rect -12960 40974 -12946 41026
rect -12894 40974 -12880 41026
rect -12960 40960 -12880 40974
rect -12800 41026 -12720 41040
rect -12800 40974 -12786 41026
rect -12734 40974 -12720 41026
rect -12800 40960 -12720 40974
rect -12640 41026 -12560 41040
rect -12640 40974 -12626 41026
rect -12574 40974 -12560 41026
rect -12640 40960 -12560 40974
rect -12480 41026 -12400 41040
rect -12480 40974 -12466 41026
rect -12414 40974 -12400 41026
rect -12480 40960 -12400 40974
rect -12320 41026 -12240 41040
rect -12320 40974 -12306 41026
rect -12254 40974 -12240 41026
rect -12320 40960 -12240 40974
rect -11360 41026 -11280 41040
rect -11360 40974 -11346 41026
rect -11294 40974 -11280 41026
rect -11360 40960 -11280 40974
rect -11200 41026 -11120 41040
rect -11200 40974 -11186 41026
rect -11134 40974 -11120 41026
rect -11200 40960 -11120 40974
rect -11040 41026 -10960 41040
rect -11040 40974 -11026 41026
rect -10974 40974 -10960 41026
rect -11040 40960 -10960 40974
rect -10880 41026 -10800 41040
rect -10880 40974 -10866 41026
rect -10814 40974 -10800 41026
rect -10880 40960 -10800 40974
rect -10720 41026 -10640 41040
rect -10720 40974 -10706 41026
rect -10654 40974 -10640 41026
rect -10720 40960 -10640 40974
rect -10560 41026 -10480 41040
rect -10560 40974 -10546 41026
rect -10494 40974 -10480 41026
rect -10560 40960 -10480 40974
rect -10400 41026 -10320 41040
rect -10400 40974 -10386 41026
rect -10334 40974 -10320 41026
rect -10400 40960 -10320 40974
rect -10240 41026 -10160 41040
rect -10240 40974 -10226 41026
rect -10174 40974 -10160 41026
rect -10240 40960 -10160 40974
rect -10080 41026 -10000 41040
rect -10080 40974 -10066 41026
rect -10014 40974 -10000 41026
rect -10080 40960 -10000 40974
rect -9920 41026 -9840 41040
rect -9920 40974 -9906 41026
rect -9854 40974 -9840 41026
rect -9920 40960 -9840 40974
rect -9760 41026 -9680 41040
rect -9760 40974 -9746 41026
rect -9694 40974 -9680 41026
rect -9760 40960 -9680 40974
rect -9600 41026 -9520 41040
rect -9600 40974 -9586 41026
rect -9534 40974 -9520 41026
rect -9600 40960 -9520 40974
rect -9440 41026 -9360 41040
rect -9440 40974 -9426 41026
rect -9374 40974 -9360 41026
rect -9440 40960 -9360 40974
rect -9280 41026 -9200 41040
rect -9280 40974 -9266 41026
rect -9214 40974 -9200 41026
rect -9280 40960 -9200 40974
rect -9120 41026 -9040 41040
rect -9120 40974 -9106 41026
rect -9054 40974 -9040 41026
rect -9120 40960 -9040 40974
rect -8960 41026 -8880 41040
rect -8960 40974 -8946 41026
rect -8894 40974 -8880 41026
rect -8960 40960 -8880 40974
rect -8800 41026 -8720 41040
rect -8800 40974 -8786 41026
rect -8734 40974 -8720 41026
rect -8800 40960 -8720 40974
rect -8640 41026 -8560 41040
rect -8640 40974 -8626 41026
rect -8574 40974 -8560 41026
rect -8640 40960 -8560 40974
rect -8480 41026 -8400 41040
rect -8480 40974 -8466 41026
rect -8414 40974 -8400 41026
rect -8480 40960 -8400 40974
rect -8320 41026 -8240 41040
rect -8320 40974 -8306 41026
rect -8254 40974 -8240 41026
rect -8320 40960 -8240 40974
rect -8160 41026 -8080 41040
rect -8160 40974 -8146 41026
rect -8094 40974 -8080 41026
rect -8160 40960 -8080 40974
rect -8000 41026 -7920 41040
rect -8000 40974 -7986 41026
rect -7934 40974 -7920 41026
rect -8000 40960 -7920 40974
rect -7840 41026 -7760 41040
rect -7840 40974 -7826 41026
rect -7774 40974 -7760 41026
rect -7840 40960 -7760 40974
rect -7680 41026 -7600 41040
rect -7680 40974 -7666 41026
rect -7614 40974 -7600 41026
rect -7680 40960 -7600 40974
rect -7520 41026 -7440 41040
rect -7520 40974 -7506 41026
rect -7454 40974 -7440 41026
rect -7520 40960 -7440 40974
rect -7360 41026 -7280 41040
rect -7360 40974 -7346 41026
rect -7294 40974 -7280 41026
rect -7360 40960 -7280 40974
rect -7200 41026 -7120 41040
rect -7200 40974 -7186 41026
rect -7134 40974 -7120 41026
rect -7200 40960 -7120 40974
rect -7040 41026 -6960 41040
rect -7040 40974 -7026 41026
rect -6974 40974 -6960 41026
rect -7040 40960 -6960 40974
rect -6880 41026 -6800 41040
rect -6880 40974 -6866 41026
rect -6814 40974 -6800 41026
rect -6880 40960 -6800 40974
rect -6720 41026 -6640 41040
rect -6720 40974 -6706 41026
rect -6654 40974 -6640 41026
rect -6720 40960 -6640 40974
rect -6560 41026 -6480 41040
rect -6560 40974 -6546 41026
rect -6494 40974 -6480 41026
rect -6560 40960 -6480 40974
rect -6400 41026 -6320 41040
rect -6400 40974 -6386 41026
rect -6334 40974 -6320 41026
rect -6400 40960 -6320 40974
rect -6240 41026 -6160 41040
rect -6240 40974 -6226 41026
rect -6174 40974 -6160 41026
rect -6240 40960 -6160 40974
rect -6080 41026 -6000 41040
rect -6080 40974 -6066 41026
rect -6014 40974 -6000 41026
rect -6080 40960 -6000 40974
rect -5920 41026 -5840 41040
rect -5920 40974 -5906 41026
rect -5854 40974 -5840 41026
rect -5920 40960 -5840 40974
rect -5760 41026 -5680 41040
rect -5760 40974 -5746 41026
rect -5694 40974 -5680 41026
rect -5760 40960 -5680 40974
rect -5600 41026 -5520 41040
rect -5600 40974 -5586 41026
rect -5534 40974 -5520 41026
rect -5600 40960 -5520 40974
rect -5440 41026 -5360 41040
rect -5440 40974 -5426 41026
rect -5374 40974 -5360 41026
rect -5440 40960 -5360 40974
rect -5280 41026 -5200 41040
rect -5280 40974 -5266 41026
rect -5214 40974 -5200 41026
rect -5280 40960 -5200 40974
rect -5120 41026 -5040 41040
rect -5120 40974 -5106 41026
rect -5054 40974 -5040 41026
rect -5120 40960 -5040 40974
rect -4960 41026 -4880 41040
rect -4960 40974 -4946 41026
rect -4894 40974 -4880 41026
rect -4960 40960 -4880 40974
rect -4800 41026 -4720 41040
rect -4800 40974 -4786 41026
rect -4734 40974 -4720 41026
rect -4800 40960 -4720 40974
rect -4640 41026 -4560 41040
rect -4640 40974 -4626 41026
rect -4574 40974 -4560 41026
rect -4640 40960 -4560 40974
rect -4480 41026 -4400 41040
rect -4480 40974 -4466 41026
rect -4414 40974 -4400 41026
rect -4480 40960 -4400 40974
rect -4320 41026 -4240 41040
rect -4320 40974 -4306 41026
rect -4254 40974 -4240 41026
rect -4320 40960 -4240 40974
rect -4160 41026 -4080 41040
rect -4160 40974 -4146 41026
rect -4094 40974 -4080 41026
rect -4160 40960 -4080 40974
rect -4000 41026 -3920 41040
rect -4000 40974 -3986 41026
rect -3934 40974 -3920 41026
rect -4000 40960 -3920 40974
rect -3840 41017 -3760 41040
rect -3840 40983 -3817 41017
rect -3783 40983 -3760 41017
rect -3840 40960 -3760 40983
rect -3680 41026 -3600 41040
rect -3680 40974 -3666 41026
rect -3614 40974 -3600 41026
rect -3680 40960 -3600 40974
rect -3520 41026 -3440 41040
rect -3520 40974 -3506 41026
rect -3454 40974 -3440 41026
rect -3520 40960 -3440 40974
rect 41040 41026 41120 41040
rect 41040 40974 41054 41026
rect 41106 40974 41120 41026
rect 41040 40960 41120 40974
rect 41200 41026 41280 41040
rect 41200 40974 41214 41026
rect 41266 40974 41280 41026
rect 41200 40960 41280 40974
rect 41360 41026 41440 41040
rect 41360 40974 41374 41026
rect 41426 40974 41440 41026
rect 41360 40960 41440 40974
rect 41520 41026 41600 41040
rect 41520 40974 41534 41026
rect 41586 40974 41600 41026
rect 41520 40960 41600 40974
rect 41680 41026 41760 41040
rect 41680 40974 41694 41026
rect 41746 40974 41760 41026
rect 41680 40960 41760 40974
rect 41840 41026 41920 41040
rect 41840 40974 41854 41026
rect 41906 40974 41920 41026
rect 41840 40960 41920 40974
rect 42000 41026 42080 41040
rect 42000 40974 42014 41026
rect 42066 40974 42080 41026
rect 42000 40960 42080 40974
rect 42160 41026 42240 41040
rect 42160 40974 42174 41026
rect 42226 40974 42240 41026
rect 42160 40960 42240 40974
rect 42320 41026 42400 41040
rect 42320 40974 42334 41026
rect 42386 40974 42400 41026
rect 42320 40960 42400 40974
rect 42480 41026 42560 41040
rect 42480 40974 42494 41026
rect 42546 40974 42560 41026
rect 42480 40960 42560 40974
rect 42640 41026 42720 41040
rect 42640 40974 42654 41026
rect 42706 40974 42720 41026
rect 42640 40960 42720 40974
rect 42800 41026 42880 41040
rect 42800 40974 42814 41026
rect 42866 40974 42880 41026
rect 42800 40960 42880 40974
rect 42960 41026 43040 41040
rect 42960 40974 42974 41026
rect 43026 40974 43040 41026
rect 42960 40960 43040 40974
rect 43120 41026 43200 41040
rect 43120 40974 43134 41026
rect 43186 40974 43200 41026
rect 43120 40960 43200 40974
rect -10560 40706 -10480 40720
rect -10560 40654 -10546 40706
rect -10494 40654 -10480 40706
rect -10560 40640 -10480 40654
rect -10240 40706 -10160 40720
rect -10240 40654 -10226 40706
rect -10174 40654 -10160 40706
rect -10240 40640 -10160 40654
rect -10080 40706 -10000 40720
rect -10080 40654 -10066 40706
rect -10014 40654 -10000 40706
rect -10080 40640 -10000 40654
rect -9920 40706 -9840 40720
rect -9920 40654 -9906 40706
rect -9854 40654 -9840 40706
rect -9920 40640 -9840 40654
rect -9760 40706 -9680 40720
rect -9760 40654 -9746 40706
rect -9694 40654 -9680 40706
rect -9760 40640 -9680 40654
rect -9600 40706 -9520 40720
rect -9600 40654 -9586 40706
rect -9534 40654 -9520 40706
rect -9600 40640 -9520 40654
rect -9440 40706 -9360 40720
rect -9440 40654 -9426 40706
rect -9374 40654 -9360 40706
rect -9440 40640 -9360 40654
rect -9280 40706 -9200 40720
rect -9280 40654 -9266 40706
rect -9214 40654 -9200 40706
rect -9280 40640 -9200 40654
rect -9120 40706 -9040 40720
rect -9120 40654 -9106 40706
rect -9054 40654 -9040 40706
rect -9120 40640 -9040 40654
rect -8960 40706 -8880 40720
rect -8960 40654 -8946 40706
rect -8894 40654 -8880 40706
rect -8960 40640 -8880 40654
rect -8800 40706 -8720 40720
rect -8800 40654 -8786 40706
rect -8734 40654 -8720 40706
rect -8800 40640 -8720 40654
rect -8640 40706 -8560 40720
rect -8640 40654 -8626 40706
rect -8574 40654 -8560 40706
rect -8640 40640 -8560 40654
rect -8480 40706 -8400 40720
rect -8480 40654 -8466 40706
rect -8414 40654 -8400 40706
rect -8480 40640 -8400 40654
rect -8320 40706 -8240 40720
rect -8320 40654 -8306 40706
rect -8254 40654 -8240 40706
rect -8320 40640 -8240 40654
rect -8160 40706 -8080 40720
rect -8160 40654 -8146 40706
rect -8094 40654 -8080 40706
rect -8160 40640 -8080 40654
rect -8000 40706 -7920 40720
rect -8000 40654 -7986 40706
rect -7934 40654 -7920 40706
rect -8000 40640 -7920 40654
rect -7840 40706 -7760 40720
rect -7840 40654 -7826 40706
rect -7774 40654 -7760 40706
rect -7840 40640 -7760 40654
rect -7680 40706 -7600 40720
rect -7680 40654 -7666 40706
rect -7614 40654 -7600 40706
rect -7680 40640 -7600 40654
rect -7520 40706 -7440 40720
rect -7520 40654 -7506 40706
rect -7454 40654 -7440 40706
rect -7520 40640 -7440 40654
rect -7360 40706 -7280 40720
rect -7360 40654 -7346 40706
rect -7294 40654 -7280 40706
rect -7360 40640 -7280 40654
rect -7200 40706 -7120 40720
rect -7200 40654 -7186 40706
rect -7134 40654 -7120 40706
rect -7200 40640 -7120 40654
rect -7040 40706 -6960 40720
rect -7040 40654 -7026 40706
rect -6974 40654 -6960 40706
rect -7040 40640 -6960 40654
rect -6880 40706 -6800 40720
rect -6880 40654 -6866 40706
rect -6814 40654 -6800 40706
rect -6880 40640 -6800 40654
rect -6720 40706 -6640 40720
rect -6720 40654 -6706 40706
rect -6654 40654 -6640 40706
rect -6720 40640 -6640 40654
rect -6560 40706 -6480 40720
rect -6560 40654 -6546 40706
rect -6494 40654 -6480 40706
rect -6560 40640 -6480 40654
rect -6400 40706 -6320 40720
rect -6400 40654 -6386 40706
rect -6334 40654 -6320 40706
rect -6400 40640 -6320 40654
rect -6240 40706 -6160 40720
rect -6240 40654 -6226 40706
rect -6174 40654 -6160 40706
rect -6240 40640 -6160 40654
rect -6080 40706 -6000 40720
rect -6080 40654 -6066 40706
rect -6014 40654 -6000 40706
rect -6080 40640 -6000 40654
rect -5920 40706 -5840 40720
rect -5920 40654 -5906 40706
rect -5854 40654 -5840 40706
rect -5920 40640 -5840 40654
rect -5760 40706 -5680 40720
rect -5760 40654 -5746 40706
rect -5694 40654 -5680 40706
rect -5760 40640 -5680 40654
rect -5600 40706 -5520 40720
rect -5600 40654 -5586 40706
rect -5534 40654 -5520 40706
rect -5600 40640 -5520 40654
rect -5440 40706 -5360 40720
rect -5440 40654 -5426 40706
rect -5374 40654 -5360 40706
rect -5440 40640 -5360 40654
rect -5280 40706 -5200 40720
rect -5280 40654 -5266 40706
rect -5214 40654 -5200 40706
rect -5280 40640 -5200 40654
rect -5120 40706 -5040 40720
rect -5120 40654 -5106 40706
rect -5054 40654 -5040 40706
rect -5120 40640 -5040 40654
rect -4960 40706 -4880 40720
rect -4960 40654 -4946 40706
rect -4894 40654 -4880 40706
rect -4960 40640 -4880 40654
rect -4800 40706 -4720 40720
rect -4800 40654 -4786 40706
rect -4734 40654 -4720 40706
rect -4800 40640 -4720 40654
rect -4640 40706 -4560 40720
rect -4640 40654 -4626 40706
rect -4574 40654 -4560 40706
rect -4640 40640 -4560 40654
rect -4480 40706 -4400 40720
rect -4480 40654 -4466 40706
rect -4414 40654 -4400 40706
rect -4480 40640 -4400 40654
rect -4320 40706 -4240 40720
rect -4320 40654 -4306 40706
rect -4254 40654 -4240 40706
rect -4320 40640 -4240 40654
rect -4160 40706 -4080 40720
rect -4160 40654 -4146 40706
rect -4094 40654 -4080 40706
rect -4160 40640 -4080 40654
rect -4000 40706 -3920 40720
rect -4000 40654 -3986 40706
rect -3934 40654 -3920 40706
rect -4000 40640 -3920 40654
rect -3680 40706 -3600 40720
rect -3680 40654 -3666 40706
rect -3614 40654 -3600 40706
rect -3680 40640 -3600 40654
rect -3520 40706 -3440 40720
rect -3520 40654 -3506 40706
rect -3454 40654 -3440 40706
rect -3520 40640 -3440 40654
rect -10560 40386 -10480 40400
rect -10560 40334 -10546 40386
rect -10494 40334 -10480 40386
rect -10560 40320 -10480 40334
rect -10240 40386 -10160 40400
rect -10240 40334 -10226 40386
rect -10174 40334 -10160 40386
rect -10240 40320 -10160 40334
rect -10080 40386 -10000 40400
rect -10080 40334 -10066 40386
rect -10014 40334 -10000 40386
rect -10080 40320 -10000 40334
rect -9920 40386 -9840 40400
rect -9920 40334 -9906 40386
rect -9854 40334 -9840 40386
rect -9920 40320 -9840 40334
rect -9760 40386 -9680 40400
rect -9760 40334 -9746 40386
rect -9694 40334 -9680 40386
rect -9760 40320 -9680 40334
rect -9600 40386 -9520 40400
rect -9600 40334 -9586 40386
rect -9534 40334 -9520 40386
rect -9600 40320 -9520 40334
rect -9440 40386 -9360 40400
rect -9440 40334 -9426 40386
rect -9374 40334 -9360 40386
rect -9440 40320 -9360 40334
rect -9280 40386 -9200 40400
rect -9280 40334 -9266 40386
rect -9214 40334 -9200 40386
rect -9280 40320 -9200 40334
rect -9120 40386 -9040 40400
rect -9120 40334 -9106 40386
rect -9054 40334 -9040 40386
rect -9120 40320 -9040 40334
rect -8960 40386 -8880 40400
rect -8960 40334 -8946 40386
rect -8894 40334 -8880 40386
rect -8960 40320 -8880 40334
rect -8800 40386 -8720 40400
rect -8800 40334 -8786 40386
rect -8734 40334 -8720 40386
rect -8800 40320 -8720 40334
rect -8640 40386 -8560 40400
rect -8640 40334 -8626 40386
rect -8574 40334 -8560 40386
rect -8640 40320 -8560 40334
rect -8480 40386 -8400 40400
rect -8480 40334 -8466 40386
rect -8414 40334 -8400 40386
rect -8480 40320 -8400 40334
rect -8320 40386 -8240 40400
rect -8320 40334 -8306 40386
rect -8254 40334 -8240 40386
rect -8320 40320 -8240 40334
rect -8160 40386 -8080 40400
rect -8160 40334 -8146 40386
rect -8094 40334 -8080 40386
rect -8160 40320 -8080 40334
rect -8000 40386 -7920 40400
rect -8000 40334 -7986 40386
rect -7934 40334 -7920 40386
rect -8000 40320 -7920 40334
rect -7840 40386 -7760 40400
rect -7840 40334 -7826 40386
rect -7774 40334 -7760 40386
rect -7840 40320 -7760 40334
rect -7680 40386 -7600 40400
rect -7680 40334 -7666 40386
rect -7614 40334 -7600 40386
rect -7680 40320 -7600 40334
rect -7520 40386 -7440 40400
rect -7520 40334 -7506 40386
rect -7454 40334 -7440 40386
rect -7520 40320 -7440 40334
rect -7360 40386 -7280 40400
rect -7360 40334 -7346 40386
rect -7294 40334 -7280 40386
rect -7360 40320 -7280 40334
rect -7200 40386 -7120 40400
rect -7200 40334 -7186 40386
rect -7134 40334 -7120 40386
rect -7200 40320 -7120 40334
rect -7040 40386 -6960 40400
rect -7040 40334 -7026 40386
rect -6974 40334 -6960 40386
rect -7040 40320 -6960 40334
rect -6880 40386 -6800 40400
rect -6880 40334 -6866 40386
rect -6814 40334 -6800 40386
rect -6880 40320 -6800 40334
rect -6720 40386 -6640 40400
rect -6720 40334 -6706 40386
rect -6654 40334 -6640 40386
rect -6720 40320 -6640 40334
rect -6560 40386 -6480 40400
rect -6560 40334 -6546 40386
rect -6494 40334 -6480 40386
rect -6560 40320 -6480 40334
rect -6400 40386 -6320 40400
rect -6400 40334 -6386 40386
rect -6334 40334 -6320 40386
rect -6400 40320 -6320 40334
rect -6240 40386 -6160 40400
rect -6240 40334 -6226 40386
rect -6174 40334 -6160 40386
rect -6240 40320 -6160 40334
rect -6080 40386 -6000 40400
rect -6080 40334 -6066 40386
rect -6014 40334 -6000 40386
rect -6080 40320 -6000 40334
rect -5920 40386 -5840 40400
rect -5920 40334 -5906 40386
rect -5854 40334 -5840 40386
rect -5920 40320 -5840 40334
rect -5760 40386 -5680 40400
rect -5760 40334 -5746 40386
rect -5694 40334 -5680 40386
rect -5760 40320 -5680 40334
rect -5600 40386 -5520 40400
rect -5600 40334 -5586 40386
rect -5534 40334 -5520 40386
rect -5600 40320 -5520 40334
rect -5440 40386 -5360 40400
rect -5440 40334 -5426 40386
rect -5374 40334 -5360 40386
rect -5440 40320 -5360 40334
rect -5280 40386 -5200 40400
rect -5280 40334 -5266 40386
rect -5214 40334 -5200 40386
rect -5280 40320 -5200 40334
rect -5120 40386 -5040 40400
rect -5120 40334 -5106 40386
rect -5054 40334 -5040 40386
rect -5120 40320 -5040 40334
rect -4960 40386 -4880 40400
rect -4960 40334 -4946 40386
rect -4894 40334 -4880 40386
rect -4960 40320 -4880 40334
rect -4800 40386 -4720 40400
rect -4800 40334 -4786 40386
rect -4734 40334 -4720 40386
rect -4800 40320 -4720 40334
rect -4640 40386 -4560 40400
rect -4640 40334 -4626 40386
rect -4574 40334 -4560 40386
rect -4640 40320 -4560 40334
rect -4480 40386 -4400 40400
rect -4480 40334 -4466 40386
rect -4414 40334 -4400 40386
rect -4480 40320 -4400 40334
rect -4320 40386 -4240 40400
rect -4320 40334 -4306 40386
rect -4254 40334 -4240 40386
rect -4320 40320 -4240 40334
rect -4160 40386 -4080 40400
rect -4160 40334 -4146 40386
rect -4094 40334 -4080 40386
rect -4160 40320 -4080 40334
rect -4000 40386 -3920 40400
rect -4000 40334 -3986 40386
rect -3934 40334 -3920 40386
rect -4000 40320 -3920 40334
rect -3680 40386 -3600 40400
rect -3680 40334 -3666 40386
rect -3614 40334 -3600 40386
rect -3680 40320 -3600 40334
rect -3520 40386 -3440 40400
rect -3520 40334 -3506 40386
rect -3454 40334 -3440 40386
rect -3520 40320 -3440 40334
rect 41040 40066 41120 40080
rect 41040 40014 41054 40066
rect 41106 40014 41120 40066
rect 41040 40000 41120 40014
rect 41200 40066 41280 40080
rect 41200 40014 41214 40066
rect 41266 40014 41280 40066
rect 41200 40000 41280 40014
rect 41360 40066 41440 40080
rect 41360 40014 41374 40066
rect 41426 40014 41440 40066
rect 41360 40000 41440 40014
rect 41520 40066 41600 40080
rect 41520 40014 41534 40066
rect 41586 40014 41600 40066
rect 41520 40000 41600 40014
rect 41680 40066 41760 40080
rect 41680 40014 41694 40066
rect 41746 40014 41760 40066
rect 41680 40000 41760 40014
rect 41840 40066 41920 40080
rect 41840 40014 41854 40066
rect 41906 40014 41920 40066
rect 41840 40000 41920 40014
rect 42000 40066 42080 40080
rect 42000 40014 42014 40066
rect 42066 40014 42080 40066
rect 42000 40000 42080 40014
rect 42160 40066 42240 40080
rect 42160 40014 42174 40066
rect 42226 40014 42240 40066
rect 42160 40000 42240 40014
rect 42320 40066 42400 40080
rect 42320 40014 42334 40066
rect 42386 40014 42400 40066
rect 42320 40000 42400 40014
rect 42480 40066 42560 40080
rect 42480 40014 42494 40066
rect 42546 40014 42560 40066
rect 42480 40000 42560 40014
rect 42640 40066 42720 40080
rect 42640 40014 42654 40066
rect 42706 40014 42720 40066
rect 42640 40000 42720 40014
rect 42800 40066 42880 40080
rect 42800 40014 42814 40066
rect 42866 40014 42880 40066
rect 42800 40000 42880 40014
rect 42960 40066 43040 40080
rect 42960 40014 42974 40066
rect 43026 40014 43040 40066
rect 42960 40000 43040 40014
rect 43120 40066 43200 40080
rect 43120 40014 43134 40066
rect 43186 40014 43200 40066
rect 43120 40000 43200 40014
rect 41040 39746 41120 39760
rect 41040 39694 41054 39746
rect 41106 39694 41120 39746
rect 41040 39680 41120 39694
rect 41200 39746 41280 39760
rect 41200 39694 41214 39746
rect 41266 39694 41280 39746
rect 41200 39680 41280 39694
rect 41360 39746 41440 39760
rect 41360 39694 41374 39746
rect 41426 39694 41440 39746
rect 41360 39680 41440 39694
rect 41520 39746 41600 39760
rect 41520 39694 41534 39746
rect 41586 39694 41600 39746
rect 41520 39680 41600 39694
rect 41680 39746 41760 39760
rect 41680 39694 41694 39746
rect 41746 39694 41760 39746
rect 41680 39680 41760 39694
rect 41840 39746 41920 39760
rect 41840 39694 41854 39746
rect 41906 39694 41920 39746
rect 41840 39680 41920 39694
rect 42000 39746 42080 39760
rect 42000 39694 42014 39746
rect 42066 39694 42080 39746
rect 42000 39680 42080 39694
rect 42160 39746 42240 39760
rect 42160 39694 42174 39746
rect 42226 39694 42240 39746
rect 42160 39680 42240 39694
rect 42320 39746 42400 39760
rect 42320 39694 42334 39746
rect 42386 39694 42400 39746
rect 42320 39680 42400 39694
rect 42480 39746 42560 39760
rect 42480 39694 42494 39746
rect 42546 39694 42560 39746
rect 42480 39680 42560 39694
rect 42640 39746 42720 39760
rect 42640 39694 42654 39746
rect 42706 39694 42720 39746
rect 42640 39680 42720 39694
rect 42800 39746 42880 39760
rect 42800 39694 42814 39746
rect 42866 39694 42880 39746
rect 42800 39680 42880 39694
rect 42960 39746 43040 39760
rect 42960 39694 42974 39746
rect 43026 39694 43040 39746
rect 42960 39680 43040 39694
rect 43120 39746 43200 39760
rect 43120 39694 43134 39746
rect 43186 39694 43200 39746
rect 43120 39680 43200 39694
rect -33120 37746 -33040 37760
rect -33120 37694 -33106 37746
rect -33054 37694 -33040 37746
rect -33120 37680 -33040 37694
rect -32960 37746 -32880 37760
rect -32960 37694 -32946 37746
rect -32894 37694 -32880 37746
rect -32960 37680 -32880 37694
rect -32800 37746 -32720 37760
rect -32800 37694 -32786 37746
rect -32734 37694 -32720 37746
rect -32800 37680 -32720 37694
rect -32640 37746 -32560 37760
rect -32640 37694 -32626 37746
rect -32574 37694 -32560 37746
rect -32640 37680 -32560 37694
rect -32480 37746 -32400 37760
rect -32480 37694 -32466 37746
rect -32414 37694 -32400 37746
rect -32480 37680 -32400 37694
rect -32320 37746 -32240 37760
rect -32320 37694 -32306 37746
rect -32254 37694 -32240 37746
rect -32320 37680 -32240 37694
rect -32160 37746 -32080 37760
rect -32160 37694 -32146 37746
rect -32094 37694 -32080 37746
rect -32160 37680 -32080 37694
rect -32000 37746 -31920 37760
rect -32000 37694 -31986 37746
rect -31934 37694 -31920 37746
rect -32000 37680 -31920 37694
rect -31840 37746 -31760 37760
rect -31840 37694 -31826 37746
rect -31774 37694 -31760 37746
rect -31840 37680 -31760 37694
rect -31680 37746 -31600 37760
rect -31680 37694 -31666 37746
rect -31614 37694 -31600 37746
rect -31680 37680 -31600 37694
rect -31520 37746 -31440 37760
rect -31520 37694 -31506 37746
rect -31454 37694 -31440 37746
rect -31520 37680 -31440 37694
rect -31360 37746 -31280 37760
rect -31360 37694 -31346 37746
rect -31294 37694 -31280 37746
rect -31360 37680 -31280 37694
rect -31200 37746 -31120 37760
rect -31200 37694 -31186 37746
rect -31134 37694 -31120 37746
rect -31200 37680 -31120 37694
rect -33120 37426 -33040 37440
rect -33120 37374 -33106 37426
rect -33054 37374 -33040 37426
rect -33120 37360 -33040 37374
rect -32960 37426 -32880 37440
rect -32960 37374 -32946 37426
rect -32894 37374 -32880 37426
rect -32960 37360 -32880 37374
rect -32800 37426 -32720 37440
rect -32800 37374 -32786 37426
rect -32734 37374 -32720 37426
rect -32800 37360 -32720 37374
rect -32640 37426 -32560 37440
rect -32640 37374 -32626 37426
rect -32574 37374 -32560 37426
rect -32640 37360 -32560 37374
rect -32480 37426 -32400 37440
rect -32480 37374 -32466 37426
rect -32414 37374 -32400 37426
rect -32480 37360 -32400 37374
rect -32320 37426 -32240 37440
rect -32320 37374 -32306 37426
rect -32254 37374 -32240 37426
rect -32320 37360 -32240 37374
rect -32160 37426 -32080 37440
rect -32160 37374 -32146 37426
rect -32094 37374 -32080 37426
rect -32160 37360 -32080 37374
rect -32000 37426 -31920 37440
rect -32000 37374 -31986 37426
rect -31934 37374 -31920 37426
rect -32000 37360 -31920 37374
rect -31840 37426 -31760 37440
rect -31840 37374 -31826 37426
rect -31774 37374 -31760 37426
rect -31840 37360 -31760 37374
rect -31680 37426 -31600 37440
rect -31680 37374 -31666 37426
rect -31614 37374 -31600 37426
rect -31680 37360 -31600 37374
rect -31520 37426 -31440 37440
rect -31520 37374 -31506 37426
rect -31454 37374 -31440 37426
rect -31520 37360 -31440 37374
rect -31360 37426 -31280 37440
rect -31360 37374 -31346 37426
rect -31294 37374 -31280 37426
rect -31360 37360 -31280 37374
rect -31200 37426 -31120 37440
rect -31200 37374 -31186 37426
rect -31134 37374 -31120 37426
rect -31200 37360 -31120 37374
rect -33120 37106 -33040 37120
rect -33120 37054 -33106 37106
rect -33054 37054 -33040 37106
rect -33120 37040 -33040 37054
rect -32960 37106 -32880 37120
rect -32960 37054 -32946 37106
rect -32894 37054 -32880 37106
rect -32960 37040 -32880 37054
rect -32800 37106 -32720 37120
rect -32800 37054 -32786 37106
rect -32734 37054 -32720 37106
rect -32800 37040 -32720 37054
rect -32640 37106 -32560 37120
rect -32640 37054 -32626 37106
rect -32574 37054 -32560 37106
rect -32640 37040 -32560 37054
rect -32480 37106 -32400 37120
rect -32480 37054 -32466 37106
rect -32414 37054 -32400 37106
rect -32480 37040 -32400 37054
rect -32320 37106 -32240 37120
rect -32320 37054 -32306 37106
rect -32254 37054 -32240 37106
rect -32320 37040 -32240 37054
rect -32160 37106 -32080 37120
rect -32160 37054 -32146 37106
rect -32094 37054 -32080 37106
rect -32160 37040 -32080 37054
rect -32000 37106 -31920 37120
rect -32000 37054 -31986 37106
rect -31934 37054 -31920 37106
rect -32000 37040 -31920 37054
rect -31840 37106 -31760 37120
rect -31840 37054 -31826 37106
rect -31774 37054 -31760 37106
rect -31840 37040 -31760 37054
rect -31680 37106 -31600 37120
rect -31680 37054 -31666 37106
rect -31614 37054 -31600 37106
rect -31680 37040 -31600 37054
rect -31520 37106 -31440 37120
rect -31520 37054 -31506 37106
rect -31454 37054 -31440 37106
rect -31520 37040 -31440 37054
rect -31360 37106 -31280 37120
rect -31360 37054 -31346 37106
rect -31294 37054 -31280 37106
rect -31360 37040 -31280 37054
rect -31200 37106 -31120 37120
rect -31200 37054 -31186 37106
rect -31134 37054 -31120 37106
rect -31200 37040 -31120 37054
rect 41040 36066 41120 36080
rect 41040 36014 41054 36066
rect 41106 36014 41120 36066
rect 41040 36000 41120 36014
rect 41200 36066 41280 36080
rect 41200 36014 41214 36066
rect 41266 36014 41280 36066
rect 41200 36000 41280 36014
rect 41360 36066 41440 36080
rect 41360 36014 41374 36066
rect 41426 36014 41440 36066
rect 41360 36000 41440 36014
rect 41520 36066 41600 36080
rect 41520 36014 41534 36066
rect 41586 36014 41600 36066
rect 41520 36000 41600 36014
rect 41680 36066 41760 36080
rect 41680 36014 41694 36066
rect 41746 36014 41760 36066
rect 41680 36000 41760 36014
rect 41840 36066 41920 36080
rect 41840 36014 41854 36066
rect 41906 36014 41920 36066
rect 41840 36000 41920 36014
rect 42000 36066 42080 36080
rect 42000 36014 42014 36066
rect 42066 36014 42080 36066
rect 42000 36000 42080 36014
rect 42160 36066 42240 36080
rect 42160 36014 42174 36066
rect 42226 36014 42240 36066
rect 42160 36000 42240 36014
rect 42320 36066 42400 36080
rect 42320 36014 42334 36066
rect 42386 36014 42400 36066
rect 42320 36000 42400 36014
rect 42480 36066 42560 36080
rect 42480 36014 42494 36066
rect 42546 36014 42560 36066
rect 42480 36000 42560 36014
rect 42640 36066 42720 36080
rect 42640 36014 42654 36066
rect 42706 36014 42720 36066
rect 42640 36000 42720 36014
rect 42800 36066 42880 36080
rect 42800 36014 42814 36066
rect 42866 36014 42880 36066
rect 42800 36000 42880 36014
rect 42960 36066 43040 36080
rect 42960 36014 42974 36066
rect 43026 36014 43040 36066
rect 42960 36000 43040 36014
rect 43120 36066 43200 36080
rect 43120 36014 43134 36066
rect 43186 36014 43200 36066
rect 43120 36000 43200 36014
rect 41040 35746 41120 35760
rect 41040 35694 41054 35746
rect 41106 35694 41120 35746
rect 41040 35680 41120 35694
rect 41200 35746 41280 35760
rect 41200 35694 41214 35746
rect 41266 35694 41280 35746
rect 41200 35680 41280 35694
rect 41360 35746 41440 35760
rect 41360 35694 41374 35746
rect 41426 35694 41440 35746
rect 41360 35680 41440 35694
rect 41520 35746 41600 35760
rect 41520 35694 41534 35746
rect 41586 35694 41600 35746
rect 41520 35680 41600 35694
rect 41680 35746 41760 35760
rect 41680 35694 41694 35746
rect 41746 35694 41760 35746
rect 41680 35680 41760 35694
rect 41840 35746 41920 35760
rect 41840 35694 41854 35746
rect 41906 35694 41920 35746
rect 41840 35680 41920 35694
rect 42000 35746 42080 35760
rect 42000 35694 42014 35746
rect 42066 35694 42080 35746
rect 42000 35680 42080 35694
rect 42160 35746 42240 35760
rect 42160 35694 42174 35746
rect 42226 35694 42240 35746
rect 42160 35680 42240 35694
rect 42320 35746 42400 35760
rect 42320 35694 42334 35746
rect 42386 35694 42400 35746
rect 42320 35680 42400 35694
rect 42480 35746 42560 35760
rect 42480 35694 42494 35746
rect 42546 35694 42560 35746
rect 42480 35680 42560 35694
rect 42640 35746 42720 35760
rect 42640 35694 42654 35746
rect 42706 35694 42720 35746
rect 42640 35680 42720 35694
rect 42800 35746 42880 35760
rect 42800 35694 42814 35746
rect 42866 35694 42880 35746
rect 42800 35680 42880 35694
rect 42960 35746 43040 35760
rect 42960 35694 42974 35746
rect 43026 35694 43040 35746
rect 42960 35680 43040 35694
rect 43120 35746 43200 35760
rect 43120 35694 43134 35746
rect 43186 35694 43200 35746
rect 43120 35680 43200 35694
rect -33120 34706 -33040 34720
rect -33120 34654 -33106 34706
rect -33054 34654 -33040 34706
rect -33120 34640 -33040 34654
rect -32960 34706 -32880 34720
rect -32960 34654 -32946 34706
rect -32894 34654 -32880 34706
rect -32960 34640 -32880 34654
rect -32800 34706 -32720 34720
rect -32800 34654 -32786 34706
rect -32734 34654 -32720 34706
rect -32800 34640 -32720 34654
rect -32640 34706 -32560 34720
rect -32640 34654 -32626 34706
rect -32574 34654 -32560 34706
rect -32640 34640 -32560 34654
rect -32480 34706 -32400 34720
rect -32480 34654 -32466 34706
rect -32414 34654 -32400 34706
rect -32480 34640 -32400 34654
rect -32320 34706 -32240 34720
rect -32320 34654 -32306 34706
rect -32254 34654 -32240 34706
rect -32320 34640 -32240 34654
rect -32160 34706 -32080 34720
rect -32160 34654 -32146 34706
rect -32094 34654 -32080 34706
rect -32160 34640 -32080 34654
rect -32000 34706 -31920 34720
rect -32000 34654 -31986 34706
rect -31934 34654 -31920 34706
rect -32000 34640 -31920 34654
rect -31840 34706 -31760 34720
rect -31840 34654 -31826 34706
rect -31774 34654 -31760 34706
rect -31840 34640 -31760 34654
rect -31680 34706 -31600 34720
rect -31680 34654 -31666 34706
rect -31614 34654 -31600 34706
rect -31680 34640 -31600 34654
rect -31520 34706 -31440 34720
rect -31520 34654 -31506 34706
rect -31454 34654 -31440 34706
rect -31520 34640 -31440 34654
rect -31360 34706 -31280 34720
rect -31360 34654 -31346 34706
rect -31294 34654 -31280 34706
rect -31360 34640 -31280 34654
rect -31200 34706 -31120 34720
rect -31200 34654 -31186 34706
rect -31134 34654 -31120 34706
rect -31200 34640 -31120 34654
rect -29920 34706 -29840 34720
rect -29920 34654 -29906 34706
rect -29854 34654 -29840 34706
rect -29920 34640 -29840 34654
rect -29760 34706 -29680 34720
rect -29760 34654 -29746 34706
rect -29694 34654 -29680 34706
rect -29760 34640 -29680 34654
rect -29600 34706 -29520 34720
rect -29600 34654 -29586 34706
rect -29534 34654 -29520 34706
rect -29600 34640 -29520 34654
rect -29440 34706 -29360 34720
rect -29440 34654 -29426 34706
rect -29374 34654 -29360 34706
rect -29440 34640 -29360 34654
rect -29280 34706 -29200 34720
rect -29280 34654 -29266 34706
rect -29214 34654 -29200 34706
rect -29280 34640 -29200 34654
rect -29120 34706 -29040 34720
rect -29120 34654 -29106 34706
rect -29054 34654 -29040 34706
rect -29120 34640 -29040 34654
rect -28960 34706 -28880 34720
rect -28960 34654 -28946 34706
rect -28894 34654 -28880 34706
rect -28960 34640 -28880 34654
rect -28800 34706 -28720 34720
rect -28800 34654 -28786 34706
rect -28734 34654 -28720 34706
rect -28800 34640 -28720 34654
rect -28640 34706 -28560 34720
rect -28640 34654 -28626 34706
rect -28574 34654 -28560 34706
rect -28640 34640 -28560 34654
rect -28480 34706 -28400 34720
rect -28480 34654 -28466 34706
rect -28414 34654 -28400 34706
rect -28480 34640 -28400 34654
rect -28320 34706 -28240 34720
rect -28320 34654 -28306 34706
rect -28254 34654 -28240 34706
rect -28320 34640 -28240 34654
rect -28160 34706 -28080 34720
rect -28160 34654 -28146 34706
rect -28094 34654 -28080 34706
rect -28160 34640 -28080 34654
rect -28000 34706 -27920 34720
rect -28000 34654 -27986 34706
rect -27934 34654 -27920 34706
rect -28000 34640 -27920 34654
rect -27840 34706 -27760 34720
rect -27840 34654 -27826 34706
rect -27774 34654 -27760 34706
rect -27840 34640 -27760 34654
rect -27680 34706 -27600 34720
rect -27680 34654 -27666 34706
rect -27614 34654 -27600 34706
rect -27680 34640 -27600 34654
rect -27520 34706 -27440 34720
rect -27520 34654 -27506 34706
rect -27454 34654 -27440 34706
rect -27520 34640 -27440 34654
rect -27360 34706 -27280 34720
rect -27360 34654 -27346 34706
rect -27294 34654 -27280 34706
rect -27360 34640 -27280 34654
rect -27200 34706 -27120 34720
rect -27200 34654 -27186 34706
rect -27134 34654 -27120 34706
rect -27200 34640 -27120 34654
rect -27040 34706 -26960 34720
rect -27040 34654 -27026 34706
rect -26974 34654 -26960 34706
rect -27040 34640 -26960 34654
rect -26880 34706 -26800 34720
rect -26880 34654 -26866 34706
rect -26814 34654 -26800 34706
rect -26880 34640 -26800 34654
rect -26720 34706 -26640 34720
rect -26720 34654 -26706 34706
rect -26654 34654 -26640 34706
rect -26720 34640 -26640 34654
rect -26560 34706 -26480 34720
rect -26560 34654 -26546 34706
rect -26494 34654 -26480 34706
rect -26560 34640 -26480 34654
rect -26400 34706 -26320 34720
rect -26400 34654 -26386 34706
rect -26334 34654 -26320 34706
rect -26400 34640 -26320 34654
rect -26240 34706 -26160 34720
rect -26240 34654 -26226 34706
rect -26174 34654 -26160 34706
rect -26240 34640 -26160 34654
rect -26080 34706 -26000 34720
rect -26080 34654 -26066 34706
rect -26014 34654 -26000 34706
rect -26080 34640 -26000 34654
rect -25920 34706 -25840 34720
rect -25920 34654 -25906 34706
rect -25854 34654 -25840 34706
rect -25920 34640 -25840 34654
rect -25760 34706 -25680 34720
rect -25760 34654 -25746 34706
rect -25694 34654 -25680 34706
rect -25760 34640 -25680 34654
rect -25600 34706 -25520 34720
rect -25600 34654 -25586 34706
rect -25534 34654 -25520 34706
rect -25600 34640 -25520 34654
rect -25440 34706 -25360 34720
rect -25440 34654 -25426 34706
rect -25374 34654 -25360 34706
rect -25440 34640 -25360 34654
rect -25280 34706 -25200 34720
rect -25280 34654 -25266 34706
rect -25214 34654 -25200 34706
rect -25280 34640 -25200 34654
rect -25120 34706 -25040 34720
rect -25120 34654 -25106 34706
rect -25054 34654 -25040 34706
rect -25120 34640 -25040 34654
rect -24960 34706 -24880 34720
rect -24960 34654 -24946 34706
rect -24894 34654 -24880 34706
rect -24960 34640 -24880 34654
rect -24800 34706 -24720 34720
rect -24800 34654 -24786 34706
rect -24734 34654 -24720 34706
rect -24800 34640 -24720 34654
rect -24640 34706 -24560 34720
rect -24640 34654 -24626 34706
rect -24574 34654 -24560 34706
rect -24640 34640 -24560 34654
rect -24480 34706 -24400 34720
rect -24480 34654 -24466 34706
rect -24414 34654 -24400 34706
rect -24480 34640 -24400 34654
rect -24320 34706 -24240 34720
rect -24320 34654 -24306 34706
rect -24254 34654 -24240 34706
rect -24320 34640 -24240 34654
rect -24160 34706 -24080 34720
rect -24160 34654 -24146 34706
rect -24094 34654 -24080 34706
rect -24160 34640 -24080 34654
rect -24000 34706 -23920 34720
rect -24000 34654 -23986 34706
rect -23934 34654 -23920 34706
rect -24000 34640 -23920 34654
rect -23840 34706 -23760 34720
rect -23840 34654 -23826 34706
rect -23774 34654 -23760 34706
rect -23840 34640 -23760 34654
rect -23680 34706 -23600 34720
rect -23680 34654 -23666 34706
rect -23614 34654 -23600 34706
rect -23680 34640 -23600 34654
rect -23520 34706 -23440 34720
rect -23520 34654 -23506 34706
rect -23454 34654 -23440 34706
rect -23520 34640 -23440 34654
rect -23360 34706 -23280 34720
rect -23360 34654 -23346 34706
rect -23294 34654 -23280 34706
rect -23360 34640 -23280 34654
rect -23200 34706 -23120 34720
rect -23200 34654 -23186 34706
rect -23134 34654 -23120 34706
rect -23200 34640 -23120 34654
rect -23040 34706 -22960 34720
rect -23040 34654 -23026 34706
rect -22974 34654 -22960 34706
rect -23040 34640 -22960 34654
rect -22880 34706 -22800 34720
rect -22880 34654 -22866 34706
rect -22814 34654 -22800 34706
rect -22880 34640 -22800 34654
rect -22720 34706 -22640 34720
rect -22720 34654 -22706 34706
rect -22654 34654 -22640 34706
rect -22720 34640 -22640 34654
rect -22560 34706 -22480 34720
rect -22560 34654 -22546 34706
rect -22494 34654 -22480 34706
rect -22560 34640 -22480 34654
rect -22400 34706 -22320 34720
rect -22400 34654 -22386 34706
rect -22334 34654 -22320 34706
rect -22400 34640 -22320 34654
rect -22240 34706 -22160 34720
rect -22240 34654 -22226 34706
rect -22174 34654 -22160 34706
rect -22240 34640 -22160 34654
rect -22080 34706 -22000 34720
rect -22080 34654 -22066 34706
rect -22014 34654 -22000 34706
rect -22080 34640 -22000 34654
rect -21920 34706 -21840 34720
rect -21920 34654 -21906 34706
rect -21854 34654 -21840 34706
rect -21920 34640 -21840 34654
rect -21760 34706 -21680 34720
rect -21760 34654 -21746 34706
rect -21694 34654 -21680 34706
rect -21760 34640 -21680 34654
rect -21600 34706 -21520 34720
rect -21600 34654 -21586 34706
rect -21534 34654 -21520 34706
rect -21600 34640 -21520 34654
rect -21440 34706 -21360 34720
rect -21440 34654 -21426 34706
rect -21374 34654 -21360 34706
rect -21440 34640 -21360 34654
rect -21280 34706 -21200 34720
rect -21280 34654 -21266 34706
rect -21214 34654 -21200 34706
rect -21280 34640 -21200 34654
rect -21120 34706 -21040 34720
rect -21120 34654 -21106 34706
rect -21054 34654 -21040 34706
rect -21120 34640 -21040 34654
rect -20960 34706 -20880 34720
rect -20960 34654 -20946 34706
rect -20894 34654 -20880 34706
rect -20960 34640 -20880 34654
rect -20800 34706 -20720 34720
rect -20800 34654 -20786 34706
rect -20734 34654 -20720 34706
rect -20800 34640 -20720 34654
rect -20640 34706 -20560 34720
rect -20640 34654 -20626 34706
rect -20574 34654 -20560 34706
rect -20640 34640 -20560 34654
rect -20480 34706 -20400 34720
rect -20480 34654 -20466 34706
rect -20414 34654 -20400 34706
rect -20480 34640 -20400 34654
rect -20320 34706 -20240 34720
rect -20320 34654 -20306 34706
rect -20254 34654 -20240 34706
rect -20320 34640 -20240 34654
rect -20160 34706 -20080 34720
rect -20160 34654 -20146 34706
rect -20094 34654 -20080 34706
rect -20160 34640 -20080 34654
rect -20000 34706 -19920 34720
rect -20000 34654 -19986 34706
rect -19934 34654 -19920 34706
rect -20000 34640 -19920 34654
rect -19840 34706 -19760 34720
rect -19840 34654 -19826 34706
rect -19774 34654 -19760 34706
rect -19840 34640 -19760 34654
rect -19680 34706 -19600 34720
rect -19680 34654 -19666 34706
rect -19614 34654 -19600 34706
rect -19680 34640 -19600 34654
rect -19520 34706 -19440 34720
rect -19520 34654 -19506 34706
rect -19454 34654 -19440 34706
rect -19520 34640 -19440 34654
rect -19360 34706 -19280 34720
rect -19360 34654 -19346 34706
rect -19294 34654 -19280 34706
rect -19360 34640 -19280 34654
rect -19200 34706 -19120 34720
rect -19200 34654 -19186 34706
rect -19134 34654 -19120 34706
rect -19200 34640 -19120 34654
rect -19040 34706 -18960 34720
rect -19040 34654 -19026 34706
rect -18974 34654 -18960 34706
rect -19040 34640 -18960 34654
rect -18880 34706 -18800 34720
rect -18880 34654 -18866 34706
rect -18814 34654 -18800 34706
rect -18880 34640 -18800 34654
rect -18720 34706 -18640 34720
rect -18720 34654 -18706 34706
rect -18654 34654 -18640 34706
rect -18720 34640 -18640 34654
rect -18560 34706 -18480 34720
rect -18560 34654 -18546 34706
rect -18494 34654 -18480 34706
rect -18560 34640 -18480 34654
rect -18400 34706 -18320 34720
rect -18400 34654 -18386 34706
rect -18334 34654 -18320 34706
rect -18400 34640 -18320 34654
rect -18240 34706 -18160 34720
rect -18240 34654 -18226 34706
rect -18174 34654 -18160 34706
rect -18240 34640 -18160 34654
rect -18080 34706 -18000 34720
rect -18080 34654 -18066 34706
rect -18014 34654 -18000 34706
rect -18080 34640 -18000 34654
rect -17920 34706 -17840 34720
rect -17920 34654 -17906 34706
rect -17854 34654 -17840 34706
rect -17920 34640 -17840 34654
rect -17760 34706 -17680 34720
rect -17760 34654 -17746 34706
rect -17694 34654 -17680 34706
rect -17760 34640 -17680 34654
rect -17600 34706 -17520 34720
rect -17600 34654 -17586 34706
rect -17534 34654 -17520 34706
rect -17600 34640 -17520 34654
rect -17440 34706 -17360 34720
rect -17440 34654 -17426 34706
rect -17374 34654 -17360 34706
rect -17440 34640 -17360 34654
rect -17280 34706 -17200 34720
rect -17280 34654 -17266 34706
rect -17214 34654 -17200 34706
rect -17280 34640 -17200 34654
rect -17120 34706 -17040 34720
rect -17120 34654 -17106 34706
rect -17054 34654 -17040 34706
rect -17120 34640 -17040 34654
rect -16960 34706 -16880 34720
rect -16960 34654 -16946 34706
rect -16894 34654 -16880 34706
rect -16960 34640 -16880 34654
rect -16800 34706 -16720 34720
rect -16800 34654 -16786 34706
rect -16734 34654 -16720 34706
rect -16800 34640 -16720 34654
rect -16640 34706 -16560 34720
rect -16640 34654 -16626 34706
rect -16574 34654 -16560 34706
rect -16640 34640 -16560 34654
rect -16480 34706 -16400 34720
rect -16480 34654 -16466 34706
rect -16414 34654 -16400 34706
rect -16480 34640 -16400 34654
rect -16320 34706 -16240 34720
rect -16320 34654 -16306 34706
rect -16254 34654 -16240 34706
rect -16320 34640 -16240 34654
rect -16160 34706 -16080 34720
rect -16160 34654 -16146 34706
rect -16094 34654 -16080 34706
rect -16160 34640 -16080 34654
rect -16000 34706 -15920 34720
rect -16000 34654 -15986 34706
rect -15934 34654 -15920 34706
rect -16000 34640 -15920 34654
rect -15840 34706 -15760 34720
rect -15840 34654 -15826 34706
rect -15774 34654 -15760 34706
rect -15840 34640 -15760 34654
rect -15680 34706 -15600 34720
rect -15680 34654 -15666 34706
rect -15614 34654 -15600 34706
rect -15680 34640 -15600 34654
rect -15520 34706 -15440 34720
rect -15520 34654 -15506 34706
rect -15454 34654 -15440 34706
rect -15520 34640 -15440 34654
rect -15360 34706 -15280 34720
rect -15360 34654 -15346 34706
rect -15294 34654 -15280 34706
rect -15360 34640 -15280 34654
rect -15200 34706 -15120 34720
rect -15200 34654 -15186 34706
rect -15134 34654 -15120 34706
rect -15200 34640 -15120 34654
rect -15040 34706 -14960 34720
rect -15040 34654 -15026 34706
rect -14974 34654 -14960 34706
rect -15040 34640 -14960 34654
rect -14880 34706 -14800 34720
rect -14880 34654 -14866 34706
rect -14814 34654 -14800 34706
rect -14880 34640 -14800 34654
rect -14720 34706 -14640 34720
rect -14720 34654 -14706 34706
rect -14654 34654 -14640 34706
rect -14720 34640 -14640 34654
rect -14560 34706 -14480 34720
rect -14560 34654 -14546 34706
rect -14494 34654 -14480 34706
rect -14560 34640 -14480 34654
rect -14400 34706 -14320 34720
rect -14400 34654 -14386 34706
rect -14334 34654 -14320 34706
rect -14400 34640 -14320 34654
rect -14240 34706 -14160 34720
rect -14240 34654 -14226 34706
rect -14174 34654 -14160 34706
rect -14240 34640 -14160 34654
rect -14080 34706 -14000 34720
rect -14080 34654 -14066 34706
rect -14014 34654 -14000 34706
rect -14080 34640 -14000 34654
rect -13920 34706 -13840 34720
rect -13920 34654 -13906 34706
rect -13854 34654 -13840 34706
rect -13920 34640 -13840 34654
rect -13760 34706 -13680 34720
rect -13760 34654 -13746 34706
rect -13694 34654 -13680 34706
rect -13760 34640 -13680 34654
rect -13600 34706 -13520 34720
rect -13600 34654 -13586 34706
rect -13534 34654 -13520 34706
rect -13600 34640 -13520 34654
rect -13440 34706 -13360 34720
rect -13440 34654 -13426 34706
rect -13374 34654 -13360 34706
rect -13440 34640 -13360 34654
rect -13280 34706 -13200 34720
rect -13280 34654 -13266 34706
rect -13214 34654 -13200 34706
rect -13280 34640 -13200 34654
rect -13120 34706 -13040 34720
rect -13120 34654 -13106 34706
rect -13054 34654 -13040 34706
rect -13120 34640 -13040 34654
rect -12960 34706 -12880 34720
rect -12960 34654 -12946 34706
rect -12894 34654 -12880 34706
rect -12960 34640 -12880 34654
rect -12800 34706 -12720 34720
rect -12800 34654 -12786 34706
rect -12734 34654 -12720 34706
rect -12800 34640 -12720 34654
rect -12640 34706 -12560 34720
rect -12640 34654 -12626 34706
rect -12574 34654 -12560 34706
rect -12640 34640 -12560 34654
rect -12480 34706 -12400 34720
rect -12480 34654 -12466 34706
rect -12414 34654 -12400 34706
rect -12480 34640 -12400 34654
rect -12320 34706 -12240 34720
rect -12320 34654 -12306 34706
rect -12254 34654 -12240 34706
rect -12320 34640 -12240 34654
rect -12160 34706 -12080 34720
rect -12160 34654 -12146 34706
rect -12094 34654 -12080 34706
rect -12160 34640 -12080 34654
rect -12000 34706 -11920 34720
rect -12000 34654 -11986 34706
rect -11934 34654 -11920 34706
rect -12000 34640 -11920 34654
rect -11840 34706 -11760 34720
rect -11840 34654 -11826 34706
rect -11774 34654 -11760 34706
rect -11840 34640 -11760 34654
rect -11680 34706 -11600 34720
rect -11680 34654 -11666 34706
rect -11614 34654 -11600 34706
rect -11680 34640 -11600 34654
rect -11520 34706 -11440 34720
rect -11520 34654 -11506 34706
rect -11454 34654 -11440 34706
rect -11520 34640 -11440 34654
rect -10880 34706 -10800 34720
rect -10880 34654 -10866 34706
rect -10814 34654 -10800 34706
rect -10880 34640 -10800 34654
rect -10560 34706 -10480 34720
rect -10560 34654 -10546 34706
rect -10494 34654 -10480 34706
rect -10560 34640 -10480 34654
rect -33120 34386 -33040 34400
rect -33120 34334 -33106 34386
rect -33054 34334 -33040 34386
rect -33120 34320 -33040 34334
rect -32960 34386 -32880 34400
rect -32960 34334 -32946 34386
rect -32894 34334 -32880 34386
rect -32960 34320 -32880 34334
rect -32800 34386 -32720 34400
rect -32800 34334 -32786 34386
rect -32734 34334 -32720 34386
rect -32800 34320 -32720 34334
rect -32640 34386 -32560 34400
rect -32640 34334 -32626 34386
rect -32574 34334 -32560 34386
rect -32640 34320 -32560 34334
rect -32480 34386 -32400 34400
rect -32480 34334 -32466 34386
rect -32414 34334 -32400 34386
rect -32480 34320 -32400 34334
rect -32320 34386 -32240 34400
rect -32320 34334 -32306 34386
rect -32254 34334 -32240 34386
rect -32320 34320 -32240 34334
rect -32160 34386 -32080 34400
rect -32160 34334 -32146 34386
rect -32094 34334 -32080 34386
rect -32160 34320 -32080 34334
rect -32000 34386 -31920 34400
rect -32000 34334 -31986 34386
rect -31934 34334 -31920 34386
rect -32000 34320 -31920 34334
rect -31840 34386 -31760 34400
rect -31840 34334 -31826 34386
rect -31774 34334 -31760 34386
rect -31840 34320 -31760 34334
rect -31680 34386 -31600 34400
rect -31680 34334 -31666 34386
rect -31614 34334 -31600 34386
rect -31680 34320 -31600 34334
rect -31520 34386 -31440 34400
rect -31520 34334 -31506 34386
rect -31454 34334 -31440 34386
rect -31520 34320 -31440 34334
rect -31360 34386 -31280 34400
rect -31360 34334 -31346 34386
rect -31294 34334 -31280 34386
rect -31360 34320 -31280 34334
rect -31200 34386 -31120 34400
rect -31200 34334 -31186 34386
rect -31134 34334 -31120 34386
rect -31200 34320 -31120 34334
rect -29920 34386 -29840 34400
rect -29920 34334 -29906 34386
rect -29854 34334 -29840 34386
rect -29920 34320 -29840 34334
rect -29760 34386 -29680 34400
rect -29760 34334 -29746 34386
rect -29694 34334 -29680 34386
rect -29760 34320 -29680 34334
rect -29600 34386 -29520 34400
rect -29600 34334 -29586 34386
rect -29534 34334 -29520 34386
rect -29600 34320 -29520 34334
rect -29440 34386 -29360 34400
rect -29440 34334 -29426 34386
rect -29374 34334 -29360 34386
rect -29440 34320 -29360 34334
rect -29280 34386 -29200 34400
rect -29280 34334 -29266 34386
rect -29214 34334 -29200 34386
rect -29280 34320 -29200 34334
rect -29120 34386 -29040 34400
rect -29120 34334 -29106 34386
rect -29054 34334 -29040 34386
rect -29120 34320 -29040 34334
rect -28960 34386 -28880 34400
rect -28960 34334 -28946 34386
rect -28894 34334 -28880 34386
rect -28960 34320 -28880 34334
rect -28800 34386 -28720 34400
rect -28800 34334 -28786 34386
rect -28734 34334 -28720 34386
rect -28800 34320 -28720 34334
rect -28640 34386 -28560 34400
rect -28640 34334 -28626 34386
rect -28574 34334 -28560 34386
rect -28640 34320 -28560 34334
rect -28480 34386 -28400 34400
rect -28480 34334 -28466 34386
rect -28414 34334 -28400 34386
rect -28480 34320 -28400 34334
rect -28320 34386 -28240 34400
rect -28320 34334 -28306 34386
rect -28254 34334 -28240 34386
rect -28320 34320 -28240 34334
rect -28160 34386 -28080 34400
rect -28160 34334 -28146 34386
rect -28094 34334 -28080 34386
rect -28160 34320 -28080 34334
rect -28000 34386 -27920 34400
rect -28000 34334 -27986 34386
rect -27934 34334 -27920 34386
rect -28000 34320 -27920 34334
rect -27840 34386 -27760 34400
rect -27840 34334 -27826 34386
rect -27774 34334 -27760 34386
rect -27840 34320 -27760 34334
rect -27680 34386 -27600 34400
rect -27680 34334 -27666 34386
rect -27614 34334 -27600 34386
rect -27680 34320 -27600 34334
rect -27520 34386 -27440 34400
rect -27520 34334 -27506 34386
rect -27454 34334 -27440 34386
rect -27520 34320 -27440 34334
rect -27360 34386 -27280 34400
rect -27360 34334 -27346 34386
rect -27294 34334 -27280 34386
rect -27360 34320 -27280 34334
rect -27200 34386 -27120 34400
rect -27200 34334 -27186 34386
rect -27134 34334 -27120 34386
rect -27200 34320 -27120 34334
rect -27040 34386 -26960 34400
rect -27040 34334 -27026 34386
rect -26974 34334 -26960 34386
rect -27040 34320 -26960 34334
rect -26880 34386 -26800 34400
rect -26880 34334 -26866 34386
rect -26814 34334 -26800 34386
rect -26880 34320 -26800 34334
rect -26720 34386 -26640 34400
rect -26720 34334 -26706 34386
rect -26654 34334 -26640 34386
rect -26720 34320 -26640 34334
rect -26560 34386 -26480 34400
rect -26560 34334 -26546 34386
rect -26494 34334 -26480 34386
rect -26560 34320 -26480 34334
rect -26400 34386 -26320 34400
rect -26400 34334 -26386 34386
rect -26334 34334 -26320 34386
rect -26400 34320 -26320 34334
rect -26240 34386 -26160 34400
rect -26240 34334 -26226 34386
rect -26174 34334 -26160 34386
rect -26240 34320 -26160 34334
rect -26080 34386 -26000 34400
rect -26080 34334 -26066 34386
rect -26014 34334 -26000 34386
rect -26080 34320 -26000 34334
rect -25920 34386 -25840 34400
rect -25920 34334 -25906 34386
rect -25854 34334 -25840 34386
rect -25920 34320 -25840 34334
rect -25760 34386 -25680 34400
rect -25760 34334 -25746 34386
rect -25694 34334 -25680 34386
rect -25760 34320 -25680 34334
rect -25600 34386 -25520 34400
rect -25600 34334 -25586 34386
rect -25534 34334 -25520 34386
rect -25600 34320 -25520 34334
rect -25440 34386 -25360 34400
rect -25440 34334 -25426 34386
rect -25374 34334 -25360 34386
rect -25440 34320 -25360 34334
rect -25280 34386 -25200 34400
rect -25280 34334 -25266 34386
rect -25214 34334 -25200 34386
rect -25280 34320 -25200 34334
rect -25120 34386 -25040 34400
rect -25120 34334 -25106 34386
rect -25054 34334 -25040 34386
rect -25120 34320 -25040 34334
rect -24960 34386 -24880 34400
rect -24960 34334 -24946 34386
rect -24894 34334 -24880 34386
rect -24960 34320 -24880 34334
rect -24800 34386 -24720 34400
rect -24800 34334 -24786 34386
rect -24734 34334 -24720 34386
rect -24800 34320 -24720 34334
rect -24640 34386 -24560 34400
rect -24640 34334 -24626 34386
rect -24574 34334 -24560 34386
rect -24640 34320 -24560 34334
rect -24480 34386 -24400 34400
rect -24480 34334 -24466 34386
rect -24414 34334 -24400 34386
rect -24480 34320 -24400 34334
rect -24320 34386 -24240 34400
rect -24320 34334 -24306 34386
rect -24254 34334 -24240 34386
rect -24320 34320 -24240 34334
rect -24160 34386 -24080 34400
rect -24160 34334 -24146 34386
rect -24094 34334 -24080 34386
rect -24160 34320 -24080 34334
rect -24000 34386 -23920 34400
rect -24000 34334 -23986 34386
rect -23934 34334 -23920 34386
rect -24000 34320 -23920 34334
rect -23840 34386 -23760 34400
rect -23840 34334 -23826 34386
rect -23774 34334 -23760 34386
rect -23840 34320 -23760 34334
rect -23680 34386 -23600 34400
rect -23680 34334 -23666 34386
rect -23614 34334 -23600 34386
rect -23680 34320 -23600 34334
rect -23520 34386 -23440 34400
rect -23520 34334 -23506 34386
rect -23454 34334 -23440 34386
rect -23520 34320 -23440 34334
rect -23360 34386 -23280 34400
rect -23360 34334 -23346 34386
rect -23294 34334 -23280 34386
rect -23360 34320 -23280 34334
rect -23200 34386 -23120 34400
rect -23200 34334 -23186 34386
rect -23134 34334 -23120 34386
rect -23200 34320 -23120 34334
rect -23040 34386 -22960 34400
rect -23040 34334 -23026 34386
rect -22974 34334 -22960 34386
rect -23040 34320 -22960 34334
rect -22880 34386 -22800 34400
rect -22880 34334 -22866 34386
rect -22814 34334 -22800 34386
rect -22880 34320 -22800 34334
rect -22720 34386 -22640 34400
rect -22720 34334 -22706 34386
rect -22654 34334 -22640 34386
rect -22720 34320 -22640 34334
rect -22560 34386 -22480 34400
rect -22560 34334 -22546 34386
rect -22494 34334 -22480 34386
rect -22560 34320 -22480 34334
rect -22400 34386 -22320 34400
rect -22400 34334 -22386 34386
rect -22334 34334 -22320 34386
rect -22400 34320 -22320 34334
rect -22240 34386 -22160 34400
rect -22240 34334 -22226 34386
rect -22174 34334 -22160 34386
rect -22240 34320 -22160 34334
rect -22080 34386 -22000 34400
rect -22080 34334 -22066 34386
rect -22014 34334 -22000 34386
rect -22080 34320 -22000 34334
rect -21920 34386 -21840 34400
rect -21920 34334 -21906 34386
rect -21854 34334 -21840 34386
rect -21920 34320 -21840 34334
rect -21760 34386 -21680 34400
rect -21760 34334 -21746 34386
rect -21694 34334 -21680 34386
rect -21760 34320 -21680 34334
rect -21600 34386 -21520 34400
rect -21600 34334 -21586 34386
rect -21534 34334 -21520 34386
rect -21600 34320 -21520 34334
rect -21440 34386 -21360 34400
rect -21440 34334 -21426 34386
rect -21374 34334 -21360 34386
rect -21440 34320 -21360 34334
rect -21280 34386 -21200 34400
rect -21280 34334 -21266 34386
rect -21214 34334 -21200 34386
rect -21280 34320 -21200 34334
rect -21120 34386 -21040 34400
rect -21120 34334 -21106 34386
rect -21054 34334 -21040 34386
rect -21120 34320 -21040 34334
rect -20960 34386 -20880 34400
rect -20960 34334 -20946 34386
rect -20894 34334 -20880 34386
rect -20960 34320 -20880 34334
rect -20800 34386 -20720 34400
rect -20800 34334 -20786 34386
rect -20734 34334 -20720 34386
rect -20800 34320 -20720 34334
rect -20640 34386 -20560 34400
rect -20640 34334 -20626 34386
rect -20574 34334 -20560 34386
rect -20640 34320 -20560 34334
rect -20480 34386 -20400 34400
rect -20480 34334 -20466 34386
rect -20414 34334 -20400 34386
rect -20480 34320 -20400 34334
rect -20320 34386 -20240 34400
rect -20320 34334 -20306 34386
rect -20254 34334 -20240 34386
rect -20320 34320 -20240 34334
rect -20160 34386 -20080 34400
rect -20160 34334 -20146 34386
rect -20094 34334 -20080 34386
rect -20160 34320 -20080 34334
rect -20000 34386 -19920 34400
rect -20000 34334 -19986 34386
rect -19934 34334 -19920 34386
rect -20000 34320 -19920 34334
rect -19840 34386 -19760 34400
rect -19840 34334 -19826 34386
rect -19774 34334 -19760 34386
rect -19840 34320 -19760 34334
rect -19680 34386 -19600 34400
rect -19680 34334 -19666 34386
rect -19614 34334 -19600 34386
rect -19680 34320 -19600 34334
rect -19520 34386 -19440 34400
rect -19520 34334 -19506 34386
rect -19454 34334 -19440 34386
rect -19520 34320 -19440 34334
rect -19360 34386 -19280 34400
rect -19360 34334 -19346 34386
rect -19294 34334 -19280 34386
rect -19360 34320 -19280 34334
rect -19200 34386 -19120 34400
rect -19200 34334 -19186 34386
rect -19134 34334 -19120 34386
rect -19200 34320 -19120 34334
rect -19040 34386 -18960 34400
rect -19040 34334 -19026 34386
rect -18974 34334 -18960 34386
rect -19040 34320 -18960 34334
rect -18880 34386 -18800 34400
rect -18880 34334 -18866 34386
rect -18814 34334 -18800 34386
rect -18880 34320 -18800 34334
rect -18720 34386 -18640 34400
rect -18720 34334 -18706 34386
rect -18654 34334 -18640 34386
rect -18720 34320 -18640 34334
rect -18560 34386 -18480 34400
rect -18560 34334 -18546 34386
rect -18494 34334 -18480 34386
rect -18560 34320 -18480 34334
rect -18400 34386 -18320 34400
rect -18400 34334 -18386 34386
rect -18334 34334 -18320 34386
rect -18400 34320 -18320 34334
rect -18240 34386 -18160 34400
rect -18240 34334 -18226 34386
rect -18174 34334 -18160 34386
rect -18240 34320 -18160 34334
rect -18080 34386 -18000 34400
rect -18080 34334 -18066 34386
rect -18014 34334 -18000 34386
rect -18080 34320 -18000 34334
rect -17920 34386 -17840 34400
rect -17920 34334 -17906 34386
rect -17854 34334 -17840 34386
rect -17920 34320 -17840 34334
rect -17760 34386 -17680 34400
rect -17760 34334 -17746 34386
rect -17694 34334 -17680 34386
rect -17760 34320 -17680 34334
rect -17600 34386 -17520 34400
rect -17600 34334 -17586 34386
rect -17534 34334 -17520 34386
rect -17600 34320 -17520 34334
rect -17440 34386 -17360 34400
rect -17440 34334 -17426 34386
rect -17374 34334 -17360 34386
rect -17440 34320 -17360 34334
rect -17280 34386 -17200 34400
rect -17280 34334 -17266 34386
rect -17214 34334 -17200 34386
rect -17280 34320 -17200 34334
rect -17120 34386 -17040 34400
rect -17120 34334 -17106 34386
rect -17054 34334 -17040 34386
rect -17120 34320 -17040 34334
rect -16960 34386 -16880 34400
rect -16960 34334 -16946 34386
rect -16894 34334 -16880 34386
rect -16960 34320 -16880 34334
rect -16800 34386 -16720 34400
rect -16800 34334 -16786 34386
rect -16734 34334 -16720 34386
rect -16800 34320 -16720 34334
rect -16640 34386 -16560 34400
rect -16640 34334 -16626 34386
rect -16574 34334 -16560 34386
rect -16640 34320 -16560 34334
rect -16480 34386 -16400 34400
rect -16480 34334 -16466 34386
rect -16414 34334 -16400 34386
rect -16480 34320 -16400 34334
rect -16320 34386 -16240 34400
rect -16320 34334 -16306 34386
rect -16254 34334 -16240 34386
rect -16320 34320 -16240 34334
rect -16160 34386 -16080 34400
rect -16160 34334 -16146 34386
rect -16094 34334 -16080 34386
rect -16160 34320 -16080 34334
rect -16000 34386 -15920 34400
rect -16000 34334 -15986 34386
rect -15934 34334 -15920 34386
rect -16000 34320 -15920 34334
rect -15840 34386 -15760 34400
rect -15840 34334 -15826 34386
rect -15774 34334 -15760 34386
rect -15840 34320 -15760 34334
rect -15680 34386 -15600 34400
rect -15680 34334 -15666 34386
rect -15614 34334 -15600 34386
rect -15680 34320 -15600 34334
rect -15520 34386 -15440 34400
rect -15520 34334 -15506 34386
rect -15454 34334 -15440 34386
rect -15520 34320 -15440 34334
rect -15360 34386 -15280 34400
rect -15360 34334 -15346 34386
rect -15294 34334 -15280 34386
rect -15360 34320 -15280 34334
rect -15200 34386 -15120 34400
rect -15200 34334 -15186 34386
rect -15134 34334 -15120 34386
rect -15200 34320 -15120 34334
rect -15040 34386 -14960 34400
rect -15040 34334 -15026 34386
rect -14974 34334 -14960 34386
rect -15040 34320 -14960 34334
rect -14880 34386 -14800 34400
rect -14880 34334 -14866 34386
rect -14814 34334 -14800 34386
rect -14880 34320 -14800 34334
rect -14720 34386 -14640 34400
rect -14720 34334 -14706 34386
rect -14654 34334 -14640 34386
rect -14720 34320 -14640 34334
rect -14560 34386 -14480 34400
rect -14560 34334 -14546 34386
rect -14494 34334 -14480 34386
rect -14560 34320 -14480 34334
rect -14400 34386 -14320 34400
rect -14400 34334 -14386 34386
rect -14334 34334 -14320 34386
rect -14400 34320 -14320 34334
rect -14240 34386 -14160 34400
rect -14240 34334 -14226 34386
rect -14174 34334 -14160 34386
rect -14240 34320 -14160 34334
rect -14080 34386 -14000 34400
rect -14080 34334 -14066 34386
rect -14014 34334 -14000 34386
rect -14080 34320 -14000 34334
rect -13920 34386 -13840 34400
rect -13920 34334 -13906 34386
rect -13854 34334 -13840 34386
rect -13920 34320 -13840 34334
rect -13760 34386 -13680 34400
rect -13760 34334 -13746 34386
rect -13694 34334 -13680 34386
rect -13760 34320 -13680 34334
rect -13600 34386 -13520 34400
rect -13600 34334 -13586 34386
rect -13534 34334 -13520 34386
rect -13600 34320 -13520 34334
rect -13440 34386 -13360 34400
rect -13440 34334 -13426 34386
rect -13374 34334 -13360 34386
rect -13440 34320 -13360 34334
rect -13280 34386 -13200 34400
rect -13280 34334 -13266 34386
rect -13214 34334 -13200 34386
rect -13280 34320 -13200 34334
rect -13120 34386 -13040 34400
rect -13120 34334 -13106 34386
rect -13054 34334 -13040 34386
rect -13120 34320 -13040 34334
rect -12960 34386 -12880 34400
rect -12960 34334 -12946 34386
rect -12894 34334 -12880 34386
rect -12960 34320 -12880 34334
rect -12800 34386 -12720 34400
rect -12800 34334 -12786 34386
rect -12734 34334 -12720 34386
rect -12800 34320 -12720 34334
rect -12640 34386 -12560 34400
rect -12640 34334 -12626 34386
rect -12574 34334 -12560 34386
rect -12640 34320 -12560 34334
rect -12480 34386 -12400 34400
rect -12480 34334 -12466 34386
rect -12414 34334 -12400 34386
rect -12480 34320 -12400 34334
rect -12320 34386 -12240 34400
rect -12320 34334 -12306 34386
rect -12254 34334 -12240 34386
rect -12320 34320 -12240 34334
rect -12160 34386 -12080 34400
rect -12160 34334 -12146 34386
rect -12094 34334 -12080 34386
rect -12160 34320 -12080 34334
rect -12000 34386 -11920 34400
rect -12000 34334 -11986 34386
rect -11934 34334 -11920 34386
rect -12000 34320 -11920 34334
rect -11840 34386 -11760 34400
rect -11840 34334 -11826 34386
rect -11774 34334 -11760 34386
rect -11840 34320 -11760 34334
rect -11680 34386 -11600 34400
rect -11680 34334 -11666 34386
rect -11614 34334 -11600 34386
rect -11680 34320 -11600 34334
rect -11520 34386 -11440 34400
rect -11520 34334 -11506 34386
rect -11454 34334 -11440 34386
rect -11520 34320 -11440 34334
rect -10880 34386 -10800 34400
rect -10880 34334 -10866 34386
rect -10814 34334 -10800 34386
rect -10880 34320 -10800 34334
rect -10560 34386 -10480 34400
rect -10560 34334 -10546 34386
rect -10494 34334 -10480 34386
rect -10560 34320 -10480 34334
rect -29920 32946 -29840 32960
rect -29920 32894 -29906 32946
rect -29854 32894 -29840 32946
rect -29920 32880 -29840 32894
rect -29760 32946 -29680 32960
rect -29760 32894 -29746 32946
rect -29694 32894 -29680 32946
rect -29760 32880 -29680 32894
rect -29600 32946 -29520 32960
rect -29600 32894 -29586 32946
rect -29534 32894 -29520 32946
rect -29600 32880 -29520 32894
rect -29440 32946 -29360 32960
rect -29440 32894 -29426 32946
rect -29374 32894 -29360 32946
rect -29440 32880 -29360 32894
rect -29280 32946 -29200 32960
rect -29280 32894 -29266 32946
rect -29214 32894 -29200 32946
rect -29280 32880 -29200 32894
rect -29120 32946 -29040 32960
rect -29120 32894 -29106 32946
rect -29054 32894 -29040 32946
rect -29120 32880 -29040 32894
rect -28960 32946 -28880 32960
rect -28960 32894 -28946 32946
rect -28894 32894 -28880 32946
rect -28960 32880 -28880 32894
rect -28800 32946 -28720 32960
rect -28800 32894 -28786 32946
rect -28734 32894 -28720 32946
rect -28800 32880 -28720 32894
rect -28640 32946 -28560 32960
rect -28640 32894 -28626 32946
rect -28574 32894 -28560 32946
rect -28640 32880 -28560 32894
rect -28480 32946 -28400 32960
rect -28480 32894 -28466 32946
rect -28414 32894 -28400 32946
rect -28480 32880 -28400 32894
rect -28320 32946 -28240 32960
rect -28320 32894 -28306 32946
rect -28254 32894 -28240 32946
rect -28320 32880 -28240 32894
rect -28160 32946 -28080 32960
rect -28160 32894 -28146 32946
rect -28094 32894 -28080 32946
rect -28160 32880 -28080 32894
rect -28000 32946 -27920 32960
rect -28000 32894 -27986 32946
rect -27934 32894 -27920 32946
rect -28000 32880 -27920 32894
rect -27840 32946 -27760 32960
rect -27840 32894 -27826 32946
rect -27774 32894 -27760 32946
rect -27840 32880 -27760 32894
rect -27680 32946 -27600 32960
rect -27680 32894 -27666 32946
rect -27614 32894 -27600 32946
rect -27680 32880 -27600 32894
rect -27520 32946 -27440 32960
rect -27520 32894 -27506 32946
rect -27454 32894 -27440 32946
rect -27520 32880 -27440 32894
rect -27360 32946 -27280 32960
rect -27360 32894 -27346 32946
rect -27294 32894 -27280 32946
rect -27360 32880 -27280 32894
rect -27200 32946 -27120 32960
rect -27200 32894 -27186 32946
rect -27134 32894 -27120 32946
rect -27200 32880 -27120 32894
rect -27040 32946 -26960 32960
rect -27040 32894 -27026 32946
rect -26974 32894 -26960 32946
rect -27040 32880 -26960 32894
rect -26880 32946 -26800 32960
rect -26880 32894 -26866 32946
rect -26814 32894 -26800 32946
rect -26880 32880 -26800 32894
rect -26720 32946 -26640 32960
rect -26720 32894 -26706 32946
rect -26654 32894 -26640 32946
rect -26720 32880 -26640 32894
rect -26560 32946 -26480 32960
rect -26560 32894 -26546 32946
rect -26494 32894 -26480 32946
rect -26560 32880 -26480 32894
rect -26400 32946 -26320 32960
rect -26400 32894 -26386 32946
rect -26334 32894 -26320 32946
rect -26400 32880 -26320 32894
rect -26240 32946 -26160 32960
rect -26240 32894 -26226 32946
rect -26174 32894 -26160 32946
rect -26240 32880 -26160 32894
rect -26080 32946 -26000 32960
rect -26080 32894 -26066 32946
rect -26014 32894 -26000 32946
rect -26080 32880 -26000 32894
rect -25920 32946 -25840 32960
rect -25920 32894 -25906 32946
rect -25854 32894 -25840 32946
rect -25920 32880 -25840 32894
rect -25760 32946 -25680 32960
rect -25760 32894 -25746 32946
rect -25694 32894 -25680 32946
rect -25760 32880 -25680 32894
rect -25600 32946 -25520 32960
rect -25600 32894 -25586 32946
rect -25534 32894 -25520 32946
rect -25600 32880 -25520 32894
rect -25440 32946 -25360 32960
rect -25440 32894 -25426 32946
rect -25374 32894 -25360 32946
rect -25440 32880 -25360 32894
rect -25280 32946 -25200 32960
rect -25280 32894 -25266 32946
rect -25214 32894 -25200 32946
rect -25280 32880 -25200 32894
rect -25120 32946 -25040 32960
rect -25120 32894 -25106 32946
rect -25054 32894 -25040 32946
rect -25120 32880 -25040 32894
rect -24960 32946 -24880 32960
rect -24960 32894 -24946 32946
rect -24894 32894 -24880 32946
rect -24960 32880 -24880 32894
rect -24800 32946 -24720 32960
rect -24800 32894 -24786 32946
rect -24734 32894 -24720 32946
rect -24800 32880 -24720 32894
rect -24640 32946 -24560 32960
rect -24640 32894 -24626 32946
rect -24574 32894 -24560 32946
rect -24640 32880 -24560 32894
rect -24480 32946 -24400 32960
rect -24480 32894 -24466 32946
rect -24414 32894 -24400 32946
rect -24480 32880 -24400 32894
rect -24320 32946 -24240 32960
rect -24320 32894 -24306 32946
rect -24254 32894 -24240 32946
rect -24320 32880 -24240 32894
rect -24160 32946 -24080 32960
rect -24160 32894 -24146 32946
rect -24094 32894 -24080 32946
rect -24160 32880 -24080 32894
rect -24000 32946 -23920 32960
rect -24000 32894 -23986 32946
rect -23934 32894 -23920 32946
rect -24000 32880 -23920 32894
rect -23840 32946 -23760 32960
rect -23840 32894 -23826 32946
rect -23774 32894 -23760 32946
rect -23840 32880 -23760 32894
rect -23680 32946 -23600 32960
rect -23680 32894 -23666 32946
rect -23614 32894 -23600 32946
rect -23680 32880 -23600 32894
rect -23520 32946 -23440 32960
rect -23520 32894 -23506 32946
rect -23454 32894 -23440 32946
rect -23520 32880 -23440 32894
rect -23360 32946 -23280 32960
rect -23360 32894 -23346 32946
rect -23294 32894 -23280 32946
rect -23360 32880 -23280 32894
rect -23200 32946 -23120 32960
rect -23200 32894 -23186 32946
rect -23134 32894 -23120 32946
rect -23200 32880 -23120 32894
rect -23040 32946 -22960 32960
rect -23040 32894 -23026 32946
rect -22974 32894 -22960 32946
rect -23040 32880 -22960 32894
rect -22880 32946 -22800 32960
rect -22880 32894 -22866 32946
rect -22814 32894 -22800 32946
rect -22880 32880 -22800 32894
rect -22720 32946 -22640 32960
rect -22720 32894 -22706 32946
rect -22654 32894 -22640 32946
rect -22720 32880 -22640 32894
rect -22560 32946 -22480 32960
rect -22560 32894 -22546 32946
rect -22494 32894 -22480 32946
rect -22560 32880 -22480 32894
rect -22400 32946 -22320 32960
rect -22400 32894 -22386 32946
rect -22334 32894 -22320 32946
rect -22400 32880 -22320 32894
rect -22240 32946 -22160 32960
rect -22240 32894 -22226 32946
rect -22174 32894 -22160 32946
rect -22240 32880 -22160 32894
rect -22080 32946 -22000 32960
rect -22080 32894 -22066 32946
rect -22014 32894 -22000 32946
rect -22080 32880 -22000 32894
rect -21920 32946 -21840 32960
rect -21920 32894 -21906 32946
rect -21854 32894 -21840 32946
rect -21920 32880 -21840 32894
rect -21760 32946 -21680 32960
rect -21760 32894 -21746 32946
rect -21694 32894 -21680 32946
rect -21760 32880 -21680 32894
rect -21600 32946 -21520 32960
rect -21600 32894 -21586 32946
rect -21534 32894 -21520 32946
rect -21600 32880 -21520 32894
rect -21440 32946 -21360 32960
rect -21440 32894 -21426 32946
rect -21374 32894 -21360 32946
rect -21440 32880 -21360 32894
rect -21280 32946 -21200 32960
rect -21280 32894 -21266 32946
rect -21214 32894 -21200 32946
rect -21280 32880 -21200 32894
rect -21120 32946 -21040 32960
rect -21120 32894 -21106 32946
rect -21054 32894 -21040 32946
rect -21120 32880 -21040 32894
rect -20960 32946 -20880 32960
rect -20960 32894 -20946 32946
rect -20894 32894 -20880 32946
rect -20960 32880 -20880 32894
rect -20800 32946 -20720 32960
rect -20800 32894 -20786 32946
rect -20734 32894 -20720 32946
rect -20800 32880 -20720 32894
rect -20640 32946 -20560 32960
rect -20640 32894 -20626 32946
rect -20574 32894 -20560 32946
rect -20640 32880 -20560 32894
rect -20480 32946 -20400 32960
rect -20480 32894 -20466 32946
rect -20414 32894 -20400 32946
rect -20480 32880 -20400 32894
rect -20320 32946 -20240 32960
rect -20320 32894 -20306 32946
rect -20254 32894 -20240 32946
rect -20320 32880 -20240 32894
rect -20160 32946 -20080 32960
rect -20160 32894 -20146 32946
rect -20094 32894 -20080 32946
rect -20160 32880 -20080 32894
rect -20000 32946 -19920 32960
rect -20000 32894 -19986 32946
rect -19934 32894 -19920 32946
rect -20000 32880 -19920 32894
rect -19840 32946 -19760 32960
rect -19840 32894 -19826 32946
rect -19774 32894 -19760 32946
rect -19840 32880 -19760 32894
rect -19680 32946 -19600 32960
rect -19680 32894 -19666 32946
rect -19614 32894 -19600 32946
rect -19680 32880 -19600 32894
rect -19520 32946 -19440 32960
rect -19520 32894 -19506 32946
rect -19454 32894 -19440 32946
rect -19520 32880 -19440 32894
rect -19360 32946 -19280 32960
rect -19360 32894 -19346 32946
rect -19294 32894 -19280 32946
rect -19360 32880 -19280 32894
rect -19200 32946 -19120 32960
rect -19200 32894 -19186 32946
rect -19134 32894 -19120 32946
rect -19200 32880 -19120 32894
rect -19040 32946 -18960 32960
rect -19040 32894 -19026 32946
rect -18974 32894 -18960 32946
rect -19040 32880 -18960 32894
rect -18880 32946 -18800 32960
rect -18880 32894 -18866 32946
rect -18814 32894 -18800 32946
rect -18880 32880 -18800 32894
rect -18720 32946 -18640 32960
rect -18720 32894 -18706 32946
rect -18654 32894 -18640 32946
rect -18720 32880 -18640 32894
rect -18560 32946 -18480 32960
rect -18560 32894 -18546 32946
rect -18494 32894 -18480 32946
rect -18560 32880 -18480 32894
rect -18400 32946 -18320 32960
rect -18400 32894 -18386 32946
rect -18334 32894 -18320 32946
rect -18400 32880 -18320 32894
rect -18240 32946 -18160 32960
rect -18240 32894 -18226 32946
rect -18174 32894 -18160 32946
rect -18240 32880 -18160 32894
rect -18080 32946 -18000 32960
rect -18080 32894 -18066 32946
rect -18014 32894 -18000 32946
rect -18080 32880 -18000 32894
rect -17920 32946 -17840 32960
rect -17920 32894 -17906 32946
rect -17854 32894 -17840 32946
rect -17920 32880 -17840 32894
rect -17760 32946 -17680 32960
rect -17760 32894 -17746 32946
rect -17694 32894 -17680 32946
rect -17760 32880 -17680 32894
rect -17600 32946 -17520 32960
rect -17600 32894 -17586 32946
rect -17534 32894 -17520 32946
rect -17600 32880 -17520 32894
rect -17440 32946 -17360 32960
rect -17440 32894 -17426 32946
rect -17374 32894 -17360 32946
rect -17440 32880 -17360 32894
rect -17280 32946 -17200 32960
rect -17280 32894 -17266 32946
rect -17214 32894 -17200 32946
rect -17280 32880 -17200 32894
rect -17120 32946 -17040 32960
rect -17120 32894 -17106 32946
rect -17054 32894 -17040 32946
rect -17120 32880 -17040 32894
rect -16960 32946 -16880 32960
rect -16960 32894 -16946 32946
rect -16894 32894 -16880 32946
rect -16960 32880 -16880 32894
rect -16800 32946 -16720 32960
rect -16800 32894 -16786 32946
rect -16734 32894 -16720 32946
rect -16800 32880 -16720 32894
rect -16640 32946 -16560 32960
rect -16640 32894 -16626 32946
rect -16574 32894 -16560 32946
rect -16640 32880 -16560 32894
rect -16480 32946 -16400 32960
rect -16480 32894 -16466 32946
rect -16414 32894 -16400 32946
rect -16480 32880 -16400 32894
rect -16320 32946 -16240 32960
rect -16320 32894 -16306 32946
rect -16254 32894 -16240 32946
rect -16320 32880 -16240 32894
rect -16160 32946 -16080 32960
rect -16160 32894 -16146 32946
rect -16094 32894 -16080 32946
rect -16160 32880 -16080 32894
rect -16000 32946 -15920 32960
rect -16000 32894 -15986 32946
rect -15934 32894 -15920 32946
rect -16000 32880 -15920 32894
rect -15840 32946 -15760 32960
rect -15840 32894 -15826 32946
rect -15774 32894 -15760 32946
rect -15840 32880 -15760 32894
rect -15680 32946 -15600 32960
rect -15680 32894 -15666 32946
rect -15614 32894 -15600 32946
rect -15680 32880 -15600 32894
rect -15520 32946 -15440 32960
rect -15520 32894 -15506 32946
rect -15454 32894 -15440 32946
rect -15520 32880 -15440 32894
rect -15360 32946 -15280 32960
rect -15360 32894 -15346 32946
rect -15294 32894 -15280 32946
rect -15360 32880 -15280 32894
rect -15200 32946 -15120 32960
rect -15200 32894 -15186 32946
rect -15134 32894 -15120 32946
rect -15200 32880 -15120 32894
rect -15040 32946 -14960 32960
rect -15040 32894 -15026 32946
rect -14974 32894 -14960 32946
rect -15040 32880 -14960 32894
rect -14880 32946 -14800 32960
rect -14880 32894 -14866 32946
rect -14814 32894 -14800 32946
rect -14880 32880 -14800 32894
rect -14720 32946 -14640 32960
rect -14720 32894 -14706 32946
rect -14654 32894 -14640 32946
rect -14720 32880 -14640 32894
rect -14560 32946 -14480 32960
rect -14560 32894 -14546 32946
rect -14494 32894 -14480 32946
rect -14560 32880 -14480 32894
rect -14400 32946 -14320 32960
rect -14400 32894 -14386 32946
rect -14334 32894 -14320 32946
rect -14400 32880 -14320 32894
rect -14240 32946 -14160 32960
rect -14240 32894 -14226 32946
rect -14174 32894 -14160 32946
rect -14240 32880 -14160 32894
rect -14080 32946 -14000 32960
rect -14080 32894 -14066 32946
rect -14014 32894 -14000 32946
rect -14080 32880 -14000 32894
rect -13920 32946 -13840 32960
rect -13920 32894 -13906 32946
rect -13854 32894 -13840 32946
rect -13920 32880 -13840 32894
rect -13760 32946 -13680 32960
rect -13760 32894 -13746 32946
rect -13694 32894 -13680 32946
rect -13760 32880 -13680 32894
rect -13600 32946 -13520 32960
rect -13600 32894 -13586 32946
rect -13534 32894 -13520 32946
rect -13600 32880 -13520 32894
rect -13440 32946 -13360 32960
rect -13440 32894 -13426 32946
rect -13374 32894 -13360 32946
rect -13440 32880 -13360 32894
rect -13280 32946 -13200 32960
rect -13280 32894 -13266 32946
rect -13214 32894 -13200 32946
rect -13280 32880 -13200 32894
rect -13120 32946 -13040 32960
rect -13120 32894 -13106 32946
rect -13054 32894 -13040 32946
rect -13120 32880 -13040 32894
rect -12960 32946 -12880 32960
rect -12960 32894 -12946 32946
rect -12894 32894 -12880 32946
rect -12960 32880 -12880 32894
rect -12800 32946 -12720 32960
rect -12800 32894 -12786 32946
rect -12734 32894 -12720 32946
rect -12800 32880 -12720 32894
rect -12640 32946 -12560 32960
rect -12640 32894 -12626 32946
rect -12574 32894 -12560 32946
rect -12640 32880 -12560 32894
rect -12480 32946 -12400 32960
rect -12480 32894 -12466 32946
rect -12414 32894 -12400 32946
rect -12480 32880 -12400 32894
rect -12320 32946 -12240 32960
rect -12320 32894 -12306 32946
rect -12254 32894 -12240 32946
rect -12320 32880 -12240 32894
rect -12160 32946 -12080 32960
rect -12160 32894 -12146 32946
rect -12094 32894 -12080 32946
rect -12160 32880 -12080 32894
rect -12000 32946 -11920 32960
rect -12000 32894 -11986 32946
rect -11934 32894 -11920 32946
rect -12000 32880 -11920 32894
rect -11840 32946 -11760 32960
rect -11840 32894 -11826 32946
rect -11774 32894 -11760 32946
rect -11840 32880 -11760 32894
rect -11680 32946 -11600 32960
rect -11680 32894 -11666 32946
rect -11614 32894 -11600 32946
rect -11680 32880 -11600 32894
rect -11520 32946 -11440 32960
rect -11520 32894 -11506 32946
rect -11454 32894 -11440 32946
rect -11520 32880 -11440 32894
rect -11200 32946 -11120 32960
rect -11200 32894 -11186 32946
rect -11134 32894 -11120 32946
rect -11200 32880 -11120 32894
rect -10880 32946 -10800 32960
rect -10880 32894 -10866 32946
rect -10814 32894 -10800 32946
rect -10880 32880 -10800 32894
rect -10720 32946 -10640 32960
rect -10720 32894 -10706 32946
rect -10654 32894 -10640 32946
rect -10720 32880 -10640 32894
rect -10560 32946 -10480 32960
rect -10560 32894 -10546 32946
rect -10494 32894 -10480 32946
rect -10560 32880 -10480 32894
rect -10400 32946 -10320 32960
rect -10400 32894 -10386 32946
rect -10334 32894 -10320 32946
rect -10400 32880 -10320 32894
rect -10240 32946 -10160 32960
rect -10240 32894 -10226 32946
rect -10174 32894 -10160 32946
rect -10240 32880 -10160 32894
rect -10080 32946 -10000 32960
rect -10080 32894 -10066 32946
rect -10014 32894 -10000 32946
rect -10080 32880 -10000 32894
rect -9920 32946 -9840 32960
rect -9920 32894 -9906 32946
rect -9854 32894 -9840 32946
rect -9920 32880 -9840 32894
rect -9760 32946 -9680 32960
rect -9760 32894 -9746 32946
rect -9694 32894 -9680 32946
rect -9760 32880 -9680 32894
rect -9600 32946 -9520 32960
rect -9600 32894 -9586 32946
rect -9534 32894 -9520 32946
rect -9600 32880 -9520 32894
rect -9440 32946 -9360 32960
rect -9440 32894 -9426 32946
rect -9374 32894 -9360 32946
rect -9440 32880 -9360 32894
rect -9280 32946 -9200 32960
rect -9280 32894 -9266 32946
rect -9214 32894 -9200 32946
rect -9280 32880 -9200 32894
rect -9120 32946 -9040 32960
rect -9120 32894 -9106 32946
rect -9054 32894 -9040 32946
rect -9120 32880 -9040 32894
rect -8960 32946 -8880 32960
rect -8960 32894 -8946 32946
rect -8894 32894 -8880 32946
rect -8960 32880 -8880 32894
rect -8800 32946 -8720 32960
rect -8800 32894 -8786 32946
rect -8734 32894 -8720 32946
rect -8800 32880 -8720 32894
rect -8640 32946 -8560 32960
rect -8640 32894 -8626 32946
rect -8574 32894 -8560 32946
rect -8640 32880 -8560 32894
rect -8480 32946 -8400 32960
rect -8480 32894 -8466 32946
rect -8414 32894 -8400 32946
rect -8480 32880 -8400 32894
rect -8320 32946 -8240 32960
rect -8320 32894 -8306 32946
rect -8254 32894 -8240 32946
rect -8320 32880 -8240 32894
rect -8160 32946 -8080 32960
rect -8160 32894 -8146 32946
rect -8094 32894 -8080 32946
rect -8160 32880 -8080 32894
rect -8000 32946 -7920 32960
rect -8000 32894 -7986 32946
rect -7934 32894 -7920 32946
rect -8000 32880 -7920 32894
rect -7840 32946 -7760 32960
rect -7840 32894 -7826 32946
rect -7774 32894 -7760 32946
rect -7840 32880 -7760 32894
rect -7680 32946 -7600 32960
rect -7680 32894 -7666 32946
rect -7614 32894 -7600 32946
rect -7680 32880 -7600 32894
rect -7520 32946 -7440 32960
rect -7520 32894 -7506 32946
rect -7454 32894 -7440 32946
rect -7520 32880 -7440 32894
rect -7360 32946 -7280 32960
rect -7360 32894 -7346 32946
rect -7294 32894 -7280 32946
rect -7360 32880 -7280 32894
rect -7200 32946 -7120 32960
rect -7200 32894 -7186 32946
rect -7134 32894 -7120 32946
rect -7200 32880 -7120 32894
rect -7040 32946 -6960 32960
rect -7040 32894 -7026 32946
rect -6974 32894 -6960 32946
rect -7040 32880 -6960 32894
rect -6880 32946 -6800 32960
rect -6880 32894 -6866 32946
rect -6814 32894 -6800 32946
rect -6880 32880 -6800 32894
rect -6720 32946 -6640 32960
rect -6720 32894 -6706 32946
rect -6654 32894 -6640 32946
rect -6720 32880 -6640 32894
rect -6560 32946 -6480 32960
rect -6560 32894 -6546 32946
rect -6494 32894 -6480 32946
rect -6560 32880 -6480 32894
rect -6400 32946 -6320 32960
rect -6400 32894 -6386 32946
rect -6334 32894 -6320 32946
rect -6400 32880 -6320 32894
rect -6240 32946 -6160 32960
rect -6240 32894 -6226 32946
rect -6174 32894 -6160 32946
rect -6240 32880 -6160 32894
rect -6080 32946 -6000 32960
rect -6080 32894 -6066 32946
rect -6014 32894 -6000 32946
rect -6080 32880 -6000 32894
rect -5920 32946 -5840 32960
rect -5920 32894 -5906 32946
rect -5854 32894 -5840 32946
rect -5920 32880 -5840 32894
rect -5760 32946 -5680 32960
rect -5760 32894 -5746 32946
rect -5694 32894 -5680 32946
rect -5760 32880 -5680 32894
rect -5600 32946 -5520 32960
rect -5600 32894 -5586 32946
rect -5534 32894 -5520 32946
rect -5600 32880 -5520 32894
rect -5440 32946 -5360 32960
rect -5440 32894 -5426 32946
rect -5374 32894 -5360 32946
rect -5440 32880 -5360 32894
rect -5280 32946 -5200 32960
rect -5280 32894 -5266 32946
rect -5214 32894 -5200 32946
rect -5280 32880 -5200 32894
rect -5120 32946 -5040 32960
rect -5120 32894 -5106 32946
rect -5054 32894 -5040 32946
rect -5120 32880 -5040 32894
rect -4960 32946 -4880 32960
rect -4960 32894 -4946 32946
rect -4894 32894 -4880 32946
rect -4960 32880 -4880 32894
rect -4800 32946 -4720 32960
rect -4800 32894 -4786 32946
rect -4734 32894 -4720 32946
rect -4800 32880 -4720 32894
rect -4640 32946 -4560 32960
rect -4640 32894 -4626 32946
rect -4574 32894 -4560 32946
rect -4640 32880 -4560 32894
rect -4480 32946 -4400 32960
rect -4480 32894 -4466 32946
rect -4414 32894 -4400 32946
rect -4480 32880 -4400 32894
rect -4320 32946 -4240 32960
rect -4320 32894 -4306 32946
rect -4254 32894 -4240 32946
rect -4320 32880 -4240 32894
rect -4160 32946 -4080 32960
rect -4160 32894 -4146 32946
rect -4094 32894 -4080 32946
rect -4160 32880 -4080 32894
rect -4000 32946 -3920 32960
rect -4000 32894 -3986 32946
rect -3934 32894 -3920 32946
rect -4000 32880 -3920 32894
rect -3680 32946 -3600 32960
rect -3680 32894 -3666 32946
rect -3614 32894 -3600 32946
rect -3680 32880 -3600 32894
rect -3520 32946 -3440 32960
rect -3520 32894 -3506 32946
rect -3454 32894 -3440 32946
rect -3520 32880 -3440 32894
rect -3360 32946 -3280 32960
rect -3360 32894 -3346 32946
rect -3294 32894 -3280 32946
rect -3360 32880 -3280 32894
rect -3200 32946 -3120 32960
rect -3200 32894 -3186 32946
rect -3134 32894 -3120 32946
rect -3200 32880 -3120 32894
rect -3040 32946 -2960 32960
rect -3040 32894 -3026 32946
rect -2974 32894 -2960 32946
rect -3040 32880 -2960 32894
rect -2880 32946 -2800 32960
rect -2880 32894 -2866 32946
rect -2814 32894 -2800 32946
rect -2880 32880 -2800 32894
rect -2720 32946 -2640 32960
rect -2720 32894 -2706 32946
rect -2654 32894 -2640 32946
rect -2720 32880 -2640 32894
rect -2400 32946 -2320 32960
rect -2400 32894 -2386 32946
rect -2334 32894 -2320 32946
rect -2400 32880 -2320 32894
rect -2080 32946 -2000 32960
rect -2080 32894 -2066 32946
rect -2014 32894 -2000 32946
rect -2080 32880 -2000 32894
rect -1760 32946 -1680 32960
rect -1760 32894 -1746 32946
rect -1694 32894 -1680 32946
rect -1760 32880 -1680 32894
rect -1440 32946 -1360 32960
rect -1440 32894 -1426 32946
rect -1374 32894 -1360 32946
rect -1440 32880 -1360 32894
rect -1120 32946 -1040 32960
rect -1120 32894 -1106 32946
rect -1054 32894 -1040 32946
rect -1120 32880 -1040 32894
rect -29920 32626 -29840 32640
rect -29920 32574 -29906 32626
rect -29854 32574 -29840 32626
rect -29920 32560 -29840 32574
rect -29760 32626 -29680 32640
rect -29760 32574 -29746 32626
rect -29694 32574 -29680 32626
rect -29760 32560 -29680 32574
rect -29600 32626 -29520 32640
rect -29600 32574 -29586 32626
rect -29534 32574 -29520 32626
rect -29600 32560 -29520 32574
rect -29440 32626 -29360 32640
rect -29440 32574 -29426 32626
rect -29374 32574 -29360 32626
rect -29440 32560 -29360 32574
rect -29280 32626 -29200 32640
rect -29280 32574 -29266 32626
rect -29214 32574 -29200 32626
rect -29280 32560 -29200 32574
rect -29120 32626 -29040 32640
rect -29120 32574 -29106 32626
rect -29054 32574 -29040 32626
rect -29120 32560 -29040 32574
rect -28960 32626 -28880 32640
rect -28960 32574 -28946 32626
rect -28894 32574 -28880 32626
rect -28960 32560 -28880 32574
rect -28800 32626 -28720 32640
rect -28800 32574 -28786 32626
rect -28734 32574 -28720 32626
rect -28800 32560 -28720 32574
rect -28640 32626 -28560 32640
rect -28640 32574 -28626 32626
rect -28574 32574 -28560 32626
rect -28640 32560 -28560 32574
rect -28480 32626 -28400 32640
rect -28480 32574 -28466 32626
rect -28414 32574 -28400 32626
rect -28480 32560 -28400 32574
rect -28320 32626 -28240 32640
rect -28320 32574 -28306 32626
rect -28254 32574 -28240 32626
rect -28320 32560 -28240 32574
rect -28160 32626 -28080 32640
rect -28160 32574 -28146 32626
rect -28094 32574 -28080 32626
rect -28160 32560 -28080 32574
rect -28000 32626 -27920 32640
rect -28000 32574 -27986 32626
rect -27934 32574 -27920 32626
rect -28000 32560 -27920 32574
rect -27840 32626 -27760 32640
rect -27840 32574 -27826 32626
rect -27774 32574 -27760 32626
rect -27840 32560 -27760 32574
rect -27680 32626 -27600 32640
rect -27680 32574 -27666 32626
rect -27614 32574 -27600 32626
rect -27680 32560 -27600 32574
rect -27520 32626 -27440 32640
rect -27520 32574 -27506 32626
rect -27454 32574 -27440 32626
rect -27520 32560 -27440 32574
rect -27360 32626 -27280 32640
rect -27360 32574 -27346 32626
rect -27294 32574 -27280 32626
rect -27360 32560 -27280 32574
rect -27200 32626 -27120 32640
rect -27200 32574 -27186 32626
rect -27134 32574 -27120 32626
rect -27200 32560 -27120 32574
rect -27040 32626 -26960 32640
rect -27040 32574 -27026 32626
rect -26974 32574 -26960 32626
rect -27040 32560 -26960 32574
rect -26880 32626 -26800 32640
rect -26880 32574 -26866 32626
rect -26814 32574 -26800 32626
rect -26880 32560 -26800 32574
rect -26720 32626 -26640 32640
rect -26720 32574 -26706 32626
rect -26654 32574 -26640 32626
rect -26720 32560 -26640 32574
rect -26560 32626 -26480 32640
rect -26560 32574 -26546 32626
rect -26494 32574 -26480 32626
rect -26560 32560 -26480 32574
rect -26400 32626 -26320 32640
rect -26400 32574 -26386 32626
rect -26334 32574 -26320 32626
rect -26400 32560 -26320 32574
rect -26240 32626 -26160 32640
rect -26240 32574 -26226 32626
rect -26174 32574 -26160 32626
rect -26240 32560 -26160 32574
rect -26080 32626 -26000 32640
rect -26080 32574 -26066 32626
rect -26014 32574 -26000 32626
rect -26080 32560 -26000 32574
rect -25920 32626 -25840 32640
rect -25920 32574 -25906 32626
rect -25854 32574 -25840 32626
rect -25920 32560 -25840 32574
rect -25760 32626 -25680 32640
rect -25760 32574 -25746 32626
rect -25694 32574 -25680 32626
rect -25760 32560 -25680 32574
rect -25600 32626 -25520 32640
rect -25600 32574 -25586 32626
rect -25534 32574 -25520 32626
rect -25600 32560 -25520 32574
rect -25440 32626 -25360 32640
rect -25440 32574 -25426 32626
rect -25374 32574 -25360 32626
rect -25440 32560 -25360 32574
rect -25280 32626 -25200 32640
rect -25280 32574 -25266 32626
rect -25214 32574 -25200 32626
rect -25280 32560 -25200 32574
rect -25120 32626 -25040 32640
rect -25120 32574 -25106 32626
rect -25054 32574 -25040 32626
rect -25120 32560 -25040 32574
rect -24960 32626 -24880 32640
rect -24960 32574 -24946 32626
rect -24894 32574 -24880 32626
rect -24960 32560 -24880 32574
rect -24800 32626 -24720 32640
rect -24800 32574 -24786 32626
rect -24734 32574 -24720 32626
rect -24800 32560 -24720 32574
rect -24640 32626 -24560 32640
rect -24640 32574 -24626 32626
rect -24574 32574 -24560 32626
rect -24640 32560 -24560 32574
rect -24480 32626 -24400 32640
rect -24480 32574 -24466 32626
rect -24414 32574 -24400 32626
rect -24480 32560 -24400 32574
rect -24320 32626 -24240 32640
rect -24320 32574 -24306 32626
rect -24254 32574 -24240 32626
rect -24320 32560 -24240 32574
rect -24160 32626 -24080 32640
rect -24160 32574 -24146 32626
rect -24094 32574 -24080 32626
rect -24160 32560 -24080 32574
rect -24000 32626 -23920 32640
rect -24000 32574 -23986 32626
rect -23934 32574 -23920 32626
rect -24000 32560 -23920 32574
rect -23840 32626 -23760 32640
rect -23840 32574 -23826 32626
rect -23774 32574 -23760 32626
rect -23840 32560 -23760 32574
rect -23680 32626 -23600 32640
rect -23680 32574 -23666 32626
rect -23614 32574 -23600 32626
rect -23680 32560 -23600 32574
rect -23520 32626 -23440 32640
rect -23520 32574 -23506 32626
rect -23454 32574 -23440 32626
rect -23520 32560 -23440 32574
rect -23360 32626 -23280 32640
rect -23360 32574 -23346 32626
rect -23294 32574 -23280 32626
rect -23360 32560 -23280 32574
rect -23200 32626 -23120 32640
rect -23200 32574 -23186 32626
rect -23134 32574 -23120 32626
rect -23200 32560 -23120 32574
rect -23040 32626 -22960 32640
rect -23040 32574 -23026 32626
rect -22974 32574 -22960 32626
rect -23040 32560 -22960 32574
rect -22880 32626 -22800 32640
rect -22880 32574 -22866 32626
rect -22814 32574 -22800 32626
rect -22880 32560 -22800 32574
rect -22720 32626 -22640 32640
rect -22720 32574 -22706 32626
rect -22654 32574 -22640 32626
rect -22720 32560 -22640 32574
rect -22560 32626 -22480 32640
rect -22560 32574 -22546 32626
rect -22494 32574 -22480 32626
rect -22560 32560 -22480 32574
rect -22400 32626 -22320 32640
rect -22400 32574 -22386 32626
rect -22334 32574 -22320 32626
rect -22400 32560 -22320 32574
rect -22240 32626 -22160 32640
rect -22240 32574 -22226 32626
rect -22174 32574 -22160 32626
rect -22240 32560 -22160 32574
rect -22080 32626 -22000 32640
rect -22080 32574 -22066 32626
rect -22014 32574 -22000 32626
rect -22080 32560 -22000 32574
rect -21920 32626 -21840 32640
rect -21920 32574 -21906 32626
rect -21854 32574 -21840 32626
rect -21920 32560 -21840 32574
rect -21760 32626 -21680 32640
rect -21760 32574 -21746 32626
rect -21694 32574 -21680 32626
rect -21760 32560 -21680 32574
rect -21600 32626 -21520 32640
rect -21600 32574 -21586 32626
rect -21534 32574 -21520 32626
rect -21600 32560 -21520 32574
rect -21440 32626 -21360 32640
rect -21440 32574 -21426 32626
rect -21374 32574 -21360 32626
rect -21440 32560 -21360 32574
rect -21280 32626 -21200 32640
rect -21280 32574 -21266 32626
rect -21214 32574 -21200 32626
rect -21280 32560 -21200 32574
rect -21120 32626 -21040 32640
rect -21120 32574 -21106 32626
rect -21054 32574 -21040 32626
rect -21120 32560 -21040 32574
rect -20960 32626 -20880 32640
rect -20960 32574 -20946 32626
rect -20894 32574 -20880 32626
rect -20960 32560 -20880 32574
rect -20800 32626 -20720 32640
rect -20800 32574 -20786 32626
rect -20734 32574 -20720 32626
rect -20800 32560 -20720 32574
rect -20640 32626 -20560 32640
rect -20640 32574 -20626 32626
rect -20574 32574 -20560 32626
rect -20640 32560 -20560 32574
rect -20480 32626 -20400 32640
rect -20480 32574 -20466 32626
rect -20414 32574 -20400 32626
rect -20480 32560 -20400 32574
rect -20320 32626 -20240 32640
rect -20320 32574 -20306 32626
rect -20254 32574 -20240 32626
rect -20320 32560 -20240 32574
rect -20160 32626 -20080 32640
rect -20160 32574 -20146 32626
rect -20094 32574 -20080 32626
rect -20160 32560 -20080 32574
rect -20000 32626 -19920 32640
rect -20000 32574 -19986 32626
rect -19934 32574 -19920 32626
rect -20000 32560 -19920 32574
rect -19840 32626 -19760 32640
rect -19840 32574 -19826 32626
rect -19774 32574 -19760 32626
rect -19840 32560 -19760 32574
rect -19680 32626 -19600 32640
rect -19680 32574 -19666 32626
rect -19614 32574 -19600 32626
rect -19680 32560 -19600 32574
rect -19520 32626 -19440 32640
rect -19520 32574 -19506 32626
rect -19454 32574 -19440 32626
rect -19520 32560 -19440 32574
rect -19360 32626 -19280 32640
rect -19360 32574 -19346 32626
rect -19294 32574 -19280 32626
rect -19360 32560 -19280 32574
rect -19200 32626 -19120 32640
rect -19200 32574 -19186 32626
rect -19134 32574 -19120 32626
rect -19200 32560 -19120 32574
rect -19040 32626 -18960 32640
rect -19040 32574 -19026 32626
rect -18974 32574 -18960 32626
rect -19040 32560 -18960 32574
rect -18880 32626 -18800 32640
rect -18880 32574 -18866 32626
rect -18814 32574 -18800 32626
rect -18880 32560 -18800 32574
rect -18720 32626 -18640 32640
rect -18720 32574 -18706 32626
rect -18654 32574 -18640 32626
rect -18720 32560 -18640 32574
rect -18560 32626 -18480 32640
rect -18560 32574 -18546 32626
rect -18494 32574 -18480 32626
rect -18560 32560 -18480 32574
rect -18400 32626 -18320 32640
rect -18400 32574 -18386 32626
rect -18334 32574 -18320 32626
rect -18400 32560 -18320 32574
rect -18240 32626 -18160 32640
rect -18240 32574 -18226 32626
rect -18174 32574 -18160 32626
rect -18240 32560 -18160 32574
rect -18080 32626 -18000 32640
rect -18080 32574 -18066 32626
rect -18014 32574 -18000 32626
rect -18080 32560 -18000 32574
rect -17920 32626 -17840 32640
rect -17920 32574 -17906 32626
rect -17854 32574 -17840 32626
rect -17920 32560 -17840 32574
rect -17760 32626 -17680 32640
rect -17760 32574 -17746 32626
rect -17694 32574 -17680 32626
rect -17760 32560 -17680 32574
rect -17600 32626 -17520 32640
rect -17600 32574 -17586 32626
rect -17534 32574 -17520 32626
rect -17600 32560 -17520 32574
rect -17440 32626 -17360 32640
rect -17440 32574 -17426 32626
rect -17374 32574 -17360 32626
rect -17440 32560 -17360 32574
rect -17280 32626 -17200 32640
rect -17280 32574 -17266 32626
rect -17214 32574 -17200 32626
rect -17280 32560 -17200 32574
rect -17120 32626 -17040 32640
rect -17120 32574 -17106 32626
rect -17054 32574 -17040 32626
rect -17120 32560 -17040 32574
rect -16960 32626 -16880 32640
rect -16960 32574 -16946 32626
rect -16894 32574 -16880 32626
rect -16960 32560 -16880 32574
rect -16800 32626 -16720 32640
rect -16800 32574 -16786 32626
rect -16734 32574 -16720 32626
rect -16800 32560 -16720 32574
rect -16640 32626 -16560 32640
rect -16640 32574 -16626 32626
rect -16574 32574 -16560 32626
rect -16640 32560 -16560 32574
rect -16480 32626 -16400 32640
rect -16480 32574 -16466 32626
rect -16414 32574 -16400 32626
rect -16480 32560 -16400 32574
rect -16320 32626 -16240 32640
rect -16320 32574 -16306 32626
rect -16254 32574 -16240 32626
rect -16320 32560 -16240 32574
rect -16160 32626 -16080 32640
rect -16160 32574 -16146 32626
rect -16094 32574 -16080 32626
rect -16160 32560 -16080 32574
rect -16000 32626 -15920 32640
rect -16000 32574 -15986 32626
rect -15934 32574 -15920 32626
rect -16000 32560 -15920 32574
rect -15840 32626 -15760 32640
rect -15840 32574 -15826 32626
rect -15774 32574 -15760 32626
rect -15840 32560 -15760 32574
rect -15680 32626 -15600 32640
rect -15680 32574 -15666 32626
rect -15614 32574 -15600 32626
rect -15680 32560 -15600 32574
rect -15520 32626 -15440 32640
rect -15520 32574 -15506 32626
rect -15454 32574 -15440 32626
rect -15520 32560 -15440 32574
rect -15360 32626 -15280 32640
rect -15360 32574 -15346 32626
rect -15294 32574 -15280 32626
rect -15360 32560 -15280 32574
rect -15200 32626 -15120 32640
rect -15200 32574 -15186 32626
rect -15134 32574 -15120 32626
rect -15200 32560 -15120 32574
rect -15040 32626 -14960 32640
rect -15040 32574 -15026 32626
rect -14974 32574 -14960 32626
rect -15040 32560 -14960 32574
rect -14880 32626 -14800 32640
rect -14880 32574 -14866 32626
rect -14814 32574 -14800 32626
rect -14880 32560 -14800 32574
rect -14720 32626 -14640 32640
rect -14720 32574 -14706 32626
rect -14654 32574 -14640 32626
rect -14720 32560 -14640 32574
rect -14560 32626 -14480 32640
rect -14560 32574 -14546 32626
rect -14494 32574 -14480 32626
rect -14560 32560 -14480 32574
rect -14400 32626 -14320 32640
rect -14400 32574 -14386 32626
rect -14334 32574 -14320 32626
rect -14400 32560 -14320 32574
rect -14240 32626 -14160 32640
rect -14240 32574 -14226 32626
rect -14174 32574 -14160 32626
rect -14240 32560 -14160 32574
rect -14080 32626 -14000 32640
rect -14080 32574 -14066 32626
rect -14014 32574 -14000 32626
rect -14080 32560 -14000 32574
rect -13920 32626 -13840 32640
rect -13920 32574 -13906 32626
rect -13854 32574 -13840 32626
rect -13920 32560 -13840 32574
rect -13760 32626 -13680 32640
rect -13760 32574 -13746 32626
rect -13694 32574 -13680 32626
rect -13760 32560 -13680 32574
rect -13600 32626 -13520 32640
rect -13600 32574 -13586 32626
rect -13534 32574 -13520 32626
rect -13600 32560 -13520 32574
rect -13440 32626 -13360 32640
rect -13440 32574 -13426 32626
rect -13374 32574 -13360 32626
rect -13440 32560 -13360 32574
rect -13280 32626 -13200 32640
rect -13280 32574 -13266 32626
rect -13214 32574 -13200 32626
rect -13280 32560 -13200 32574
rect -13120 32626 -13040 32640
rect -13120 32574 -13106 32626
rect -13054 32574 -13040 32626
rect -13120 32560 -13040 32574
rect -12960 32626 -12880 32640
rect -12960 32574 -12946 32626
rect -12894 32574 -12880 32626
rect -12960 32560 -12880 32574
rect -12800 32626 -12720 32640
rect -12800 32574 -12786 32626
rect -12734 32574 -12720 32626
rect -12800 32560 -12720 32574
rect -12640 32626 -12560 32640
rect -12640 32574 -12626 32626
rect -12574 32574 -12560 32626
rect -12640 32560 -12560 32574
rect -12480 32626 -12400 32640
rect -12480 32574 -12466 32626
rect -12414 32574 -12400 32626
rect -12480 32560 -12400 32574
rect -12320 32626 -12240 32640
rect -12320 32574 -12306 32626
rect -12254 32574 -12240 32626
rect -12320 32560 -12240 32574
rect -12160 32626 -12080 32640
rect -12160 32574 -12146 32626
rect -12094 32574 -12080 32626
rect -12160 32560 -12080 32574
rect -12000 32626 -11920 32640
rect -12000 32574 -11986 32626
rect -11934 32574 -11920 32626
rect -12000 32560 -11920 32574
rect -11840 32626 -11760 32640
rect -11840 32574 -11826 32626
rect -11774 32574 -11760 32626
rect -11840 32560 -11760 32574
rect -11680 32626 -11600 32640
rect -11680 32574 -11666 32626
rect -11614 32574 -11600 32626
rect -11680 32560 -11600 32574
rect -11520 32626 -11440 32640
rect -11520 32574 -11506 32626
rect -11454 32574 -11440 32626
rect -11520 32560 -11440 32574
rect -11200 32626 -11120 32640
rect -11200 32574 -11186 32626
rect -11134 32574 -11120 32626
rect -11200 32560 -11120 32574
rect -10880 32626 -10800 32640
rect -10880 32574 -10866 32626
rect -10814 32574 -10800 32626
rect -10880 32560 -10800 32574
rect -10720 32626 -10640 32640
rect -10720 32574 -10706 32626
rect -10654 32574 -10640 32626
rect -10720 32560 -10640 32574
rect -10560 32626 -10480 32640
rect -10560 32574 -10546 32626
rect -10494 32574 -10480 32626
rect -10560 32560 -10480 32574
rect -10400 32626 -10320 32640
rect -10400 32574 -10386 32626
rect -10334 32574 -10320 32626
rect -10400 32560 -10320 32574
rect -10240 32626 -10160 32640
rect -10240 32574 -10226 32626
rect -10174 32574 -10160 32626
rect -10240 32560 -10160 32574
rect -10080 32626 -10000 32640
rect -10080 32574 -10066 32626
rect -10014 32574 -10000 32626
rect -10080 32560 -10000 32574
rect -9920 32626 -9840 32640
rect -9920 32574 -9906 32626
rect -9854 32574 -9840 32626
rect -9920 32560 -9840 32574
rect -9760 32626 -9680 32640
rect -9760 32574 -9746 32626
rect -9694 32574 -9680 32626
rect -9760 32560 -9680 32574
rect -9600 32626 -9520 32640
rect -9600 32574 -9586 32626
rect -9534 32574 -9520 32626
rect -9600 32560 -9520 32574
rect -9440 32626 -9360 32640
rect -9440 32574 -9426 32626
rect -9374 32574 -9360 32626
rect -9440 32560 -9360 32574
rect -9280 32626 -9200 32640
rect -9280 32574 -9266 32626
rect -9214 32574 -9200 32626
rect -9280 32560 -9200 32574
rect -9120 32626 -9040 32640
rect -9120 32574 -9106 32626
rect -9054 32574 -9040 32626
rect -9120 32560 -9040 32574
rect -8960 32626 -8880 32640
rect -8960 32574 -8946 32626
rect -8894 32574 -8880 32626
rect -8960 32560 -8880 32574
rect -8800 32626 -8720 32640
rect -8800 32574 -8786 32626
rect -8734 32574 -8720 32626
rect -8800 32560 -8720 32574
rect -8640 32626 -8560 32640
rect -8640 32574 -8626 32626
rect -8574 32574 -8560 32626
rect -8640 32560 -8560 32574
rect -8480 32626 -8400 32640
rect -8480 32574 -8466 32626
rect -8414 32574 -8400 32626
rect -8480 32560 -8400 32574
rect -8320 32626 -8240 32640
rect -8320 32574 -8306 32626
rect -8254 32574 -8240 32626
rect -8320 32560 -8240 32574
rect -8160 32626 -8080 32640
rect -8160 32574 -8146 32626
rect -8094 32574 -8080 32626
rect -8160 32560 -8080 32574
rect -8000 32626 -7920 32640
rect -8000 32574 -7986 32626
rect -7934 32574 -7920 32626
rect -8000 32560 -7920 32574
rect -7840 32626 -7760 32640
rect -7840 32574 -7826 32626
rect -7774 32574 -7760 32626
rect -7840 32560 -7760 32574
rect -7680 32626 -7600 32640
rect -7680 32574 -7666 32626
rect -7614 32574 -7600 32626
rect -7680 32560 -7600 32574
rect -7520 32626 -7440 32640
rect -7520 32574 -7506 32626
rect -7454 32574 -7440 32626
rect -7520 32560 -7440 32574
rect -7360 32626 -7280 32640
rect -7360 32574 -7346 32626
rect -7294 32574 -7280 32626
rect -7360 32560 -7280 32574
rect -7200 32626 -7120 32640
rect -7200 32574 -7186 32626
rect -7134 32574 -7120 32626
rect -7200 32560 -7120 32574
rect -7040 32626 -6960 32640
rect -7040 32574 -7026 32626
rect -6974 32574 -6960 32626
rect -7040 32560 -6960 32574
rect -6880 32626 -6800 32640
rect -6880 32574 -6866 32626
rect -6814 32574 -6800 32626
rect -6880 32560 -6800 32574
rect -6720 32626 -6640 32640
rect -6720 32574 -6706 32626
rect -6654 32574 -6640 32626
rect -6720 32560 -6640 32574
rect -6560 32626 -6480 32640
rect -6560 32574 -6546 32626
rect -6494 32574 -6480 32626
rect -6560 32560 -6480 32574
rect -6400 32626 -6320 32640
rect -6400 32574 -6386 32626
rect -6334 32574 -6320 32626
rect -6400 32560 -6320 32574
rect -6240 32626 -6160 32640
rect -6240 32574 -6226 32626
rect -6174 32574 -6160 32626
rect -6240 32560 -6160 32574
rect -6080 32626 -6000 32640
rect -6080 32574 -6066 32626
rect -6014 32574 -6000 32626
rect -6080 32560 -6000 32574
rect -5920 32626 -5840 32640
rect -5920 32574 -5906 32626
rect -5854 32574 -5840 32626
rect -5920 32560 -5840 32574
rect -5760 32626 -5680 32640
rect -5760 32574 -5746 32626
rect -5694 32574 -5680 32626
rect -5760 32560 -5680 32574
rect -5600 32626 -5520 32640
rect -5600 32574 -5586 32626
rect -5534 32574 -5520 32626
rect -5600 32560 -5520 32574
rect -5440 32626 -5360 32640
rect -5440 32574 -5426 32626
rect -5374 32574 -5360 32626
rect -5440 32560 -5360 32574
rect -5280 32626 -5200 32640
rect -5280 32574 -5266 32626
rect -5214 32574 -5200 32626
rect -5280 32560 -5200 32574
rect -5120 32626 -5040 32640
rect -5120 32574 -5106 32626
rect -5054 32574 -5040 32626
rect -5120 32560 -5040 32574
rect -4960 32626 -4880 32640
rect -4960 32574 -4946 32626
rect -4894 32574 -4880 32626
rect -4960 32560 -4880 32574
rect -4800 32626 -4720 32640
rect -4800 32574 -4786 32626
rect -4734 32574 -4720 32626
rect -4800 32560 -4720 32574
rect -4640 32626 -4560 32640
rect -4640 32574 -4626 32626
rect -4574 32574 -4560 32626
rect -4640 32560 -4560 32574
rect -4480 32626 -4400 32640
rect -4480 32574 -4466 32626
rect -4414 32574 -4400 32626
rect -4480 32560 -4400 32574
rect -4320 32626 -4240 32640
rect -4320 32574 -4306 32626
rect -4254 32574 -4240 32626
rect -4320 32560 -4240 32574
rect -4160 32626 -4080 32640
rect -4160 32574 -4146 32626
rect -4094 32574 -4080 32626
rect -4160 32560 -4080 32574
rect -4000 32626 -3920 32640
rect -4000 32574 -3986 32626
rect -3934 32574 -3920 32626
rect -4000 32560 -3920 32574
rect -3680 32626 -3600 32640
rect -3680 32574 -3666 32626
rect -3614 32574 -3600 32626
rect -3680 32560 -3600 32574
rect -3520 32626 -3440 32640
rect -3520 32574 -3506 32626
rect -3454 32574 -3440 32626
rect -3520 32560 -3440 32574
rect -3360 32626 -3280 32640
rect -3360 32574 -3346 32626
rect -3294 32574 -3280 32626
rect -3360 32560 -3280 32574
rect -3200 32626 -3120 32640
rect -3200 32574 -3186 32626
rect -3134 32574 -3120 32626
rect -3200 32560 -3120 32574
rect -3040 32626 -2960 32640
rect -3040 32574 -3026 32626
rect -2974 32574 -2960 32626
rect -3040 32560 -2960 32574
rect -2880 32626 -2800 32640
rect -2880 32574 -2866 32626
rect -2814 32574 -2800 32626
rect -2880 32560 -2800 32574
rect -2720 32626 -2640 32640
rect -2720 32574 -2706 32626
rect -2654 32574 -2640 32626
rect -2720 32560 -2640 32574
rect -2400 32626 -2320 32640
rect -2400 32574 -2386 32626
rect -2334 32574 -2320 32626
rect -2400 32560 -2320 32574
rect -2080 32626 -2000 32640
rect -2080 32574 -2066 32626
rect -2014 32574 -2000 32626
rect -2080 32560 -2000 32574
rect -1760 32626 -1680 32640
rect -1760 32574 -1746 32626
rect -1694 32574 -1680 32626
rect -1760 32560 -1680 32574
rect -1440 32626 -1360 32640
rect -1440 32574 -1426 32626
rect -1374 32574 -1360 32626
rect -1440 32560 -1360 32574
rect -1120 32626 -1040 32640
rect -1120 32574 -1106 32626
rect -1054 32574 -1040 32626
rect -1120 32560 -1040 32574
rect -29920 32306 -29840 32320
rect -29920 32254 -29906 32306
rect -29854 32254 -29840 32306
rect -29920 32240 -29840 32254
rect -29760 32306 -29680 32320
rect -29760 32254 -29746 32306
rect -29694 32254 -29680 32306
rect -29760 32240 -29680 32254
rect -29600 32306 -29520 32320
rect -29600 32254 -29586 32306
rect -29534 32254 -29520 32306
rect -29600 32240 -29520 32254
rect -29440 32306 -29360 32320
rect -29440 32254 -29426 32306
rect -29374 32254 -29360 32306
rect -29440 32240 -29360 32254
rect -29280 32306 -29200 32320
rect -29280 32254 -29266 32306
rect -29214 32254 -29200 32306
rect -29280 32240 -29200 32254
rect -29120 32306 -29040 32320
rect -29120 32254 -29106 32306
rect -29054 32254 -29040 32306
rect -29120 32240 -29040 32254
rect -28960 32306 -28880 32320
rect -28960 32254 -28946 32306
rect -28894 32254 -28880 32306
rect -28960 32240 -28880 32254
rect -28800 32306 -28720 32320
rect -28800 32254 -28786 32306
rect -28734 32254 -28720 32306
rect -28800 32240 -28720 32254
rect -28640 32306 -28560 32320
rect -28640 32254 -28626 32306
rect -28574 32254 -28560 32306
rect -28640 32240 -28560 32254
rect -28480 32306 -28400 32320
rect -28480 32254 -28466 32306
rect -28414 32254 -28400 32306
rect -28480 32240 -28400 32254
rect -28320 32306 -28240 32320
rect -28320 32254 -28306 32306
rect -28254 32254 -28240 32306
rect -28320 32240 -28240 32254
rect -28160 32306 -28080 32320
rect -28160 32254 -28146 32306
rect -28094 32254 -28080 32306
rect -28160 32240 -28080 32254
rect -28000 32306 -27920 32320
rect -28000 32254 -27986 32306
rect -27934 32254 -27920 32306
rect -28000 32240 -27920 32254
rect -27840 32306 -27760 32320
rect -27840 32254 -27826 32306
rect -27774 32254 -27760 32306
rect -27840 32240 -27760 32254
rect -27680 32306 -27600 32320
rect -27680 32254 -27666 32306
rect -27614 32254 -27600 32306
rect -27680 32240 -27600 32254
rect -27520 32306 -27440 32320
rect -27520 32254 -27506 32306
rect -27454 32254 -27440 32306
rect -27520 32240 -27440 32254
rect -27360 32306 -27280 32320
rect -27360 32254 -27346 32306
rect -27294 32254 -27280 32306
rect -27360 32240 -27280 32254
rect -27200 32306 -27120 32320
rect -27200 32254 -27186 32306
rect -27134 32254 -27120 32306
rect -27200 32240 -27120 32254
rect -27040 32306 -26960 32320
rect -27040 32254 -27026 32306
rect -26974 32254 -26960 32306
rect -27040 32240 -26960 32254
rect -26880 32306 -26800 32320
rect -26880 32254 -26866 32306
rect -26814 32254 -26800 32306
rect -26880 32240 -26800 32254
rect -26720 32306 -26640 32320
rect -26720 32254 -26706 32306
rect -26654 32254 -26640 32306
rect -26720 32240 -26640 32254
rect -26560 32306 -26480 32320
rect -26560 32254 -26546 32306
rect -26494 32254 -26480 32306
rect -26560 32240 -26480 32254
rect -26400 32306 -26320 32320
rect -26400 32254 -26386 32306
rect -26334 32254 -26320 32306
rect -26400 32240 -26320 32254
rect -26240 32306 -26160 32320
rect -26240 32254 -26226 32306
rect -26174 32254 -26160 32306
rect -26240 32240 -26160 32254
rect -26080 32306 -26000 32320
rect -26080 32254 -26066 32306
rect -26014 32254 -26000 32306
rect -26080 32240 -26000 32254
rect -25920 32306 -25840 32320
rect -25920 32254 -25906 32306
rect -25854 32254 -25840 32306
rect -25920 32240 -25840 32254
rect -25760 32306 -25680 32320
rect -25760 32254 -25746 32306
rect -25694 32254 -25680 32306
rect -25760 32240 -25680 32254
rect -25600 32306 -25520 32320
rect -25600 32254 -25586 32306
rect -25534 32254 -25520 32306
rect -25600 32240 -25520 32254
rect -25440 32306 -25360 32320
rect -25440 32254 -25426 32306
rect -25374 32254 -25360 32306
rect -25440 32240 -25360 32254
rect -25280 32306 -25200 32320
rect -25280 32254 -25266 32306
rect -25214 32254 -25200 32306
rect -25280 32240 -25200 32254
rect -25120 32306 -25040 32320
rect -25120 32254 -25106 32306
rect -25054 32254 -25040 32306
rect -25120 32240 -25040 32254
rect -24960 32306 -24880 32320
rect -24960 32254 -24946 32306
rect -24894 32254 -24880 32306
rect -24960 32240 -24880 32254
rect -24800 32306 -24720 32320
rect -24800 32254 -24786 32306
rect -24734 32254 -24720 32306
rect -24800 32240 -24720 32254
rect -24640 32306 -24560 32320
rect -24640 32254 -24626 32306
rect -24574 32254 -24560 32306
rect -24640 32240 -24560 32254
rect -24480 32306 -24400 32320
rect -24480 32254 -24466 32306
rect -24414 32254 -24400 32306
rect -24480 32240 -24400 32254
rect -24320 32306 -24240 32320
rect -24320 32254 -24306 32306
rect -24254 32254 -24240 32306
rect -24320 32240 -24240 32254
rect -24160 32306 -24080 32320
rect -24160 32254 -24146 32306
rect -24094 32254 -24080 32306
rect -24160 32240 -24080 32254
rect -24000 32306 -23920 32320
rect -24000 32254 -23986 32306
rect -23934 32254 -23920 32306
rect -24000 32240 -23920 32254
rect -23840 32306 -23760 32320
rect -23840 32254 -23826 32306
rect -23774 32254 -23760 32306
rect -23840 32240 -23760 32254
rect -23680 32306 -23600 32320
rect -23680 32254 -23666 32306
rect -23614 32254 -23600 32306
rect -23680 32240 -23600 32254
rect -23520 32306 -23440 32320
rect -23520 32254 -23506 32306
rect -23454 32254 -23440 32306
rect -23520 32240 -23440 32254
rect -23360 32306 -23280 32320
rect -23360 32254 -23346 32306
rect -23294 32254 -23280 32306
rect -23360 32240 -23280 32254
rect -23200 32306 -23120 32320
rect -23200 32254 -23186 32306
rect -23134 32254 -23120 32306
rect -23200 32240 -23120 32254
rect -23040 32306 -22960 32320
rect -23040 32254 -23026 32306
rect -22974 32254 -22960 32306
rect -23040 32240 -22960 32254
rect -22880 32306 -22800 32320
rect -22880 32254 -22866 32306
rect -22814 32254 -22800 32306
rect -22880 32240 -22800 32254
rect -22720 32306 -22640 32320
rect -22720 32254 -22706 32306
rect -22654 32254 -22640 32306
rect -22720 32240 -22640 32254
rect -22560 32306 -22480 32320
rect -22560 32254 -22546 32306
rect -22494 32254 -22480 32306
rect -22560 32240 -22480 32254
rect -22400 32306 -22320 32320
rect -22400 32254 -22386 32306
rect -22334 32254 -22320 32306
rect -22400 32240 -22320 32254
rect -22240 32306 -22160 32320
rect -22240 32254 -22226 32306
rect -22174 32254 -22160 32306
rect -22240 32240 -22160 32254
rect -22080 32306 -22000 32320
rect -22080 32254 -22066 32306
rect -22014 32254 -22000 32306
rect -22080 32240 -22000 32254
rect -21920 32306 -21840 32320
rect -21920 32254 -21906 32306
rect -21854 32254 -21840 32306
rect -21920 32240 -21840 32254
rect -21760 32306 -21680 32320
rect -21760 32254 -21746 32306
rect -21694 32254 -21680 32306
rect -21760 32240 -21680 32254
rect -21600 32306 -21520 32320
rect -21600 32254 -21586 32306
rect -21534 32254 -21520 32306
rect -21600 32240 -21520 32254
rect -21440 32306 -21360 32320
rect -21440 32254 -21426 32306
rect -21374 32254 -21360 32306
rect -21440 32240 -21360 32254
rect -21280 32306 -21200 32320
rect -21280 32254 -21266 32306
rect -21214 32254 -21200 32306
rect -21280 32240 -21200 32254
rect -21120 32306 -21040 32320
rect -21120 32254 -21106 32306
rect -21054 32254 -21040 32306
rect -21120 32240 -21040 32254
rect -20960 32306 -20880 32320
rect -20960 32254 -20946 32306
rect -20894 32254 -20880 32306
rect -20960 32240 -20880 32254
rect -20800 32306 -20720 32320
rect -20800 32254 -20786 32306
rect -20734 32254 -20720 32306
rect -20800 32240 -20720 32254
rect -20640 32306 -20560 32320
rect -20640 32254 -20626 32306
rect -20574 32254 -20560 32306
rect -20640 32240 -20560 32254
rect -20480 32306 -20400 32320
rect -20480 32254 -20466 32306
rect -20414 32254 -20400 32306
rect -20480 32240 -20400 32254
rect -20320 32306 -20240 32320
rect -20320 32254 -20306 32306
rect -20254 32254 -20240 32306
rect -20320 32240 -20240 32254
rect -20160 32306 -20080 32320
rect -20160 32254 -20146 32306
rect -20094 32254 -20080 32306
rect -20160 32240 -20080 32254
rect -20000 32306 -19920 32320
rect -20000 32254 -19986 32306
rect -19934 32254 -19920 32306
rect -20000 32240 -19920 32254
rect -19840 32306 -19760 32320
rect -19840 32254 -19826 32306
rect -19774 32254 -19760 32306
rect -19840 32240 -19760 32254
rect -19680 32306 -19600 32320
rect -19680 32254 -19666 32306
rect -19614 32254 -19600 32306
rect -19680 32240 -19600 32254
rect -19520 32306 -19440 32320
rect -19520 32254 -19506 32306
rect -19454 32254 -19440 32306
rect -19520 32240 -19440 32254
rect -19360 32306 -19280 32320
rect -19360 32254 -19346 32306
rect -19294 32254 -19280 32306
rect -19360 32240 -19280 32254
rect -19200 32306 -19120 32320
rect -19200 32254 -19186 32306
rect -19134 32254 -19120 32306
rect -19200 32240 -19120 32254
rect -19040 32306 -18960 32320
rect -19040 32254 -19026 32306
rect -18974 32254 -18960 32306
rect -19040 32240 -18960 32254
rect -18880 32306 -18800 32320
rect -18880 32254 -18866 32306
rect -18814 32254 -18800 32306
rect -18880 32240 -18800 32254
rect -18720 32306 -18640 32320
rect -18720 32254 -18706 32306
rect -18654 32254 -18640 32306
rect -18720 32240 -18640 32254
rect -18560 32306 -18480 32320
rect -18560 32254 -18546 32306
rect -18494 32254 -18480 32306
rect -18560 32240 -18480 32254
rect -18400 32306 -18320 32320
rect -18400 32254 -18386 32306
rect -18334 32254 -18320 32306
rect -18400 32240 -18320 32254
rect -18240 32306 -18160 32320
rect -18240 32254 -18226 32306
rect -18174 32254 -18160 32306
rect -18240 32240 -18160 32254
rect -18080 32306 -18000 32320
rect -18080 32254 -18066 32306
rect -18014 32254 -18000 32306
rect -18080 32240 -18000 32254
rect -17920 32306 -17840 32320
rect -17920 32254 -17906 32306
rect -17854 32254 -17840 32306
rect -17920 32240 -17840 32254
rect -17760 32306 -17680 32320
rect -17760 32254 -17746 32306
rect -17694 32254 -17680 32306
rect -17760 32240 -17680 32254
rect -17600 32306 -17520 32320
rect -17600 32254 -17586 32306
rect -17534 32254 -17520 32306
rect -17600 32240 -17520 32254
rect -17440 32306 -17360 32320
rect -17440 32254 -17426 32306
rect -17374 32254 -17360 32306
rect -17440 32240 -17360 32254
rect -17280 32306 -17200 32320
rect -17280 32254 -17266 32306
rect -17214 32254 -17200 32306
rect -17280 32240 -17200 32254
rect -17120 32306 -17040 32320
rect -17120 32254 -17106 32306
rect -17054 32254 -17040 32306
rect -17120 32240 -17040 32254
rect -16960 32306 -16880 32320
rect -16960 32254 -16946 32306
rect -16894 32254 -16880 32306
rect -16960 32240 -16880 32254
rect -16800 32306 -16720 32320
rect -16800 32254 -16786 32306
rect -16734 32254 -16720 32306
rect -16800 32240 -16720 32254
rect -16640 32306 -16560 32320
rect -16640 32254 -16626 32306
rect -16574 32254 -16560 32306
rect -16640 32240 -16560 32254
rect -16480 32306 -16400 32320
rect -16480 32254 -16466 32306
rect -16414 32254 -16400 32306
rect -16480 32240 -16400 32254
rect -16320 32306 -16240 32320
rect -16320 32254 -16306 32306
rect -16254 32254 -16240 32306
rect -16320 32240 -16240 32254
rect -16160 32306 -16080 32320
rect -16160 32254 -16146 32306
rect -16094 32254 -16080 32306
rect -16160 32240 -16080 32254
rect -16000 32306 -15920 32320
rect -16000 32254 -15986 32306
rect -15934 32254 -15920 32306
rect -16000 32240 -15920 32254
rect -15840 32306 -15760 32320
rect -15840 32254 -15826 32306
rect -15774 32254 -15760 32306
rect -15840 32240 -15760 32254
rect -15680 32306 -15600 32320
rect -15680 32254 -15666 32306
rect -15614 32254 -15600 32306
rect -15680 32240 -15600 32254
rect -15520 32306 -15440 32320
rect -15520 32254 -15506 32306
rect -15454 32254 -15440 32306
rect -15520 32240 -15440 32254
rect -15360 32306 -15280 32320
rect -15360 32254 -15346 32306
rect -15294 32254 -15280 32306
rect -15360 32240 -15280 32254
rect -15200 32306 -15120 32320
rect -15200 32254 -15186 32306
rect -15134 32254 -15120 32306
rect -15200 32240 -15120 32254
rect -15040 32306 -14960 32320
rect -15040 32254 -15026 32306
rect -14974 32254 -14960 32306
rect -15040 32240 -14960 32254
rect -14880 32306 -14800 32320
rect -14880 32254 -14866 32306
rect -14814 32254 -14800 32306
rect -14880 32240 -14800 32254
rect -14720 32306 -14640 32320
rect -14720 32254 -14706 32306
rect -14654 32254 -14640 32306
rect -14720 32240 -14640 32254
rect -14560 32306 -14480 32320
rect -14560 32254 -14546 32306
rect -14494 32254 -14480 32306
rect -14560 32240 -14480 32254
rect -14400 32306 -14320 32320
rect -14400 32254 -14386 32306
rect -14334 32254 -14320 32306
rect -14400 32240 -14320 32254
rect -14240 32306 -14160 32320
rect -14240 32254 -14226 32306
rect -14174 32254 -14160 32306
rect -14240 32240 -14160 32254
rect -14080 32306 -14000 32320
rect -14080 32254 -14066 32306
rect -14014 32254 -14000 32306
rect -14080 32240 -14000 32254
rect -13920 32306 -13840 32320
rect -13920 32254 -13906 32306
rect -13854 32254 -13840 32306
rect -13920 32240 -13840 32254
rect -13760 32306 -13680 32320
rect -13760 32254 -13746 32306
rect -13694 32254 -13680 32306
rect -13760 32240 -13680 32254
rect -13600 32306 -13520 32320
rect -13600 32254 -13586 32306
rect -13534 32254 -13520 32306
rect -13600 32240 -13520 32254
rect -13440 32306 -13360 32320
rect -13440 32254 -13426 32306
rect -13374 32254 -13360 32306
rect -13440 32240 -13360 32254
rect -13280 32306 -13200 32320
rect -13280 32254 -13266 32306
rect -13214 32254 -13200 32306
rect -13280 32240 -13200 32254
rect -13120 32306 -13040 32320
rect -13120 32254 -13106 32306
rect -13054 32254 -13040 32306
rect -13120 32240 -13040 32254
rect -12960 32306 -12880 32320
rect -12960 32254 -12946 32306
rect -12894 32254 -12880 32306
rect -12960 32240 -12880 32254
rect -12800 32306 -12720 32320
rect -12800 32254 -12786 32306
rect -12734 32254 -12720 32306
rect -12800 32240 -12720 32254
rect -12640 32306 -12560 32320
rect -12640 32254 -12626 32306
rect -12574 32254 -12560 32306
rect -12640 32240 -12560 32254
rect -12480 32306 -12400 32320
rect -12480 32254 -12466 32306
rect -12414 32254 -12400 32306
rect -12480 32240 -12400 32254
rect -12320 32306 -12240 32320
rect -12320 32254 -12306 32306
rect -12254 32254 -12240 32306
rect -12320 32240 -12240 32254
rect -12160 32306 -12080 32320
rect -12160 32254 -12146 32306
rect -12094 32254 -12080 32306
rect -12160 32240 -12080 32254
rect -12000 32306 -11920 32320
rect -12000 32254 -11986 32306
rect -11934 32254 -11920 32306
rect -12000 32240 -11920 32254
rect -11840 32306 -11760 32320
rect -11840 32254 -11826 32306
rect -11774 32254 -11760 32306
rect -11840 32240 -11760 32254
rect -11680 32306 -11600 32320
rect -11680 32254 -11666 32306
rect -11614 32254 -11600 32306
rect -11680 32240 -11600 32254
rect -11520 32306 -11440 32320
rect -11520 32254 -11506 32306
rect -11454 32254 -11440 32306
rect -11520 32240 -11440 32254
rect -11360 32306 -11280 32320
rect -11360 32254 -11346 32306
rect -11294 32254 -11280 32306
rect -11360 32240 -11280 32254
rect -11200 32306 -11120 32320
rect -11200 32254 -11186 32306
rect -11134 32254 -11120 32306
rect -11200 32240 -11120 32254
rect -10880 32306 -10800 32320
rect -10880 32254 -10866 32306
rect -10814 32254 -10800 32306
rect -10880 32240 -10800 32254
rect -10720 32306 -10640 32320
rect -10720 32254 -10706 32306
rect -10654 32254 -10640 32306
rect -10720 32240 -10640 32254
rect -10560 32306 -10480 32320
rect -10560 32254 -10546 32306
rect -10494 32254 -10480 32306
rect -10560 32240 -10480 32254
rect -10400 32306 -10320 32320
rect -10400 32254 -10386 32306
rect -10334 32254 -10320 32306
rect -10400 32240 -10320 32254
rect -10240 32306 -10160 32320
rect -10240 32254 -10226 32306
rect -10174 32254 -10160 32306
rect -10240 32240 -10160 32254
rect -10080 32306 -10000 32320
rect -10080 32254 -10066 32306
rect -10014 32254 -10000 32306
rect -10080 32240 -10000 32254
rect -9920 32306 -9840 32320
rect -9920 32254 -9906 32306
rect -9854 32254 -9840 32306
rect -9920 32240 -9840 32254
rect -9760 32306 -9680 32320
rect -9760 32254 -9746 32306
rect -9694 32254 -9680 32306
rect -9760 32240 -9680 32254
rect -9600 32306 -9520 32320
rect -9600 32254 -9586 32306
rect -9534 32254 -9520 32306
rect -9600 32240 -9520 32254
rect -9440 32306 -9360 32320
rect -9440 32254 -9426 32306
rect -9374 32254 -9360 32306
rect -9440 32240 -9360 32254
rect -9280 32306 -9200 32320
rect -9280 32254 -9266 32306
rect -9214 32254 -9200 32306
rect -9280 32240 -9200 32254
rect -9120 32306 -9040 32320
rect -9120 32254 -9106 32306
rect -9054 32254 -9040 32306
rect -9120 32240 -9040 32254
rect -8960 32306 -8880 32320
rect -8960 32254 -8946 32306
rect -8894 32254 -8880 32306
rect -8960 32240 -8880 32254
rect -8800 32306 -8720 32320
rect -8800 32254 -8786 32306
rect -8734 32254 -8720 32306
rect -8800 32240 -8720 32254
rect -8640 32306 -8560 32320
rect -8640 32254 -8626 32306
rect -8574 32254 -8560 32306
rect -8640 32240 -8560 32254
rect -8480 32306 -8400 32320
rect -8480 32254 -8466 32306
rect -8414 32254 -8400 32306
rect -8480 32240 -8400 32254
rect -8320 32306 -8240 32320
rect -8320 32254 -8306 32306
rect -8254 32254 -8240 32306
rect -8320 32240 -8240 32254
rect -8160 32306 -8080 32320
rect -8160 32254 -8146 32306
rect -8094 32254 -8080 32306
rect -8160 32240 -8080 32254
rect -8000 32306 -7920 32320
rect -8000 32254 -7986 32306
rect -7934 32254 -7920 32306
rect -8000 32240 -7920 32254
rect -7840 32306 -7760 32320
rect -7840 32254 -7826 32306
rect -7774 32254 -7760 32306
rect -7840 32240 -7760 32254
rect -7680 32306 -7600 32320
rect -7680 32254 -7666 32306
rect -7614 32254 -7600 32306
rect -7680 32240 -7600 32254
rect -7520 32306 -7440 32320
rect -7520 32254 -7506 32306
rect -7454 32254 -7440 32306
rect -7520 32240 -7440 32254
rect -7360 32306 -7280 32320
rect -7360 32254 -7346 32306
rect -7294 32254 -7280 32306
rect -7360 32240 -7280 32254
rect -7200 32306 -7120 32320
rect -7200 32254 -7186 32306
rect -7134 32254 -7120 32306
rect -7200 32240 -7120 32254
rect -7040 32306 -6960 32320
rect -7040 32254 -7026 32306
rect -6974 32254 -6960 32306
rect -7040 32240 -6960 32254
rect -6880 32306 -6800 32320
rect -6880 32254 -6866 32306
rect -6814 32254 -6800 32306
rect -6880 32240 -6800 32254
rect -6720 32306 -6640 32320
rect -6720 32254 -6706 32306
rect -6654 32254 -6640 32306
rect -6720 32240 -6640 32254
rect -6560 32306 -6480 32320
rect -6560 32254 -6546 32306
rect -6494 32254 -6480 32306
rect -6560 32240 -6480 32254
rect -6400 32306 -6320 32320
rect -6400 32254 -6386 32306
rect -6334 32254 -6320 32306
rect -6400 32240 -6320 32254
rect -6240 32306 -6160 32320
rect -6240 32254 -6226 32306
rect -6174 32254 -6160 32306
rect -6240 32240 -6160 32254
rect -6080 32306 -6000 32320
rect -6080 32254 -6066 32306
rect -6014 32254 -6000 32306
rect -6080 32240 -6000 32254
rect -5920 32306 -5840 32320
rect -5920 32254 -5906 32306
rect -5854 32254 -5840 32306
rect -5920 32240 -5840 32254
rect -5760 32306 -5680 32320
rect -5760 32254 -5746 32306
rect -5694 32254 -5680 32306
rect -5760 32240 -5680 32254
rect -5600 32306 -5520 32320
rect -5600 32254 -5586 32306
rect -5534 32254 -5520 32306
rect -5600 32240 -5520 32254
rect -5440 32306 -5360 32320
rect -5440 32254 -5426 32306
rect -5374 32254 -5360 32306
rect -5440 32240 -5360 32254
rect -5280 32306 -5200 32320
rect -5280 32254 -5266 32306
rect -5214 32254 -5200 32306
rect -5280 32240 -5200 32254
rect -5120 32306 -5040 32320
rect -5120 32254 -5106 32306
rect -5054 32254 -5040 32306
rect -5120 32240 -5040 32254
rect -4960 32306 -4880 32320
rect -4960 32254 -4946 32306
rect -4894 32254 -4880 32306
rect -4960 32240 -4880 32254
rect -4800 32306 -4720 32320
rect -4800 32254 -4786 32306
rect -4734 32254 -4720 32306
rect -4800 32240 -4720 32254
rect -4640 32306 -4560 32320
rect -4640 32254 -4626 32306
rect -4574 32254 -4560 32306
rect -4640 32240 -4560 32254
rect -4480 32306 -4400 32320
rect -4480 32254 -4466 32306
rect -4414 32254 -4400 32306
rect -4480 32240 -4400 32254
rect -4320 32306 -4240 32320
rect -4320 32254 -4306 32306
rect -4254 32254 -4240 32306
rect -4320 32240 -4240 32254
rect -4160 32306 -4080 32320
rect -4160 32254 -4146 32306
rect -4094 32254 -4080 32306
rect -4160 32240 -4080 32254
rect -4000 32306 -3920 32320
rect -4000 32254 -3986 32306
rect -3934 32254 -3920 32306
rect -4000 32240 -3920 32254
rect -3680 32306 -3600 32320
rect -3680 32254 -3666 32306
rect -3614 32254 -3600 32306
rect -3680 32240 -3600 32254
rect -3520 32306 -3440 32320
rect -3520 32254 -3506 32306
rect -3454 32254 -3440 32306
rect -3520 32240 -3440 32254
rect -3360 32306 -3280 32320
rect -3360 32254 -3346 32306
rect -3294 32254 -3280 32306
rect -3360 32240 -3280 32254
rect -3200 32306 -3120 32320
rect -3200 32254 -3186 32306
rect -3134 32254 -3120 32306
rect -3200 32240 -3120 32254
rect -3040 32306 -2960 32320
rect -3040 32254 -3026 32306
rect -2974 32254 -2960 32306
rect -3040 32240 -2960 32254
rect -2880 32306 -2800 32320
rect -2880 32254 -2866 32306
rect -2814 32254 -2800 32306
rect -2880 32240 -2800 32254
rect -2720 32306 -2640 32320
rect -2720 32254 -2706 32306
rect -2654 32254 -2640 32306
rect -2720 32240 -2640 32254
rect -2400 32306 -2320 32320
rect -2400 32254 -2386 32306
rect -2334 32254 -2320 32306
rect -2400 32240 -2320 32254
rect -2080 32306 -2000 32320
rect -2080 32254 -2066 32306
rect -2014 32254 -2000 32306
rect -2080 32240 -2000 32254
rect -1760 32306 -1680 32320
rect -1760 32254 -1746 32306
rect -1694 32254 -1680 32306
rect -1760 32240 -1680 32254
rect -1440 32306 -1360 32320
rect -1440 32254 -1426 32306
rect -1374 32254 -1360 32306
rect -1440 32240 -1360 32254
rect -1120 32306 -1040 32320
rect -1120 32254 -1106 32306
rect -1054 32254 -1040 32306
rect -1120 32240 -1040 32254
rect -11040 32080 -10960 32160
rect -29920 31986 -29840 32000
rect -29920 31934 -29906 31986
rect -29854 31934 -29840 31986
rect -29920 31920 -29840 31934
rect -29760 31986 -29680 32000
rect -29760 31934 -29746 31986
rect -29694 31934 -29680 31986
rect -29760 31920 -29680 31934
rect -29600 31986 -29520 32000
rect -29600 31934 -29586 31986
rect -29534 31934 -29520 31986
rect -29600 31920 -29520 31934
rect -29440 31986 -29360 32000
rect -29440 31934 -29426 31986
rect -29374 31934 -29360 31986
rect -29440 31920 -29360 31934
rect -29280 31986 -29200 32000
rect -29280 31934 -29266 31986
rect -29214 31934 -29200 31986
rect -29280 31920 -29200 31934
rect -29120 31986 -29040 32000
rect -29120 31934 -29106 31986
rect -29054 31934 -29040 31986
rect -29120 31920 -29040 31934
rect -28960 31986 -28880 32000
rect -28960 31934 -28946 31986
rect -28894 31934 -28880 31986
rect -28960 31920 -28880 31934
rect -28800 31986 -28720 32000
rect -28800 31934 -28786 31986
rect -28734 31934 -28720 31986
rect -28800 31920 -28720 31934
rect -28640 31986 -28560 32000
rect -28640 31934 -28626 31986
rect -28574 31934 -28560 31986
rect -28640 31920 -28560 31934
rect -28480 31986 -28400 32000
rect -28480 31934 -28466 31986
rect -28414 31934 -28400 31986
rect -28480 31920 -28400 31934
rect -28320 31986 -28240 32000
rect -28320 31934 -28306 31986
rect -28254 31934 -28240 31986
rect -28320 31920 -28240 31934
rect -28160 31986 -28080 32000
rect -28160 31934 -28146 31986
rect -28094 31934 -28080 31986
rect -28160 31920 -28080 31934
rect -28000 31986 -27920 32000
rect -28000 31934 -27986 31986
rect -27934 31934 -27920 31986
rect -28000 31920 -27920 31934
rect -27840 31986 -27760 32000
rect -27840 31934 -27826 31986
rect -27774 31934 -27760 31986
rect -27840 31920 -27760 31934
rect -27680 31986 -27600 32000
rect -27680 31934 -27666 31986
rect -27614 31934 -27600 31986
rect -27680 31920 -27600 31934
rect -27520 31986 -27440 32000
rect -27520 31934 -27506 31986
rect -27454 31934 -27440 31986
rect -27520 31920 -27440 31934
rect -27360 31986 -27280 32000
rect -27360 31934 -27346 31986
rect -27294 31934 -27280 31986
rect -27360 31920 -27280 31934
rect -27200 31986 -27120 32000
rect -27200 31934 -27186 31986
rect -27134 31934 -27120 31986
rect -27200 31920 -27120 31934
rect -27040 31986 -26960 32000
rect -27040 31934 -27026 31986
rect -26974 31934 -26960 31986
rect -27040 31920 -26960 31934
rect -26880 31986 -26800 32000
rect -26880 31934 -26866 31986
rect -26814 31934 -26800 31986
rect -26880 31920 -26800 31934
rect -26720 31986 -26640 32000
rect -26720 31934 -26706 31986
rect -26654 31934 -26640 31986
rect -26720 31920 -26640 31934
rect -26560 31986 -26480 32000
rect -26560 31934 -26546 31986
rect -26494 31934 -26480 31986
rect -26560 31920 -26480 31934
rect -26400 31986 -26320 32000
rect -26400 31934 -26386 31986
rect -26334 31934 -26320 31986
rect -26400 31920 -26320 31934
rect -26240 31986 -26160 32000
rect -26240 31934 -26226 31986
rect -26174 31934 -26160 31986
rect -26240 31920 -26160 31934
rect -26080 31986 -26000 32000
rect -26080 31934 -26066 31986
rect -26014 31934 -26000 31986
rect -26080 31920 -26000 31934
rect -25920 31986 -25840 32000
rect -25920 31934 -25906 31986
rect -25854 31934 -25840 31986
rect -25920 31920 -25840 31934
rect -25760 31986 -25680 32000
rect -25760 31934 -25746 31986
rect -25694 31934 -25680 31986
rect -25760 31920 -25680 31934
rect -25600 31986 -25520 32000
rect -25600 31934 -25586 31986
rect -25534 31934 -25520 31986
rect -25600 31920 -25520 31934
rect -25440 31986 -25360 32000
rect -25440 31934 -25426 31986
rect -25374 31934 -25360 31986
rect -25440 31920 -25360 31934
rect -25280 31986 -25200 32000
rect -25280 31934 -25266 31986
rect -25214 31934 -25200 31986
rect -25280 31920 -25200 31934
rect -25120 31986 -25040 32000
rect -25120 31934 -25106 31986
rect -25054 31934 -25040 31986
rect -25120 31920 -25040 31934
rect -24960 31986 -24880 32000
rect -24960 31934 -24946 31986
rect -24894 31934 -24880 31986
rect -24960 31920 -24880 31934
rect -24800 31986 -24720 32000
rect -24800 31934 -24786 31986
rect -24734 31934 -24720 31986
rect -24800 31920 -24720 31934
rect -24640 31986 -24560 32000
rect -24640 31934 -24626 31986
rect -24574 31934 -24560 31986
rect -24640 31920 -24560 31934
rect -24480 31986 -24400 32000
rect -24480 31934 -24466 31986
rect -24414 31934 -24400 31986
rect -24480 31920 -24400 31934
rect -24320 31986 -24240 32000
rect -24320 31934 -24306 31986
rect -24254 31934 -24240 31986
rect -24320 31920 -24240 31934
rect -24160 31986 -24080 32000
rect -24160 31934 -24146 31986
rect -24094 31934 -24080 31986
rect -24160 31920 -24080 31934
rect -24000 31986 -23920 32000
rect -24000 31934 -23986 31986
rect -23934 31934 -23920 31986
rect -24000 31920 -23920 31934
rect -23840 31986 -23760 32000
rect -23840 31934 -23826 31986
rect -23774 31934 -23760 31986
rect -23840 31920 -23760 31934
rect -23680 31986 -23600 32000
rect -23680 31934 -23666 31986
rect -23614 31934 -23600 31986
rect -23680 31920 -23600 31934
rect -23520 31986 -23440 32000
rect -23520 31934 -23506 31986
rect -23454 31934 -23440 31986
rect -23520 31920 -23440 31934
rect -23360 31986 -23280 32000
rect -23360 31934 -23346 31986
rect -23294 31934 -23280 31986
rect -23360 31920 -23280 31934
rect -23200 31986 -23120 32000
rect -23200 31934 -23186 31986
rect -23134 31934 -23120 31986
rect -23200 31920 -23120 31934
rect -23040 31986 -22960 32000
rect -23040 31934 -23026 31986
rect -22974 31934 -22960 31986
rect -23040 31920 -22960 31934
rect -22880 31986 -22800 32000
rect -22880 31934 -22866 31986
rect -22814 31934 -22800 31986
rect -22880 31920 -22800 31934
rect -22720 31986 -22640 32000
rect -22720 31934 -22706 31986
rect -22654 31934 -22640 31986
rect -22720 31920 -22640 31934
rect -22560 31986 -22480 32000
rect -22560 31934 -22546 31986
rect -22494 31934 -22480 31986
rect -22560 31920 -22480 31934
rect -22400 31986 -22320 32000
rect -22400 31934 -22386 31986
rect -22334 31934 -22320 31986
rect -22400 31920 -22320 31934
rect -22240 31986 -22160 32000
rect -22240 31934 -22226 31986
rect -22174 31934 -22160 31986
rect -22240 31920 -22160 31934
rect -22080 31986 -22000 32000
rect -22080 31934 -22066 31986
rect -22014 31934 -22000 31986
rect -22080 31920 -22000 31934
rect -21920 31986 -21840 32000
rect -21920 31934 -21906 31986
rect -21854 31934 -21840 31986
rect -21920 31920 -21840 31934
rect -21760 31986 -21680 32000
rect -21760 31934 -21746 31986
rect -21694 31934 -21680 31986
rect -21760 31920 -21680 31934
rect -21600 31986 -21520 32000
rect -21600 31934 -21586 31986
rect -21534 31934 -21520 31986
rect -21600 31920 -21520 31934
rect -21440 31986 -21360 32000
rect -21440 31934 -21426 31986
rect -21374 31934 -21360 31986
rect -21440 31920 -21360 31934
rect -21280 31986 -21200 32000
rect -21280 31934 -21266 31986
rect -21214 31934 -21200 31986
rect -21280 31920 -21200 31934
rect -21120 31986 -21040 32000
rect -21120 31934 -21106 31986
rect -21054 31934 -21040 31986
rect -21120 31920 -21040 31934
rect -20960 31986 -20880 32000
rect -20960 31934 -20946 31986
rect -20894 31934 -20880 31986
rect -20960 31920 -20880 31934
rect -20800 31986 -20720 32000
rect -20800 31934 -20786 31986
rect -20734 31934 -20720 31986
rect -20800 31920 -20720 31934
rect -20640 31986 -20560 32000
rect -20640 31934 -20626 31986
rect -20574 31934 -20560 31986
rect -20640 31920 -20560 31934
rect -20480 31986 -20400 32000
rect -20480 31934 -20466 31986
rect -20414 31934 -20400 31986
rect -20480 31920 -20400 31934
rect -20320 31986 -20240 32000
rect -20320 31934 -20306 31986
rect -20254 31934 -20240 31986
rect -20320 31920 -20240 31934
rect -20160 31986 -20080 32000
rect -20160 31934 -20146 31986
rect -20094 31934 -20080 31986
rect -20160 31920 -20080 31934
rect -20000 31986 -19920 32000
rect -20000 31934 -19986 31986
rect -19934 31934 -19920 31986
rect -20000 31920 -19920 31934
rect -19840 31986 -19760 32000
rect -19840 31934 -19826 31986
rect -19774 31934 -19760 31986
rect -19840 31920 -19760 31934
rect -19680 31986 -19600 32000
rect -19680 31934 -19666 31986
rect -19614 31934 -19600 31986
rect -19680 31920 -19600 31934
rect -19520 31986 -19440 32000
rect -19520 31934 -19506 31986
rect -19454 31934 -19440 31986
rect -19520 31920 -19440 31934
rect -19360 31986 -19280 32000
rect -19360 31934 -19346 31986
rect -19294 31934 -19280 31986
rect -19360 31920 -19280 31934
rect -19200 31986 -19120 32000
rect -19200 31934 -19186 31986
rect -19134 31934 -19120 31986
rect -19200 31920 -19120 31934
rect -19040 31986 -18960 32000
rect -19040 31934 -19026 31986
rect -18974 31934 -18960 31986
rect -19040 31920 -18960 31934
rect -18880 31986 -18800 32000
rect -18880 31934 -18866 31986
rect -18814 31934 -18800 31986
rect -18880 31920 -18800 31934
rect -18720 31986 -18640 32000
rect -18720 31934 -18706 31986
rect -18654 31934 -18640 31986
rect -18720 31920 -18640 31934
rect -18560 31986 -18480 32000
rect -18560 31934 -18546 31986
rect -18494 31934 -18480 31986
rect -18560 31920 -18480 31934
rect -18400 31986 -18320 32000
rect -18400 31934 -18386 31986
rect -18334 31934 -18320 31986
rect -18400 31920 -18320 31934
rect -18240 31986 -18160 32000
rect -18240 31934 -18226 31986
rect -18174 31934 -18160 31986
rect -18240 31920 -18160 31934
rect -18080 31986 -18000 32000
rect -18080 31934 -18066 31986
rect -18014 31934 -18000 31986
rect -18080 31920 -18000 31934
rect -17920 31986 -17840 32000
rect -17920 31934 -17906 31986
rect -17854 31934 -17840 31986
rect -17920 31920 -17840 31934
rect -17760 31986 -17680 32000
rect -17760 31934 -17746 31986
rect -17694 31934 -17680 31986
rect -17760 31920 -17680 31934
rect -17600 31986 -17520 32000
rect -17600 31934 -17586 31986
rect -17534 31934 -17520 31986
rect -17600 31920 -17520 31934
rect -17440 31986 -17360 32000
rect -17440 31934 -17426 31986
rect -17374 31934 -17360 31986
rect -17440 31920 -17360 31934
rect -17280 31986 -17200 32000
rect -17280 31934 -17266 31986
rect -17214 31934 -17200 31986
rect -17280 31920 -17200 31934
rect -17120 31986 -17040 32000
rect -17120 31934 -17106 31986
rect -17054 31934 -17040 31986
rect -17120 31920 -17040 31934
rect -16960 31986 -16880 32000
rect -16960 31934 -16946 31986
rect -16894 31934 -16880 31986
rect -16960 31920 -16880 31934
rect -16800 31986 -16720 32000
rect -16800 31934 -16786 31986
rect -16734 31934 -16720 31986
rect -16800 31920 -16720 31934
rect -16640 31986 -16560 32000
rect -16640 31934 -16626 31986
rect -16574 31934 -16560 31986
rect -16640 31920 -16560 31934
rect -16480 31986 -16400 32000
rect -16480 31934 -16466 31986
rect -16414 31934 -16400 31986
rect -16480 31920 -16400 31934
rect -16320 31986 -16240 32000
rect -16320 31934 -16306 31986
rect -16254 31934 -16240 31986
rect -16320 31920 -16240 31934
rect -16160 31986 -16080 32000
rect -16160 31934 -16146 31986
rect -16094 31934 -16080 31986
rect -16160 31920 -16080 31934
rect -16000 31986 -15920 32000
rect -16000 31934 -15986 31986
rect -15934 31934 -15920 31986
rect -16000 31920 -15920 31934
rect -15840 31986 -15760 32000
rect -15840 31934 -15826 31986
rect -15774 31934 -15760 31986
rect -15840 31920 -15760 31934
rect -15680 31986 -15600 32000
rect -15680 31934 -15666 31986
rect -15614 31934 -15600 31986
rect -15680 31920 -15600 31934
rect -15520 31986 -15440 32000
rect -15520 31934 -15506 31986
rect -15454 31934 -15440 31986
rect -15520 31920 -15440 31934
rect -15360 31986 -15280 32000
rect -15360 31934 -15346 31986
rect -15294 31934 -15280 31986
rect -15360 31920 -15280 31934
rect -15200 31986 -15120 32000
rect -15200 31934 -15186 31986
rect -15134 31934 -15120 31986
rect -15200 31920 -15120 31934
rect -15040 31986 -14960 32000
rect -15040 31934 -15026 31986
rect -14974 31934 -14960 31986
rect -15040 31920 -14960 31934
rect -14880 31986 -14800 32000
rect -14880 31934 -14866 31986
rect -14814 31934 -14800 31986
rect -14880 31920 -14800 31934
rect -14720 31986 -14640 32000
rect -14720 31934 -14706 31986
rect -14654 31934 -14640 31986
rect -14720 31920 -14640 31934
rect -14560 31986 -14480 32000
rect -14560 31934 -14546 31986
rect -14494 31934 -14480 31986
rect -14560 31920 -14480 31934
rect -14400 31986 -14320 32000
rect -14400 31934 -14386 31986
rect -14334 31934 -14320 31986
rect -14400 31920 -14320 31934
rect -14240 31986 -14160 32000
rect -14240 31934 -14226 31986
rect -14174 31934 -14160 31986
rect -14240 31920 -14160 31934
rect -14080 31986 -14000 32000
rect -14080 31934 -14066 31986
rect -14014 31934 -14000 31986
rect -14080 31920 -14000 31934
rect -13920 31986 -13840 32000
rect -13920 31934 -13906 31986
rect -13854 31934 -13840 31986
rect -13920 31920 -13840 31934
rect -13760 31986 -13680 32000
rect -13760 31934 -13746 31986
rect -13694 31934 -13680 31986
rect -13760 31920 -13680 31934
rect -13600 31986 -13520 32000
rect -13600 31934 -13586 31986
rect -13534 31934 -13520 31986
rect -13600 31920 -13520 31934
rect -13440 31986 -13360 32000
rect -13440 31934 -13426 31986
rect -13374 31934 -13360 31986
rect -13440 31920 -13360 31934
rect -13280 31986 -13200 32000
rect -13280 31934 -13266 31986
rect -13214 31934 -13200 31986
rect -13280 31920 -13200 31934
rect -13120 31986 -13040 32000
rect -13120 31934 -13106 31986
rect -13054 31934 -13040 31986
rect -13120 31920 -13040 31934
rect -12960 31986 -12880 32000
rect -12960 31934 -12946 31986
rect -12894 31934 -12880 31986
rect -12960 31920 -12880 31934
rect -12800 31986 -12720 32000
rect -12800 31934 -12786 31986
rect -12734 31934 -12720 31986
rect -12800 31920 -12720 31934
rect -12640 31986 -12560 32000
rect -12640 31934 -12626 31986
rect -12574 31934 -12560 31986
rect -12640 31920 -12560 31934
rect -12480 31986 -12400 32000
rect -12480 31934 -12466 31986
rect -12414 31934 -12400 31986
rect -12480 31920 -12400 31934
rect -12320 31986 -12240 32000
rect -12320 31934 -12306 31986
rect -12254 31934 -12240 31986
rect -12320 31920 -12240 31934
rect -12160 31986 -12080 32000
rect -12160 31934 -12146 31986
rect -12094 31934 -12080 31986
rect -12160 31920 -12080 31934
rect -12000 31986 -11920 32000
rect -12000 31934 -11986 31986
rect -11934 31934 -11920 31986
rect -12000 31920 -11920 31934
rect -11840 31986 -11760 32000
rect -11840 31934 -11826 31986
rect -11774 31934 -11760 31986
rect -11840 31920 -11760 31934
rect -11680 31986 -11600 32000
rect -11680 31934 -11666 31986
rect -11614 31934 -11600 31986
rect -11680 31920 -11600 31934
rect -11520 31986 -11440 32000
rect -11520 31934 -11506 31986
rect -11454 31934 -11440 31986
rect -11520 31920 -11440 31934
rect -11360 31986 -11280 32000
rect -11360 31934 -11346 31986
rect -11294 31934 -11280 31986
rect -11360 31920 -11280 31934
rect -11200 31986 -11120 32000
rect -11200 31934 -11186 31986
rect -11134 31934 -11120 31986
rect -11200 31920 -11120 31934
rect -10880 31986 -10800 32000
rect -10880 31934 -10866 31986
rect -10814 31934 -10800 31986
rect -10880 31920 -10800 31934
rect -10720 31986 -10640 32000
rect -10720 31934 -10706 31986
rect -10654 31934 -10640 31986
rect -10720 31920 -10640 31934
rect -10560 31986 -10480 32000
rect -10560 31934 -10546 31986
rect -10494 31934 -10480 31986
rect -10560 31920 -10480 31934
rect -10400 31986 -10320 32000
rect -10400 31934 -10386 31986
rect -10334 31934 -10320 31986
rect -10400 31920 -10320 31934
rect -10240 31986 -10160 32000
rect -10240 31934 -10226 31986
rect -10174 31934 -10160 31986
rect -10240 31920 -10160 31934
rect -10080 31986 -10000 32000
rect -10080 31934 -10066 31986
rect -10014 31934 -10000 31986
rect -10080 31920 -10000 31934
rect -9920 31986 -9840 32000
rect -9920 31934 -9906 31986
rect -9854 31934 -9840 31986
rect -9920 31920 -9840 31934
rect -9760 31986 -9680 32000
rect -9760 31934 -9746 31986
rect -9694 31934 -9680 31986
rect -9760 31920 -9680 31934
rect -9600 31986 -9520 32000
rect -9600 31934 -9586 31986
rect -9534 31934 -9520 31986
rect -9600 31920 -9520 31934
rect -9440 31986 -9360 32000
rect -9440 31934 -9426 31986
rect -9374 31934 -9360 31986
rect -9440 31920 -9360 31934
rect -9280 31986 -9200 32000
rect -9280 31934 -9266 31986
rect -9214 31934 -9200 31986
rect -9280 31920 -9200 31934
rect -9120 31986 -9040 32000
rect -9120 31934 -9106 31986
rect -9054 31934 -9040 31986
rect -9120 31920 -9040 31934
rect -8960 31986 -8880 32000
rect -8960 31934 -8946 31986
rect -8894 31934 -8880 31986
rect -8960 31920 -8880 31934
rect -8800 31986 -8720 32000
rect -8800 31934 -8786 31986
rect -8734 31934 -8720 31986
rect -8800 31920 -8720 31934
rect -8640 31986 -8560 32000
rect -8640 31934 -8626 31986
rect -8574 31934 -8560 31986
rect -8640 31920 -8560 31934
rect -8480 31986 -8400 32000
rect -8480 31934 -8466 31986
rect -8414 31934 -8400 31986
rect -8480 31920 -8400 31934
rect -8320 31986 -8240 32000
rect -8320 31934 -8306 31986
rect -8254 31934 -8240 31986
rect -8320 31920 -8240 31934
rect -8160 31986 -8080 32000
rect -8160 31934 -8146 31986
rect -8094 31934 -8080 31986
rect -8160 31920 -8080 31934
rect -8000 31986 -7920 32000
rect -8000 31934 -7986 31986
rect -7934 31934 -7920 31986
rect -8000 31920 -7920 31934
rect -7840 31986 -7760 32000
rect -7840 31934 -7826 31986
rect -7774 31934 -7760 31986
rect -7840 31920 -7760 31934
rect -7680 31986 -7600 32000
rect -7680 31934 -7666 31986
rect -7614 31934 -7600 31986
rect -7680 31920 -7600 31934
rect -7520 31986 -7440 32000
rect -7520 31934 -7506 31986
rect -7454 31934 -7440 31986
rect -7520 31920 -7440 31934
rect -7360 31986 -7280 32000
rect -7360 31934 -7346 31986
rect -7294 31934 -7280 31986
rect -7360 31920 -7280 31934
rect -7200 31986 -7120 32000
rect -7200 31934 -7186 31986
rect -7134 31934 -7120 31986
rect -7200 31920 -7120 31934
rect -7040 31986 -6960 32000
rect -7040 31934 -7026 31986
rect -6974 31934 -6960 31986
rect -7040 31920 -6960 31934
rect -6880 31986 -6800 32000
rect -6880 31934 -6866 31986
rect -6814 31934 -6800 31986
rect -6880 31920 -6800 31934
rect -6720 31986 -6640 32000
rect -6720 31934 -6706 31986
rect -6654 31934 -6640 31986
rect -6720 31920 -6640 31934
rect -6560 31986 -6480 32000
rect -6560 31934 -6546 31986
rect -6494 31934 -6480 31986
rect -6560 31920 -6480 31934
rect -6400 31986 -6320 32000
rect -6400 31934 -6386 31986
rect -6334 31934 -6320 31986
rect -6400 31920 -6320 31934
rect -6240 31986 -6160 32000
rect -6240 31934 -6226 31986
rect -6174 31934 -6160 31986
rect -6240 31920 -6160 31934
rect -6080 31986 -6000 32000
rect -6080 31934 -6066 31986
rect -6014 31934 -6000 31986
rect -6080 31920 -6000 31934
rect -5920 31986 -5840 32000
rect -5920 31934 -5906 31986
rect -5854 31934 -5840 31986
rect -5920 31920 -5840 31934
rect -5760 31986 -5680 32000
rect -5760 31934 -5746 31986
rect -5694 31934 -5680 31986
rect -5760 31920 -5680 31934
rect -5600 31986 -5520 32000
rect -5600 31934 -5586 31986
rect -5534 31934 -5520 31986
rect -5600 31920 -5520 31934
rect -5440 31986 -5360 32000
rect -5440 31934 -5426 31986
rect -5374 31934 -5360 31986
rect -5440 31920 -5360 31934
rect -5280 31986 -5200 32000
rect -5280 31934 -5266 31986
rect -5214 31934 -5200 31986
rect -5280 31920 -5200 31934
rect -5120 31986 -5040 32000
rect -5120 31934 -5106 31986
rect -5054 31934 -5040 31986
rect -5120 31920 -5040 31934
rect -4960 31986 -4880 32000
rect -4960 31934 -4946 31986
rect -4894 31934 -4880 31986
rect -4960 31920 -4880 31934
rect -4800 31986 -4720 32000
rect -4800 31934 -4786 31986
rect -4734 31934 -4720 31986
rect -4800 31920 -4720 31934
rect -4640 31986 -4560 32000
rect -4640 31934 -4626 31986
rect -4574 31934 -4560 31986
rect -4640 31920 -4560 31934
rect -4480 31986 -4400 32000
rect -4480 31934 -4466 31986
rect -4414 31934 -4400 31986
rect -4480 31920 -4400 31934
rect -4320 31986 -4240 32000
rect -4320 31934 -4306 31986
rect -4254 31934 -4240 31986
rect -4320 31920 -4240 31934
rect -4160 31986 -4080 32000
rect -4160 31934 -4146 31986
rect -4094 31934 -4080 31986
rect -4160 31920 -4080 31934
rect -4000 31986 -3920 32000
rect -4000 31934 -3986 31986
rect -3934 31934 -3920 31986
rect -4000 31920 -3920 31934
rect -3680 31986 -3600 32000
rect -3680 31934 -3666 31986
rect -3614 31934 -3600 31986
rect -3680 31920 -3600 31934
rect -3520 31986 -3440 32000
rect -3520 31934 -3506 31986
rect -3454 31934 -3440 31986
rect -3520 31920 -3440 31934
rect -3360 31986 -3280 32000
rect -3360 31934 -3346 31986
rect -3294 31934 -3280 31986
rect -3360 31920 -3280 31934
rect -3200 31986 -3120 32000
rect -3200 31934 -3186 31986
rect -3134 31934 -3120 31986
rect -3200 31920 -3120 31934
rect -3040 31986 -2960 32000
rect -3040 31934 -3026 31986
rect -2974 31934 -2960 31986
rect -3040 31920 -2960 31934
rect -2880 31986 -2800 32000
rect -2880 31934 -2866 31986
rect -2814 31934 -2800 31986
rect -2880 31920 -2800 31934
rect -2720 31986 -2640 32000
rect -2720 31934 -2706 31986
rect -2654 31934 -2640 31986
rect -2720 31920 -2640 31934
rect -2400 31986 -2320 32000
rect -2400 31934 -2386 31986
rect -2334 31934 -2320 31986
rect -2400 31920 -2320 31934
rect -2080 31986 -2000 32000
rect -2080 31934 -2066 31986
rect -2014 31934 -2000 31986
rect -2080 31920 -2000 31934
rect -1760 31986 -1680 32000
rect -1760 31934 -1746 31986
rect -1694 31934 -1680 31986
rect -1760 31920 -1680 31934
rect -1440 31986 -1360 32000
rect -1440 31934 -1426 31986
rect -1374 31934 -1360 31986
rect -1440 31920 -1360 31934
rect -1120 31986 -1040 32000
rect -1120 31934 -1106 31986
rect -1054 31934 -1040 31986
rect -1120 31920 -1040 31934
<< via1 >>
rect -29906 42857 -29854 42866
rect -29906 42823 -29897 42857
rect -29897 42823 -29863 42857
rect -29863 42823 -29854 42857
rect -29906 42814 -29854 42823
rect -29746 42857 -29694 42866
rect -29746 42823 -29737 42857
rect -29737 42823 -29703 42857
rect -29703 42823 -29694 42857
rect -29746 42814 -29694 42823
rect -29586 42857 -29534 42866
rect -29586 42823 -29577 42857
rect -29577 42823 -29543 42857
rect -29543 42823 -29534 42857
rect -29586 42814 -29534 42823
rect -29426 42857 -29374 42866
rect -29426 42823 -29417 42857
rect -29417 42823 -29383 42857
rect -29383 42823 -29374 42857
rect -29426 42814 -29374 42823
rect -29266 42857 -29214 42866
rect -29266 42823 -29257 42857
rect -29257 42823 -29223 42857
rect -29223 42823 -29214 42857
rect -29266 42814 -29214 42823
rect -29106 42857 -29054 42866
rect -29106 42823 -29097 42857
rect -29097 42823 -29063 42857
rect -29063 42823 -29054 42857
rect -29106 42814 -29054 42823
rect -28946 42857 -28894 42866
rect -28946 42823 -28937 42857
rect -28937 42823 -28903 42857
rect -28903 42823 -28894 42857
rect -28946 42814 -28894 42823
rect -28786 42857 -28734 42866
rect -28786 42823 -28777 42857
rect -28777 42823 -28743 42857
rect -28743 42823 -28734 42857
rect -28786 42814 -28734 42823
rect -28626 42857 -28574 42866
rect -28626 42823 -28617 42857
rect -28617 42823 -28583 42857
rect -28583 42823 -28574 42857
rect -28626 42814 -28574 42823
rect -28466 42857 -28414 42866
rect -28466 42823 -28457 42857
rect -28457 42823 -28423 42857
rect -28423 42823 -28414 42857
rect -28466 42814 -28414 42823
rect -28306 42857 -28254 42866
rect -28306 42823 -28297 42857
rect -28297 42823 -28263 42857
rect -28263 42823 -28254 42857
rect -28306 42814 -28254 42823
rect -28146 42857 -28094 42866
rect -28146 42823 -28137 42857
rect -28137 42823 -28103 42857
rect -28103 42823 -28094 42857
rect -28146 42814 -28094 42823
rect -27986 42857 -27934 42866
rect -27986 42823 -27977 42857
rect -27977 42823 -27943 42857
rect -27943 42823 -27934 42857
rect -27986 42814 -27934 42823
rect -27826 42857 -27774 42866
rect -27826 42823 -27817 42857
rect -27817 42823 -27783 42857
rect -27783 42823 -27774 42857
rect -27826 42814 -27774 42823
rect -27666 42857 -27614 42866
rect -27666 42823 -27657 42857
rect -27657 42823 -27623 42857
rect -27623 42823 -27614 42857
rect -27666 42814 -27614 42823
rect -27506 42857 -27454 42866
rect -27506 42823 -27497 42857
rect -27497 42823 -27463 42857
rect -27463 42823 -27454 42857
rect -27506 42814 -27454 42823
rect -27346 42857 -27294 42866
rect -27346 42823 -27337 42857
rect -27337 42823 -27303 42857
rect -27303 42823 -27294 42857
rect -27346 42814 -27294 42823
rect -27186 42857 -27134 42866
rect -27186 42823 -27177 42857
rect -27177 42823 -27143 42857
rect -27143 42823 -27134 42857
rect -27186 42814 -27134 42823
rect -27026 42857 -26974 42866
rect -27026 42823 -27017 42857
rect -27017 42823 -26983 42857
rect -26983 42823 -26974 42857
rect -27026 42814 -26974 42823
rect -26866 42857 -26814 42866
rect -26866 42823 -26857 42857
rect -26857 42823 -26823 42857
rect -26823 42823 -26814 42857
rect -26866 42814 -26814 42823
rect -26706 42857 -26654 42866
rect -26706 42823 -26697 42857
rect -26697 42823 -26663 42857
rect -26663 42823 -26654 42857
rect -26706 42814 -26654 42823
rect -26546 42857 -26494 42866
rect -26546 42823 -26537 42857
rect -26537 42823 -26503 42857
rect -26503 42823 -26494 42857
rect -26546 42814 -26494 42823
rect -26386 42857 -26334 42866
rect -26386 42823 -26377 42857
rect -26377 42823 -26343 42857
rect -26343 42823 -26334 42857
rect -26386 42814 -26334 42823
rect -26226 42857 -26174 42866
rect -26226 42823 -26217 42857
rect -26217 42823 -26183 42857
rect -26183 42823 -26174 42857
rect -26226 42814 -26174 42823
rect -26066 42857 -26014 42866
rect -26066 42823 -26057 42857
rect -26057 42823 -26023 42857
rect -26023 42823 -26014 42857
rect -26066 42814 -26014 42823
rect -25906 42857 -25854 42866
rect -25906 42823 -25897 42857
rect -25897 42823 -25863 42857
rect -25863 42823 -25854 42857
rect -25906 42814 -25854 42823
rect -25746 42857 -25694 42866
rect -25746 42823 -25737 42857
rect -25737 42823 -25703 42857
rect -25703 42823 -25694 42857
rect -25746 42814 -25694 42823
rect -25586 42857 -25534 42866
rect -25586 42823 -25577 42857
rect -25577 42823 -25543 42857
rect -25543 42823 -25534 42857
rect -25586 42814 -25534 42823
rect -25426 42857 -25374 42866
rect -25426 42823 -25417 42857
rect -25417 42823 -25383 42857
rect -25383 42823 -25374 42857
rect -25426 42814 -25374 42823
rect -25266 42857 -25214 42866
rect -25266 42823 -25257 42857
rect -25257 42823 -25223 42857
rect -25223 42823 -25214 42857
rect -25266 42814 -25214 42823
rect -25106 42857 -25054 42866
rect -25106 42823 -25097 42857
rect -25097 42823 -25063 42857
rect -25063 42823 -25054 42857
rect -25106 42814 -25054 42823
rect -24946 42857 -24894 42866
rect -24946 42823 -24937 42857
rect -24937 42823 -24903 42857
rect -24903 42823 -24894 42857
rect -24946 42814 -24894 42823
rect -24786 42857 -24734 42866
rect -24786 42823 -24777 42857
rect -24777 42823 -24743 42857
rect -24743 42823 -24734 42857
rect -24786 42814 -24734 42823
rect -24626 42857 -24574 42866
rect -24626 42823 -24617 42857
rect -24617 42823 -24583 42857
rect -24583 42823 -24574 42857
rect -24626 42814 -24574 42823
rect -24466 42857 -24414 42866
rect -24466 42823 -24457 42857
rect -24457 42823 -24423 42857
rect -24423 42823 -24414 42857
rect -24466 42814 -24414 42823
rect -24306 42857 -24254 42866
rect -24306 42823 -24297 42857
rect -24297 42823 -24263 42857
rect -24263 42823 -24254 42857
rect -24306 42814 -24254 42823
rect -24146 42857 -24094 42866
rect -24146 42823 -24137 42857
rect -24137 42823 -24103 42857
rect -24103 42823 -24094 42857
rect -24146 42814 -24094 42823
rect -23986 42857 -23934 42866
rect -23986 42823 -23977 42857
rect -23977 42823 -23943 42857
rect -23943 42823 -23934 42857
rect -23986 42814 -23934 42823
rect -23826 42857 -23774 42866
rect -23826 42823 -23817 42857
rect -23817 42823 -23783 42857
rect -23783 42823 -23774 42857
rect -23826 42814 -23774 42823
rect -23666 42857 -23614 42866
rect -23666 42823 -23657 42857
rect -23657 42823 -23623 42857
rect -23623 42823 -23614 42857
rect -23666 42814 -23614 42823
rect -23506 42857 -23454 42866
rect -23506 42823 -23497 42857
rect -23497 42823 -23463 42857
rect -23463 42823 -23454 42857
rect -23506 42814 -23454 42823
rect -23346 42857 -23294 42866
rect -23346 42823 -23337 42857
rect -23337 42823 -23303 42857
rect -23303 42823 -23294 42857
rect -23346 42814 -23294 42823
rect -23186 42857 -23134 42866
rect -23186 42823 -23177 42857
rect -23177 42823 -23143 42857
rect -23143 42823 -23134 42857
rect -23186 42814 -23134 42823
rect -23026 42857 -22974 42866
rect -23026 42823 -23017 42857
rect -23017 42823 -22983 42857
rect -22983 42823 -22974 42857
rect -23026 42814 -22974 42823
rect -22866 42857 -22814 42866
rect -22866 42823 -22857 42857
rect -22857 42823 -22823 42857
rect -22823 42823 -22814 42857
rect -22866 42814 -22814 42823
rect -22706 42857 -22654 42866
rect -22706 42823 -22697 42857
rect -22697 42823 -22663 42857
rect -22663 42823 -22654 42857
rect -22706 42814 -22654 42823
rect -22546 42857 -22494 42866
rect -22546 42823 -22537 42857
rect -22537 42823 -22503 42857
rect -22503 42823 -22494 42857
rect -22546 42814 -22494 42823
rect -22386 42857 -22334 42866
rect -22386 42823 -22377 42857
rect -22377 42823 -22343 42857
rect -22343 42823 -22334 42857
rect -22386 42814 -22334 42823
rect -22226 42857 -22174 42866
rect -22226 42823 -22217 42857
rect -22217 42823 -22183 42857
rect -22183 42823 -22174 42857
rect -22226 42814 -22174 42823
rect -22066 42857 -22014 42866
rect -22066 42823 -22057 42857
rect -22057 42823 -22023 42857
rect -22023 42823 -22014 42857
rect -22066 42814 -22014 42823
rect -21906 42857 -21854 42866
rect -21906 42823 -21897 42857
rect -21897 42823 -21863 42857
rect -21863 42823 -21854 42857
rect -21906 42814 -21854 42823
rect -21746 42857 -21694 42866
rect -21746 42823 -21737 42857
rect -21737 42823 -21703 42857
rect -21703 42823 -21694 42857
rect -21746 42814 -21694 42823
rect -21586 42857 -21534 42866
rect -21586 42823 -21577 42857
rect -21577 42823 -21543 42857
rect -21543 42823 -21534 42857
rect -21586 42814 -21534 42823
rect -21426 42857 -21374 42866
rect -21426 42823 -21417 42857
rect -21417 42823 -21383 42857
rect -21383 42823 -21374 42857
rect -21426 42814 -21374 42823
rect -21266 42857 -21214 42866
rect -21266 42823 -21257 42857
rect -21257 42823 -21223 42857
rect -21223 42823 -21214 42857
rect -21266 42814 -21214 42823
rect -21106 42857 -21054 42866
rect -21106 42823 -21097 42857
rect -21097 42823 -21063 42857
rect -21063 42823 -21054 42857
rect -21106 42814 -21054 42823
rect -20946 42857 -20894 42866
rect -20946 42823 -20937 42857
rect -20937 42823 -20903 42857
rect -20903 42823 -20894 42857
rect -20946 42814 -20894 42823
rect -20786 42857 -20734 42866
rect -20786 42823 -20777 42857
rect -20777 42823 -20743 42857
rect -20743 42823 -20734 42857
rect -20786 42814 -20734 42823
rect -20626 42857 -20574 42866
rect -20626 42823 -20617 42857
rect -20617 42823 -20583 42857
rect -20583 42823 -20574 42857
rect -20626 42814 -20574 42823
rect -20466 42857 -20414 42866
rect -20466 42823 -20457 42857
rect -20457 42823 -20423 42857
rect -20423 42823 -20414 42857
rect -20466 42814 -20414 42823
rect -20306 42857 -20254 42866
rect -20306 42823 -20297 42857
rect -20297 42823 -20263 42857
rect -20263 42823 -20254 42857
rect -20306 42814 -20254 42823
rect -20146 42857 -20094 42866
rect -20146 42823 -20137 42857
rect -20137 42823 -20103 42857
rect -20103 42823 -20094 42857
rect -20146 42814 -20094 42823
rect -19986 42857 -19934 42866
rect -19986 42823 -19977 42857
rect -19977 42823 -19943 42857
rect -19943 42823 -19934 42857
rect -19986 42814 -19934 42823
rect -19826 42857 -19774 42866
rect -19826 42823 -19817 42857
rect -19817 42823 -19783 42857
rect -19783 42823 -19774 42857
rect -19826 42814 -19774 42823
rect -19666 42857 -19614 42866
rect -19666 42823 -19657 42857
rect -19657 42823 -19623 42857
rect -19623 42823 -19614 42857
rect -19666 42814 -19614 42823
rect -19506 42857 -19454 42866
rect -19506 42823 -19497 42857
rect -19497 42823 -19463 42857
rect -19463 42823 -19454 42857
rect -19506 42814 -19454 42823
rect -19346 42857 -19294 42866
rect -19346 42823 -19337 42857
rect -19337 42823 -19303 42857
rect -19303 42823 -19294 42857
rect -19346 42814 -19294 42823
rect -19186 42857 -19134 42866
rect -19186 42823 -19177 42857
rect -19177 42823 -19143 42857
rect -19143 42823 -19134 42857
rect -19186 42814 -19134 42823
rect -19026 42857 -18974 42866
rect -19026 42823 -19017 42857
rect -19017 42823 -18983 42857
rect -18983 42823 -18974 42857
rect -19026 42814 -18974 42823
rect -18866 42857 -18814 42866
rect -18866 42823 -18857 42857
rect -18857 42823 -18823 42857
rect -18823 42823 -18814 42857
rect -18866 42814 -18814 42823
rect -18706 42857 -18654 42866
rect -18706 42823 -18697 42857
rect -18697 42823 -18663 42857
rect -18663 42823 -18654 42857
rect -18706 42814 -18654 42823
rect -18546 42857 -18494 42866
rect -18546 42823 -18537 42857
rect -18537 42823 -18503 42857
rect -18503 42823 -18494 42857
rect -18546 42814 -18494 42823
rect -18386 42857 -18334 42866
rect -18386 42823 -18377 42857
rect -18377 42823 -18343 42857
rect -18343 42823 -18334 42857
rect -18386 42814 -18334 42823
rect -18226 42857 -18174 42866
rect -18226 42823 -18217 42857
rect -18217 42823 -18183 42857
rect -18183 42823 -18174 42857
rect -18226 42814 -18174 42823
rect -18066 42857 -18014 42866
rect -18066 42823 -18057 42857
rect -18057 42823 -18023 42857
rect -18023 42823 -18014 42857
rect -18066 42814 -18014 42823
rect -17906 42857 -17854 42866
rect -17906 42823 -17897 42857
rect -17897 42823 -17863 42857
rect -17863 42823 -17854 42857
rect -17906 42814 -17854 42823
rect -17746 42857 -17694 42866
rect -17746 42823 -17737 42857
rect -17737 42823 -17703 42857
rect -17703 42823 -17694 42857
rect -17746 42814 -17694 42823
rect -17586 42857 -17534 42866
rect -17586 42823 -17577 42857
rect -17577 42823 -17543 42857
rect -17543 42823 -17534 42857
rect -17586 42814 -17534 42823
rect -17426 42857 -17374 42866
rect -17426 42823 -17417 42857
rect -17417 42823 -17383 42857
rect -17383 42823 -17374 42857
rect -17426 42814 -17374 42823
rect -17266 42857 -17214 42866
rect -17266 42823 -17257 42857
rect -17257 42823 -17223 42857
rect -17223 42823 -17214 42857
rect -17266 42814 -17214 42823
rect -17106 42857 -17054 42866
rect -17106 42823 -17097 42857
rect -17097 42823 -17063 42857
rect -17063 42823 -17054 42857
rect -17106 42814 -17054 42823
rect -16946 42857 -16894 42866
rect -16946 42823 -16937 42857
rect -16937 42823 -16903 42857
rect -16903 42823 -16894 42857
rect -16946 42814 -16894 42823
rect -16786 42857 -16734 42866
rect -16786 42823 -16777 42857
rect -16777 42823 -16743 42857
rect -16743 42823 -16734 42857
rect -16786 42814 -16734 42823
rect -16626 42857 -16574 42866
rect -16626 42823 -16617 42857
rect -16617 42823 -16583 42857
rect -16583 42823 -16574 42857
rect -16626 42814 -16574 42823
rect -16466 42857 -16414 42866
rect -16466 42823 -16457 42857
rect -16457 42823 -16423 42857
rect -16423 42823 -16414 42857
rect -16466 42814 -16414 42823
rect -16306 42857 -16254 42866
rect -16306 42823 -16297 42857
rect -16297 42823 -16263 42857
rect -16263 42823 -16254 42857
rect -16306 42814 -16254 42823
rect -16146 42857 -16094 42866
rect -16146 42823 -16137 42857
rect -16137 42823 -16103 42857
rect -16103 42823 -16094 42857
rect -16146 42814 -16094 42823
rect -15986 42857 -15934 42866
rect -15986 42823 -15977 42857
rect -15977 42823 -15943 42857
rect -15943 42823 -15934 42857
rect -15986 42814 -15934 42823
rect -15826 42857 -15774 42866
rect -15826 42823 -15817 42857
rect -15817 42823 -15783 42857
rect -15783 42823 -15774 42857
rect -15826 42814 -15774 42823
rect -15666 42857 -15614 42866
rect -15666 42823 -15657 42857
rect -15657 42823 -15623 42857
rect -15623 42823 -15614 42857
rect -15666 42814 -15614 42823
rect -15506 42857 -15454 42866
rect -15506 42823 -15497 42857
rect -15497 42823 -15463 42857
rect -15463 42823 -15454 42857
rect -15506 42814 -15454 42823
rect -15346 42857 -15294 42866
rect -15346 42823 -15337 42857
rect -15337 42823 -15303 42857
rect -15303 42823 -15294 42857
rect -15346 42814 -15294 42823
rect -15186 42857 -15134 42866
rect -15186 42823 -15177 42857
rect -15177 42823 -15143 42857
rect -15143 42823 -15134 42857
rect -15186 42814 -15134 42823
rect -15026 42857 -14974 42866
rect -15026 42823 -15017 42857
rect -15017 42823 -14983 42857
rect -14983 42823 -14974 42857
rect -15026 42814 -14974 42823
rect -14866 42857 -14814 42866
rect -14866 42823 -14857 42857
rect -14857 42823 -14823 42857
rect -14823 42823 -14814 42857
rect -14866 42814 -14814 42823
rect -14706 42857 -14654 42866
rect -14706 42823 -14697 42857
rect -14697 42823 -14663 42857
rect -14663 42823 -14654 42857
rect -14706 42814 -14654 42823
rect -14546 42857 -14494 42866
rect -14546 42823 -14537 42857
rect -14537 42823 -14503 42857
rect -14503 42823 -14494 42857
rect -14546 42814 -14494 42823
rect -14386 42857 -14334 42866
rect -14386 42823 -14377 42857
rect -14377 42823 -14343 42857
rect -14343 42823 -14334 42857
rect -14386 42814 -14334 42823
rect -14226 42857 -14174 42866
rect -14226 42823 -14217 42857
rect -14217 42823 -14183 42857
rect -14183 42823 -14174 42857
rect -14226 42814 -14174 42823
rect -14066 42857 -14014 42866
rect -14066 42823 -14057 42857
rect -14057 42823 -14023 42857
rect -14023 42823 -14014 42857
rect -14066 42814 -14014 42823
rect -13906 42857 -13854 42866
rect -13906 42823 -13897 42857
rect -13897 42823 -13863 42857
rect -13863 42823 -13854 42857
rect -13906 42814 -13854 42823
rect -13746 42857 -13694 42866
rect -13746 42823 -13737 42857
rect -13737 42823 -13703 42857
rect -13703 42823 -13694 42857
rect -13746 42814 -13694 42823
rect -13586 42857 -13534 42866
rect -13586 42823 -13577 42857
rect -13577 42823 -13543 42857
rect -13543 42823 -13534 42857
rect -13586 42814 -13534 42823
rect -13426 42857 -13374 42866
rect -13426 42823 -13417 42857
rect -13417 42823 -13383 42857
rect -13383 42823 -13374 42857
rect -13426 42814 -13374 42823
rect -13266 42857 -13214 42866
rect -13266 42823 -13257 42857
rect -13257 42823 -13223 42857
rect -13223 42823 -13214 42857
rect -13266 42814 -13214 42823
rect -13106 42857 -13054 42866
rect -13106 42823 -13097 42857
rect -13097 42823 -13063 42857
rect -13063 42823 -13054 42857
rect -13106 42814 -13054 42823
rect -12946 42857 -12894 42866
rect -12946 42823 -12937 42857
rect -12937 42823 -12903 42857
rect -12903 42823 -12894 42857
rect -12946 42814 -12894 42823
rect -12786 42857 -12734 42866
rect -12786 42823 -12777 42857
rect -12777 42823 -12743 42857
rect -12743 42823 -12734 42857
rect -12786 42814 -12734 42823
rect -12626 42857 -12574 42866
rect -12626 42823 -12617 42857
rect -12617 42823 -12583 42857
rect -12583 42823 -12574 42857
rect -12626 42814 -12574 42823
rect -12466 42857 -12414 42866
rect -12466 42823 -12457 42857
rect -12457 42823 -12423 42857
rect -12423 42823 -12414 42857
rect -12466 42814 -12414 42823
rect -12306 42857 -12254 42866
rect -12306 42823 -12297 42857
rect -12297 42823 -12263 42857
rect -12263 42823 -12254 42857
rect -12306 42814 -12254 42823
rect -11346 42857 -11294 42866
rect -11346 42823 -11337 42857
rect -11337 42823 -11303 42857
rect -11303 42823 -11294 42857
rect -11346 42814 -11294 42823
rect -11186 42857 -11134 42866
rect -11186 42823 -11177 42857
rect -11177 42823 -11143 42857
rect -11143 42823 -11134 42857
rect -11186 42814 -11134 42823
rect -11026 42857 -10974 42866
rect -11026 42823 -11017 42857
rect -11017 42823 -10983 42857
rect -10983 42823 -10974 42857
rect -11026 42814 -10974 42823
rect -10866 42857 -10814 42866
rect -10866 42823 -10857 42857
rect -10857 42823 -10823 42857
rect -10823 42823 -10814 42857
rect -10866 42814 -10814 42823
rect -10706 42857 -10654 42866
rect -10706 42823 -10697 42857
rect -10697 42823 -10663 42857
rect -10663 42823 -10654 42857
rect -10706 42814 -10654 42823
rect -10546 42857 -10494 42866
rect -10546 42823 -10537 42857
rect -10537 42823 -10503 42857
rect -10503 42823 -10494 42857
rect -10546 42814 -10494 42823
rect -10386 42857 -10334 42866
rect -10386 42823 -10377 42857
rect -10377 42823 -10343 42857
rect -10343 42823 -10334 42857
rect -10386 42814 -10334 42823
rect -10226 42857 -10174 42866
rect -10226 42823 -10217 42857
rect -10217 42823 -10183 42857
rect -10183 42823 -10174 42857
rect -10226 42814 -10174 42823
rect -10066 42857 -10014 42866
rect -10066 42823 -10057 42857
rect -10057 42823 -10023 42857
rect -10023 42823 -10014 42857
rect -10066 42814 -10014 42823
rect -9906 42857 -9854 42866
rect -9906 42823 -9897 42857
rect -9897 42823 -9863 42857
rect -9863 42823 -9854 42857
rect -9906 42814 -9854 42823
rect -9746 42857 -9694 42866
rect -9746 42823 -9737 42857
rect -9737 42823 -9703 42857
rect -9703 42823 -9694 42857
rect -9746 42814 -9694 42823
rect -9586 42857 -9534 42866
rect -9586 42823 -9577 42857
rect -9577 42823 -9543 42857
rect -9543 42823 -9534 42857
rect -9586 42814 -9534 42823
rect -9426 42857 -9374 42866
rect -9426 42823 -9417 42857
rect -9417 42823 -9383 42857
rect -9383 42823 -9374 42857
rect -9426 42814 -9374 42823
rect -9266 42857 -9214 42866
rect -9266 42823 -9257 42857
rect -9257 42823 -9223 42857
rect -9223 42823 -9214 42857
rect -9266 42814 -9214 42823
rect -9106 42857 -9054 42866
rect -9106 42823 -9097 42857
rect -9097 42823 -9063 42857
rect -9063 42823 -9054 42857
rect -9106 42814 -9054 42823
rect -8946 42857 -8894 42866
rect -8946 42823 -8937 42857
rect -8937 42823 -8903 42857
rect -8903 42823 -8894 42857
rect -8946 42814 -8894 42823
rect -8786 42857 -8734 42866
rect -8786 42823 -8777 42857
rect -8777 42823 -8743 42857
rect -8743 42823 -8734 42857
rect -8786 42814 -8734 42823
rect -8626 42857 -8574 42866
rect -8626 42823 -8617 42857
rect -8617 42823 -8583 42857
rect -8583 42823 -8574 42857
rect -8626 42814 -8574 42823
rect -8466 42857 -8414 42866
rect -8466 42823 -8457 42857
rect -8457 42823 -8423 42857
rect -8423 42823 -8414 42857
rect -8466 42814 -8414 42823
rect -8306 42857 -8254 42866
rect -8306 42823 -8297 42857
rect -8297 42823 -8263 42857
rect -8263 42823 -8254 42857
rect -8306 42814 -8254 42823
rect -8146 42857 -8094 42866
rect -8146 42823 -8137 42857
rect -8137 42823 -8103 42857
rect -8103 42823 -8094 42857
rect -8146 42814 -8094 42823
rect -7986 42857 -7934 42866
rect -7986 42823 -7977 42857
rect -7977 42823 -7943 42857
rect -7943 42823 -7934 42857
rect -7986 42814 -7934 42823
rect -7826 42857 -7774 42866
rect -7826 42823 -7817 42857
rect -7817 42823 -7783 42857
rect -7783 42823 -7774 42857
rect -7826 42814 -7774 42823
rect -7666 42857 -7614 42866
rect -7666 42823 -7657 42857
rect -7657 42823 -7623 42857
rect -7623 42823 -7614 42857
rect -7666 42814 -7614 42823
rect -7506 42857 -7454 42866
rect -7506 42823 -7497 42857
rect -7497 42823 -7463 42857
rect -7463 42823 -7454 42857
rect -7506 42814 -7454 42823
rect -7346 42857 -7294 42866
rect -7346 42823 -7337 42857
rect -7337 42823 -7303 42857
rect -7303 42823 -7294 42857
rect -7346 42814 -7294 42823
rect -7186 42857 -7134 42866
rect -7186 42823 -7177 42857
rect -7177 42823 -7143 42857
rect -7143 42823 -7134 42857
rect -7186 42814 -7134 42823
rect -7026 42857 -6974 42866
rect -7026 42823 -7017 42857
rect -7017 42823 -6983 42857
rect -6983 42823 -6974 42857
rect -7026 42814 -6974 42823
rect -6866 42857 -6814 42866
rect -6866 42823 -6857 42857
rect -6857 42823 -6823 42857
rect -6823 42823 -6814 42857
rect -6866 42814 -6814 42823
rect -6706 42857 -6654 42866
rect -6706 42823 -6697 42857
rect -6697 42823 -6663 42857
rect -6663 42823 -6654 42857
rect -6706 42814 -6654 42823
rect -6546 42857 -6494 42866
rect -6546 42823 -6537 42857
rect -6537 42823 -6503 42857
rect -6503 42823 -6494 42857
rect -6546 42814 -6494 42823
rect -6386 42857 -6334 42866
rect -6386 42823 -6377 42857
rect -6377 42823 -6343 42857
rect -6343 42823 -6334 42857
rect -6386 42814 -6334 42823
rect -6226 42857 -6174 42866
rect -6226 42823 -6217 42857
rect -6217 42823 -6183 42857
rect -6183 42823 -6174 42857
rect -6226 42814 -6174 42823
rect -6066 42857 -6014 42866
rect -6066 42823 -6057 42857
rect -6057 42823 -6023 42857
rect -6023 42823 -6014 42857
rect -6066 42814 -6014 42823
rect -5906 42857 -5854 42866
rect -5906 42823 -5897 42857
rect -5897 42823 -5863 42857
rect -5863 42823 -5854 42857
rect -5906 42814 -5854 42823
rect -5746 42857 -5694 42866
rect -5746 42823 -5737 42857
rect -5737 42823 -5703 42857
rect -5703 42823 -5694 42857
rect -5746 42814 -5694 42823
rect -5586 42857 -5534 42866
rect -5586 42823 -5577 42857
rect -5577 42823 -5543 42857
rect -5543 42823 -5534 42857
rect -5586 42814 -5534 42823
rect -5426 42857 -5374 42866
rect -5426 42823 -5417 42857
rect -5417 42823 -5383 42857
rect -5383 42823 -5374 42857
rect -5426 42814 -5374 42823
rect -5266 42857 -5214 42866
rect -5266 42823 -5257 42857
rect -5257 42823 -5223 42857
rect -5223 42823 -5214 42857
rect -5266 42814 -5214 42823
rect -5106 42857 -5054 42866
rect -5106 42823 -5097 42857
rect -5097 42823 -5063 42857
rect -5063 42823 -5054 42857
rect -5106 42814 -5054 42823
rect -4946 42857 -4894 42866
rect -4946 42823 -4937 42857
rect -4937 42823 -4903 42857
rect -4903 42823 -4894 42857
rect -4946 42814 -4894 42823
rect -4786 42857 -4734 42866
rect -4786 42823 -4777 42857
rect -4777 42823 -4743 42857
rect -4743 42823 -4734 42857
rect -4786 42814 -4734 42823
rect -4626 42857 -4574 42866
rect -4626 42823 -4617 42857
rect -4617 42823 -4583 42857
rect -4583 42823 -4574 42857
rect -4626 42814 -4574 42823
rect -4466 42857 -4414 42866
rect -4466 42823 -4457 42857
rect -4457 42823 -4423 42857
rect -4423 42823 -4414 42857
rect -4466 42814 -4414 42823
rect -4306 42857 -4254 42866
rect -4306 42823 -4297 42857
rect -4297 42823 -4263 42857
rect -4263 42823 -4254 42857
rect -4306 42814 -4254 42823
rect -4146 42857 -4094 42866
rect -4146 42823 -4137 42857
rect -4137 42823 -4103 42857
rect -4103 42823 -4094 42857
rect -4146 42814 -4094 42823
rect -3986 42857 -3934 42866
rect -3986 42823 -3977 42857
rect -3977 42823 -3943 42857
rect -3943 42823 -3934 42857
rect -3986 42814 -3934 42823
rect -3666 42857 -3614 42866
rect -3666 42823 -3657 42857
rect -3657 42823 -3623 42857
rect -3623 42823 -3614 42857
rect -3666 42814 -3614 42823
rect -3506 42857 -3454 42866
rect -3506 42823 -3497 42857
rect -3497 42823 -3463 42857
rect -3463 42823 -3454 42857
rect -3506 42814 -3454 42823
rect -3346 42857 -3294 42866
rect -3346 42823 -3337 42857
rect -3337 42823 -3303 42857
rect -3303 42823 -3294 42857
rect -3346 42814 -3294 42823
rect -3026 42857 -2974 42866
rect -3026 42823 -3017 42857
rect -3017 42823 -2983 42857
rect -2983 42823 -2974 42857
rect -3026 42814 -2974 42823
rect -2706 42857 -2654 42866
rect -2706 42823 -2697 42857
rect -2697 42823 -2663 42857
rect -2663 42823 -2654 42857
rect -2706 42814 -2654 42823
rect -2546 42857 -2494 42866
rect -2546 42823 -2537 42857
rect -2537 42823 -2503 42857
rect -2503 42823 -2494 42857
rect -2546 42814 -2494 42823
rect -2386 42857 -2334 42866
rect -2386 42823 -2377 42857
rect -2377 42823 -2343 42857
rect -2343 42823 -2334 42857
rect -2386 42814 -2334 42823
rect -2226 42857 -2174 42866
rect -2226 42823 -2217 42857
rect -2217 42823 -2183 42857
rect -2183 42823 -2174 42857
rect -2226 42814 -2174 42823
rect -2066 42857 -2014 42866
rect -2066 42823 -2057 42857
rect -2057 42823 -2023 42857
rect -2023 42823 -2014 42857
rect -2066 42814 -2014 42823
rect -1746 42857 -1694 42866
rect -1746 42823 -1737 42857
rect -1737 42823 -1703 42857
rect -1703 42823 -1694 42857
rect -1746 42814 -1694 42823
rect -1426 42857 -1374 42866
rect -1426 42823 -1417 42857
rect -1417 42823 -1383 42857
rect -1383 42823 -1374 42857
rect -1426 42814 -1374 42823
rect -1106 42857 -1054 42866
rect -1106 42823 -1097 42857
rect -1097 42823 -1063 42857
rect -1063 42823 -1054 42857
rect -1106 42814 -1054 42823
rect -29906 42537 -29854 42546
rect -29906 42503 -29897 42537
rect -29897 42503 -29863 42537
rect -29863 42503 -29854 42537
rect -29906 42494 -29854 42503
rect -29746 42537 -29694 42546
rect -29746 42503 -29737 42537
rect -29737 42503 -29703 42537
rect -29703 42503 -29694 42537
rect -29746 42494 -29694 42503
rect -29586 42537 -29534 42546
rect -29586 42503 -29577 42537
rect -29577 42503 -29543 42537
rect -29543 42503 -29534 42537
rect -29586 42494 -29534 42503
rect -29426 42537 -29374 42546
rect -29426 42503 -29417 42537
rect -29417 42503 -29383 42537
rect -29383 42503 -29374 42537
rect -29426 42494 -29374 42503
rect -29266 42537 -29214 42546
rect -29266 42503 -29257 42537
rect -29257 42503 -29223 42537
rect -29223 42503 -29214 42537
rect -29266 42494 -29214 42503
rect -29106 42537 -29054 42546
rect -29106 42503 -29097 42537
rect -29097 42503 -29063 42537
rect -29063 42503 -29054 42537
rect -29106 42494 -29054 42503
rect -28946 42537 -28894 42546
rect -28946 42503 -28937 42537
rect -28937 42503 -28903 42537
rect -28903 42503 -28894 42537
rect -28946 42494 -28894 42503
rect -28786 42537 -28734 42546
rect -28786 42503 -28777 42537
rect -28777 42503 -28743 42537
rect -28743 42503 -28734 42537
rect -28786 42494 -28734 42503
rect -28626 42537 -28574 42546
rect -28626 42503 -28617 42537
rect -28617 42503 -28583 42537
rect -28583 42503 -28574 42537
rect -28626 42494 -28574 42503
rect -28466 42537 -28414 42546
rect -28466 42503 -28457 42537
rect -28457 42503 -28423 42537
rect -28423 42503 -28414 42537
rect -28466 42494 -28414 42503
rect -28306 42537 -28254 42546
rect -28306 42503 -28297 42537
rect -28297 42503 -28263 42537
rect -28263 42503 -28254 42537
rect -28306 42494 -28254 42503
rect -28146 42537 -28094 42546
rect -28146 42503 -28137 42537
rect -28137 42503 -28103 42537
rect -28103 42503 -28094 42537
rect -28146 42494 -28094 42503
rect -27986 42537 -27934 42546
rect -27986 42503 -27977 42537
rect -27977 42503 -27943 42537
rect -27943 42503 -27934 42537
rect -27986 42494 -27934 42503
rect -27826 42537 -27774 42546
rect -27826 42503 -27817 42537
rect -27817 42503 -27783 42537
rect -27783 42503 -27774 42537
rect -27826 42494 -27774 42503
rect -27666 42537 -27614 42546
rect -27666 42503 -27657 42537
rect -27657 42503 -27623 42537
rect -27623 42503 -27614 42537
rect -27666 42494 -27614 42503
rect -27506 42537 -27454 42546
rect -27506 42503 -27497 42537
rect -27497 42503 -27463 42537
rect -27463 42503 -27454 42537
rect -27506 42494 -27454 42503
rect -27346 42537 -27294 42546
rect -27346 42503 -27337 42537
rect -27337 42503 -27303 42537
rect -27303 42503 -27294 42537
rect -27346 42494 -27294 42503
rect -27186 42537 -27134 42546
rect -27186 42503 -27177 42537
rect -27177 42503 -27143 42537
rect -27143 42503 -27134 42537
rect -27186 42494 -27134 42503
rect -27026 42537 -26974 42546
rect -27026 42503 -27017 42537
rect -27017 42503 -26983 42537
rect -26983 42503 -26974 42537
rect -27026 42494 -26974 42503
rect -26866 42537 -26814 42546
rect -26866 42503 -26857 42537
rect -26857 42503 -26823 42537
rect -26823 42503 -26814 42537
rect -26866 42494 -26814 42503
rect -26706 42537 -26654 42546
rect -26706 42503 -26697 42537
rect -26697 42503 -26663 42537
rect -26663 42503 -26654 42537
rect -26706 42494 -26654 42503
rect -26546 42537 -26494 42546
rect -26546 42503 -26537 42537
rect -26537 42503 -26503 42537
rect -26503 42503 -26494 42537
rect -26546 42494 -26494 42503
rect -26386 42537 -26334 42546
rect -26386 42503 -26377 42537
rect -26377 42503 -26343 42537
rect -26343 42503 -26334 42537
rect -26386 42494 -26334 42503
rect -26226 42537 -26174 42546
rect -26226 42503 -26217 42537
rect -26217 42503 -26183 42537
rect -26183 42503 -26174 42537
rect -26226 42494 -26174 42503
rect -26066 42537 -26014 42546
rect -26066 42503 -26057 42537
rect -26057 42503 -26023 42537
rect -26023 42503 -26014 42537
rect -26066 42494 -26014 42503
rect -25906 42537 -25854 42546
rect -25906 42503 -25897 42537
rect -25897 42503 -25863 42537
rect -25863 42503 -25854 42537
rect -25906 42494 -25854 42503
rect -25746 42537 -25694 42546
rect -25746 42503 -25737 42537
rect -25737 42503 -25703 42537
rect -25703 42503 -25694 42537
rect -25746 42494 -25694 42503
rect -25586 42537 -25534 42546
rect -25586 42503 -25577 42537
rect -25577 42503 -25543 42537
rect -25543 42503 -25534 42537
rect -25586 42494 -25534 42503
rect -25426 42537 -25374 42546
rect -25426 42503 -25417 42537
rect -25417 42503 -25383 42537
rect -25383 42503 -25374 42537
rect -25426 42494 -25374 42503
rect -25266 42537 -25214 42546
rect -25266 42503 -25257 42537
rect -25257 42503 -25223 42537
rect -25223 42503 -25214 42537
rect -25266 42494 -25214 42503
rect -25106 42537 -25054 42546
rect -25106 42503 -25097 42537
rect -25097 42503 -25063 42537
rect -25063 42503 -25054 42537
rect -25106 42494 -25054 42503
rect -24946 42537 -24894 42546
rect -24946 42503 -24937 42537
rect -24937 42503 -24903 42537
rect -24903 42503 -24894 42537
rect -24946 42494 -24894 42503
rect -24786 42537 -24734 42546
rect -24786 42503 -24777 42537
rect -24777 42503 -24743 42537
rect -24743 42503 -24734 42537
rect -24786 42494 -24734 42503
rect -24626 42537 -24574 42546
rect -24626 42503 -24617 42537
rect -24617 42503 -24583 42537
rect -24583 42503 -24574 42537
rect -24626 42494 -24574 42503
rect -24466 42537 -24414 42546
rect -24466 42503 -24457 42537
rect -24457 42503 -24423 42537
rect -24423 42503 -24414 42537
rect -24466 42494 -24414 42503
rect -24306 42537 -24254 42546
rect -24306 42503 -24297 42537
rect -24297 42503 -24263 42537
rect -24263 42503 -24254 42537
rect -24306 42494 -24254 42503
rect -24146 42537 -24094 42546
rect -24146 42503 -24137 42537
rect -24137 42503 -24103 42537
rect -24103 42503 -24094 42537
rect -24146 42494 -24094 42503
rect -23986 42537 -23934 42546
rect -23986 42503 -23977 42537
rect -23977 42503 -23943 42537
rect -23943 42503 -23934 42537
rect -23986 42494 -23934 42503
rect -23826 42537 -23774 42546
rect -23826 42503 -23817 42537
rect -23817 42503 -23783 42537
rect -23783 42503 -23774 42537
rect -23826 42494 -23774 42503
rect -23666 42537 -23614 42546
rect -23666 42503 -23657 42537
rect -23657 42503 -23623 42537
rect -23623 42503 -23614 42537
rect -23666 42494 -23614 42503
rect -23506 42537 -23454 42546
rect -23506 42503 -23497 42537
rect -23497 42503 -23463 42537
rect -23463 42503 -23454 42537
rect -23506 42494 -23454 42503
rect -23346 42537 -23294 42546
rect -23346 42503 -23337 42537
rect -23337 42503 -23303 42537
rect -23303 42503 -23294 42537
rect -23346 42494 -23294 42503
rect -23186 42537 -23134 42546
rect -23186 42503 -23177 42537
rect -23177 42503 -23143 42537
rect -23143 42503 -23134 42537
rect -23186 42494 -23134 42503
rect -23026 42537 -22974 42546
rect -23026 42503 -23017 42537
rect -23017 42503 -22983 42537
rect -22983 42503 -22974 42537
rect -23026 42494 -22974 42503
rect -22866 42537 -22814 42546
rect -22866 42503 -22857 42537
rect -22857 42503 -22823 42537
rect -22823 42503 -22814 42537
rect -22866 42494 -22814 42503
rect -22706 42537 -22654 42546
rect -22706 42503 -22697 42537
rect -22697 42503 -22663 42537
rect -22663 42503 -22654 42537
rect -22706 42494 -22654 42503
rect -22546 42537 -22494 42546
rect -22546 42503 -22537 42537
rect -22537 42503 -22503 42537
rect -22503 42503 -22494 42537
rect -22546 42494 -22494 42503
rect -22386 42537 -22334 42546
rect -22386 42503 -22377 42537
rect -22377 42503 -22343 42537
rect -22343 42503 -22334 42537
rect -22386 42494 -22334 42503
rect -22226 42537 -22174 42546
rect -22226 42503 -22217 42537
rect -22217 42503 -22183 42537
rect -22183 42503 -22174 42537
rect -22226 42494 -22174 42503
rect -22066 42537 -22014 42546
rect -22066 42503 -22057 42537
rect -22057 42503 -22023 42537
rect -22023 42503 -22014 42537
rect -22066 42494 -22014 42503
rect -21906 42537 -21854 42546
rect -21906 42503 -21897 42537
rect -21897 42503 -21863 42537
rect -21863 42503 -21854 42537
rect -21906 42494 -21854 42503
rect -21746 42537 -21694 42546
rect -21746 42503 -21737 42537
rect -21737 42503 -21703 42537
rect -21703 42503 -21694 42537
rect -21746 42494 -21694 42503
rect -21586 42537 -21534 42546
rect -21586 42503 -21577 42537
rect -21577 42503 -21543 42537
rect -21543 42503 -21534 42537
rect -21586 42494 -21534 42503
rect -21426 42537 -21374 42546
rect -21426 42503 -21417 42537
rect -21417 42503 -21383 42537
rect -21383 42503 -21374 42537
rect -21426 42494 -21374 42503
rect -21266 42537 -21214 42546
rect -21266 42503 -21257 42537
rect -21257 42503 -21223 42537
rect -21223 42503 -21214 42537
rect -21266 42494 -21214 42503
rect -21106 42537 -21054 42546
rect -21106 42503 -21097 42537
rect -21097 42503 -21063 42537
rect -21063 42503 -21054 42537
rect -21106 42494 -21054 42503
rect -20946 42537 -20894 42546
rect -20946 42503 -20937 42537
rect -20937 42503 -20903 42537
rect -20903 42503 -20894 42537
rect -20946 42494 -20894 42503
rect -20786 42537 -20734 42546
rect -20786 42503 -20777 42537
rect -20777 42503 -20743 42537
rect -20743 42503 -20734 42537
rect -20786 42494 -20734 42503
rect -20626 42537 -20574 42546
rect -20626 42503 -20617 42537
rect -20617 42503 -20583 42537
rect -20583 42503 -20574 42537
rect -20626 42494 -20574 42503
rect -20466 42537 -20414 42546
rect -20466 42503 -20457 42537
rect -20457 42503 -20423 42537
rect -20423 42503 -20414 42537
rect -20466 42494 -20414 42503
rect -20306 42537 -20254 42546
rect -20306 42503 -20297 42537
rect -20297 42503 -20263 42537
rect -20263 42503 -20254 42537
rect -20306 42494 -20254 42503
rect -20146 42537 -20094 42546
rect -20146 42503 -20137 42537
rect -20137 42503 -20103 42537
rect -20103 42503 -20094 42537
rect -20146 42494 -20094 42503
rect -19986 42537 -19934 42546
rect -19986 42503 -19977 42537
rect -19977 42503 -19943 42537
rect -19943 42503 -19934 42537
rect -19986 42494 -19934 42503
rect -19826 42537 -19774 42546
rect -19826 42503 -19817 42537
rect -19817 42503 -19783 42537
rect -19783 42503 -19774 42537
rect -19826 42494 -19774 42503
rect -19666 42537 -19614 42546
rect -19666 42503 -19657 42537
rect -19657 42503 -19623 42537
rect -19623 42503 -19614 42537
rect -19666 42494 -19614 42503
rect -19506 42537 -19454 42546
rect -19506 42503 -19497 42537
rect -19497 42503 -19463 42537
rect -19463 42503 -19454 42537
rect -19506 42494 -19454 42503
rect -19346 42537 -19294 42546
rect -19346 42503 -19337 42537
rect -19337 42503 -19303 42537
rect -19303 42503 -19294 42537
rect -19346 42494 -19294 42503
rect -19186 42537 -19134 42546
rect -19186 42503 -19177 42537
rect -19177 42503 -19143 42537
rect -19143 42503 -19134 42537
rect -19186 42494 -19134 42503
rect -19026 42537 -18974 42546
rect -19026 42503 -19017 42537
rect -19017 42503 -18983 42537
rect -18983 42503 -18974 42537
rect -19026 42494 -18974 42503
rect -18866 42537 -18814 42546
rect -18866 42503 -18857 42537
rect -18857 42503 -18823 42537
rect -18823 42503 -18814 42537
rect -18866 42494 -18814 42503
rect -18706 42537 -18654 42546
rect -18706 42503 -18697 42537
rect -18697 42503 -18663 42537
rect -18663 42503 -18654 42537
rect -18706 42494 -18654 42503
rect -18546 42537 -18494 42546
rect -18546 42503 -18537 42537
rect -18537 42503 -18503 42537
rect -18503 42503 -18494 42537
rect -18546 42494 -18494 42503
rect -18386 42537 -18334 42546
rect -18386 42503 -18377 42537
rect -18377 42503 -18343 42537
rect -18343 42503 -18334 42537
rect -18386 42494 -18334 42503
rect -18226 42537 -18174 42546
rect -18226 42503 -18217 42537
rect -18217 42503 -18183 42537
rect -18183 42503 -18174 42537
rect -18226 42494 -18174 42503
rect -18066 42537 -18014 42546
rect -18066 42503 -18057 42537
rect -18057 42503 -18023 42537
rect -18023 42503 -18014 42537
rect -18066 42494 -18014 42503
rect -17906 42537 -17854 42546
rect -17906 42503 -17897 42537
rect -17897 42503 -17863 42537
rect -17863 42503 -17854 42537
rect -17906 42494 -17854 42503
rect -17746 42537 -17694 42546
rect -17746 42503 -17737 42537
rect -17737 42503 -17703 42537
rect -17703 42503 -17694 42537
rect -17746 42494 -17694 42503
rect -17586 42537 -17534 42546
rect -17586 42503 -17577 42537
rect -17577 42503 -17543 42537
rect -17543 42503 -17534 42537
rect -17586 42494 -17534 42503
rect -17426 42537 -17374 42546
rect -17426 42503 -17417 42537
rect -17417 42503 -17383 42537
rect -17383 42503 -17374 42537
rect -17426 42494 -17374 42503
rect -17266 42537 -17214 42546
rect -17266 42503 -17257 42537
rect -17257 42503 -17223 42537
rect -17223 42503 -17214 42537
rect -17266 42494 -17214 42503
rect -17106 42537 -17054 42546
rect -17106 42503 -17097 42537
rect -17097 42503 -17063 42537
rect -17063 42503 -17054 42537
rect -17106 42494 -17054 42503
rect -16946 42537 -16894 42546
rect -16946 42503 -16937 42537
rect -16937 42503 -16903 42537
rect -16903 42503 -16894 42537
rect -16946 42494 -16894 42503
rect -16786 42537 -16734 42546
rect -16786 42503 -16777 42537
rect -16777 42503 -16743 42537
rect -16743 42503 -16734 42537
rect -16786 42494 -16734 42503
rect -16626 42537 -16574 42546
rect -16626 42503 -16617 42537
rect -16617 42503 -16583 42537
rect -16583 42503 -16574 42537
rect -16626 42494 -16574 42503
rect -16466 42537 -16414 42546
rect -16466 42503 -16457 42537
rect -16457 42503 -16423 42537
rect -16423 42503 -16414 42537
rect -16466 42494 -16414 42503
rect -16306 42537 -16254 42546
rect -16306 42503 -16297 42537
rect -16297 42503 -16263 42537
rect -16263 42503 -16254 42537
rect -16306 42494 -16254 42503
rect -16146 42537 -16094 42546
rect -16146 42503 -16137 42537
rect -16137 42503 -16103 42537
rect -16103 42503 -16094 42537
rect -16146 42494 -16094 42503
rect -15986 42537 -15934 42546
rect -15986 42503 -15977 42537
rect -15977 42503 -15943 42537
rect -15943 42503 -15934 42537
rect -15986 42494 -15934 42503
rect -15826 42537 -15774 42546
rect -15826 42503 -15817 42537
rect -15817 42503 -15783 42537
rect -15783 42503 -15774 42537
rect -15826 42494 -15774 42503
rect -15666 42537 -15614 42546
rect -15666 42503 -15657 42537
rect -15657 42503 -15623 42537
rect -15623 42503 -15614 42537
rect -15666 42494 -15614 42503
rect -15506 42537 -15454 42546
rect -15506 42503 -15497 42537
rect -15497 42503 -15463 42537
rect -15463 42503 -15454 42537
rect -15506 42494 -15454 42503
rect -15346 42537 -15294 42546
rect -15346 42503 -15337 42537
rect -15337 42503 -15303 42537
rect -15303 42503 -15294 42537
rect -15346 42494 -15294 42503
rect -15186 42537 -15134 42546
rect -15186 42503 -15177 42537
rect -15177 42503 -15143 42537
rect -15143 42503 -15134 42537
rect -15186 42494 -15134 42503
rect -15026 42537 -14974 42546
rect -15026 42503 -15017 42537
rect -15017 42503 -14983 42537
rect -14983 42503 -14974 42537
rect -15026 42494 -14974 42503
rect -14866 42537 -14814 42546
rect -14866 42503 -14857 42537
rect -14857 42503 -14823 42537
rect -14823 42503 -14814 42537
rect -14866 42494 -14814 42503
rect -14706 42537 -14654 42546
rect -14706 42503 -14697 42537
rect -14697 42503 -14663 42537
rect -14663 42503 -14654 42537
rect -14706 42494 -14654 42503
rect -14546 42537 -14494 42546
rect -14546 42503 -14537 42537
rect -14537 42503 -14503 42537
rect -14503 42503 -14494 42537
rect -14546 42494 -14494 42503
rect -14386 42537 -14334 42546
rect -14386 42503 -14377 42537
rect -14377 42503 -14343 42537
rect -14343 42503 -14334 42537
rect -14386 42494 -14334 42503
rect -14226 42537 -14174 42546
rect -14226 42503 -14217 42537
rect -14217 42503 -14183 42537
rect -14183 42503 -14174 42537
rect -14226 42494 -14174 42503
rect -14066 42537 -14014 42546
rect -14066 42503 -14057 42537
rect -14057 42503 -14023 42537
rect -14023 42503 -14014 42537
rect -14066 42494 -14014 42503
rect -13906 42537 -13854 42546
rect -13906 42503 -13897 42537
rect -13897 42503 -13863 42537
rect -13863 42503 -13854 42537
rect -13906 42494 -13854 42503
rect -13746 42537 -13694 42546
rect -13746 42503 -13737 42537
rect -13737 42503 -13703 42537
rect -13703 42503 -13694 42537
rect -13746 42494 -13694 42503
rect -13586 42537 -13534 42546
rect -13586 42503 -13577 42537
rect -13577 42503 -13543 42537
rect -13543 42503 -13534 42537
rect -13586 42494 -13534 42503
rect -13426 42537 -13374 42546
rect -13426 42503 -13417 42537
rect -13417 42503 -13383 42537
rect -13383 42503 -13374 42537
rect -13426 42494 -13374 42503
rect -13266 42537 -13214 42546
rect -13266 42503 -13257 42537
rect -13257 42503 -13223 42537
rect -13223 42503 -13214 42537
rect -13266 42494 -13214 42503
rect -13106 42537 -13054 42546
rect -13106 42503 -13097 42537
rect -13097 42503 -13063 42537
rect -13063 42503 -13054 42537
rect -13106 42494 -13054 42503
rect -12946 42537 -12894 42546
rect -12946 42503 -12937 42537
rect -12937 42503 -12903 42537
rect -12903 42503 -12894 42537
rect -12946 42494 -12894 42503
rect -12786 42537 -12734 42546
rect -12786 42503 -12777 42537
rect -12777 42503 -12743 42537
rect -12743 42503 -12734 42537
rect -12786 42494 -12734 42503
rect -12626 42537 -12574 42546
rect -12626 42503 -12617 42537
rect -12617 42503 -12583 42537
rect -12583 42503 -12574 42537
rect -12626 42494 -12574 42503
rect -12466 42537 -12414 42546
rect -12466 42503 -12457 42537
rect -12457 42503 -12423 42537
rect -12423 42503 -12414 42537
rect -12466 42494 -12414 42503
rect -12306 42537 -12254 42546
rect -12306 42503 -12297 42537
rect -12297 42503 -12263 42537
rect -12263 42503 -12254 42537
rect -12306 42494 -12254 42503
rect -11346 42537 -11294 42546
rect -11346 42503 -11337 42537
rect -11337 42503 -11303 42537
rect -11303 42503 -11294 42537
rect -11346 42494 -11294 42503
rect -11186 42537 -11134 42546
rect -11186 42503 -11177 42537
rect -11177 42503 -11143 42537
rect -11143 42503 -11134 42537
rect -11186 42494 -11134 42503
rect -11026 42537 -10974 42546
rect -11026 42503 -11017 42537
rect -11017 42503 -10983 42537
rect -10983 42503 -10974 42537
rect -11026 42494 -10974 42503
rect -10866 42537 -10814 42546
rect -10866 42503 -10857 42537
rect -10857 42503 -10823 42537
rect -10823 42503 -10814 42537
rect -10866 42494 -10814 42503
rect -10706 42537 -10654 42546
rect -10706 42503 -10697 42537
rect -10697 42503 -10663 42537
rect -10663 42503 -10654 42537
rect -10706 42494 -10654 42503
rect -10546 42537 -10494 42546
rect -10546 42503 -10537 42537
rect -10537 42503 -10503 42537
rect -10503 42503 -10494 42537
rect -10546 42494 -10494 42503
rect -10386 42537 -10334 42546
rect -10386 42503 -10377 42537
rect -10377 42503 -10343 42537
rect -10343 42503 -10334 42537
rect -10386 42494 -10334 42503
rect -10226 42537 -10174 42546
rect -10226 42503 -10217 42537
rect -10217 42503 -10183 42537
rect -10183 42503 -10174 42537
rect -10226 42494 -10174 42503
rect -10066 42537 -10014 42546
rect -10066 42503 -10057 42537
rect -10057 42503 -10023 42537
rect -10023 42503 -10014 42537
rect -10066 42494 -10014 42503
rect -9906 42537 -9854 42546
rect -9906 42503 -9897 42537
rect -9897 42503 -9863 42537
rect -9863 42503 -9854 42537
rect -9906 42494 -9854 42503
rect -9746 42537 -9694 42546
rect -9746 42503 -9737 42537
rect -9737 42503 -9703 42537
rect -9703 42503 -9694 42537
rect -9746 42494 -9694 42503
rect -9586 42537 -9534 42546
rect -9586 42503 -9577 42537
rect -9577 42503 -9543 42537
rect -9543 42503 -9534 42537
rect -9586 42494 -9534 42503
rect -9426 42537 -9374 42546
rect -9426 42503 -9417 42537
rect -9417 42503 -9383 42537
rect -9383 42503 -9374 42537
rect -9426 42494 -9374 42503
rect -9266 42537 -9214 42546
rect -9266 42503 -9257 42537
rect -9257 42503 -9223 42537
rect -9223 42503 -9214 42537
rect -9266 42494 -9214 42503
rect -9106 42537 -9054 42546
rect -9106 42503 -9097 42537
rect -9097 42503 -9063 42537
rect -9063 42503 -9054 42537
rect -9106 42494 -9054 42503
rect -8946 42537 -8894 42546
rect -8946 42503 -8937 42537
rect -8937 42503 -8903 42537
rect -8903 42503 -8894 42537
rect -8946 42494 -8894 42503
rect -8786 42537 -8734 42546
rect -8786 42503 -8777 42537
rect -8777 42503 -8743 42537
rect -8743 42503 -8734 42537
rect -8786 42494 -8734 42503
rect -8626 42537 -8574 42546
rect -8626 42503 -8617 42537
rect -8617 42503 -8583 42537
rect -8583 42503 -8574 42537
rect -8626 42494 -8574 42503
rect -8466 42537 -8414 42546
rect -8466 42503 -8457 42537
rect -8457 42503 -8423 42537
rect -8423 42503 -8414 42537
rect -8466 42494 -8414 42503
rect -8306 42537 -8254 42546
rect -8306 42503 -8297 42537
rect -8297 42503 -8263 42537
rect -8263 42503 -8254 42537
rect -8306 42494 -8254 42503
rect -8146 42537 -8094 42546
rect -8146 42503 -8137 42537
rect -8137 42503 -8103 42537
rect -8103 42503 -8094 42537
rect -8146 42494 -8094 42503
rect -7986 42537 -7934 42546
rect -7986 42503 -7977 42537
rect -7977 42503 -7943 42537
rect -7943 42503 -7934 42537
rect -7986 42494 -7934 42503
rect -7826 42537 -7774 42546
rect -7826 42503 -7817 42537
rect -7817 42503 -7783 42537
rect -7783 42503 -7774 42537
rect -7826 42494 -7774 42503
rect -7666 42537 -7614 42546
rect -7666 42503 -7657 42537
rect -7657 42503 -7623 42537
rect -7623 42503 -7614 42537
rect -7666 42494 -7614 42503
rect -7506 42537 -7454 42546
rect -7506 42503 -7497 42537
rect -7497 42503 -7463 42537
rect -7463 42503 -7454 42537
rect -7506 42494 -7454 42503
rect -7346 42537 -7294 42546
rect -7346 42503 -7337 42537
rect -7337 42503 -7303 42537
rect -7303 42503 -7294 42537
rect -7346 42494 -7294 42503
rect -7186 42537 -7134 42546
rect -7186 42503 -7177 42537
rect -7177 42503 -7143 42537
rect -7143 42503 -7134 42537
rect -7186 42494 -7134 42503
rect -7026 42537 -6974 42546
rect -7026 42503 -7017 42537
rect -7017 42503 -6983 42537
rect -6983 42503 -6974 42537
rect -7026 42494 -6974 42503
rect -6866 42537 -6814 42546
rect -6866 42503 -6857 42537
rect -6857 42503 -6823 42537
rect -6823 42503 -6814 42537
rect -6866 42494 -6814 42503
rect -6706 42537 -6654 42546
rect -6706 42503 -6697 42537
rect -6697 42503 -6663 42537
rect -6663 42503 -6654 42537
rect -6706 42494 -6654 42503
rect -6546 42537 -6494 42546
rect -6546 42503 -6537 42537
rect -6537 42503 -6503 42537
rect -6503 42503 -6494 42537
rect -6546 42494 -6494 42503
rect -6386 42537 -6334 42546
rect -6386 42503 -6377 42537
rect -6377 42503 -6343 42537
rect -6343 42503 -6334 42537
rect -6386 42494 -6334 42503
rect -6226 42537 -6174 42546
rect -6226 42503 -6217 42537
rect -6217 42503 -6183 42537
rect -6183 42503 -6174 42537
rect -6226 42494 -6174 42503
rect -6066 42537 -6014 42546
rect -6066 42503 -6057 42537
rect -6057 42503 -6023 42537
rect -6023 42503 -6014 42537
rect -6066 42494 -6014 42503
rect -5906 42537 -5854 42546
rect -5906 42503 -5897 42537
rect -5897 42503 -5863 42537
rect -5863 42503 -5854 42537
rect -5906 42494 -5854 42503
rect -5746 42537 -5694 42546
rect -5746 42503 -5737 42537
rect -5737 42503 -5703 42537
rect -5703 42503 -5694 42537
rect -5746 42494 -5694 42503
rect -5586 42537 -5534 42546
rect -5586 42503 -5577 42537
rect -5577 42503 -5543 42537
rect -5543 42503 -5534 42537
rect -5586 42494 -5534 42503
rect -5426 42537 -5374 42546
rect -5426 42503 -5417 42537
rect -5417 42503 -5383 42537
rect -5383 42503 -5374 42537
rect -5426 42494 -5374 42503
rect -5266 42537 -5214 42546
rect -5266 42503 -5257 42537
rect -5257 42503 -5223 42537
rect -5223 42503 -5214 42537
rect -5266 42494 -5214 42503
rect -5106 42537 -5054 42546
rect -5106 42503 -5097 42537
rect -5097 42503 -5063 42537
rect -5063 42503 -5054 42537
rect -5106 42494 -5054 42503
rect -4946 42537 -4894 42546
rect -4946 42503 -4937 42537
rect -4937 42503 -4903 42537
rect -4903 42503 -4894 42537
rect -4946 42494 -4894 42503
rect -4786 42537 -4734 42546
rect -4786 42503 -4777 42537
rect -4777 42503 -4743 42537
rect -4743 42503 -4734 42537
rect -4786 42494 -4734 42503
rect -4626 42537 -4574 42546
rect -4626 42503 -4617 42537
rect -4617 42503 -4583 42537
rect -4583 42503 -4574 42537
rect -4626 42494 -4574 42503
rect -4466 42537 -4414 42546
rect -4466 42503 -4457 42537
rect -4457 42503 -4423 42537
rect -4423 42503 -4414 42537
rect -4466 42494 -4414 42503
rect -4306 42537 -4254 42546
rect -4306 42503 -4297 42537
rect -4297 42503 -4263 42537
rect -4263 42503 -4254 42537
rect -4306 42494 -4254 42503
rect -4146 42537 -4094 42546
rect -4146 42503 -4137 42537
rect -4137 42503 -4103 42537
rect -4103 42503 -4094 42537
rect -4146 42494 -4094 42503
rect -3986 42537 -3934 42546
rect -3986 42503 -3977 42537
rect -3977 42503 -3943 42537
rect -3943 42503 -3934 42537
rect -3986 42494 -3934 42503
rect -3666 42537 -3614 42546
rect -3666 42503 -3657 42537
rect -3657 42503 -3623 42537
rect -3623 42503 -3614 42537
rect -3666 42494 -3614 42503
rect -3506 42537 -3454 42546
rect -3506 42503 -3497 42537
rect -3497 42503 -3463 42537
rect -3463 42503 -3454 42537
rect -3506 42494 -3454 42503
rect -3346 42537 -3294 42546
rect -3346 42503 -3337 42537
rect -3337 42503 -3303 42537
rect -3303 42503 -3294 42537
rect -3346 42494 -3294 42503
rect -3026 42537 -2974 42546
rect -3026 42503 -3017 42537
rect -3017 42503 -2983 42537
rect -2983 42503 -2974 42537
rect -3026 42494 -2974 42503
rect -2706 42537 -2654 42546
rect -2706 42503 -2697 42537
rect -2697 42503 -2663 42537
rect -2663 42503 -2654 42537
rect -2706 42494 -2654 42503
rect -2546 42537 -2494 42546
rect -2546 42503 -2537 42537
rect -2537 42503 -2503 42537
rect -2503 42503 -2494 42537
rect -2546 42494 -2494 42503
rect -2386 42537 -2334 42546
rect -2386 42503 -2377 42537
rect -2377 42503 -2343 42537
rect -2343 42503 -2334 42537
rect -2386 42494 -2334 42503
rect -2226 42537 -2174 42546
rect -2226 42503 -2217 42537
rect -2217 42503 -2183 42537
rect -2183 42503 -2174 42537
rect -2226 42494 -2174 42503
rect -2066 42537 -2014 42546
rect -2066 42503 -2057 42537
rect -2057 42503 -2023 42537
rect -2023 42503 -2014 42537
rect -2066 42494 -2014 42503
rect -1746 42537 -1694 42546
rect -1746 42503 -1737 42537
rect -1737 42503 -1703 42537
rect -1703 42503 -1694 42537
rect -1746 42494 -1694 42503
rect -1426 42537 -1374 42546
rect -1426 42503 -1417 42537
rect -1417 42503 -1383 42537
rect -1383 42503 -1374 42537
rect -1426 42494 -1374 42503
rect -1106 42537 -1054 42546
rect -1106 42503 -1097 42537
rect -1097 42503 -1063 42537
rect -1063 42503 -1054 42537
rect -1106 42494 -1054 42503
rect -29906 42217 -29854 42226
rect -29906 42183 -29897 42217
rect -29897 42183 -29863 42217
rect -29863 42183 -29854 42217
rect -29906 42174 -29854 42183
rect -29746 42217 -29694 42226
rect -29746 42183 -29737 42217
rect -29737 42183 -29703 42217
rect -29703 42183 -29694 42217
rect -29746 42174 -29694 42183
rect -29586 42217 -29534 42226
rect -29586 42183 -29577 42217
rect -29577 42183 -29543 42217
rect -29543 42183 -29534 42217
rect -29586 42174 -29534 42183
rect -29426 42217 -29374 42226
rect -29426 42183 -29417 42217
rect -29417 42183 -29383 42217
rect -29383 42183 -29374 42217
rect -29426 42174 -29374 42183
rect -29266 42217 -29214 42226
rect -29266 42183 -29257 42217
rect -29257 42183 -29223 42217
rect -29223 42183 -29214 42217
rect -29266 42174 -29214 42183
rect -29106 42217 -29054 42226
rect -29106 42183 -29097 42217
rect -29097 42183 -29063 42217
rect -29063 42183 -29054 42217
rect -29106 42174 -29054 42183
rect -28946 42217 -28894 42226
rect -28946 42183 -28937 42217
rect -28937 42183 -28903 42217
rect -28903 42183 -28894 42217
rect -28946 42174 -28894 42183
rect -28786 42217 -28734 42226
rect -28786 42183 -28777 42217
rect -28777 42183 -28743 42217
rect -28743 42183 -28734 42217
rect -28786 42174 -28734 42183
rect -28626 42217 -28574 42226
rect -28626 42183 -28617 42217
rect -28617 42183 -28583 42217
rect -28583 42183 -28574 42217
rect -28626 42174 -28574 42183
rect -28466 42217 -28414 42226
rect -28466 42183 -28457 42217
rect -28457 42183 -28423 42217
rect -28423 42183 -28414 42217
rect -28466 42174 -28414 42183
rect -28306 42217 -28254 42226
rect -28306 42183 -28297 42217
rect -28297 42183 -28263 42217
rect -28263 42183 -28254 42217
rect -28306 42174 -28254 42183
rect -28146 42217 -28094 42226
rect -28146 42183 -28137 42217
rect -28137 42183 -28103 42217
rect -28103 42183 -28094 42217
rect -28146 42174 -28094 42183
rect -27986 42217 -27934 42226
rect -27986 42183 -27977 42217
rect -27977 42183 -27943 42217
rect -27943 42183 -27934 42217
rect -27986 42174 -27934 42183
rect -27826 42217 -27774 42226
rect -27826 42183 -27817 42217
rect -27817 42183 -27783 42217
rect -27783 42183 -27774 42217
rect -27826 42174 -27774 42183
rect -27666 42217 -27614 42226
rect -27666 42183 -27657 42217
rect -27657 42183 -27623 42217
rect -27623 42183 -27614 42217
rect -27666 42174 -27614 42183
rect -27506 42217 -27454 42226
rect -27506 42183 -27497 42217
rect -27497 42183 -27463 42217
rect -27463 42183 -27454 42217
rect -27506 42174 -27454 42183
rect -27346 42217 -27294 42226
rect -27346 42183 -27337 42217
rect -27337 42183 -27303 42217
rect -27303 42183 -27294 42217
rect -27346 42174 -27294 42183
rect -27186 42217 -27134 42226
rect -27186 42183 -27177 42217
rect -27177 42183 -27143 42217
rect -27143 42183 -27134 42217
rect -27186 42174 -27134 42183
rect -27026 42217 -26974 42226
rect -27026 42183 -27017 42217
rect -27017 42183 -26983 42217
rect -26983 42183 -26974 42217
rect -27026 42174 -26974 42183
rect -26866 42217 -26814 42226
rect -26866 42183 -26857 42217
rect -26857 42183 -26823 42217
rect -26823 42183 -26814 42217
rect -26866 42174 -26814 42183
rect -26706 42217 -26654 42226
rect -26706 42183 -26697 42217
rect -26697 42183 -26663 42217
rect -26663 42183 -26654 42217
rect -26706 42174 -26654 42183
rect -26546 42217 -26494 42226
rect -26546 42183 -26537 42217
rect -26537 42183 -26503 42217
rect -26503 42183 -26494 42217
rect -26546 42174 -26494 42183
rect -26386 42217 -26334 42226
rect -26386 42183 -26377 42217
rect -26377 42183 -26343 42217
rect -26343 42183 -26334 42217
rect -26386 42174 -26334 42183
rect -26226 42217 -26174 42226
rect -26226 42183 -26217 42217
rect -26217 42183 -26183 42217
rect -26183 42183 -26174 42217
rect -26226 42174 -26174 42183
rect -26066 42217 -26014 42226
rect -26066 42183 -26057 42217
rect -26057 42183 -26023 42217
rect -26023 42183 -26014 42217
rect -26066 42174 -26014 42183
rect -25906 42217 -25854 42226
rect -25906 42183 -25897 42217
rect -25897 42183 -25863 42217
rect -25863 42183 -25854 42217
rect -25906 42174 -25854 42183
rect -25746 42217 -25694 42226
rect -25746 42183 -25737 42217
rect -25737 42183 -25703 42217
rect -25703 42183 -25694 42217
rect -25746 42174 -25694 42183
rect -25586 42217 -25534 42226
rect -25586 42183 -25577 42217
rect -25577 42183 -25543 42217
rect -25543 42183 -25534 42217
rect -25586 42174 -25534 42183
rect -25426 42217 -25374 42226
rect -25426 42183 -25417 42217
rect -25417 42183 -25383 42217
rect -25383 42183 -25374 42217
rect -25426 42174 -25374 42183
rect -25266 42217 -25214 42226
rect -25266 42183 -25257 42217
rect -25257 42183 -25223 42217
rect -25223 42183 -25214 42217
rect -25266 42174 -25214 42183
rect -25106 42217 -25054 42226
rect -25106 42183 -25097 42217
rect -25097 42183 -25063 42217
rect -25063 42183 -25054 42217
rect -25106 42174 -25054 42183
rect -24946 42217 -24894 42226
rect -24946 42183 -24937 42217
rect -24937 42183 -24903 42217
rect -24903 42183 -24894 42217
rect -24946 42174 -24894 42183
rect -24786 42217 -24734 42226
rect -24786 42183 -24777 42217
rect -24777 42183 -24743 42217
rect -24743 42183 -24734 42217
rect -24786 42174 -24734 42183
rect -24626 42217 -24574 42226
rect -24626 42183 -24617 42217
rect -24617 42183 -24583 42217
rect -24583 42183 -24574 42217
rect -24626 42174 -24574 42183
rect -24466 42217 -24414 42226
rect -24466 42183 -24457 42217
rect -24457 42183 -24423 42217
rect -24423 42183 -24414 42217
rect -24466 42174 -24414 42183
rect -24306 42217 -24254 42226
rect -24306 42183 -24297 42217
rect -24297 42183 -24263 42217
rect -24263 42183 -24254 42217
rect -24306 42174 -24254 42183
rect -24146 42217 -24094 42226
rect -24146 42183 -24137 42217
rect -24137 42183 -24103 42217
rect -24103 42183 -24094 42217
rect -24146 42174 -24094 42183
rect -23986 42217 -23934 42226
rect -23986 42183 -23977 42217
rect -23977 42183 -23943 42217
rect -23943 42183 -23934 42217
rect -23986 42174 -23934 42183
rect -23826 42217 -23774 42226
rect -23826 42183 -23817 42217
rect -23817 42183 -23783 42217
rect -23783 42183 -23774 42217
rect -23826 42174 -23774 42183
rect -23666 42217 -23614 42226
rect -23666 42183 -23657 42217
rect -23657 42183 -23623 42217
rect -23623 42183 -23614 42217
rect -23666 42174 -23614 42183
rect -23506 42217 -23454 42226
rect -23506 42183 -23497 42217
rect -23497 42183 -23463 42217
rect -23463 42183 -23454 42217
rect -23506 42174 -23454 42183
rect -23346 42217 -23294 42226
rect -23346 42183 -23337 42217
rect -23337 42183 -23303 42217
rect -23303 42183 -23294 42217
rect -23346 42174 -23294 42183
rect -23186 42217 -23134 42226
rect -23186 42183 -23177 42217
rect -23177 42183 -23143 42217
rect -23143 42183 -23134 42217
rect -23186 42174 -23134 42183
rect -23026 42217 -22974 42226
rect -23026 42183 -23017 42217
rect -23017 42183 -22983 42217
rect -22983 42183 -22974 42217
rect -23026 42174 -22974 42183
rect -22866 42217 -22814 42226
rect -22866 42183 -22857 42217
rect -22857 42183 -22823 42217
rect -22823 42183 -22814 42217
rect -22866 42174 -22814 42183
rect -22706 42217 -22654 42226
rect -22706 42183 -22697 42217
rect -22697 42183 -22663 42217
rect -22663 42183 -22654 42217
rect -22706 42174 -22654 42183
rect -22546 42217 -22494 42226
rect -22546 42183 -22537 42217
rect -22537 42183 -22503 42217
rect -22503 42183 -22494 42217
rect -22546 42174 -22494 42183
rect -22386 42217 -22334 42226
rect -22386 42183 -22377 42217
rect -22377 42183 -22343 42217
rect -22343 42183 -22334 42217
rect -22386 42174 -22334 42183
rect -22226 42217 -22174 42226
rect -22226 42183 -22217 42217
rect -22217 42183 -22183 42217
rect -22183 42183 -22174 42217
rect -22226 42174 -22174 42183
rect -22066 42217 -22014 42226
rect -22066 42183 -22057 42217
rect -22057 42183 -22023 42217
rect -22023 42183 -22014 42217
rect -22066 42174 -22014 42183
rect -21906 42217 -21854 42226
rect -21906 42183 -21897 42217
rect -21897 42183 -21863 42217
rect -21863 42183 -21854 42217
rect -21906 42174 -21854 42183
rect -21746 42217 -21694 42226
rect -21746 42183 -21737 42217
rect -21737 42183 -21703 42217
rect -21703 42183 -21694 42217
rect -21746 42174 -21694 42183
rect -21586 42217 -21534 42226
rect -21586 42183 -21577 42217
rect -21577 42183 -21543 42217
rect -21543 42183 -21534 42217
rect -21586 42174 -21534 42183
rect -21426 42217 -21374 42226
rect -21426 42183 -21417 42217
rect -21417 42183 -21383 42217
rect -21383 42183 -21374 42217
rect -21426 42174 -21374 42183
rect -21266 42217 -21214 42226
rect -21266 42183 -21257 42217
rect -21257 42183 -21223 42217
rect -21223 42183 -21214 42217
rect -21266 42174 -21214 42183
rect -21106 42217 -21054 42226
rect -21106 42183 -21097 42217
rect -21097 42183 -21063 42217
rect -21063 42183 -21054 42217
rect -21106 42174 -21054 42183
rect -20946 42217 -20894 42226
rect -20946 42183 -20937 42217
rect -20937 42183 -20903 42217
rect -20903 42183 -20894 42217
rect -20946 42174 -20894 42183
rect -20786 42217 -20734 42226
rect -20786 42183 -20777 42217
rect -20777 42183 -20743 42217
rect -20743 42183 -20734 42217
rect -20786 42174 -20734 42183
rect -20626 42217 -20574 42226
rect -20626 42183 -20617 42217
rect -20617 42183 -20583 42217
rect -20583 42183 -20574 42217
rect -20626 42174 -20574 42183
rect -20466 42217 -20414 42226
rect -20466 42183 -20457 42217
rect -20457 42183 -20423 42217
rect -20423 42183 -20414 42217
rect -20466 42174 -20414 42183
rect -20306 42217 -20254 42226
rect -20306 42183 -20297 42217
rect -20297 42183 -20263 42217
rect -20263 42183 -20254 42217
rect -20306 42174 -20254 42183
rect -20146 42217 -20094 42226
rect -20146 42183 -20137 42217
rect -20137 42183 -20103 42217
rect -20103 42183 -20094 42217
rect -20146 42174 -20094 42183
rect -19986 42217 -19934 42226
rect -19986 42183 -19977 42217
rect -19977 42183 -19943 42217
rect -19943 42183 -19934 42217
rect -19986 42174 -19934 42183
rect -19826 42217 -19774 42226
rect -19826 42183 -19817 42217
rect -19817 42183 -19783 42217
rect -19783 42183 -19774 42217
rect -19826 42174 -19774 42183
rect -19666 42217 -19614 42226
rect -19666 42183 -19657 42217
rect -19657 42183 -19623 42217
rect -19623 42183 -19614 42217
rect -19666 42174 -19614 42183
rect -19506 42217 -19454 42226
rect -19506 42183 -19497 42217
rect -19497 42183 -19463 42217
rect -19463 42183 -19454 42217
rect -19506 42174 -19454 42183
rect -19346 42217 -19294 42226
rect -19346 42183 -19337 42217
rect -19337 42183 -19303 42217
rect -19303 42183 -19294 42217
rect -19346 42174 -19294 42183
rect -19186 42217 -19134 42226
rect -19186 42183 -19177 42217
rect -19177 42183 -19143 42217
rect -19143 42183 -19134 42217
rect -19186 42174 -19134 42183
rect -19026 42217 -18974 42226
rect -19026 42183 -19017 42217
rect -19017 42183 -18983 42217
rect -18983 42183 -18974 42217
rect -19026 42174 -18974 42183
rect -18866 42217 -18814 42226
rect -18866 42183 -18857 42217
rect -18857 42183 -18823 42217
rect -18823 42183 -18814 42217
rect -18866 42174 -18814 42183
rect -18706 42217 -18654 42226
rect -18706 42183 -18697 42217
rect -18697 42183 -18663 42217
rect -18663 42183 -18654 42217
rect -18706 42174 -18654 42183
rect -18546 42217 -18494 42226
rect -18546 42183 -18537 42217
rect -18537 42183 -18503 42217
rect -18503 42183 -18494 42217
rect -18546 42174 -18494 42183
rect -18386 42217 -18334 42226
rect -18386 42183 -18377 42217
rect -18377 42183 -18343 42217
rect -18343 42183 -18334 42217
rect -18386 42174 -18334 42183
rect -18226 42217 -18174 42226
rect -18226 42183 -18217 42217
rect -18217 42183 -18183 42217
rect -18183 42183 -18174 42217
rect -18226 42174 -18174 42183
rect -18066 42217 -18014 42226
rect -18066 42183 -18057 42217
rect -18057 42183 -18023 42217
rect -18023 42183 -18014 42217
rect -18066 42174 -18014 42183
rect -17906 42217 -17854 42226
rect -17906 42183 -17897 42217
rect -17897 42183 -17863 42217
rect -17863 42183 -17854 42217
rect -17906 42174 -17854 42183
rect -17746 42217 -17694 42226
rect -17746 42183 -17737 42217
rect -17737 42183 -17703 42217
rect -17703 42183 -17694 42217
rect -17746 42174 -17694 42183
rect -17586 42217 -17534 42226
rect -17586 42183 -17577 42217
rect -17577 42183 -17543 42217
rect -17543 42183 -17534 42217
rect -17586 42174 -17534 42183
rect -17426 42217 -17374 42226
rect -17426 42183 -17417 42217
rect -17417 42183 -17383 42217
rect -17383 42183 -17374 42217
rect -17426 42174 -17374 42183
rect -17266 42217 -17214 42226
rect -17266 42183 -17257 42217
rect -17257 42183 -17223 42217
rect -17223 42183 -17214 42217
rect -17266 42174 -17214 42183
rect -17106 42217 -17054 42226
rect -17106 42183 -17097 42217
rect -17097 42183 -17063 42217
rect -17063 42183 -17054 42217
rect -17106 42174 -17054 42183
rect -16946 42217 -16894 42226
rect -16946 42183 -16937 42217
rect -16937 42183 -16903 42217
rect -16903 42183 -16894 42217
rect -16946 42174 -16894 42183
rect -16786 42217 -16734 42226
rect -16786 42183 -16777 42217
rect -16777 42183 -16743 42217
rect -16743 42183 -16734 42217
rect -16786 42174 -16734 42183
rect -16626 42217 -16574 42226
rect -16626 42183 -16617 42217
rect -16617 42183 -16583 42217
rect -16583 42183 -16574 42217
rect -16626 42174 -16574 42183
rect -16466 42217 -16414 42226
rect -16466 42183 -16457 42217
rect -16457 42183 -16423 42217
rect -16423 42183 -16414 42217
rect -16466 42174 -16414 42183
rect -16306 42217 -16254 42226
rect -16306 42183 -16297 42217
rect -16297 42183 -16263 42217
rect -16263 42183 -16254 42217
rect -16306 42174 -16254 42183
rect -16146 42217 -16094 42226
rect -16146 42183 -16137 42217
rect -16137 42183 -16103 42217
rect -16103 42183 -16094 42217
rect -16146 42174 -16094 42183
rect -15986 42217 -15934 42226
rect -15986 42183 -15977 42217
rect -15977 42183 -15943 42217
rect -15943 42183 -15934 42217
rect -15986 42174 -15934 42183
rect -15826 42217 -15774 42226
rect -15826 42183 -15817 42217
rect -15817 42183 -15783 42217
rect -15783 42183 -15774 42217
rect -15826 42174 -15774 42183
rect -15666 42217 -15614 42226
rect -15666 42183 -15657 42217
rect -15657 42183 -15623 42217
rect -15623 42183 -15614 42217
rect -15666 42174 -15614 42183
rect -15506 42217 -15454 42226
rect -15506 42183 -15497 42217
rect -15497 42183 -15463 42217
rect -15463 42183 -15454 42217
rect -15506 42174 -15454 42183
rect -15346 42217 -15294 42226
rect -15346 42183 -15337 42217
rect -15337 42183 -15303 42217
rect -15303 42183 -15294 42217
rect -15346 42174 -15294 42183
rect -15186 42217 -15134 42226
rect -15186 42183 -15177 42217
rect -15177 42183 -15143 42217
rect -15143 42183 -15134 42217
rect -15186 42174 -15134 42183
rect -15026 42217 -14974 42226
rect -15026 42183 -15017 42217
rect -15017 42183 -14983 42217
rect -14983 42183 -14974 42217
rect -15026 42174 -14974 42183
rect -14866 42217 -14814 42226
rect -14866 42183 -14857 42217
rect -14857 42183 -14823 42217
rect -14823 42183 -14814 42217
rect -14866 42174 -14814 42183
rect -14706 42217 -14654 42226
rect -14706 42183 -14697 42217
rect -14697 42183 -14663 42217
rect -14663 42183 -14654 42217
rect -14706 42174 -14654 42183
rect -14546 42217 -14494 42226
rect -14546 42183 -14537 42217
rect -14537 42183 -14503 42217
rect -14503 42183 -14494 42217
rect -14546 42174 -14494 42183
rect -14386 42217 -14334 42226
rect -14386 42183 -14377 42217
rect -14377 42183 -14343 42217
rect -14343 42183 -14334 42217
rect -14386 42174 -14334 42183
rect -14226 42217 -14174 42226
rect -14226 42183 -14217 42217
rect -14217 42183 -14183 42217
rect -14183 42183 -14174 42217
rect -14226 42174 -14174 42183
rect -14066 42217 -14014 42226
rect -14066 42183 -14057 42217
rect -14057 42183 -14023 42217
rect -14023 42183 -14014 42217
rect -14066 42174 -14014 42183
rect -13906 42217 -13854 42226
rect -13906 42183 -13897 42217
rect -13897 42183 -13863 42217
rect -13863 42183 -13854 42217
rect -13906 42174 -13854 42183
rect -13746 42217 -13694 42226
rect -13746 42183 -13737 42217
rect -13737 42183 -13703 42217
rect -13703 42183 -13694 42217
rect -13746 42174 -13694 42183
rect -13586 42217 -13534 42226
rect -13586 42183 -13577 42217
rect -13577 42183 -13543 42217
rect -13543 42183 -13534 42217
rect -13586 42174 -13534 42183
rect -13426 42217 -13374 42226
rect -13426 42183 -13417 42217
rect -13417 42183 -13383 42217
rect -13383 42183 -13374 42217
rect -13426 42174 -13374 42183
rect -13266 42217 -13214 42226
rect -13266 42183 -13257 42217
rect -13257 42183 -13223 42217
rect -13223 42183 -13214 42217
rect -13266 42174 -13214 42183
rect -13106 42217 -13054 42226
rect -13106 42183 -13097 42217
rect -13097 42183 -13063 42217
rect -13063 42183 -13054 42217
rect -13106 42174 -13054 42183
rect -12946 42217 -12894 42226
rect -12946 42183 -12937 42217
rect -12937 42183 -12903 42217
rect -12903 42183 -12894 42217
rect -12946 42174 -12894 42183
rect -12786 42217 -12734 42226
rect -12786 42183 -12777 42217
rect -12777 42183 -12743 42217
rect -12743 42183 -12734 42217
rect -12786 42174 -12734 42183
rect -12626 42217 -12574 42226
rect -12626 42183 -12617 42217
rect -12617 42183 -12583 42217
rect -12583 42183 -12574 42217
rect -12626 42174 -12574 42183
rect -12466 42217 -12414 42226
rect -12466 42183 -12457 42217
rect -12457 42183 -12423 42217
rect -12423 42183 -12414 42217
rect -12466 42174 -12414 42183
rect -12306 42217 -12254 42226
rect -12306 42183 -12297 42217
rect -12297 42183 -12263 42217
rect -12263 42183 -12254 42217
rect -12306 42174 -12254 42183
rect -11346 42217 -11294 42226
rect -11346 42183 -11337 42217
rect -11337 42183 -11303 42217
rect -11303 42183 -11294 42217
rect -11346 42174 -11294 42183
rect -11186 42217 -11134 42226
rect -11186 42183 -11177 42217
rect -11177 42183 -11143 42217
rect -11143 42183 -11134 42217
rect -11186 42174 -11134 42183
rect -11026 42217 -10974 42226
rect -11026 42183 -11017 42217
rect -11017 42183 -10983 42217
rect -10983 42183 -10974 42217
rect -11026 42174 -10974 42183
rect -10866 42217 -10814 42226
rect -10866 42183 -10857 42217
rect -10857 42183 -10823 42217
rect -10823 42183 -10814 42217
rect -10866 42174 -10814 42183
rect -10706 42217 -10654 42226
rect -10706 42183 -10697 42217
rect -10697 42183 -10663 42217
rect -10663 42183 -10654 42217
rect -10706 42174 -10654 42183
rect -10546 42217 -10494 42226
rect -10546 42183 -10537 42217
rect -10537 42183 -10503 42217
rect -10503 42183 -10494 42217
rect -10546 42174 -10494 42183
rect -10386 42217 -10334 42226
rect -10386 42183 -10377 42217
rect -10377 42183 -10343 42217
rect -10343 42183 -10334 42217
rect -10386 42174 -10334 42183
rect -10226 42217 -10174 42226
rect -10226 42183 -10217 42217
rect -10217 42183 -10183 42217
rect -10183 42183 -10174 42217
rect -10226 42174 -10174 42183
rect -10066 42217 -10014 42226
rect -10066 42183 -10057 42217
rect -10057 42183 -10023 42217
rect -10023 42183 -10014 42217
rect -10066 42174 -10014 42183
rect -9906 42217 -9854 42226
rect -9906 42183 -9897 42217
rect -9897 42183 -9863 42217
rect -9863 42183 -9854 42217
rect -9906 42174 -9854 42183
rect -9746 42217 -9694 42226
rect -9746 42183 -9737 42217
rect -9737 42183 -9703 42217
rect -9703 42183 -9694 42217
rect -9746 42174 -9694 42183
rect -9586 42217 -9534 42226
rect -9586 42183 -9577 42217
rect -9577 42183 -9543 42217
rect -9543 42183 -9534 42217
rect -9586 42174 -9534 42183
rect -9426 42217 -9374 42226
rect -9426 42183 -9417 42217
rect -9417 42183 -9383 42217
rect -9383 42183 -9374 42217
rect -9426 42174 -9374 42183
rect -9266 42217 -9214 42226
rect -9266 42183 -9257 42217
rect -9257 42183 -9223 42217
rect -9223 42183 -9214 42217
rect -9266 42174 -9214 42183
rect -9106 42217 -9054 42226
rect -9106 42183 -9097 42217
rect -9097 42183 -9063 42217
rect -9063 42183 -9054 42217
rect -9106 42174 -9054 42183
rect -8946 42217 -8894 42226
rect -8946 42183 -8937 42217
rect -8937 42183 -8903 42217
rect -8903 42183 -8894 42217
rect -8946 42174 -8894 42183
rect -8786 42217 -8734 42226
rect -8786 42183 -8777 42217
rect -8777 42183 -8743 42217
rect -8743 42183 -8734 42217
rect -8786 42174 -8734 42183
rect -8626 42217 -8574 42226
rect -8626 42183 -8617 42217
rect -8617 42183 -8583 42217
rect -8583 42183 -8574 42217
rect -8626 42174 -8574 42183
rect -8466 42217 -8414 42226
rect -8466 42183 -8457 42217
rect -8457 42183 -8423 42217
rect -8423 42183 -8414 42217
rect -8466 42174 -8414 42183
rect -8306 42217 -8254 42226
rect -8306 42183 -8297 42217
rect -8297 42183 -8263 42217
rect -8263 42183 -8254 42217
rect -8306 42174 -8254 42183
rect -8146 42217 -8094 42226
rect -8146 42183 -8137 42217
rect -8137 42183 -8103 42217
rect -8103 42183 -8094 42217
rect -8146 42174 -8094 42183
rect -7986 42217 -7934 42226
rect -7986 42183 -7977 42217
rect -7977 42183 -7943 42217
rect -7943 42183 -7934 42217
rect -7986 42174 -7934 42183
rect -7826 42217 -7774 42226
rect -7826 42183 -7817 42217
rect -7817 42183 -7783 42217
rect -7783 42183 -7774 42217
rect -7826 42174 -7774 42183
rect -7666 42217 -7614 42226
rect -7666 42183 -7657 42217
rect -7657 42183 -7623 42217
rect -7623 42183 -7614 42217
rect -7666 42174 -7614 42183
rect -7506 42217 -7454 42226
rect -7506 42183 -7497 42217
rect -7497 42183 -7463 42217
rect -7463 42183 -7454 42217
rect -7506 42174 -7454 42183
rect -7346 42217 -7294 42226
rect -7346 42183 -7337 42217
rect -7337 42183 -7303 42217
rect -7303 42183 -7294 42217
rect -7346 42174 -7294 42183
rect -7186 42217 -7134 42226
rect -7186 42183 -7177 42217
rect -7177 42183 -7143 42217
rect -7143 42183 -7134 42217
rect -7186 42174 -7134 42183
rect -7026 42217 -6974 42226
rect -7026 42183 -7017 42217
rect -7017 42183 -6983 42217
rect -6983 42183 -6974 42217
rect -7026 42174 -6974 42183
rect -6866 42217 -6814 42226
rect -6866 42183 -6857 42217
rect -6857 42183 -6823 42217
rect -6823 42183 -6814 42217
rect -6866 42174 -6814 42183
rect -6706 42217 -6654 42226
rect -6706 42183 -6697 42217
rect -6697 42183 -6663 42217
rect -6663 42183 -6654 42217
rect -6706 42174 -6654 42183
rect -6546 42217 -6494 42226
rect -6546 42183 -6537 42217
rect -6537 42183 -6503 42217
rect -6503 42183 -6494 42217
rect -6546 42174 -6494 42183
rect -6386 42217 -6334 42226
rect -6386 42183 -6377 42217
rect -6377 42183 -6343 42217
rect -6343 42183 -6334 42217
rect -6386 42174 -6334 42183
rect -6226 42217 -6174 42226
rect -6226 42183 -6217 42217
rect -6217 42183 -6183 42217
rect -6183 42183 -6174 42217
rect -6226 42174 -6174 42183
rect -6066 42217 -6014 42226
rect -6066 42183 -6057 42217
rect -6057 42183 -6023 42217
rect -6023 42183 -6014 42217
rect -6066 42174 -6014 42183
rect -5906 42217 -5854 42226
rect -5906 42183 -5897 42217
rect -5897 42183 -5863 42217
rect -5863 42183 -5854 42217
rect -5906 42174 -5854 42183
rect -5746 42217 -5694 42226
rect -5746 42183 -5737 42217
rect -5737 42183 -5703 42217
rect -5703 42183 -5694 42217
rect -5746 42174 -5694 42183
rect -5586 42217 -5534 42226
rect -5586 42183 -5577 42217
rect -5577 42183 -5543 42217
rect -5543 42183 -5534 42217
rect -5586 42174 -5534 42183
rect -5426 42217 -5374 42226
rect -5426 42183 -5417 42217
rect -5417 42183 -5383 42217
rect -5383 42183 -5374 42217
rect -5426 42174 -5374 42183
rect -5266 42217 -5214 42226
rect -5266 42183 -5257 42217
rect -5257 42183 -5223 42217
rect -5223 42183 -5214 42217
rect -5266 42174 -5214 42183
rect -5106 42217 -5054 42226
rect -5106 42183 -5097 42217
rect -5097 42183 -5063 42217
rect -5063 42183 -5054 42217
rect -5106 42174 -5054 42183
rect -4946 42217 -4894 42226
rect -4946 42183 -4937 42217
rect -4937 42183 -4903 42217
rect -4903 42183 -4894 42217
rect -4946 42174 -4894 42183
rect -4786 42217 -4734 42226
rect -4786 42183 -4777 42217
rect -4777 42183 -4743 42217
rect -4743 42183 -4734 42217
rect -4786 42174 -4734 42183
rect -4626 42217 -4574 42226
rect -4626 42183 -4617 42217
rect -4617 42183 -4583 42217
rect -4583 42183 -4574 42217
rect -4626 42174 -4574 42183
rect -4466 42217 -4414 42226
rect -4466 42183 -4457 42217
rect -4457 42183 -4423 42217
rect -4423 42183 -4414 42217
rect -4466 42174 -4414 42183
rect -4306 42217 -4254 42226
rect -4306 42183 -4297 42217
rect -4297 42183 -4263 42217
rect -4263 42183 -4254 42217
rect -4306 42174 -4254 42183
rect -4146 42217 -4094 42226
rect -4146 42183 -4137 42217
rect -4137 42183 -4103 42217
rect -4103 42183 -4094 42217
rect -4146 42174 -4094 42183
rect -3986 42217 -3934 42226
rect -3986 42183 -3977 42217
rect -3977 42183 -3943 42217
rect -3943 42183 -3934 42217
rect -3986 42174 -3934 42183
rect -3666 42217 -3614 42226
rect -3666 42183 -3657 42217
rect -3657 42183 -3623 42217
rect -3623 42183 -3614 42217
rect -3666 42174 -3614 42183
rect -3506 42217 -3454 42226
rect -3506 42183 -3497 42217
rect -3497 42183 -3463 42217
rect -3463 42183 -3454 42217
rect -3506 42174 -3454 42183
rect -3346 42217 -3294 42226
rect -3346 42183 -3337 42217
rect -3337 42183 -3303 42217
rect -3303 42183 -3294 42217
rect -3346 42174 -3294 42183
rect -3026 42217 -2974 42226
rect -3026 42183 -3017 42217
rect -3017 42183 -2983 42217
rect -2983 42183 -2974 42217
rect -3026 42174 -2974 42183
rect -2706 42217 -2654 42226
rect -2706 42183 -2697 42217
rect -2697 42183 -2663 42217
rect -2663 42183 -2654 42217
rect -2706 42174 -2654 42183
rect -2546 42217 -2494 42226
rect -2546 42183 -2537 42217
rect -2537 42183 -2503 42217
rect -2503 42183 -2494 42217
rect -2546 42174 -2494 42183
rect -2386 42217 -2334 42226
rect -2386 42183 -2377 42217
rect -2377 42183 -2343 42217
rect -2343 42183 -2334 42217
rect -2386 42174 -2334 42183
rect -2226 42217 -2174 42226
rect -2226 42183 -2217 42217
rect -2217 42183 -2183 42217
rect -2183 42183 -2174 42217
rect -2226 42174 -2174 42183
rect -2066 42217 -2014 42226
rect -2066 42183 -2057 42217
rect -2057 42183 -2023 42217
rect -2023 42183 -2014 42217
rect -2066 42174 -2014 42183
rect -1746 42217 -1694 42226
rect -1746 42183 -1737 42217
rect -1737 42183 -1703 42217
rect -1703 42183 -1694 42217
rect -1746 42174 -1694 42183
rect -1426 42217 -1374 42226
rect -1426 42183 -1417 42217
rect -1417 42183 -1383 42217
rect -1383 42183 -1374 42217
rect -1426 42174 -1374 42183
rect -1106 42217 -1054 42226
rect -1106 42183 -1097 42217
rect -1097 42183 -1063 42217
rect -1063 42183 -1054 42217
rect -1106 42174 -1054 42183
rect -29906 41897 -29854 41906
rect -29906 41863 -29897 41897
rect -29897 41863 -29863 41897
rect -29863 41863 -29854 41897
rect -29906 41854 -29854 41863
rect -29746 41897 -29694 41906
rect -29746 41863 -29737 41897
rect -29737 41863 -29703 41897
rect -29703 41863 -29694 41897
rect -29746 41854 -29694 41863
rect -29586 41897 -29534 41906
rect -29586 41863 -29577 41897
rect -29577 41863 -29543 41897
rect -29543 41863 -29534 41897
rect -29586 41854 -29534 41863
rect -29426 41897 -29374 41906
rect -29426 41863 -29417 41897
rect -29417 41863 -29383 41897
rect -29383 41863 -29374 41897
rect -29426 41854 -29374 41863
rect -29266 41897 -29214 41906
rect -29266 41863 -29257 41897
rect -29257 41863 -29223 41897
rect -29223 41863 -29214 41897
rect -29266 41854 -29214 41863
rect -29106 41897 -29054 41906
rect -29106 41863 -29097 41897
rect -29097 41863 -29063 41897
rect -29063 41863 -29054 41897
rect -29106 41854 -29054 41863
rect -28946 41897 -28894 41906
rect -28946 41863 -28937 41897
rect -28937 41863 -28903 41897
rect -28903 41863 -28894 41897
rect -28946 41854 -28894 41863
rect -28786 41897 -28734 41906
rect -28786 41863 -28777 41897
rect -28777 41863 -28743 41897
rect -28743 41863 -28734 41897
rect -28786 41854 -28734 41863
rect -28626 41897 -28574 41906
rect -28626 41863 -28617 41897
rect -28617 41863 -28583 41897
rect -28583 41863 -28574 41897
rect -28626 41854 -28574 41863
rect -28466 41897 -28414 41906
rect -28466 41863 -28457 41897
rect -28457 41863 -28423 41897
rect -28423 41863 -28414 41897
rect -28466 41854 -28414 41863
rect -28306 41897 -28254 41906
rect -28306 41863 -28297 41897
rect -28297 41863 -28263 41897
rect -28263 41863 -28254 41897
rect -28306 41854 -28254 41863
rect -28146 41897 -28094 41906
rect -28146 41863 -28137 41897
rect -28137 41863 -28103 41897
rect -28103 41863 -28094 41897
rect -28146 41854 -28094 41863
rect -27986 41897 -27934 41906
rect -27986 41863 -27977 41897
rect -27977 41863 -27943 41897
rect -27943 41863 -27934 41897
rect -27986 41854 -27934 41863
rect -27826 41897 -27774 41906
rect -27826 41863 -27817 41897
rect -27817 41863 -27783 41897
rect -27783 41863 -27774 41897
rect -27826 41854 -27774 41863
rect -27666 41897 -27614 41906
rect -27666 41863 -27657 41897
rect -27657 41863 -27623 41897
rect -27623 41863 -27614 41897
rect -27666 41854 -27614 41863
rect -27506 41897 -27454 41906
rect -27506 41863 -27497 41897
rect -27497 41863 -27463 41897
rect -27463 41863 -27454 41897
rect -27506 41854 -27454 41863
rect -27346 41897 -27294 41906
rect -27346 41863 -27337 41897
rect -27337 41863 -27303 41897
rect -27303 41863 -27294 41897
rect -27346 41854 -27294 41863
rect -27186 41897 -27134 41906
rect -27186 41863 -27177 41897
rect -27177 41863 -27143 41897
rect -27143 41863 -27134 41897
rect -27186 41854 -27134 41863
rect -27026 41897 -26974 41906
rect -27026 41863 -27017 41897
rect -27017 41863 -26983 41897
rect -26983 41863 -26974 41897
rect -27026 41854 -26974 41863
rect -26866 41897 -26814 41906
rect -26866 41863 -26857 41897
rect -26857 41863 -26823 41897
rect -26823 41863 -26814 41897
rect -26866 41854 -26814 41863
rect -26706 41897 -26654 41906
rect -26706 41863 -26697 41897
rect -26697 41863 -26663 41897
rect -26663 41863 -26654 41897
rect -26706 41854 -26654 41863
rect -26546 41897 -26494 41906
rect -26546 41863 -26537 41897
rect -26537 41863 -26503 41897
rect -26503 41863 -26494 41897
rect -26546 41854 -26494 41863
rect -26386 41897 -26334 41906
rect -26386 41863 -26377 41897
rect -26377 41863 -26343 41897
rect -26343 41863 -26334 41897
rect -26386 41854 -26334 41863
rect -26226 41897 -26174 41906
rect -26226 41863 -26217 41897
rect -26217 41863 -26183 41897
rect -26183 41863 -26174 41897
rect -26226 41854 -26174 41863
rect -26066 41897 -26014 41906
rect -26066 41863 -26057 41897
rect -26057 41863 -26023 41897
rect -26023 41863 -26014 41897
rect -26066 41854 -26014 41863
rect -25906 41897 -25854 41906
rect -25906 41863 -25897 41897
rect -25897 41863 -25863 41897
rect -25863 41863 -25854 41897
rect -25906 41854 -25854 41863
rect -25746 41897 -25694 41906
rect -25746 41863 -25737 41897
rect -25737 41863 -25703 41897
rect -25703 41863 -25694 41897
rect -25746 41854 -25694 41863
rect -25586 41897 -25534 41906
rect -25586 41863 -25577 41897
rect -25577 41863 -25543 41897
rect -25543 41863 -25534 41897
rect -25586 41854 -25534 41863
rect -25426 41897 -25374 41906
rect -25426 41863 -25417 41897
rect -25417 41863 -25383 41897
rect -25383 41863 -25374 41897
rect -25426 41854 -25374 41863
rect -25266 41897 -25214 41906
rect -25266 41863 -25257 41897
rect -25257 41863 -25223 41897
rect -25223 41863 -25214 41897
rect -25266 41854 -25214 41863
rect -25106 41897 -25054 41906
rect -25106 41863 -25097 41897
rect -25097 41863 -25063 41897
rect -25063 41863 -25054 41897
rect -25106 41854 -25054 41863
rect -24946 41897 -24894 41906
rect -24946 41863 -24937 41897
rect -24937 41863 -24903 41897
rect -24903 41863 -24894 41897
rect -24946 41854 -24894 41863
rect -24786 41897 -24734 41906
rect -24786 41863 -24777 41897
rect -24777 41863 -24743 41897
rect -24743 41863 -24734 41897
rect -24786 41854 -24734 41863
rect -24626 41897 -24574 41906
rect -24626 41863 -24617 41897
rect -24617 41863 -24583 41897
rect -24583 41863 -24574 41897
rect -24626 41854 -24574 41863
rect -24466 41897 -24414 41906
rect -24466 41863 -24457 41897
rect -24457 41863 -24423 41897
rect -24423 41863 -24414 41897
rect -24466 41854 -24414 41863
rect -24306 41897 -24254 41906
rect -24306 41863 -24297 41897
rect -24297 41863 -24263 41897
rect -24263 41863 -24254 41897
rect -24306 41854 -24254 41863
rect -24146 41897 -24094 41906
rect -24146 41863 -24137 41897
rect -24137 41863 -24103 41897
rect -24103 41863 -24094 41897
rect -24146 41854 -24094 41863
rect -23986 41897 -23934 41906
rect -23986 41863 -23977 41897
rect -23977 41863 -23943 41897
rect -23943 41863 -23934 41897
rect -23986 41854 -23934 41863
rect -23826 41897 -23774 41906
rect -23826 41863 -23817 41897
rect -23817 41863 -23783 41897
rect -23783 41863 -23774 41897
rect -23826 41854 -23774 41863
rect -23666 41897 -23614 41906
rect -23666 41863 -23657 41897
rect -23657 41863 -23623 41897
rect -23623 41863 -23614 41897
rect -23666 41854 -23614 41863
rect -23506 41897 -23454 41906
rect -23506 41863 -23497 41897
rect -23497 41863 -23463 41897
rect -23463 41863 -23454 41897
rect -23506 41854 -23454 41863
rect -23346 41897 -23294 41906
rect -23346 41863 -23337 41897
rect -23337 41863 -23303 41897
rect -23303 41863 -23294 41897
rect -23346 41854 -23294 41863
rect -23186 41897 -23134 41906
rect -23186 41863 -23177 41897
rect -23177 41863 -23143 41897
rect -23143 41863 -23134 41897
rect -23186 41854 -23134 41863
rect -23026 41897 -22974 41906
rect -23026 41863 -23017 41897
rect -23017 41863 -22983 41897
rect -22983 41863 -22974 41897
rect -23026 41854 -22974 41863
rect -22866 41897 -22814 41906
rect -22866 41863 -22857 41897
rect -22857 41863 -22823 41897
rect -22823 41863 -22814 41897
rect -22866 41854 -22814 41863
rect -22706 41897 -22654 41906
rect -22706 41863 -22697 41897
rect -22697 41863 -22663 41897
rect -22663 41863 -22654 41897
rect -22706 41854 -22654 41863
rect -22546 41897 -22494 41906
rect -22546 41863 -22537 41897
rect -22537 41863 -22503 41897
rect -22503 41863 -22494 41897
rect -22546 41854 -22494 41863
rect -22386 41897 -22334 41906
rect -22386 41863 -22377 41897
rect -22377 41863 -22343 41897
rect -22343 41863 -22334 41897
rect -22386 41854 -22334 41863
rect -22226 41897 -22174 41906
rect -22226 41863 -22217 41897
rect -22217 41863 -22183 41897
rect -22183 41863 -22174 41897
rect -22226 41854 -22174 41863
rect -22066 41897 -22014 41906
rect -22066 41863 -22057 41897
rect -22057 41863 -22023 41897
rect -22023 41863 -22014 41897
rect -22066 41854 -22014 41863
rect -21906 41897 -21854 41906
rect -21906 41863 -21897 41897
rect -21897 41863 -21863 41897
rect -21863 41863 -21854 41897
rect -21906 41854 -21854 41863
rect -21746 41897 -21694 41906
rect -21746 41863 -21737 41897
rect -21737 41863 -21703 41897
rect -21703 41863 -21694 41897
rect -21746 41854 -21694 41863
rect -21586 41897 -21534 41906
rect -21586 41863 -21577 41897
rect -21577 41863 -21543 41897
rect -21543 41863 -21534 41897
rect -21586 41854 -21534 41863
rect -21426 41897 -21374 41906
rect -21426 41863 -21417 41897
rect -21417 41863 -21383 41897
rect -21383 41863 -21374 41897
rect -21426 41854 -21374 41863
rect -21266 41897 -21214 41906
rect -21266 41863 -21257 41897
rect -21257 41863 -21223 41897
rect -21223 41863 -21214 41897
rect -21266 41854 -21214 41863
rect -21106 41897 -21054 41906
rect -21106 41863 -21097 41897
rect -21097 41863 -21063 41897
rect -21063 41863 -21054 41897
rect -21106 41854 -21054 41863
rect -20946 41897 -20894 41906
rect -20946 41863 -20937 41897
rect -20937 41863 -20903 41897
rect -20903 41863 -20894 41897
rect -20946 41854 -20894 41863
rect -20786 41897 -20734 41906
rect -20786 41863 -20777 41897
rect -20777 41863 -20743 41897
rect -20743 41863 -20734 41897
rect -20786 41854 -20734 41863
rect -20626 41897 -20574 41906
rect -20626 41863 -20617 41897
rect -20617 41863 -20583 41897
rect -20583 41863 -20574 41897
rect -20626 41854 -20574 41863
rect -20466 41897 -20414 41906
rect -20466 41863 -20457 41897
rect -20457 41863 -20423 41897
rect -20423 41863 -20414 41897
rect -20466 41854 -20414 41863
rect -20306 41897 -20254 41906
rect -20306 41863 -20297 41897
rect -20297 41863 -20263 41897
rect -20263 41863 -20254 41897
rect -20306 41854 -20254 41863
rect -20146 41897 -20094 41906
rect -20146 41863 -20137 41897
rect -20137 41863 -20103 41897
rect -20103 41863 -20094 41897
rect -20146 41854 -20094 41863
rect -19986 41897 -19934 41906
rect -19986 41863 -19977 41897
rect -19977 41863 -19943 41897
rect -19943 41863 -19934 41897
rect -19986 41854 -19934 41863
rect -19826 41897 -19774 41906
rect -19826 41863 -19817 41897
rect -19817 41863 -19783 41897
rect -19783 41863 -19774 41897
rect -19826 41854 -19774 41863
rect -19666 41897 -19614 41906
rect -19666 41863 -19657 41897
rect -19657 41863 -19623 41897
rect -19623 41863 -19614 41897
rect -19666 41854 -19614 41863
rect -19506 41897 -19454 41906
rect -19506 41863 -19497 41897
rect -19497 41863 -19463 41897
rect -19463 41863 -19454 41897
rect -19506 41854 -19454 41863
rect -19346 41897 -19294 41906
rect -19346 41863 -19337 41897
rect -19337 41863 -19303 41897
rect -19303 41863 -19294 41897
rect -19346 41854 -19294 41863
rect -19186 41897 -19134 41906
rect -19186 41863 -19177 41897
rect -19177 41863 -19143 41897
rect -19143 41863 -19134 41897
rect -19186 41854 -19134 41863
rect -19026 41897 -18974 41906
rect -19026 41863 -19017 41897
rect -19017 41863 -18983 41897
rect -18983 41863 -18974 41897
rect -19026 41854 -18974 41863
rect -18866 41897 -18814 41906
rect -18866 41863 -18857 41897
rect -18857 41863 -18823 41897
rect -18823 41863 -18814 41897
rect -18866 41854 -18814 41863
rect -18706 41897 -18654 41906
rect -18706 41863 -18697 41897
rect -18697 41863 -18663 41897
rect -18663 41863 -18654 41897
rect -18706 41854 -18654 41863
rect -18546 41897 -18494 41906
rect -18546 41863 -18537 41897
rect -18537 41863 -18503 41897
rect -18503 41863 -18494 41897
rect -18546 41854 -18494 41863
rect -18386 41897 -18334 41906
rect -18386 41863 -18377 41897
rect -18377 41863 -18343 41897
rect -18343 41863 -18334 41897
rect -18386 41854 -18334 41863
rect -18226 41897 -18174 41906
rect -18226 41863 -18217 41897
rect -18217 41863 -18183 41897
rect -18183 41863 -18174 41897
rect -18226 41854 -18174 41863
rect -18066 41897 -18014 41906
rect -18066 41863 -18057 41897
rect -18057 41863 -18023 41897
rect -18023 41863 -18014 41897
rect -18066 41854 -18014 41863
rect -17906 41897 -17854 41906
rect -17906 41863 -17897 41897
rect -17897 41863 -17863 41897
rect -17863 41863 -17854 41897
rect -17906 41854 -17854 41863
rect -17746 41897 -17694 41906
rect -17746 41863 -17737 41897
rect -17737 41863 -17703 41897
rect -17703 41863 -17694 41897
rect -17746 41854 -17694 41863
rect -17586 41897 -17534 41906
rect -17586 41863 -17577 41897
rect -17577 41863 -17543 41897
rect -17543 41863 -17534 41897
rect -17586 41854 -17534 41863
rect -17426 41897 -17374 41906
rect -17426 41863 -17417 41897
rect -17417 41863 -17383 41897
rect -17383 41863 -17374 41897
rect -17426 41854 -17374 41863
rect -17266 41897 -17214 41906
rect -17266 41863 -17257 41897
rect -17257 41863 -17223 41897
rect -17223 41863 -17214 41897
rect -17266 41854 -17214 41863
rect -17106 41897 -17054 41906
rect -17106 41863 -17097 41897
rect -17097 41863 -17063 41897
rect -17063 41863 -17054 41897
rect -17106 41854 -17054 41863
rect -16946 41897 -16894 41906
rect -16946 41863 -16937 41897
rect -16937 41863 -16903 41897
rect -16903 41863 -16894 41897
rect -16946 41854 -16894 41863
rect -16786 41897 -16734 41906
rect -16786 41863 -16777 41897
rect -16777 41863 -16743 41897
rect -16743 41863 -16734 41897
rect -16786 41854 -16734 41863
rect -16626 41897 -16574 41906
rect -16626 41863 -16617 41897
rect -16617 41863 -16583 41897
rect -16583 41863 -16574 41897
rect -16626 41854 -16574 41863
rect -16466 41897 -16414 41906
rect -16466 41863 -16457 41897
rect -16457 41863 -16423 41897
rect -16423 41863 -16414 41897
rect -16466 41854 -16414 41863
rect -16306 41897 -16254 41906
rect -16306 41863 -16297 41897
rect -16297 41863 -16263 41897
rect -16263 41863 -16254 41897
rect -16306 41854 -16254 41863
rect -16146 41897 -16094 41906
rect -16146 41863 -16137 41897
rect -16137 41863 -16103 41897
rect -16103 41863 -16094 41897
rect -16146 41854 -16094 41863
rect -15986 41897 -15934 41906
rect -15986 41863 -15977 41897
rect -15977 41863 -15943 41897
rect -15943 41863 -15934 41897
rect -15986 41854 -15934 41863
rect -15826 41897 -15774 41906
rect -15826 41863 -15817 41897
rect -15817 41863 -15783 41897
rect -15783 41863 -15774 41897
rect -15826 41854 -15774 41863
rect -15666 41897 -15614 41906
rect -15666 41863 -15657 41897
rect -15657 41863 -15623 41897
rect -15623 41863 -15614 41897
rect -15666 41854 -15614 41863
rect -15506 41897 -15454 41906
rect -15506 41863 -15497 41897
rect -15497 41863 -15463 41897
rect -15463 41863 -15454 41897
rect -15506 41854 -15454 41863
rect -15346 41897 -15294 41906
rect -15346 41863 -15337 41897
rect -15337 41863 -15303 41897
rect -15303 41863 -15294 41897
rect -15346 41854 -15294 41863
rect -15186 41897 -15134 41906
rect -15186 41863 -15177 41897
rect -15177 41863 -15143 41897
rect -15143 41863 -15134 41897
rect -15186 41854 -15134 41863
rect -15026 41897 -14974 41906
rect -15026 41863 -15017 41897
rect -15017 41863 -14983 41897
rect -14983 41863 -14974 41897
rect -15026 41854 -14974 41863
rect -14866 41897 -14814 41906
rect -14866 41863 -14857 41897
rect -14857 41863 -14823 41897
rect -14823 41863 -14814 41897
rect -14866 41854 -14814 41863
rect -14706 41897 -14654 41906
rect -14706 41863 -14697 41897
rect -14697 41863 -14663 41897
rect -14663 41863 -14654 41897
rect -14706 41854 -14654 41863
rect -14546 41897 -14494 41906
rect -14546 41863 -14537 41897
rect -14537 41863 -14503 41897
rect -14503 41863 -14494 41897
rect -14546 41854 -14494 41863
rect -14386 41897 -14334 41906
rect -14386 41863 -14377 41897
rect -14377 41863 -14343 41897
rect -14343 41863 -14334 41897
rect -14386 41854 -14334 41863
rect -14226 41897 -14174 41906
rect -14226 41863 -14217 41897
rect -14217 41863 -14183 41897
rect -14183 41863 -14174 41897
rect -14226 41854 -14174 41863
rect -14066 41897 -14014 41906
rect -14066 41863 -14057 41897
rect -14057 41863 -14023 41897
rect -14023 41863 -14014 41897
rect -14066 41854 -14014 41863
rect -13906 41897 -13854 41906
rect -13906 41863 -13897 41897
rect -13897 41863 -13863 41897
rect -13863 41863 -13854 41897
rect -13906 41854 -13854 41863
rect -13746 41897 -13694 41906
rect -13746 41863 -13737 41897
rect -13737 41863 -13703 41897
rect -13703 41863 -13694 41897
rect -13746 41854 -13694 41863
rect -13586 41897 -13534 41906
rect -13586 41863 -13577 41897
rect -13577 41863 -13543 41897
rect -13543 41863 -13534 41897
rect -13586 41854 -13534 41863
rect -13426 41897 -13374 41906
rect -13426 41863 -13417 41897
rect -13417 41863 -13383 41897
rect -13383 41863 -13374 41897
rect -13426 41854 -13374 41863
rect -13266 41897 -13214 41906
rect -13266 41863 -13257 41897
rect -13257 41863 -13223 41897
rect -13223 41863 -13214 41897
rect -13266 41854 -13214 41863
rect -13106 41897 -13054 41906
rect -13106 41863 -13097 41897
rect -13097 41863 -13063 41897
rect -13063 41863 -13054 41897
rect -13106 41854 -13054 41863
rect -12946 41897 -12894 41906
rect -12946 41863 -12937 41897
rect -12937 41863 -12903 41897
rect -12903 41863 -12894 41897
rect -12946 41854 -12894 41863
rect -12786 41897 -12734 41906
rect -12786 41863 -12777 41897
rect -12777 41863 -12743 41897
rect -12743 41863 -12734 41897
rect -12786 41854 -12734 41863
rect -12626 41897 -12574 41906
rect -12626 41863 -12617 41897
rect -12617 41863 -12583 41897
rect -12583 41863 -12574 41897
rect -12626 41854 -12574 41863
rect -12466 41897 -12414 41906
rect -12466 41863 -12457 41897
rect -12457 41863 -12423 41897
rect -12423 41863 -12414 41897
rect -12466 41854 -12414 41863
rect -12306 41897 -12254 41906
rect -12306 41863 -12297 41897
rect -12297 41863 -12263 41897
rect -12263 41863 -12254 41897
rect -12306 41854 -12254 41863
rect -11346 41897 -11294 41906
rect -11346 41863 -11337 41897
rect -11337 41863 -11303 41897
rect -11303 41863 -11294 41897
rect -11346 41854 -11294 41863
rect -11186 41897 -11134 41906
rect -11186 41863 -11177 41897
rect -11177 41863 -11143 41897
rect -11143 41863 -11134 41897
rect -11186 41854 -11134 41863
rect -11026 41897 -10974 41906
rect -11026 41863 -11017 41897
rect -11017 41863 -10983 41897
rect -10983 41863 -10974 41897
rect -11026 41854 -10974 41863
rect -10866 41897 -10814 41906
rect -10866 41863 -10857 41897
rect -10857 41863 -10823 41897
rect -10823 41863 -10814 41897
rect -10866 41854 -10814 41863
rect -10706 41897 -10654 41906
rect -10706 41863 -10697 41897
rect -10697 41863 -10663 41897
rect -10663 41863 -10654 41897
rect -10706 41854 -10654 41863
rect -10546 41897 -10494 41906
rect -10546 41863 -10537 41897
rect -10537 41863 -10503 41897
rect -10503 41863 -10494 41897
rect -10546 41854 -10494 41863
rect -10386 41897 -10334 41906
rect -10386 41863 -10377 41897
rect -10377 41863 -10343 41897
rect -10343 41863 -10334 41897
rect -10386 41854 -10334 41863
rect -10226 41897 -10174 41906
rect -10226 41863 -10217 41897
rect -10217 41863 -10183 41897
rect -10183 41863 -10174 41897
rect -10226 41854 -10174 41863
rect -10066 41897 -10014 41906
rect -10066 41863 -10057 41897
rect -10057 41863 -10023 41897
rect -10023 41863 -10014 41897
rect -10066 41854 -10014 41863
rect -9906 41897 -9854 41906
rect -9906 41863 -9897 41897
rect -9897 41863 -9863 41897
rect -9863 41863 -9854 41897
rect -9906 41854 -9854 41863
rect -9746 41897 -9694 41906
rect -9746 41863 -9737 41897
rect -9737 41863 -9703 41897
rect -9703 41863 -9694 41897
rect -9746 41854 -9694 41863
rect -9586 41897 -9534 41906
rect -9586 41863 -9577 41897
rect -9577 41863 -9543 41897
rect -9543 41863 -9534 41897
rect -9586 41854 -9534 41863
rect -9426 41897 -9374 41906
rect -9426 41863 -9417 41897
rect -9417 41863 -9383 41897
rect -9383 41863 -9374 41897
rect -9426 41854 -9374 41863
rect -9266 41897 -9214 41906
rect -9266 41863 -9257 41897
rect -9257 41863 -9223 41897
rect -9223 41863 -9214 41897
rect -9266 41854 -9214 41863
rect -9106 41897 -9054 41906
rect -9106 41863 -9097 41897
rect -9097 41863 -9063 41897
rect -9063 41863 -9054 41897
rect -9106 41854 -9054 41863
rect -8946 41897 -8894 41906
rect -8946 41863 -8937 41897
rect -8937 41863 -8903 41897
rect -8903 41863 -8894 41897
rect -8946 41854 -8894 41863
rect -8786 41897 -8734 41906
rect -8786 41863 -8777 41897
rect -8777 41863 -8743 41897
rect -8743 41863 -8734 41897
rect -8786 41854 -8734 41863
rect -8626 41897 -8574 41906
rect -8626 41863 -8617 41897
rect -8617 41863 -8583 41897
rect -8583 41863 -8574 41897
rect -8626 41854 -8574 41863
rect -8466 41897 -8414 41906
rect -8466 41863 -8457 41897
rect -8457 41863 -8423 41897
rect -8423 41863 -8414 41897
rect -8466 41854 -8414 41863
rect -8306 41897 -8254 41906
rect -8306 41863 -8297 41897
rect -8297 41863 -8263 41897
rect -8263 41863 -8254 41897
rect -8306 41854 -8254 41863
rect -8146 41897 -8094 41906
rect -8146 41863 -8137 41897
rect -8137 41863 -8103 41897
rect -8103 41863 -8094 41897
rect -8146 41854 -8094 41863
rect -7986 41897 -7934 41906
rect -7986 41863 -7977 41897
rect -7977 41863 -7943 41897
rect -7943 41863 -7934 41897
rect -7986 41854 -7934 41863
rect -7826 41897 -7774 41906
rect -7826 41863 -7817 41897
rect -7817 41863 -7783 41897
rect -7783 41863 -7774 41897
rect -7826 41854 -7774 41863
rect -7666 41897 -7614 41906
rect -7666 41863 -7657 41897
rect -7657 41863 -7623 41897
rect -7623 41863 -7614 41897
rect -7666 41854 -7614 41863
rect -7506 41897 -7454 41906
rect -7506 41863 -7497 41897
rect -7497 41863 -7463 41897
rect -7463 41863 -7454 41897
rect -7506 41854 -7454 41863
rect -7346 41897 -7294 41906
rect -7346 41863 -7337 41897
rect -7337 41863 -7303 41897
rect -7303 41863 -7294 41897
rect -7346 41854 -7294 41863
rect -7186 41897 -7134 41906
rect -7186 41863 -7177 41897
rect -7177 41863 -7143 41897
rect -7143 41863 -7134 41897
rect -7186 41854 -7134 41863
rect -7026 41897 -6974 41906
rect -7026 41863 -7017 41897
rect -7017 41863 -6983 41897
rect -6983 41863 -6974 41897
rect -7026 41854 -6974 41863
rect -6866 41897 -6814 41906
rect -6866 41863 -6857 41897
rect -6857 41863 -6823 41897
rect -6823 41863 -6814 41897
rect -6866 41854 -6814 41863
rect -6706 41897 -6654 41906
rect -6706 41863 -6697 41897
rect -6697 41863 -6663 41897
rect -6663 41863 -6654 41897
rect -6706 41854 -6654 41863
rect -6546 41897 -6494 41906
rect -6546 41863 -6537 41897
rect -6537 41863 -6503 41897
rect -6503 41863 -6494 41897
rect -6546 41854 -6494 41863
rect -6386 41897 -6334 41906
rect -6386 41863 -6377 41897
rect -6377 41863 -6343 41897
rect -6343 41863 -6334 41897
rect -6386 41854 -6334 41863
rect -6226 41897 -6174 41906
rect -6226 41863 -6217 41897
rect -6217 41863 -6183 41897
rect -6183 41863 -6174 41897
rect -6226 41854 -6174 41863
rect -6066 41897 -6014 41906
rect -6066 41863 -6057 41897
rect -6057 41863 -6023 41897
rect -6023 41863 -6014 41897
rect -6066 41854 -6014 41863
rect -5906 41897 -5854 41906
rect -5906 41863 -5897 41897
rect -5897 41863 -5863 41897
rect -5863 41863 -5854 41897
rect -5906 41854 -5854 41863
rect -5746 41897 -5694 41906
rect -5746 41863 -5737 41897
rect -5737 41863 -5703 41897
rect -5703 41863 -5694 41897
rect -5746 41854 -5694 41863
rect -5586 41897 -5534 41906
rect -5586 41863 -5577 41897
rect -5577 41863 -5543 41897
rect -5543 41863 -5534 41897
rect -5586 41854 -5534 41863
rect -5426 41897 -5374 41906
rect -5426 41863 -5417 41897
rect -5417 41863 -5383 41897
rect -5383 41863 -5374 41897
rect -5426 41854 -5374 41863
rect -5266 41897 -5214 41906
rect -5266 41863 -5257 41897
rect -5257 41863 -5223 41897
rect -5223 41863 -5214 41897
rect -5266 41854 -5214 41863
rect -5106 41897 -5054 41906
rect -5106 41863 -5097 41897
rect -5097 41863 -5063 41897
rect -5063 41863 -5054 41897
rect -5106 41854 -5054 41863
rect -4946 41897 -4894 41906
rect -4946 41863 -4937 41897
rect -4937 41863 -4903 41897
rect -4903 41863 -4894 41897
rect -4946 41854 -4894 41863
rect -4786 41897 -4734 41906
rect -4786 41863 -4777 41897
rect -4777 41863 -4743 41897
rect -4743 41863 -4734 41897
rect -4786 41854 -4734 41863
rect -4626 41897 -4574 41906
rect -4626 41863 -4617 41897
rect -4617 41863 -4583 41897
rect -4583 41863 -4574 41897
rect -4626 41854 -4574 41863
rect -4466 41897 -4414 41906
rect -4466 41863 -4457 41897
rect -4457 41863 -4423 41897
rect -4423 41863 -4414 41897
rect -4466 41854 -4414 41863
rect -4306 41897 -4254 41906
rect -4306 41863 -4297 41897
rect -4297 41863 -4263 41897
rect -4263 41863 -4254 41897
rect -4306 41854 -4254 41863
rect -4146 41897 -4094 41906
rect -4146 41863 -4137 41897
rect -4137 41863 -4103 41897
rect -4103 41863 -4094 41897
rect -4146 41854 -4094 41863
rect -3986 41897 -3934 41906
rect -3986 41863 -3977 41897
rect -3977 41863 -3943 41897
rect -3943 41863 -3934 41897
rect -3986 41854 -3934 41863
rect -3666 41897 -3614 41906
rect -3666 41863 -3657 41897
rect -3657 41863 -3623 41897
rect -3623 41863 -3614 41897
rect -3666 41854 -3614 41863
rect -3506 41897 -3454 41906
rect -3506 41863 -3497 41897
rect -3497 41863 -3463 41897
rect -3463 41863 -3454 41897
rect -3506 41854 -3454 41863
rect -3346 41897 -3294 41906
rect -3346 41863 -3337 41897
rect -3337 41863 -3303 41897
rect -3303 41863 -3294 41897
rect -3346 41854 -3294 41863
rect -3026 41897 -2974 41906
rect -3026 41863 -3017 41897
rect -3017 41863 -2983 41897
rect -2983 41863 -2974 41897
rect -3026 41854 -2974 41863
rect -2706 41897 -2654 41906
rect -2706 41863 -2697 41897
rect -2697 41863 -2663 41897
rect -2663 41863 -2654 41897
rect -2706 41854 -2654 41863
rect -2546 41897 -2494 41906
rect -2546 41863 -2537 41897
rect -2537 41863 -2503 41897
rect -2503 41863 -2494 41897
rect -2546 41854 -2494 41863
rect -2386 41897 -2334 41906
rect -2386 41863 -2377 41897
rect -2377 41863 -2343 41897
rect -2343 41863 -2334 41897
rect -2386 41854 -2334 41863
rect -2226 41897 -2174 41906
rect -2226 41863 -2217 41897
rect -2217 41863 -2183 41897
rect -2183 41863 -2174 41897
rect -2226 41854 -2174 41863
rect -2066 41897 -2014 41906
rect -2066 41863 -2057 41897
rect -2057 41863 -2023 41897
rect -2023 41863 -2014 41897
rect -2066 41854 -2014 41863
rect -1746 41897 -1694 41906
rect -1746 41863 -1737 41897
rect -1737 41863 -1703 41897
rect -1703 41863 -1694 41897
rect -1746 41854 -1694 41863
rect -1426 41897 -1374 41906
rect -1426 41863 -1417 41897
rect -1417 41863 -1383 41897
rect -1383 41863 -1374 41897
rect -1426 41854 -1374 41863
rect -1106 41897 -1054 41906
rect -1106 41863 -1097 41897
rect -1097 41863 -1063 41897
rect -1063 41863 -1054 41897
rect -1106 41854 -1054 41863
rect -33106 41337 -33054 41346
rect -33106 41303 -33097 41337
rect -33097 41303 -33063 41337
rect -33063 41303 -33054 41337
rect -33106 41294 -33054 41303
rect -32946 41337 -32894 41346
rect -32946 41303 -32937 41337
rect -32937 41303 -32903 41337
rect -32903 41303 -32894 41337
rect -32946 41294 -32894 41303
rect -32786 41337 -32734 41346
rect -32786 41303 -32777 41337
rect -32777 41303 -32743 41337
rect -32743 41303 -32734 41337
rect -32786 41294 -32734 41303
rect -32626 41337 -32574 41346
rect -32626 41303 -32617 41337
rect -32617 41303 -32583 41337
rect -32583 41303 -32574 41337
rect -32626 41294 -32574 41303
rect -32466 41337 -32414 41346
rect -32466 41303 -32457 41337
rect -32457 41303 -32423 41337
rect -32423 41303 -32414 41337
rect -32466 41294 -32414 41303
rect -32306 41337 -32254 41346
rect -32306 41303 -32297 41337
rect -32297 41303 -32263 41337
rect -32263 41303 -32254 41337
rect -32306 41294 -32254 41303
rect -32146 41337 -32094 41346
rect -32146 41303 -32137 41337
rect -32137 41303 -32103 41337
rect -32103 41303 -32094 41337
rect -32146 41294 -32094 41303
rect -31986 41337 -31934 41346
rect -31986 41303 -31977 41337
rect -31977 41303 -31943 41337
rect -31943 41303 -31934 41337
rect -31986 41294 -31934 41303
rect -31826 41337 -31774 41346
rect -31826 41303 -31817 41337
rect -31817 41303 -31783 41337
rect -31783 41303 -31774 41337
rect -31826 41294 -31774 41303
rect -31666 41337 -31614 41346
rect -31666 41303 -31657 41337
rect -31657 41303 -31623 41337
rect -31623 41303 -31614 41337
rect -31666 41294 -31614 41303
rect -31506 41337 -31454 41346
rect -31506 41303 -31497 41337
rect -31497 41303 -31463 41337
rect -31463 41303 -31454 41337
rect -31506 41294 -31454 41303
rect -31346 41337 -31294 41346
rect -31346 41303 -31337 41337
rect -31337 41303 -31303 41337
rect -31303 41303 -31294 41337
rect -31346 41294 -31294 41303
rect -31186 41337 -31134 41346
rect -31186 41303 -31177 41337
rect -31177 41303 -31143 41337
rect -31143 41303 -31134 41337
rect -31186 41294 -31134 41303
rect -29906 41337 -29854 41346
rect -29906 41303 -29897 41337
rect -29897 41303 -29863 41337
rect -29863 41303 -29854 41337
rect -29906 41294 -29854 41303
rect -29746 41337 -29694 41346
rect -29746 41303 -29737 41337
rect -29737 41303 -29703 41337
rect -29703 41303 -29694 41337
rect -29746 41294 -29694 41303
rect -29586 41337 -29534 41346
rect -29586 41303 -29577 41337
rect -29577 41303 -29543 41337
rect -29543 41303 -29534 41337
rect -29586 41294 -29534 41303
rect -29426 41337 -29374 41346
rect -29426 41303 -29417 41337
rect -29417 41303 -29383 41337
rect -29383 41303 -29374 41337
rect -29426 41294 -29374 41303
rect -29266 41337 -29214 41346
rect -29266 41303 -29257 41337
rect -29257 41303 -29223 41337
rect -29223 41303 -29214 41337
rect -29266 41294 -29214 41303
rect -29106 41337 -29054 41346
rect -29106 41303 -29097 41337
rect -29097 41303 -29063 41337
rect -29063 41303 -29054 41337
rect -29106 41294 -29054 41303
rect -28946 41337 -28894 41346
rect -28946 41303 -28937 41337
rect -28937 41303 -28903 41337
rect -28903 41303 -28894 41337
rect -28946 41294 -28894 41303
rect -28786 41337 -28734 41346
rect -28786 41303 -28777 41337
rect -28777 41303 -28743 41337
rect -28743 41303 -28734 41337
rect -28786 41294 -28734 41303
rect -28626 41337 -28574 41346
rect -28626 41303 -28617 41337
rect -28617 41303 -28583 41337
rect -28583 41303 -28574 41337
rect -28626 41294 -28574 41303
rect -28466 41337 -28414 41346
rect -28466 41303 -28457 41337
rect -28457 41303 -28423 41337
rect -28423 41303 -28414 41337
rect -28466 41294 -28414 41303
rect -28306 41337 -28254 41346
rect -28306 41303 -28297 41337
rect -28297 41303 -28263 41337
rect -28263 41303 -28254 41337
rect -28306 41294 -28254 41303
rect -28146 41337 -28094 41346
rect -28146 41303 -28137 41337
rect -28137 41303 -28103 41337
rect -28103 41303 -28094 41337
rect -28146 41294 -28094 41303
rect -27986 41337 -27934 41346
rect -27986 41303 -27977 41337
rect -27977 41303 -27943 41337
rect -27943 41303 -27934 41337
rect -27986 41294 -27934 41303
rect -27826 41337 -27774 41346
rect -27826 41303 -27817 41337
rect -27817 41303 -27783 41337
rect -27783 41303 -27774 41337
rect -27826 41294 -27774 41303
rect -27666 41337 -27614 41346
rect -27666 41303 -27657 41337
rect -27657 41303 -27623 41337
rect -27623 41303 -27614 41337
rect -27666 41294 -27614 41303
rect -27506 41337 -27454 41346
rect -27506 41303 -27497 41337
rect -27497 41303 -27463 41337
rect -27463 41303 -27454 41337
rect -27506 41294 -27454 41303
rect -27346 41337 -27294 41346
rect -27346 41303 -27337 41337
rect -27337 41303 -27303 41337
rect -27303 41303 -27294 41337
rect -27346 41294 -27294 41303
rect -27186 41337 -27134 41346
rect -27186 41303 -27177 41337
rect -27177 41303 -27143 41337
rect -27143 41303 -27134 41337
rect -27186 41294 -27134 41303
rect -27026 41337 -26974 41346
rect -27026 41303 -27017 41337
rect -27017 41303 -26983 41337
rect -26983 41303 -26974 41337
rect -27026 41294 -26974 41303
rect -26866 41337 -26814 41346
rect -26866 41303 -26857 41337
rect -26857 41303 -26823 41337
rect -26823 41303 -26814 41337
rect -26866 41294 -26814 41303
rect -26706 41337 -26654 41346
rect -26706 41303 -26697 41337
rect -26697 41303 -26663 41337
rect -26663 41303 -26654 41337
rect -26706 41294 -26654 41303
rect -26546 41337 -26494 41346
rect -26546 41303 -26537 41337
rect -26537 41303 -26503 41337
rect -26503 41303 -26494 41337
rect -26546 41294 -26494 41303
rect -26386 41337 -26334 41346
rect -26386 41303 -26377 41337
rect -26377 41303 -26343 41337
rect -26343 41303 -26334 41337
rect -26386 41294 -26334 41303
rect -26226 41337 -26174 41346
rect -26226 41303 -26217 41337
rect -26217 41303 -26183 41337
rect -26183 41303 -26174 41337
rect -26226 41294 -26174 41303
rect -26066 41337 -26014 41346
rect -26066 41303 -26057 41337
rect -26057 41303 -26023 41337
rect -26023 41303 -26014 41337
rect -26066 41294 -26014 41303
rect -25906 41337 -25854 41346
rect -25906 41303 -25897 41337
rect -25897 41303 -25863 41337
rect -25863 41303 -25854 41337
rect -25906 41294 -25854 41303
rect -25746 41337 -25694 41346
rect -25746 41303 -25737 41337
rect -25737 41303 -25703 41337
rect -25703 41303 -25694 41337
rect -25746 41294 -25694 41303
rect -25586 41337 -25534 41346
rect -25586 41303 -25577 41337
rect -25577 41303 -25543 41337
rect -25543 41303 -25534 41337
rect -25586 41294 -25534 41303
rect -25426 41337 -25374 41346
rect -25426 41303 -25417 41337
rect -25417 41303 -25383 41337
rect -25383 41303 -25374 41337
rect -25426 41294 -25374 41303
rect -25266 41337 -25214 41346
rect -25266 41303 -25257 41337
rect -25257 41303 -25223 41337
rect -25223 41303 -25214 41337
rect -25266 41294 -25214 41303
rect -25106 41337 -25054 41346
rect -25106 41303 -25097 41337
rect -25097 41303 -25063 41337
rect -25063 41303 -25054 41337
rect -25106 41294 -25054 41303
rect -24946 41337 -24894 41346
rect -24946 41303 -24937 41337
rect -24937 41303 -24903 41337
rect -24903 41303 -24894 41337
rect -24946 41294 -24894 41303
rect -24786 41337 -24734 41346
rect -24786 41303 -24777 41337
rect -24777 41303 -24743 41337
rect -24743 41303 -24734 41337
rect -24786 41294 -24734 41303
rect -24626 41337 -24574 41346
rect -24626 41303 -24617 41337
rect -24617 41303 -24583 41337
rect -24583 41303 -24574 41337
rect -24626 41294 -24574 41303
rect -24466 41337 -24414 41346
rect -24466 41303 -24457 41337
rect -24457 41303 -24423 41337
rect -24423 41303 -24414 41337
rect -24466 41294 -24414 41303
rect -24306 41337 -24254 41346
rect -24306 41303 -24297 41337
rect -24297 41303 -24263 41337
rect -24263 41303 -24254 41337
rect -24306 41294 -24254 41303
rect -24146 41337 -24094 41346
rect -24146 41303 -24137 41337
rect -24137 41303 -24103 41337
rect -24103 41303 -24094 41337
rect -24146 41294 -24094 41303
rect -23986 41337 -23934 41346
rect -23986 41303 -23977 41337
rect -23977 41303 -23943 41337
rect -23943 41303 -23934 41337
rect -23986 41294 -23934 41303
rect -23826 41337 -23774 41346
rect -23826 41303 -23817 41337
rect -23817 41303 -23783 41337
rect -23783 41303 -23774 41337
rect -23826 41294 -23774 41303
rect -23666 41337 -23614 41346
rect -23666 41303 -23657 41337
rect -23657 41303 -23623 41337
rect -23623 41303 -23614 41337
rect -23666 41294 -23614 41303
rect -23506 41337 -23454 41346
rect -23506 41303 -23497 41337
rect -23497 41303 -23463 41337
rect -23463 41303 -23454 41337
rect -23506 41294 -23454 41303
rect -23346 41337 -23294 41346
rect -23346 41303 -23337 41337
rect -23337 41303 -23303 41337
rect -23303 41303 -23294 41337
rect -23346 41294 -23294 41303
rect -23186 41337 -23134 41346
rect -23186 41303 -23177 41337
rect -23177 41303 -23143 41337
rect -23143 41303 -23134 41337
rect -23186 41294 -23134 41303
rect -23026 41337 -22974 41346
rect -23026 41303 -23017 41337
rect -23017 41303 -22983 41337
rect -22983 41303 -22974 41337
rect -23026 41294 -22974 41303
rect -22866 41337 -22814 41346
rect -22866 41303 -22857 41337
rect -22857 41303 -22823 41337
rect -22823 41303 -22814 41337
rect -22866 41294 -22814 41303
rect -22706 41337 -22654 41346
rect -22706 41303 -22697 41337
rect -22697 41303 -22663 41337
rect -22663 41303 -22654 41337
rect -22706 41294 -22654 41303
rect -22546 41337 -22494 41346
rect -22546 41303 -22537 41337
rect -22537 41303 -22503 41337
rect -22503 41303 -22494 41337
rect -22546 41294 -22494 41303
rect -22386 41337 -22334 41346
rect -22386 41303 -22377 41337
rect -22377 41303 -22343 41337
rect -22343 41303 -22334 41337
rect -22386 41294 -22334 41303
rect -22226 41337 -22174 41346
rect -22226 41303 -22217 41337
rect -22217 41303 -22183 41337
rect -22183 41303 -22174 41337
rect -22226 41294 -22174 41303
rect -22066 41337 -22014 41346
rect -22066 41303 -22057 41337
rect -22057 41303 -22023 41337
rect -22023 41303 -22014 41337
rect -22066 41294 -22014 41303
rect -21906 41337 -21854 41346
rect -21906 41303 -21897 41337
rect -21897 41303 -21863 41337
rect -21863 41303 -21854 41337
rect -21906 41294 -21854 41303
rect -21746 41337 -21694 41346
rect -21746 41303 -21737 41337
rect -21737 41303 -21703 41337
rect -21703 41303 -21694 41337
rect -21746 41294 -21694 41303
rect -21586 41337 -21534 41346
rect -21586 41303 -21577 41337
rect -21577 41303 -21543 41337
rect -21543 41303 -21534 41337
rect -21586 41294 -21534 41303
rect -21426 41337 -21374 41346
rect -21426 41303 -21417 41337
rect -21417 41303 -21383 41337
rect -21383 41303 -21374 41337
rect -21426 41294 -21374 41303
rect -21266 41337 -21214 41346
rect -21266 41303 -21257 41337
rect -21257 41303 -21223 41337
rect -21223 41303 -21214 41337
rect -21266 41294 -21214 41303
rect -21106 41337 -21054 41346
rect -21106 41303 -21097 41337
rect -21097 41303 -21063 41337
rect -21063 41303 -21054 41337
rect -21106 41294 -21054 41303
rect -20946 41337 -20894 41346
rect -20946 41303 -20937 41337
rect -20937 41303 -20903 41337
rect -20903 41303 -20894 41337
rect -20946 41294 -20894 41303
rect -20786 41337 -20734 41346
rect -20786 41303 -20777 41337
rect -20777 41303 -20743 41337
rect -20743 41303 -20734 41337
rect -20786 41294 -20734 41303
rect -20626 41337 -20574 41346
rect -20626 41303 -20617 41337
rect -20617 41303 -20583 41337
rect -20583 41303 -20574 41337
rect -20626 41294 -20574 41303
rect -20466 41337 -20414 41346
rect -20466 41303 -20457 41337
rect -20457 41303 -20423 41337
rect -20423 41303 -20414 41337
rect -20466 41294 -20414 41303
rect -20306 41337 -20254 41346
rect -20306 41303 -20297 41337
rect -20297 41303 -20263 41337
rect -20263 41303 -20254 41337
rect -20306 41294 -20254 41303
rect -20146 41337 -20094 41346
rect -20146 41303 -20137 41337
rect -20137 41303 -20103 41337
rect -20103 41303 -20094 41337
rect -20146 41294 -20094 41303
rect -19986 41337 -19934 41346
rect -19986 41303 -19977 41337
rect -19977 41303 -19943 41337
rect -19943 41303 -19934 41337
rect -19986 41294 -19934 41303
rect -19826 41337 -19774 41346
rect -19826 41303 -19817 41337
rect -19817 41303 -19783 41337
rect -19783 41303 -19774 41337
rect -19826 41294 -19774 41303
rect -19666 41337 -19614 41346
rect -19666 41303 -19657 41337
rect -19657 41303 -19623 41337
rect -19623 41303 -19614 41337
rect -19666 41294 -19614 41303
rect -19506 41337 -19454 41346
rect -19506 41303 -19497 41337
rect -19497 41303 -19463 41337
rect -19463 41303 -19454 41337
rect -19506 41294 -19454 41303
rect -19346 41337 -19294 41346
rect -19346 41303 -19337 41337
rect -19337 41303 -19303 41337
rect -19303 41303 -19294 41337
rect -19346 41294 -19294 41303
rect -19186 41337 -19134 41346
rect -19186 41303 -19177 41337
rect -19177 41303 -19143 41337
rect -19143 41303 -19134 41337
rect -19186 41294 -19134 41303
rect -19026 41337 -18974 41346
rect -19026 41303 -19017 41337
rect -19017 41303 -18983 41337
rect -18983 41303 -18974 41337
rect -19026 41294 -18974 41303
rect -18866 41337 -18814 41346
rect -18866 41303 -18857 41337
rect -18857 41303 -18823 41337
rect -18823 41303 -18814 41337
rect -18866 41294 -18814 41303
rect -18706 41337 -18654 41346
rect -18706 41303 -18697 41337
rect -18697 41303 -18663 41337
rect -18663 41303 -18654 41337
rect -18706 41294 -18654 41303
rect -18546 41337 -18494 41346
rect -18546 41303 -18537 41337
rect -18537 41303 -18503 41337
rect -18503 41303 -18494 41337
rect -18546 41294 -18494 41303
rect -18386 41337 -18334 41346
rect -18386 41303 -18377 41337
rect -18377 41303 -18343 41337
rect -18343 41303 -18334 41337
rect -18386 41294 -18334 41303
rect -18226 41337 -18174 41346
rect -18226 41303 -18217 41337
rect -18217 41303 -18183 41337
rect -18183 41303 -18174 41337
rect -18226 41294 -18174 41303
rect -18066 41337 -18014 41346
rect -18066 41303 -18057 41337
rect -18057 41303 -18023 41337
rect -18023 41303 -18014 41337
rect -18066 41294 -18014 41303
rect -17906 41337 -17854 41346
rect -17906 41303 -17897 41337
rect -17897 41303 -17863 41337
rect -17863 41303 -17854 41337
rect -17906 41294 -17854 41303
rect -17746 41337 -17694 41346
rect -17746 41303 -17737 41337
rect -17737 41303 -17703 41337
rect -17703 41303 -17694 41337
rect -17746 41294 -17694 41303
rect -17586 41337 -17534 41346
rect -17586 41303 -17577 41337
rect -17577 41303 -17543 41337
rect -17543 41303 -17534 41337
rect -17586 41294 -17534 41303
rect -17426 41337 -17374 41346
rect -17426 41303 -17417 41337
rect -17417 41303 -17383 41337
rect -17383 41303 -17374 41337
rect -17426 41294 -17374 41303
rect -17266 41337 -17214 41346
rect -17266 41303 -17257 41337
rect -17257 41303 -17223 41337
rect -17223 41303 -17214 41337
rect -17266 41294 -17214 41303
rect -17106 41337 -17054 41346
rect -17106 41303 -17097 41337
rect -17097 41303 -17063 41337
rect -17063 41303 -17054 41337
rect -17106 41294 -17054 41303
rect -16946 41337 -16894 41346
rect -16946 41303 -16937 41337
rect -16937 41303 -16903 41337
rect -16903 41303 -16894 41337
rect -16946 41294 -16894 41303
rect -16786 41337 -16734 41346
rect -16786 41303 -16777 41337
rect -16777 41303 -16743 41337
rect -16743 41303 -16734 41337
rect -16786 41294 -16734 41303
rect -16626 41337 -16574 41346
rect -16626 41303 -16617 41337
rect -16617 41303 -16583 41337
rect -16583 41303 -16574 41337
rect -16626 41294 -16574 41303
rect -16466 41337 -16414 41346
rect -16466 41303 -16457 41337
rect -16457 41303 -16423 41337
rect -16423 41303 -16414 41337
rect -16466 41294 -16414 41303
rect -16306 41337 -16254 41346
rect -16306 41303 -16297 41337
rect -16297 41303 -16263 41337
rect -16263 41303 -16254 41337
rect -16306 41294 -16254 41303
rect -16146 41337 -16094 41346
rect -16146 41303 -16137 41337
rect -16137 41303 -16103 41337
rect -16103 41303 -16094 41337
rect -16146 41294 -16094 41303
rect -15986 41337 -15934 41346
rect -15986 41303 -15977 41337
rect -15977 41303 -15943 41337
rect -15943 41303 -15934 41337
rect -15986 41294 -15934 41303
rect -15826 41337 -15774 41346
rect -15826 41303 -15817 41337
rect -15817 41303 -15783 41337
rect -15783 41303 -15774 41337
rect -15826 41294 -15774 41303
rect -15666 41337 -15614 41346
rect -15666 41303 -15657 41337
rect -15657 41303 -15623 41337
rect -15623 41303 -15614 41337
rect -15666 41294 -15614 41303
rect -15506 41337 -15454 41346
rect -15506 41303 -15497 41337
rect -15497 41303 -15463 41337
rect -15463 41303 -15454 41337
rect -15506 41294 -15454 41303
rect -15346 41337 -15294 41346
rect -15346 41303 -15337 41337
rect -15337 41303 -15303 41337
rect -15303 41303 -15294 41337
rect -15346 41294 -15294 41303
rect -15186 41337 -15134 41346
rect -15186 41303 -15177 41337
rect -15177 41303 -15143 41337
rect -15143 41303 -15134 41337
rect -15186 41294 -15134 41303
rect -15026 41337 -14974 41346
rect -15026 41303 -15017 41337
rect -15017 41303 -14983 41337
rect -14983 41303 -14974 41337
rect -15026 41294 -14974 41303
rect -14866 41337 -14814 41346
rect -14866 41303 -14857 41337
rect -14857 41303 -14823 41337
rect -14823 41303 -14814 41337
rect -14866 41294 -14814 41303
rect -14706 41337 -14654 41346
rect -14706 41303 -14697 41337
rect -14697 41303 -14663 41337
rect -14663 41303 -14654 41337
rect -14706 41294 -14654 41303
rect -14546 41337 -14494 41346
rect -14546 41303 -14537 41337
rect -14537 41303 -14503 41337
rect -14503 41303 -14494 41337
rect -14546 41294 -14494 41303
rect -14386 41337 -14334 41346
rect -14386 41303 -14377 41337
rect -14377 41303 -14343 41337
rect -14343 41303 -14334 41337
rect -14386 41294 -14334 41303
rect -14226 41337 -14174 41346
rect -14226 41303 -14217 41337
rect -14217 41303 -14183 41337
rect -14183 41303 -14174 41337
rect -14226 41294 -14174 41303
rect -14066 41337 -14014 41346
rect -14066 41303 -14057 41337
rect -14057 41303 -14023 41337
rect -14023 41303 -14014 41337
rect -14066 41294 -14014 41303
rect -13906 41337 -13854 41346
rect -13906 41303 -13897 41337
rect -13897 41303 -13863 41337
rect -13863 41303 -13854 41337
rect -13906 41294 -13854 41303
rect -13746 41337 -13694 41346
rect -13746 41303 -13737 41337
rect -13737 41303 -13703 41337
rect -13703 41303 -13694 41337
rect -13746 41294 -13694 41303
rect -13586 41337 -13534 41346
rect -13586 41303 -13577 41337
rect -13577 41303 -13543 41337
rect -13543 41303 -13534 41337
rect -13586 41294 -13534 41303
rect -13426 41337 -13374 41346
rect -13426 41303 -13417 41337
rect -13417 41303 -13383 41337
rect -13383 41303 -13374 41337
rect -13426 41294 -13374 41303
rect -13266 41337 -13214 41346
rect -13266 41303 -13257 41337
rect -13257 41303 -13223 41337
rect -13223 41303 -13214 41337
rect -13266 41294 -13214 41303
rect -13106 41337 -13054 41346
rect -13106 41303 -13097 41337
rect -13097 41303 -13063 41337
rect -13063 41303 -13054 41337
rect -13106 41294 -13054 41303
rect -12946 41337 -12894 41346
rect -12946 41303 -12937 41337
rect -12937 41303 -12903 41337
rect -12903 41303 -12894 41337
rect -12946 41294 -12894 41303
rect -12786 41337 -12734 41346
rect -12786 41303 -12777 41337
rect -12777 41303 -12743 41337
rect -12743 41303 -12734 41337
rect -12786 41294 -12734 41303
rect -12626 41337 -12574 41346
rect -12626 41303 -12617 41337
rect -12617 41303 -12583 41337
rect -12583 41303 -12574 41337
rect -12626 41294 -12574 41303
rect -12466 41337 -12414 41346
rect -12466 41303 -12457 41337
rect -12457 41303 -12423 41337
rect -12423 41303 -12414 41337
rect -12466 41294 -12414 41303
rect -12306 41337 -12254 41346
rect -12306 41303 -12297 41337
rect -12297 41303 -12263 41337
rect -12263 41303 -12254 41337
rect -12306 41294 -12254 41303
rect -11346 41337 -11294 41346
rect -11346 41303 -11337 41337
rect -11337 41303 -11303 41337
rect -11303 41303 -11294 41337
rect -11346 41294 -11294 41303
rect -11186 41337 -11134 41346
rect -11186 41303 -11177 41337
rect -11177 41303 -11143 41337
rect -11143 41303 -11134 41337
rect -11186 41294 -11134 41303
rect -11026 41337 -10974 41346
rect -11026 41303 -11017 41337
rect -11017 41303 -10983 41337
rect -10983 41303 -10974 41337
rect -11026 41294 -10974 41303
rect -10866 41337 -10814 41346
rect -10866 41303 -10857 41337
rect -10857 41303 -10823 41337
rect -10823 41303 -10814 41337
rect -10866 41294 -10814 41303
rect -10706 41337 -10654 41346
rect -10706 41303 -10697 41337
rect -10697 41303 -10663 41337
rect -10663 41303 -10654 41337
rect -10706 41294 -10654 41303
rect -10546 41337 -10494 41346
rect -10546 41303 -10537 41337
rect -10537 41303 -10503 41337
rect -10503 41303 -10494 41337
rect -10546 41294 -10494 41303
rect -10386 41337 -10334 41346
rect -10386 41303 -10377 41337
rect -10377 41303 -10343 41337
rect -10343 41303 -10334 41337
rect -10386 41294 -10334 41303
rect -10226 41337 -10174 41346
rect -10226 41303 -10217 41337
rect -10217 41303 -10183 41337
rect -10183 41303 -10174 41337
rect -10226 41294 -10174 41303
rect -10066 41337 -10014 41346
rect -10066 41303 -10057 41337
rect -10057 41303 -10023 41337
rect -10023 41303 -10014 41337
rect -10066 41294 -10014 41303
rect -9906 41337 -9854 41346
rect -9906 41303 -9897 41337
rect -9897 41303 -9863 41337
rect -9863 41303 -9854 41337
rect -9906 41294 -9854 41303
rect -9746 41337 -9694 41346
rect -9746 41303 -9737 41337
rect -9737 41303 -9703 41337
rect -9703 41303 -9694 41337
rect -9746 41294 -9694 41303
rect -9586 41337 -9534 41346
rect -9586 41303 -9577 41337
rect -9577 41303 -9543 41337
rect -9543 41303 -9534 41337
rect -9586 41294 -9534 41303
rect -9426 41337 -9374 41346
rect -9426 41303 -9417 41337
rect -9417 41303 -9383 41337
rect -9383 41303 -9374 41337
rect -9426 41294 -9374 41303
rect -9266 41337 -9214 41346
rect -9266 41303 -9257 41337
rect -9257 41303 -9223 41337
rect -9223 41303 -9214 41337
rect -9266 41294 -9214 41303
rect -9106 41337 -9054 41346
rect -9106 41303 -9097 41337
rect -9097 41303 -9063 41337
rect -9063 41303 -9054 41337
rect -9106 41294 -9054 41303
rect -8946 41337 -8894 41346
rect -8946 41303 -8937 41337
rect -8937 41303 -8903 41337
rect -8903 41303 -8894 41337
rect -8946 41294 -8894 41303
rect -8786 41337 -8734 41346
rect -8786 41303 -8777 41337
rect -8777 41303 -8743 41337
rect -8743 41303 -8734 41337
rect -8786 41294 -8734 41303
rect -8626 41337 -8574 41346
rect -8626 41303 -8617 41337
rect -8617 41303 -8583 41337
rect -8583 41303 -8574 41337
rect -8626 41294 -8574 41303
rect -8466 41337 -8414 41346
rect -8466 41303 -8457 41337
rect -8457 41303 -8423 41337
rect -8423 41303 -8414 41337
rect -8466 41294 -8414 41303
rect -8306 41337 -8254 41346
rect -8306 41303 -8297 41337
rect -8297 41303 -8263 41337
rect -8263 41303 -8254 41337
rect -8306 41294 -8254 41303
rect -8146 41337 -8094 41346
rect -8146 41303 -8137 41337
rect -8137 41303 -8103 41337
rect -8103 41303 -8094 41337
rect -8146 41294 -8094 41303
rect -7986 41337 -7934 41346
rect -7986 41303 -7977 41337
rect -7977 41303 -7943 41337
rect -7943 41303 -7934 41337
rect -7986 41294 -7934 41303
rect -7826 41337 -7774 41346
rect -7826 41303 -7817 41337
rect -7817 41303 -7783 41337
rect -7783 41303 -7774 41337
rect -7826 41294 -7774 41303
rect -7666 41337 -7614 41346
rect -7666 41303 -7657 41337
rect -7657 41303 -7623 41337
rect -7623 41303 -7614 41337
rect -7666 41294 -7614 41303
rect -7506 41337 -7454 41346
rect -7506 41303 -7497 41337
rect -7497 41303 -7463 41337
rect -7463 41303 -7454 41337
rect -7506 41294 -7454 41303
rect -7346 41337 -7294 41346
rect -7346 41303 -7337 41337
rect -7337 41303 -7303 41337
rect -7303 41303 -7294 41337
rect -7346 41294 -7294 41303
rect -7186 41337 -7134 41346
rect -7186 41303 -7177 41337
rect -7177 41303 -7143 41337
rect -7143 41303 -7134 41337
rect -7186 41294 -7134 41303
rect -7026 41337 -6974 41346
rect -7026 41303 -7017 41337
rect -7017 41303 -6983 41337
rect -6983 41303 -6974 41337
rect -7026 41294 -6974 41303
rect -6866 41337 -6814 41346
rect -6866 41303 -6857 41337
rect -6857 41303 -6823 41337
rect -6823 41303 -6814 41337
rect -6866 41294 -6814 41303
rect -6706 41337 -6654 41346
rect -6706 41303 -6697 41337
rect -6697 41303 -6663 41337
rect -6663 41303 -6654 41337
rect -6706 41294 -6654 41303
rect -6546 41337 -6494 41346
rect -6546 41303 -6537 41337
rect -6537 41303 -6503 41337
rect -6503 41303 -6494 41337
rect -6546 41294 -6494 41303
rect -6386 41337 -6334 41346
rect -6386 41303 -6377 41337
rect -6377 41303 -6343 41337
rect -6343 41303 -6334 41337
rect -6386 41294 -6334 41303
rect -6226 41337 -6174 41346
rect -6226 41303 -6217 41337
rect -6217 41303 -6183 41337
rect -6183 41303 -6174 41337
rect -6226 41294 -6174 41303
rect -6066 41337 -6014 41346
rect -6066 41303 -6057 41337
rect -6057 41303 -6023 41337
rect -6023 41303 -6014 41337
rect -6066 41294 -6014 41303
rect -5906 41337 -5854 41346
rect -5906 41303 -5897 41337
rect -5897 41303 -5863 41337
rect -5863 41303 -5854 41337
rect -5906 41294 -5854 41303
rect -5746 41337 -5694 41346
rect -5746 41303 -5737 41337
rect -5737 41303 -5703 41337
rect -5703 41303 -5694 41337
rect -5746 41294 -5694 41303
rect -5586 41337 -5534 41346
rect -5586 41303 -5577 41337
rect -5577 41303 -5543 41337
rect -5543 41303 -5534 41337
rect -5586 41294 -5534 41303
rect -5426 41337 -5374 41346
rect -5426 41303 -5417 41337
rect -5417 41303 -5383 41337
rect -5383 41303 -5374 41337
rect -5426 41294 -5374 41303
rect -5266 41337 -5214 41346
rect -5266 41303 -5257 41337
rect -5257 41303 -5223 41337
rect -5223 41303 -5214 41337
rect -5266 41294 -5214 41303
rect -5106 41337 -5054 41346
rect -5106 41303 -5097 41337
rect -5097 41303 -5063 41337
rect -5063 41303 -5054 41337
rect -5106 41294 -5054 41303
rect -4946 41337 -4894 41346
rect -4946 41303 -4937 41337
rect -4937 41303 -4903 41337
rect -4903 41303 -4894 41337
rect -4946 41294 -4894 41303
rect -4786 41337 -4734 41346
rect -4786 41303 -4777 41337
rect -4777 41303 -4743 41337
rect -4743 41303 -4734 41337
rect -4786 41294 -4734 41303
rect -4626 41337 -4574 41346
rect -4626 41303 -4617 41337
rect -4617 41303 -4583 41337
rect -4583 41303 -4574 41337
rect -4626 41294 -4574 41303
rect -4466 41337 -4414 41346
rect -4466 41303 -4457 41337
rect -4457 41303 -4423 41337
rect -4423 41303 -4414 41337
rect -4466 41294 -4414 41303
rect -4306 41337 -4254 41346
rect -4306 41303 -4297 41337
rect -4297 41303 -4263 41337
rect -4263 41303 -4254 41337
rect -4306 41294 -4254 41303
rect -4146 41337 -4094 41346
rect -4146 41303 -4137 41337
rect -4137 41303 -4103 41337
rect -4103 41303 -4094 41337
rect -4146 41294 -4094 41303
rect -3986 41337 -3934 41346
rect -3986 41303 -3977 41337
rect -3977 41303 -3943 41337
rect -3943 41303 -3934 41337
rect -3986 41294 -3934 41303
rect -3666 41337 -3614 41346
rect -3666 41303 -3657 41337
rect -3657 41303 -3623 41337
rect -3623 41303 -3614 41337
rect -3666 41294 -3614 41303
rect -3506 41337 -3454 41346
rect -3506 41303 -3497 41337
rect -3497 41303 -3463 41337
rect -3463 41303 -3454 41337
rect -3506 41294 -3454 41303
rect 41054 41337 41106 41346
rect 41054 41303 41063 41337
rect 41063 41303 41097 41337
rect 41097 41303 41106 41337
rect 41054 41294 41106 41303
rect 41214 41337 41266 41346
rect 41214 41303 41223 41337
rect 41223 41303 41257 41337
rect 41257 41303 41266 41337
rect 41214 41294 41266 41303
rect 41374 41337 41426 41346
rect 41374 41303 41383 41337
rect 41383 41303 41417 41337
rect 41417 41303 41426 41337
rect 41374 41294 41426 41303
rect 41534 41337 41586 41346
rect 41534 41303 41543 41337
rect 41543 41303 41577 41337
rect 41577 41303 41586 41337
rect 41534 41294 41586 41303
rect 41694 41337 41746 41346
rect 41694 41303 41703 41337
rect 41703 41303 41737 41337
rect 41737 41303 41746 41337
rect 41694 41294 41746 41303
rect 41854 41337 41906 41346
rect 41854 41303 41863 41337
rect 41863 41303 41897 41337
rect 41897 41303 41906 41337
rect 41854 41294 41906 41303
rect 42014 41337 42066 41346
rect 42014 41303 42023 41337
rect 42023 41303 42057 41337
rect 42057 41303 42066 41337
rect 42014 41294 42066 41303
rect 42174 41337 42226 41346
rect 42174 41303 42183 41337
rect 42183 41303 42217 41337
rect 42217 41303 42226 41337
rect 42174 41294 42226 41303
rect 42334 41337 42386 41346
rect 42334 41303 42343 41337
rect 42343 41303 42377 41337
rect 42377 41303 42386 41337
rect 42334 41294 42386 41303
rect 42494 41337 42546 41346
rect 42494 41303 42503 41337
rect 42503 41303 42537 41337
rect 42537 41303 42546 41337
rect 42494 41294 42546 41303
rect 42654 41337 42706 41346
rect 42654 41303 42663 41337
rect 42663 41303 42697 41337
rect 42697 41303 42706 41337
rect 42654 41294 42706 41303
rect 42814 41337 42866 41346
rect 42814 41303 42823 41337
rect 42823 41303 42857 41337
rect 42857 41303 42866 41337
rect 42814 41294 42866 41303
rect 42974 41337 43026 41346
rect 42974 41303 42983 41337
rect 42983 41303 43017 41337
rect 43017 41303 43026 41337
rect 42974 41294 43026 41303
rect 43134 41337 43186 41346
rect 43134 41303 43143 41337
rect 43143 41303 43177 41337
rect 43177 41303 43186 41337
rect 43134 41294 43186 41303
rect -33106 41017 -33054 41026
rect -33106 40983 -33097 41017
rect -33097 40983 -33063 41017
rect -33063 40983 -33054 41017
rect -33106 40974 -33054 40983
rect -32946 41017 -32894 41026
rect -32946 40983 -32937 41017
rect -32937 40983 -32903 41017
rect -32903 40983 -32894 41017
rect -32946 40974 -32894 40983
rect -32786 41017 -32734 41026
rect -32786 40983 -32777 41017
rect -32777 40983 -32743 41017
rect -32743 40983 -32734 41017
rect -32786 40974 -32734 40983
rect -32626 41017 -32574 41026
rect -32626 40983 -32617 41017
rect -32617 40983 -32583 41017
rect -32583 40983 -32574 41017
rect -32626 40974 -32574 40983
rect -32466 41017 -32414 41026
rect -32466 40983 -32457 41017
rect -32457 40983 -32423 41017
rect -32423 40983 -32414 41017
rect -32466 40974 -32414 40983
rect -32306 41017 -32254 41026
rect -32306 40983 -32297 41017
rect -32297 40983 -32263 41017
rect -32263 40983 -32254 41017
rect -32306 40974 -32254 40983
rect -32146 41017 -32094 41026
rect -32146 40983 -32137 41017
rect -32137 40983 -32103 41017
rect -32103 40983 -32094 41017
rect -32146 40974 -32094 40983
rect -31986 41017 -31934 41026
rect -31986 40983 -31977 41017
rect -31977 40983 -31943 41017
rect -31943 40983 -31934 41017
rect -31986 40974 -31934 40983
rect -31826 41017 -31774 41026
rect -31826 40983 -31817 41017
rect -31817 40983 -31783 41017
rect -31783 40983 -31774 41017
rect -31826 40974 -31774 40983
rect -31666 41017 -31614 41026
rect -31666 40983 -31657 41017
rect -31657 40983 -31623 41017
rect -31623 40983 -31614 41017
rect -31666 40974 -31614 40983
rect -31506 41017 -31454 41026
rect -31506 40983 -31497 41017
rect -31497 40983 -31463 41017
rect -31463 40983 -31454 41017
rect -31506 40974 -31454 40983
rect -31346 41017 -31294 41026
rect -31346 40983 -31337 41017
rect -31337 40983 -31303 41017
rect -31303 40983 -31294 41017
rect -31346 40974 -31294 40983
rect -31186 41017 -31134 41026
rect -31186 40983 -31177 41017
rect -31177 40983 -31143 41017
rect -31143 40983 -31134 41017
rect -31186 40974 -31134 40983
rect -29906 41017 -29854 41026
rect -29906 40983 -29897 41017
rect -29897 40983 -29863 41017
rect -29863 40983 -29854 41017
rect -29906 40974 -29854 40983
rect -29746 41017 -29694 41026
rect -29746 40983 -29737 41017
rect -29737 40983 -29703 41017
rect -29703 40983 -29694 41017
rect -29746 40974 -29694 40983
rect -29586 41017 -29534 41026
rect -29586 40983 -29577 41017
rect -29577 40983 -29543 41017
rect -29543 40983 -29534 41017
rect -29586 40974 -29534 40983
rect -29426 41017 -29374 41026
rect -29426 40983 -29417 41017
rect -29417 40983 -29383 41017
rect -29383 40983 -29374 41017
rect -29426 40974 -29374 40983
rect -29266 41017 -29214 41026
rect -29266 40983 -29257 41017
rect -29257 40983 -29223 41017
rect -29223 40983 -29214 41017
rect -29266 40974 -29214 40983
rect -29106 41017 -29054 41026
rect -29106 40983 -29097 41017
rect -29097 40983 -29063 41017
rect -29063 40983 -29054 41017
rect -29106 40974 -29054 40983
rect -28946 41017 -28894 41026
rect -28946 40983 -28937 41017
rect -28937 40983 -28903 41017
rect -28903 40983 -28894 41017
rect -28946 40974 -28894 40983
rect -28786 41017 -28734 41026
rect -28786 40983 -28777 41017
rect -28777 40983 -28743 41017
rect -28743 40983 -28734 41017
rect -28786 40974 -28734 40983
rect -28626 41017 -28574 41026
rect -28626 40983 -28617 41017
rect -28617 40983 -28583 41017
rect -28583 40983 -28574 41017
rect -28626 40974 -28574 40983
rect -28466 41017 -28414 41026
rect -28466 40983 -28457 41017
rect -28457 40983 -28423 41017
rect -28423 40983 -28414 41017
rect -28466 40974 -28414 40983
rect -28306 41017 -28254 41026
rect -28306 40983 -28297 41017
rect -28297 40983 -28263 41017
rect -28263 40983 -28254 41017
rect -28306 40974 -28254 40983
rect -28146 41017 -28094 41026
rect -28146 40983 -28137 41017
rect -28137 40983 -28103 41017
rect -28103 40983 -28094 41017
rect -28146 40974 -28094 40983
rect -27986 41017 -27934 41026
rect -27986 40983 -27977 41017
rect -27977 40983 -27943 41017
rect -27943 40983 -27934 41017
rect -27986 40974 -27934 40983
rect -27826 41017 -27774 41026
rect -27826 40983 -27817 41017
rect -27817 40983 -27783 41017
rect -27783 40983 -27774 41017
rect -27826 40974 -27774 40983
rect -27666 41017 -27614 41026
rect -27666 40983 -27657 41017
rect -27657 40983 -27623 41017
rect -27623 40983 -27614 41017
rect -27666 40974 -27614 40983
rect -27506 41017 -27454 41026
rect -27506 40983 -27497 41017
rect -27497 40983 -27463 41017
rect -27463 40983 -27454 41017
rect -27506 40974 -27454 40983
rect -27346 41017 -27294 41026
rect -27346 40983 -27337 41017
rect -27337 40983 -27303 41017
rect -27303 40983 -27294 41017
rect -27346 40974 -27294 40983
rect -27186 41017 -27134 41026
rect -27186 40983 -27177 41017
rect -27177 40983 -27143 41017
rect -27143 40983 -27134 41017
rect -27186 40974 -27134 40983
rect -27026 41017 -26974 41026
rect -27026 40983 -27017 41017
rect -27017 40983 -26983 41017
rect -26983 40983 -26974 41017
rect -27026 40974 -26974 40983
rect -26866 41017 -26814 41026
rect -26866 40983 -26857 41017
rect -26857 40983 -26823 41017
rect -26823 40983 -26814 41017
rect -26866 40974 -26814 40983
rect -26706 41017 -26654 41026
rect -26706 40983 -26697 41017
rect -26697 40983 -26663 41017
rect -26663 40983 -26654 41017
rect -26706 40974 -26654 40983
rect -26546 41017 -26494 41026
rect -26546 40983 -26537 41017
rect -26537 40983 -26503 41017
rect -26503 40983 -26494 41017
rect -26546 40974 -26494 40983
rect -26386 41017 -26334 41026
rect -26386 40983 -26377 41017
rect -26377 40983 -26343 41017
rect -26343 40983 -26334 41017
rect -26386 40974 -26334 40983
rect -26226 41017 -26174 41026
rect -26226 40983 -26217 41017
rect -26217 40983 -26183 41017
rect -26183 40983 -26174 41017
rect -26226 40974 -26174 40983
rect -26066 41017 -26014 41026
rect -26066 40983 -26057 41017
rect -26057 40983 -26023 41017
rect -26023 40983 -26014 41017
rect -26066 40974 -26014 40983
rect -25906 41017 -25854 41026
rect -25906 40983 -25897 41017
rect -25897 40983 -25863 41017
rect -25863 40983 -25854 41017
rect -25906 40974 -25854 40983
rect -25746 41017 -25694 41026
rect -25746 40983 -25737 41017
rect -25737 40983 -25703 41017
rect -25703 40983 -25694 41017
rect -25746 40974 -25694 40983
rect -25586 41017 -25534 41026
rect -25586 40983 -25577 41017
rect -25577 40983 -25543 41017
rect -25543 40983 -25534 41017
rect -25586 40974 -25534 40983
rect -25426 41017 -25374 41026
rect -25426 40983 -25417 41017
rect -25417 40983 -25383 41017
rect -25383 40983 -25374 41017
rect -25426 40974 -25374 40983
rect -25266 41017 -25214 41026
rect -25266 40983 -25257 41017
rect -25257 40983 -25223 41017
rect -25223 40983 -25214 41017
rect -25266 40974 -25214 40983
rect -25106 41017 -25054 41026
rect -25106 40983 -25097 41017
rect -25097 40983 -25063 41017
rect -25063 40983 -25054 41017
rect -25106 40974 -25054 40983
rect -24946 41017 -24894 41026
rect -24946 40983 -24937 41017
rect -24937 40983 -24903 41017
rect -24903 40983 -24894 41017
rect -24946 40974 -24894 40983
rect -24786 41017 -24734 41026
rect -24786 40983 -24777 41017
rect -24777 40983 -24743 41017
rect -24743 40983 -24734 41017
rect -24786 40974 -24734 40983
rect -24626 41017 -24574 41026
rect -24626 40983 -24617 41017
rect -24617 40983 -24583 41017
rect -24583 40983 -24574 41017
rect -24626 40974 -24574 40983
rect -24466 41017 -24414 41026
rect -24466 40983 -24457 41017
rect -24457 40983 -24423 41017
rect -24423 40983 -24414 41017
rect -24466 40974 -24414 40983
rect -24306 41017 -24254 41026
rect -24306 40983 -24297 41017
rect -24297 40983 -24263 41017
rect -24263 40983 -24254 41017
rect -24306 40974 -24254 40983
rect -24146 41017 -24094 41026
rect -24146 40983 -24137 41017
rect -24137 40983 -24103 41017
rect -24103 40983 -24094 41017
rect -24146 40974 -24094 40983
rect -23986 41017 -23934 41026
rect -23986 40983 -23977 41017
rect -23977 40983 -23943 41017
rect -23943 40983 -23934 41017
rect -23986 40974 -23934 40983
rect -23826 41017 -23774 41026
rect -23826 40983 -23817 41017
rect -23817 40983 -23783 41017
rect -23783 40983 -23774 41017
rect -23826 40974 -23774 40983
rect -23666 41017 -23614 41026
rect -23666 40983 -23657 41017
rect -23657 40983 -23623 41017
rect -23623 40983 -23614 41017
rect -23666 40974 -23614 40983
rect -23506 41017 -23454 41026
rect -23506 40983 -23497 41017
rect -23497 40983 -23463 41017
rect -23463 40983 -23454 41017
rect -23506 40974 -23454 40983
rect -23346 41017 -23294 41026
rect -23346 40983 -23337 41017
rect -23337 40983 -23303 41017
rect -23303 40983 -23294 41017
rect -23346 40974 -23294 40983
rect -23186 41017 -23134 41026
rect -23186 40983 -23177 41017
rect -23177 40983 -23143 41017
rect -23143 40983 -23134 41017
rect -23186 40974 -23134 40983
rect -23026 41017 -22974 41026
rect -23026 40983 -23017 41017
rect -23017 40983 -22983 41017
rect -22983 40983 -22974 41017
rect -23026 40974 -22974 40983
rect -22866 41017 -22814 41026
rect -22866 40983 -22857 41017
rect -22857 40983 -22823 41017
rect -22823 40983 -22814 41017
rect -22866 40974 -22814 40983
rect -22706 41017 -22654 41026
rect -22706 40983 -22697 41017
rect -22697 40983 -22663 41017
rect -22663 40983 -22654 41017
rect -22706 40974 -22654 40983
rect -22546 41017 -22494 41026
rect -22546 40983 -22537 41017
rect -22537 40983 -22503 41017
rect -22503 40983 -22494 41017
rect -22546 40974 -22494 40983
rect -22386 41017 -22334 41026
rect -22386 40983 -22377 41017
rect -22377 40983 -22343 41017
rect -22343 40983 -22334 41017
rect -22386 40974 -22334 40983
rect -22226 41017 -22174 41026
rect -22226 40983 -22217 41017
rect -22217 40983 -22183 41017
rect -22183 40983 -22174 41017
rect -22226 40974 -22174 40983
rect -22066 41017 -22014 41026
rect -22066 40983 -22057 41017
rect -22057 40983 -22023 41017
rect -22023 40983 -22014 41017
rect -22066 40974 -22014 40983
rect -21906 41017 -21854 41026
rect -21906 40983 -21897 41017
rect -21897 40983 -21863 41017
rect -21863 40983 -21854 41017
rect -21906 40974 -21854 40983
rect -21746 41017 -21694 41026
rect -21746 40983 -21737 41017
rect -21737 40983 -21703 41017
rect -21703 40983 -21694 41017
rect -21746 40974 -21694 40983
rect -21586 41017 -21534 41026
rect -21586 40983 -21577 41017
rect -21577 40983 -21543 41017
rect -21543 40983 -21534 41017
rect -21586 40974 -21534 40983
rect -21426 41017 -21374 41026
rect -21426 40983 -21417 41017
rect -21417 40983 -21383 41017
rect -21383 40983 -21374 41017
rect -21426 40974 -21374 40983
rect -21266 41017 -21214 41026
rect -21266 40983 -21257 41017
rect -21257 40983 -21223 41017
rect -21223 40983 -21214 41017
rect -21266 40974 -21214 40983
rect -21106 41017 -21054 41026
rect -21106 40983 -21097 41017
rect -21097 40983 -21063 41017
rect -21063 40983 -21054 41017
rect -21106 40974 -21054 40983
rect -20946 41017 -20894 41026
rect -20946 40983 -20937 41017
rect -20937 40983 -20903 41017
rect -20903 40983 -20894 41017
rect -20946 40974 -20894 40983
rect -20786 41017 -20734 41026
rect -20786 40983 -20777 41017
rect -20777 40983 -20743 41017
rect -20743 40983 -20734 41017
rect -20786 40974 -20734 40983
rect -20626 41017 -20574 41026
rect -20626 40983 -20617 41017
rect -20617 40983 -20583 41017
rect -20583 40983 -20574 41017
rect -20626 40974 -20574 40983
rect -20466 41017 -20414 41026
rect -20466 40983 -20457 41017
rect -20457 40983 -20423 41017
rect -20423 40983 -20414 41017
rect -20466 40974 -20414 40983
rect -20306 41017 -20254 41026
rect -20306 40983 -20297 41017
rect -20297 40983 -20263 41017
rect -20263 40983 -20254 41017
rect -20306 40974 -20254 40983
rect -20146 41017 -20094 41026
rect -20146 40983 -20137 41017
rect -20137 40983 -20103 41017
rect -20103 40983 -20094 41017
rect -20146 40974 -20094 40983
rect -19986 41017 -19934 41026
rect -19986 40983 -19977 41017
rect -19977 40983 -19943 41017
rect -19943 40983 -19934 41017
rect -19986 40974 -19934 40983
rect -19826 41017 -19774 41026
rect -19826 40983 -19817 41017
rect -19817 40983 -19783 41017
rect -19783 40983 -19774 41017
rect -19826 40974 -19774 40983
rect -19666 41017 -19614 41026
rect -19666 40983 -19657 41017
rect -19657 40983 -19623 41017
rect -19623 40983 -19614 41017
rect -19666 40974 -19614 40983
rect -19506 41017 -19454 41026
rect -19506 40983 -19497 41017
rect -19497 40983 -19463 41017
rect -19463 40983 -19454 41017
rect -19506 40974 -19454 40983
rect -19346 41017 -19294 41026
rect -19346 40983 -19337 41017
rect -19337 40983 -19303 41017
rect -19303 40983 -19294 41017
rect -19346 40974 -19294 40983
rect -19186 41017 -19134 41026
rect -19186 40983 -19177 41017
rect -19177 40983 -19143 41017
rect -19143 40983 -19134 41017
rect -19186 40974 -19134 40983
rect -19026 41017 -18974 41026
rect -19026 40983 -19017 41017
rect -19017 40983 -18983 41017
rect -18983 40983 -18974 41017
rect -19026 40974 -18974 40983
rect -18866 41017 -18814 41026
rect -18866 40983 -18857 41017
rect -18857 40983 -18823 41017
rect -18823 40983 -18814 41017
rect -18866 40974 -18814 40983
rect -18706 41017 -18654 41026
rect -18706 40983 -18697 41017
rect -18697 40983 -18663 41017
rect -18663 40983 -18654 41017
rect -18706 40974 -18654 40983
rect -18546 41017 -18494 41026
rect -18546 40983 -18537 41017
rect -18537 40983 -18503 41017
rect -18503 40983 -18494 41017
rect -18546 40974 -18494 40983
rect -18386 41017 -18334 41026
rect -18386 40983 -18377 41017
rect -18377 40983 -18343 41017
rect -18343 40983 -18334 41017
rect -18386 40974 -18334 40983
rect -18226 41017 -18174 41026
rect -18226 40983 -18217 41017
rect -18217 40983 -18183 41017
rect -18183 40983 -18174 41017
rect -18226 40974 -18174 40983
rect -18066 41017 -18014 41026
rect -18066 40983 -18057 41017
rect -18057 40983 -18023 41017
rect -18023 40983 -18014 41017
rect -18066 40974 -18014 40983
rect -17906 41017 -17854 41026
rect -17906 40983 -17897 41017
rect -17897 40983 -17863 41017
rect -17863 40983 -17854 41017
rect -17906 40974 -17854 40983
rect -17746 41017 -17694 41026
rect -17746 40983 -17737 41017
rect -17737 40983 -17703 41017
rect -17703 40983 -17694 41017
rect -17746 40974 -17694 40983
rect -17586 41017 -17534 41026
rect -17586 40983 -17577 41017
rect -17577 40983 -17543 41017
rect -17543 40983 -17534 41017
rect -17586 40974 -17534 40983
rect -17426 41017 -17374 41026
rect -17426 40983 -17417 41017
rect -17417 40983 -17383 41017
rect -17383 40983 -17374 41017
rect -17426 40974 -17374 40983
rect -17266 41017 -17214 41026
rect -17266 40983 -17257 41017
rect -17257 40983 -17223 41017
rect -17223 40983 -17214 41017
rect -17266 40974 -17214 40983
rect -17106 41017 -17054 41026
rect -17106 40983 -17097 41017
rect -17097 40983 -17063 41017
rect -17063 40983 -17054 41017
rect -17106 40974 -17054 40983
rect -16946 41017 -16894 41026
rect -16946 40983 -16937 41017
rect -16937 40983 -16903 41017
rect -16903 40983 -16894 41017
rect -16946 40974 -16894 40983
rect -16786 41017 -16734 41026
rect -16786 40983 -16777 41017
rect -16777 40983 -16743 41017
rect -16743 40983 -16734 41017
rect -16786 40974 -16734 40983
rect -16626 41017 -16574 41026
rect -16626 40983 -16617 41017
rect -16617 40983 -16583 41017
rect -16583 40983 -16574 41017
rect -16626 40974 -16574 40983
rect -16466 41017 -16414 41026
rect -16466 40983 -16457 41017
rect -16457 40983 -16423 41017
rect -16423 40983 -16414 41017
rect -16466 40974 -16414 40983
rect -16306 41017 -16254 41026
rect -16306 40983 -16297 41017
rect -16297 40983 -16263 41017
rect -16263 40983 -16254 41017
rect -16306 40974 -16254 40983
rect -16146 41017 -16094 41026
rect -16146 40983 -16137 41017
rect -16137 40983 -16103 41017
rect -16103 40983 -16094 41017
rect -16146 40974 -16094 40983
rect -15986 41017 -15934 41026
rect -15986 40983 -15977 41017
rect -15977 40983 -15943 41017
rect -15943 40983 -15934 41017
rect -15986 40974 -15934 40983
rect -15826 41017 -15774 41026
rect -15826 40983 -15817 41017
rect -15817 40983 -15783 41017
rect -15783 40983 -15774 41017
rect -15826 40974 -15774 40983
rect -15666 41017 -15614 41026
rect -15666 40983 -15657 41017
rect -15657 40983 -15623 41017
rect -15623 40983 -15614 41017
rect -15666 40974 -15614 40983
rect -15506 41017 -15454 41026
rect -15506 40983 -15497 41017
rect -15497 40983 -15463 41017
rect -15463 40983 -15454 41017
rect -15506 40974 -15454 40983
rect -15346 41017 -15294 41026
rect -15346 40983 -15337 41017
rect -15337 40983 -15303 41017
rect -15303 40983 -15294 41017
rect -15346 40974 -15294 40983
rect -15186 41017 -15134 41026
rect -15186 40983 -15177 41017
rect -15177 40983 -15143 41017
rect -15143 40983 -15134 41017
rect -15186 40974 -15134 40983
rect -15026 41017 -14974 41026
rect -15026 40983 -15017 41017
rect -15017 40983 -14983 41017
rect -14983 40983 -14974 41017
rect -15026 40974 -14974 40983
rect -14866 41017 -14814 41026
rect -14866 40983 -14857 41017
rect -14857 40983 -14823 41017
rect -14823 40983 -14814 41017
rect -14866 40974 -14814 40983
rect -14706 41017 -14654 41026
rect -14706 40983 -14697 41017
rect -14697 40983 -14663 41017
rect -14663 40983 -14654 41017
rect -14706 40974 -14654 40983
rect -14546 41017 -14494 41026
rect -14546 40983 -14537 41017
rect -14537 40983 -14503 41017
rect -14503 40983 -14494 41017
rect -14546 40974 -14494 40983
rect -14386 41017 -14334 41026
rect -14386 40983 -14377 41017
rect -14377 40983 -14343 41017
rect -14343 40983 -14334 41017
rect -14386 40974 -14334 40983
rect -14226 41017 -14174 41026
rect -14226 40983 -14217 41017
rect -14217 40983 -14183 41017
rect -14183 40983 -14174 41017
rect -14226 40974 -14174 40983
rect -14066 41017 -14014 41026
rect -14066 40983 -14057 41017
rect -14057 40983 -14023 41017
rect -14023 40983 -14014 41017
rect -14066 40974 -14014 40983
rect -13906 41017 -13854 41026
rect -13906 40983 -13897 41017
rect -13897 40983 -13863 41017
rect -13863 40983 -13854 41017
rect -13906 40974 -13854 40983
rect -13746 41017 -13694 41026
rect -13746 40983 -13737 41017
rect -13737 40983 -13703 41017
rect -13703 40983 -13694 41017
rect -13746 40974 -13694 40983
rect -13586 41017 -13534 41026
rect -13586 40983 -13577 41017
rect -13577 40983 -13543 41017
rect -13543 40983 -13534 41017
rect -13586 40974 -13534 40983
rect -13426 41017 -13374 41026
rect -13426 40983 -13417 41017
rect -13417 40983 -13383 41017
rect -13383 40983 -13374 41017
rect -13426 40974 -13374 40983
rect -13266 41017 -13214 41026
rect -13266 40983 -13257 41017
rect -13257 40983 -13223 41017
rect -13223 40983 -13214 41017
rect -13266 40974 -13214 40983
rect -13106 41017 -13054 41026
rect -13106 40983 -13097 41017
rect -13097 40983 -13063 41017
rect -13063 40983 -13054 41017
rect -13106 40974 -13054 40983
rect -12946 41017 -12894 41026
rect -12946 40983 -12937 41017
rect -12937 40983 -12903 41017
rect -12903 40983 -12894 41017
rect -12946 40974 -12894 40983
rect -12786 41017 -12734 41026
rect -12786 40983 -12777 41017
rect -12777 40983 -12743 41017
rect -12743 40983 -12734 41017
rect -12786 40974 -12734 40983
rect -12626 41017 -12574 41026
rect -12626 40983 -12617 41017
rect -12617 40983 -12583 41017
rect -12583 40983 -12574 41017
rect -12626 40974 -12574 40983
rect -12466 41017 -12414 41026
rect -12466 40983 -12457 41017
rect -12457 40983 -12423 41017
rect -12423 40983 -12414 41017
rect -12466 40974 -12414 40983
rect -12306 41017 -12254 41026
rect -12306 40983 -12297 41017
rect -12297 40983 -12263 41017
rect -12263 40983 -12254 41017
rect -12306 40974 -12254 40983
rect -11346 41017 -11294 41026
rect -11346 40983 -11337 41017
rect -11337 40983 -11303 41017
rect -11303 40983 -11294 41017
rect -11346 40974 -11294 40983
rect -11186 41017 -11134 41026
rect -11186 40983 -11177 41017
rect -11177 40983 -11143 41017
rect -11143 40983 -11134 41017
rect -11186 40974 -11134 40983
rect -11026 41017 -10974 41026
rect -11026 40983 -11017 41017
rect -11017 40983 -10983 41017
rect -10983 40983 -10974 41017
rect -11026 40974 -10974 40983
rect -10866 41017 -10814 41026
rect -10866 40983 -10857 41017
rect -10857 40983 -10823 41017
rect -10823 40983 -10814 41017
rect -10866 40974 -10814 40983
rect -10706 41017 -10654 41026
rect -10706 40983 -10697 41017
rect -10697 40983 -10663 41017
rect -10663 40983 -10654 41017
rect -10706 40974 -10654 40983
rect -10546 41017 -10494 41026
rect -10546 40983 -10537 41017
rect -10537 40983 -10503 41017
rect -10503 40983 -10494 41017
rect -10546 40974 -10494 40983
rect -10386 41017 -10334 41026
rect -10386 40983 -10377 41017
rect -10377 40983 -10343 41017
rect -10343 40983 -10334 41017
rect -10386 40974 -10334 40983
rect -10226 41017 -10174 41026
rect -10226 40983 -10217 41017
rect -10217 40983 -10183 41017
rect -10183 40983 -10174 41017
rect -10226 40974 -10174 40983
rect -10066 41017 -10014 41026
rect -10066 40983 -10057 41017
rect -10057 40983 -10023 41017
rect -10023 40983 -10014 41017
rect -10066 40974 -10014 40983
rect -9906 41017 -9854 41026
rect -9906 40983 -9897 41017
rect -9897 40983 -9863 41017
rect -9863 40983 -9854 41017
rect -9906 40974 -9854 40983
rect -9746 41017 -9694 41026
rect -9746 40983 -9737 41017
rect -9737 40983 -9703 41017
rect -9703 40983 -9694 41017
rect -9746 40974 -9694 40983
rect -9586 41017 -9534 41026
rect -9586 40983 -9577 41017
rect -9577 40983 -9543 41017
rect -9543 40983 -9534 41017
rect -9586 40974 -9534 40983
rect -9426 41017 -9374 41026
rect -9426 40983 -9417 41017
rect -9417 40983 -9383 41017
rect -9383 40983 -9374 41017
rect -9426 40974 -9374 40983
rect -9266 41017 -9214 41026
rect -9266 40983 -9257 41017
rect -9257 40983 -9223 41017
rect -9223 40983 -9214 41017
rect -9266 40974 -9214 40983
rect -9106 41017 -9054 41026
rect -9106 40983 -9097 41017
rect -9097 40983 -9063 41017
rect -9063 40983 -9054 41017
rect -9106 40974 -9054 40983
rect -8946 41017 -8894 41026
rect -8946 40983 -8937 41017
rect -8937 40983 -8903 41017
rect -8903 40983 -8894 41017
rect -8946 40974 -8894 40983
rect -8786 41017 -8734 41026
rect -8786 40983 -8777 41017
rect -8777 40983 -8743 41017
rect -8743 40983 -8734 41017
rect -8786 40974 -8734 40983
rect -8626 41017 -8574 41026
rect -8626 40983 -8617 41017
rect -8617 40983 -8583 41017
rect -8583 40983 -8574 41017
rect -8626 40974 -8574 40983
rect -8466 41017 -8414 41026
rect -8466 40983 -8457 41017
rect -8457 40983 -8423 41017
rect -8423 40983 -8414 41017
rect -8466 40974 -8414 40983
rect -8306 41017 -8254 41026
rect -8306 40983 -8297 41017
rect -8297 40983 -8263 41017
rect -8263 40983 -8254 41017
rect -8306 40974 -8254 40983
rect -8146 41017 -8094 41026
rect -8146 40983 -8137 41017
rect -8137 40983 -8103 41017
rect -8103 40983 -8094 41017
rect -8146 40974 -8094 40983
rect -7986 41017 -7934 41026
rect -7986 40983 -7977 41017
rect -7977 40983 -7943 41017
rect -7943 40983 -7934 41017
rect -7986 40974 -7934 40983
rect -7826 41017 -7774 41026
rect -7826 40983 -7817 41017
rect -7817 40983 -7783 41017
rect -7783 40983 -7774 41017
rect -7826 40974 -7774 40983
rect -7666 41017 -7614 41026
rect -7666 40983 -7657 41017
rect -7657 40983 -7623 41017
rect -7623 40983 -7614 41017
rect -7666 40974 -7614 40983
rect -7506 41017 -7454 41026
rect -7506 40983 -7497 41017
rect -7497 40983 -7463 41017
rect -7463 40983 -7454 41017
rect -7506 40974 -7454 40983
rect -7346 41017 -7294 41026
rect -7346 40983 -7337 41017
rect -7337 40983 -7303 41017
rect -7303 40983 -7294 41017
rect -7346 40974 -7294 40983
rect -7186 41017 -7134 41026
rect -7186 40983 -7177 41017
rect -7177 40983 -7143 41017
rect -7143 40983 -7134 41017
rect -7186 40974 -7134 40983
rect -7026 41017 -6974 41026
rect -7026 40983 -7017 41017
rect -7017 40983 -6983 41017
rect -6983 40983 -6974 41017
rect -7026 40974 -6974 40983
rect -6866 41017 -6814 41026
rect -6866 40983 -6857 41017
rect -6857 40983 -6823 41017
rect -6823 40983 -6814 41017
rect -6866 40974 -6814 40983
rect -6706 41017 -6654 41026
rect -6706 40983 -6697 41017
rect -6697 40983 -6663 41017
rect -6663 40983 -6654 41017
rect -6706 40974 -6654 40983
rect -6546 41017 -6494 41026
rect -6546 40983 -6537 41017
rect -6537 40983 -6503 41017
rect -6503 40983 -6494 41017
rect -6546 40974 -6494 40983
rect -6386 41017 -6334 41026
rect -6386 40983 -6377 41017
rect -6377 40983 -6343 41017
rect -6343 40983 -6334 41017
rect -6386 40974 -6334 40983
rect -6226 41017 -6174 41026
rect -6226 40983 -6217 41017
rect -6217 40983 -6183 41017
rect -6183 40983 -6174 41017
rect -6226 40974 -6174 40983
rect -6066 41017 -6014 41026
rect -6066 40983 -6057 41017
rect -6057 40983 -6023 41017
rect -6023 40983 -6014 41017
rect -6066 40974 -6014 40983
rect -5906 41017 -5854 41026
rect -5906 40983 -5897 41017
rect -5897 40983 -5863 41017
rect -5863 40983 -5854 41017
rect -5906 40974 -5854 40983
rect -5746 41017 -5694 41026
rect -5746 40983 -5737 41017
rect -5737 40983 -5703 41017
rect -5703 40983 -5694 41017
rect -5746 40974 -5694 40983
rect -5586 41017 -5534 41026
rect -5586 40983 -5577 41017
rect -5577 40983 -5543 41017
rect -5543 40983 -5534 41017
rect -5586 40974 -5534 40983
rect -5426 41017 -5374 41026
rect -5426 40983 -5417 41017
rect -5417 40983 -5383 41017
rect -5383 40983 -5374 41017
rect -5426 40974 -5374 40983
rect -5266 41017 -5214 41026
rect -5266 40983 -5257 41017
rect -5257 40983 -5223 41017
rect -5223 40983 -5214 41017
rect -5266 40974 -5214 40983
rect -5106 41017 -5054 41026
rect -5106 40983 -5097 41017
rect -5097 40983 -5063 41017
rect -5063 40983 -5054 41017
rect -5106 40974 -5054 40983
rect -4946 41017 -4894 41026
rect -4946 40983 -4937 41017
rect -4937 40983 -4903 41017
rect -4903 40983 -4894 41017
rect -4946 40974 -4894 40983
rect -4786 41017 -4734 41026
rect -4786 40983 -4777 41017
rect -4777 40983 -4743 41017
rect -4743 40983 -4734 41017
rect -4786 40974 -4734 40983
rect -4626 41017 -4574 41026
rect -4626 40983 -4617 41017
rect -4617 40983 -4583 41017
rect -4583 40983 -4574 41017
rect -4626 40974 -4574 40983
rect -4466 41017 -4414 41026
rect -4466 40983 -4457 41017
rect -4457 40983 -4423 41017
rect -4423 40983 -4414 41017
rect -4466 40974 -4414 40983
rect -4306 41017 -4254 41026
rect -4306 40983 -4297 41017
rect -4297 40983 -4263 41017
rect -4263 40983 -4254 41017
rect -4306 40974 -4254 40983
rect -4146 41017 -4094 41026
rect -4146 40983 -4137 41017
rect -4137 40983 -4103 41017
rect -4103 40983 -4094 41017
rect -4146 40974 -4094 40983
rect -3986 41017 -3934 41026
rect -3986 40983 -3977 41017
rect -3977 40983 -3943 41017
rect -3943 40983 -3934 41017
rect -3986 40974 -3934 40983
rect -3666 41017 -3614 41026
rect -3666 40983 -3657 41017
rect -3657 40983 -3623 41017
rect -3623 40983 -3614 41017
rect -3666 40974 -3614 40983
rect -3506 41017 -3454 41026
rect -3506 40983 -3497 41017
rect -3497 40983 -3463 41017
rect -3463 40983 -3454 41017
rect -3506 40974 -3454 40983
rect 41054 41017 41106 41026
rect 41054 40983 41063 41017
rect 41063 40983 41097 41017
rect 41097 40983 41106 41017
rect 41054 40974 41106 40983
rect 41214 41017 41266 41026
rect 41214 40983 41223 41017
rect 41223 40983 41257 41017
rect 41257 40983 41266 41017
rect 41214 40974 41266 40983
rect 41374 41017 41426 41026
rect 41374 40983 41383 41017
rect 41383 40983 41417 41017
rect 41417 40983 41426 41017
rect 41374 40974 41426 40983
rect 41534 41017 41586 41026
rect 41534 40983 41543 41017
rect 41543 40983 41577 41017
rect 41577 40983 41586 41017
rect 41534 40974 41586 40983
rect 41694 41017 41746 41026
rect 41694 40983 41703 41017
rect 41703 40983 41737 41017
rect 41737 40983 41746 41017
rect 41694 40974 41746 40983
rect 41854 41017 41906 41026
rect 41854 40983 41863 41017
rect 41863 40983 41897 41017
rect 41897 40983 41906 41017
rect 41854 40974 41906 40983
rect 42014 41017 42066 41026
rect 42014 40983 42023 41017
rect 42023 40983 42057 41017
rect 42057 40983 42066 41017
rect 42014 40974 42066 40983
rect 42174 41017 42226 41026
rect 42174 40983 42183 41017
rect 42183 40983 42217 41017
rect 42217 40983 42226 41017
rect 42174 40974 42226 40983
rect 42334 41017 42386 41026
rect 42334 40983 42343 41017
rect 42343 40983 42377 41017
rect 42377 40983 42386 41017
rect 42334 40974 42386 40983
rect 42494 41017 42546 41026
rect 42494 40983 42503 41017
rect 42503 40983 42537 41017
rect 42537 40983 42546 41017
rect 42494 40974 42546 40983
rect 42654 41017 42706 41026
rect 42654 40983 42663 41017
rect 42663 40983 42697 41017
rect 42697 40983 42706 41017
rect 42654 40974 42706 40983
rect 42814 41017 42866 41026
rect 42814 40983 42823 41017
rect 42823 40983 42857 41017
rect 42857 40983 42866 41017
rect 42814 40974 42866 40983
rect 42974 41017 43026 41026
rect 42974 40983 42983 41017
rect 42983 40983 43017 41017
rect 43017 40983 43026 41017
rect 42974 40974 43026 40983
rect 43134 41017 43186 41026
rect 43134 40983 43143 41017
rect 43143 40983 43177 41017
rect 43177 40983 43186 41017
rect 43134 40974 43186 40983
rect -10546 40697 -10494 40706
rect -10546 40663 -10537 40697
rect -10537 40663 -10503 40697
rect -10503 40663 -10494 40697
rect -10546 40654 -10494 40663
rect -10226 40697 -10174 40706
rect -10226 40663 -10217 40697
rect -10217 40663 -10183 40697
rect -10183 40663 -10174 40697
rect -10226 40654 -10174 40663
rect -10066 40697 -10014 40706
rect -10066 40663 -10057 40697
rect -10057 40663 -10023 40697
rect -10023 40663 -10014 40697
rect -10066 40654 -10014 40663
rect -9906 40697 -9854 40706
rect -9906 40663 -9897 40697
rect -9897 40663 -9863 40697
rect -9863 40663 -9854 40697
rect -9906 40654 -9854 40663
rect -9746 40697 -9694 40706
rect -9746 40663 -9737 40697
rect -9737 40663 -9703 40697
rect -9703 40663 -9694 40697
rect -9746 40654 -9694 40663
rect -9586 40697 -9534 40706
rect -9586 40663 -9577 40697
rect -9577 40663 -9543 40697
rect -9543 40663 -9534 40697
rect -9586 40654 -9534 40663
rect -9426 40697 -9374 40706
rect -9426 40663 -9417 40697
rect -9417 40663 -9383 40697
rect -9383 40663 -9374 40697
rect -9426 40654 -9374 40663
rect -9266 40697 -9214 40706
rect -9266 40663 -9257 40697
rect -9257 40663 -9223 40697
rect -9223 40663 -9214 40697
rect -9266 40654 -9214 40663
rect -9106 40697 -9054 40706
rect -9106 40663 -9097 40697
rect -9097 40663 -9063 40697
rect -9063 40663 -9054 40697
rect -9106 40654 -9054 40663
rect -8946 40697 -8894 40706
rect -8946 40663 -8937 40697
rect -8937 40663 -8903 40697
rect -8903 40663 -8894 40697
rect -8946 40654 -8894 40663
rect -8786 40697 -8734 40706
rect -8786 40663 -8777 40697
rect -8777 40663 -8743 40697
rect -8743 40663 -8734 40697
rect -8786 40654 -8734 40663
rect -8626 40697 -8574 40706
rect -8626 40663 -8617 40697
rect -8617 40663 -8583 40697
rect -8583 40663 -8574 40697
rect -8626 40654 -8574 40663
rect -8466 40697 -8414 40706
rect -8466 40663 -8457 40697
rect -8457 40663 -8423 40697
rect -8423 40663 -8414 40697
rect -8466 40654 -8414 40663
rect -8306 40697 -8254 40706
rect -8306 40663 -8297 40697
rect -8297 40663 -8263 40697
rect -8263 40663 -8254 40697
rect -8306 40654 -8254 40663
rect -8146 40697 -8094 40706
rect -8146 40663 -8137 40697
rect -8137 40663 -8103 40697
rect -8103 40663 -8094 40697
rect -8146 40654 -8094 40663
rect -7986 40697 -7934 40706
rect -7986 40663 -7977 40697
rect -7977 40663 -7943 40697
rect -7943 40663 -7934 40697
rect -7986 40654 -7934 40663
rect -7826 40697 -7774 40706
rect -7826 40663 -7817 40697
rect -7817 40663 -7783 40697
rect -7783 40663 -7774 40697
rect -7826 40654 -7774 40663
rect -7666 40697 -7614 40706
rect -7666 40663 -7657 40697
rect -7657 40663 -7623 40697
rect -7623 40663 -7614 40697
rect -7666 40654 -7614 40663
rect -7506 40697 -7454 40706
rect -7506 40663 -7497 40697
rect -7497 40663 -7463 40697
rect -7463 40663 -7454 40697
rect -7506 40654 -7454 40663
rect -7346 40697 -7294 40706
rect -7346 40663 -7337 40697
rect -7337 40663 -7303 40697
rect -7303 40663 -7294 40697
rect -7346 40654 -7294 40663
rect -7186 40697 -7134 40706
rect -7186 40663 -7177 40697
rect -7177 40663 -7143 40697
rect -7143 40663 -7134 40697
rect -7186 40654 -7134 40663
rect -7026 40697 -6974 40706
rect -7026 40663 -7017 40697
rect -7017 40663 -6983 40697
rect -6983 40663 -6974 40697
rect -7026 40654 -6974 40663
rect -6866 40697 -6814 40706
rect -6866 40663 -6857 40697
rect -6857 40663 -6823 40697
rect -6823 40663 -6814 40697
rect -6866 40654 -6814 40663
rect -6706 40697 -6654 40706
rect -6706 40663 -6697 40697
rect -6697 40663 -6663 40697
rect -6663 40663 -6654 40697
rect -6706 40654 -6654 40663
rect -6546 40697 -6494 40706
rect -6546 40663 -6537 40697
rect -6537 40663 -6503 40697
rect -6503 40663 -6494 40697
rect -6546 40654 -6494 40663
rect -6386 40697 -6334 40706
rect -6386 40663 -6377 40697
rect -6377 40663 -6343 40697
rect -6343 40663 -6334 40697
rect -6386 40654 -6334 40663
rect -6226 40697 -6174 40706
rect -6226 40663 -6217 40697
rect -6217 40663 -6183 40697
rect -6183 40663 -6174 40697
rect -6226 40654 -6174 40663
rect -6066 40697 -6014 40706
rect -6066 40663 -6057 40697
rect -6057 40663 -6023 40697
rect -6023 40663 -6014 40697
rect -6066 40654 -6014 40663
rect -5906 40697 -5854 40706
rect -5906 40663 -5897 40697
rect -5897 40663 -5863 40697
rect -5863 40663 -5854 40697
rect -5906 40654 -5854 40663
rect -5746 40697 -5694 40706
rect -5746 40663 -5737 40697
rect -5737 40663 -5703 40697
rect -5703 40663 -5694 40697
rect -5746 40654 -5694 40663
rect -5586 40697 -5534 40706
rect -5586 40663 -5577 40697
rect -5577 40663 -5543 40697
rect -5543 40663 -5534 40697
rect -5586 40654 -5534 40663
rect -5426 40697 -5374 40706
rect -5426 40663 -5417 40697
rect -5417 40663 -5383 40697
rect -5383 40663 -5374 40697
rect -5426 40654 -5374 40663
rect -5266 40697 -5214 40706
rect -5266 40663 -5257 40697
rect -5257 40663 -5223 40697
rect -5223 40663 -5214 40697
rect -5266 40654 -5214 40663
rect -5106 40697 -5054 40706
rect -5106 40663 -5097 40697
rect -5097 40663 -5063 40697
rect -5063 40663 -5054 40697
rect -5106 40654 -5054 40663
rect -4946 40697 -4894 40706
rect -4946 40663 -4937 40697
rect -4937 40663 -4903 40697
rect -4903 40663 -4894 40697
rect -4946 40654 -4894 40663
rect -4786 40697 -4734 40706
rect -4786 40663 -4777 40697
rect -4777 40663 -4743 40697
rect -4743 40663 -4734 40697
rect -4786 40654 -4734 40663
rect -4626 40697 -4574 40706
rect -4626 40663 -4617 40697
rect -4617 40663 -4583 40697
rect -4583 40663 -4574 40697
rect -4626 40654 -4574 40663
rect -4466 40697 -4414 40706
rect -4466 40663 -4457 40697
rect -4457 40663 -4423 40697
rect -4423 40663 -4414 40697
rect -4466 40654 -4414 40663
rect -4306 40697 -4254 40706
rect -4306 40663 -4297 40697
rect -4297 40663 -4263 40697
rect -4263 40663 -4254 40697
rect -4306 40654 -4254 40663
rect -4146 40697 -4094 40706
rect -4146 40663 -4137 40697
rect -4137 40663 -4103 40697
rect -4103 40663 -4094 40697
rect -4146 40654 -4094 40663
rect -3986 40697 -3934 40706
rect -3986 40663 -3977 40697
rect -3977 40663 -3943 40697
rect -3943 40663 -3934 40697
rect -3986 40654 -3934 40663
rect -3666 40697 -3614 40706
rect -3666 40663 -3657 40697
rect -3657 40663 -3623 40697
rect -3623 40663 -3614 40697
rect -3666 40654 -3614 40663
rect -3506 40697 -3454 40706
rect -3506 40663 -3497 40697
rect -3497 40663 -3463 40697
rect -3463 40663 -3454 40697
rect -3506 40654 -3454 40663
rect -10546 40377 -10494 40386
rect -10546 40343 -10537 40377
rect -10537 40343 -10503 40377
rect -10503 40343 -10494 40377
rect -10546 40334 -10494 40343
rect -10226 40377 -10174 40386
rect -10226 40343 -10217 40377
rect -10217 40343 -10183 40377
rect -10183 40343 -10174 40377
rect -10226 40334 -10174 40343
rect -10066 40377 -10014 40386
rect -10066 40343 -10057 40377
rect -10057 40343 -10023 40377
rect -10023 40343 -10014 40377
rect -10066 40334 -10014 40343
rect -9906 40377 -9854 40386
rect -9906 40343 -9897 40377
rect -9897 40343 -9863 40377
rect -9863 40343 -9854 40377
rect -9906 40334 -9854 40343
rect -9746 40377 -9694 40386
rect -9746 40343 -9737 40377
rect -9737 40343 -9703 40377
rect -9703 40343 -9694 40377
rect -9746 40334 -9694 40343
rect -9586 40377 -9534 40386
rect -9586 40343 -9577 40377
rect -9577 40343 -9543 40377
rect -9543 40343 -9534 40377
rect -9586 40334 -9534 40343
rect -9426 40377 -9374 40386
rect -9426 40343 -9417 40377
rect -9417 40343 -9383 40377
rect -9383 40343 -9374 40377
rect -9426 40334 -9374 40343
rect -9266 40377 -9214 40386
rect -9266 40343 -9257 40377
rect -9257 40343 -9223 40377
rect -9223 40343 -9214 40377
rect -9266 40334 -9214 40343
rect -9106 40377 -9054 40386
rect -9106 40343 -9097 40377
rect -9097 40343 -9063 40377
rect -9063 40343 -9054 40377
rect -9106 40334 -9054 40343
rect -8946 40377 -8894 40386
rect -8946 40343 -8937 40377
rect -8937 40343 -8903 40377
rect -8903 40343 -8894 40377
rect -8946 40334 -8894 40343
rect -8786 40377 -8734 40386
rect -8786 40343 -8777 40377
rect -8777 40343 -8743 40377
rect -8743 40343 -8734 40377
rect -8786 40334 -8734 40343
rect -8626 40377 -8574 40386
rect -8626 40343 -8617 40377
rect -8617 40343 -8583 40377
rect -8583 40343 -8574 40377
rect -8626 40334 -8574 40343
rect -8466 40377 -8414 40386
rect -8466 40343 -8457 40377
rect -8457 40343 -8423 40377
rect -8423 40343 -8414 40377
rect -8466 40334 -8414 40343
rect -8306 40377 -8254 40386
rect -8306 40343 -8297 40377
rect -8297 40343 -8263 40377
rect -8263 40343 -8254 40377
rect -8306 40334 -8254 40343
rect -8146 40377 -8094 40386
rect -8146 40343 -8137 40377
rect -8137 40343 -8103 40377
rect -8103 40343 -8094 40377
rect -8146 40334 -8094 40343
rect -7986 40377 -7934 40386
rect -7986 40343 -7977 40377
rect -7977 40343 -7943 40377
rect -7943 40343 -7934 40377
rect -7986 40334 -7934 40343
rect -7826 40377 -7774 40386
rect -7826 40343 -7817 40377
rect -7817 40343 -7783 40377
rect -7783 40343 -7774 40377
rect -7826 40334 -7774 40343
rect -7666 40377 -7614 40386
rect -7666 40343 -7657 40377
rect -7657 40343 -7623 40377
rect -7623 40343 -7614 40377
rect -7666 40334 -7614 40343
rect -7506 40377 -7454 40386
rect -7506 40343 -7497 40377
rect -7497 40343 -7463 40377
rect -7463 40343 -7454 40377
rect -7506 40334 -7454 40343
rect -7346 40377 -7294 40386
rect -7346 40343 -7337 40377
rect -7337 40343 -7303 40377
rect -7303 40343 -7294 40377
rect -7346 40334 -7294 40343
rect -7186 40377 -7134 40386
rect -7186 40343 -7177 40377
rect -7177 40343 -7143 40377
rect -7143 40343 -7134 40377
rect -7186 40334 -7134 40343
rect -7026 40377 -6974 40386
rect -7026 40343 -7017 40377
rect -7017 40343 -6983 40377
rect -6983 40343 -6974 40377
rect -7026 40334 -6974 40343
rect -6866 40377 -6814 40386
rect -6866 40343 -6857 40377
rect -6857 40343 -6823 40377
rect -6823 40343 -6814 40377
rect -6866 40334 -6814 40343
rect -6706 40377 -6654 40386
rect -6706 40343 -6697 40377
rect -6697 40343 -6663 40377
rect -6663 40343 -6654 40377
rect -6706 40334 -6654 40343
rect -6546 40377 -6494 40386
rect -6546 40343 -6537 40377
rect -6537 40343 -6503 40377
rect -6503 40343 -6494 40377
rect -6546 40334 -6494 40343
rect -6386 40377 -6334 40386
rect -6386 40343 -6377 40377
rect -6377 40343 -6343 40377
rect -6343 40343 -6334 40377
rect -6386 40334 -6334 40343
rect -6226 40377 -6174 40386
rect -6226 40343 -6217 40377
rect -6217 40343 -6183 40377
rect -6183 40343 -6174 40377
rect -6226 40334 -6174 40343
rect -6066 40377 -6014 40386
rect -6066 40343 -6057 40377
rect -6057 40343 -6023 40377
rect -6023 40343 -6014 40377
rect -6066 40334 -6014 40343
rect -5906 40377 -5854 40386
rect -5906 40343 -5897 40377
rect -5897 40343 -5863 40377
rect -5863 40343 -5854 40377
rect -5906 40334 -5854 40343
rect -5746 40377 -5694 40386
rect -5746 40343 -5737 40377
rect -5737 40343 -5703 40377
rect -5703 40343 -5694 40377
rect -5746 40334 -5694 40343
rect -5586 40377 -5534 40386
rect -5586 40343 -5577 40377
rect -5577 40343 -5543 40377
rect -5543 40343 -5534 40377
rect -5586 40334 -5534 40343
rect -5426 40377 -5374 40386
rect -5426 40343 -5417 40377
rect -5417 40343 -5383 40377
rect -5383 40343 -5374 40377
rect -5426 40334 -5374 40343
rect -5266 40377 -5214 40386
rect -5266 40343 -5257 40377
rect -5257 40343 -5223 40377
rect -5223 40343 -5214 40377
rect -5266 40334 -5214 40343
rect -5106 40377 -5054 40386
rect -5106 40343 -5097 40377
rect -5097 40343 -5063 40377
rect -5063 40343 -5054 40377
rect -5106 40334 -5054 40343
rect -4946 40377 -4894 40386
rect -4946 40343 -4937 40377
rect -4937 40343 -4903 40377
rect -4903 40343 -4894 40377
rect -4946 40334 -4894 40343
rect -4786 40377 -4734 40386
rect -4786 40343 -4777 40377
rect -4777 40343 -4743 40377
rect -4743 40343 -4734 40377
rect -4786 40334 -4734 40343
rect -4626 40377 -4574 40386
rect -4626 40343 -4617 40377
rect -4617 40343 -4583 40377
rect -4583 40343 -4574 40377
rect -4626 40334 -4574 40343
rect -4466 40377 -4414 40386
rect -4466 40343 -4457 40377
rect -4457 40343 -4423 40377
rect -4423 40343 -4414 40377
rect -4466 40334 -4414 40343
rect -4306 40377 -4254 40386
rect -4306 40343 -4297 40377
rect -4297 40343 -4263 40377
rect -4263 40343 -4254 40377
rect -4306 40334 -4254 40343
rect -4146 40377 -4094 40386
rect -4146 40343 -4137 40377
rect -4137 40343 -4103 40377
rect -4103 40343 -4094 40377
rect -4146 40334 -4094 40343
rect -3986 40377 -3934 40386
rect -3986 40343 -3977 40377
rect -3977 40343 -3943 40377
rect -3943 40343 -3934 40377
rect -3986 40334 -3934 40343
rect -3666 40377 -3614 40386
rect -3666 40343 -3657 40377
rect -3657 40343 -3623 40377
rect -3623 40343 -3614 40377
rect -3666 40334 -3614 40343
rect -3506 40377 -3454 40386
rect -3506 40343 -3497 40377
rect -3497 40343 -3463 40377
rect -3463 40343 -3454 40377
rect -3506 40334 -3454 40343
rect 41054 40057 41106 40066
rect 41054 40023 41063 40057
rect 41063 40023 41097 40057
rect 41097 40023 41106 40057
rect 41054 40014 41106 40023
rect 41214 40057 41266 40066
rect 41214 40023 41223 40057
rect 41223 40023 41257 40057
rect 41257 40023 41266 40057
rect 41214 40014 41266 40023
rect 41374 40057 41426 40066
rect 41374 40023 41383 40057
rect 41383 40023 41417 40057
rect 41417 40023 41426 40057
rect 41374 40014 41426 40023
rect 41534 40057 41586 40066
rect 41534 40023 41543 40057
rect 41543 40023 41577 40057
rect 41577 40023 41586 40057
rect 41534 40014 41586 40023
rect 41694 40057 41746 40066
rect 41694 40023 41703 40057
rect 41703 40023 41737 40057
rect 41737 40023 41746 40057
rect 41694 40014 41746 40023
rect 41854 40057 41906 40066
rect 41854 40023 41863 40057
rect 41863 40023 41897 40057
rect 41897 40023 41906 40057
rect 41854 40014 41906 40023
rect 42014 40057 42066 40066
rect 42014 40023 42023 40057
rect 42023 40023 42057 40057
rect 42057 40023 42066 40057
rect 42014 40014 42066 40023
rect 42174 40057 42226 40066
rect 42174 40023 42183 40057
rect 42183 40023 42217 40057
rect 42217 40023 42226 40057
rect 42174 40014 42226 40023
rect 42334 40057 42386 40066
rect 42334 40023 42343 40057
rect 42343 40023 42377 40057
rect 42377 40023 42386 40057
rect 42334 40014 42386 40023
rect 42494 40057 42546 40066
rect 42494 40023 42503 40057
rect 42503 40023 42537 40057
rect 42537 40023 42546 40057
rect 42494 40014 42546 40023
rect 42654 40057 42706 40066
rect 42654 40023 42663 40057
rect 42663 40023 42697 40057
rect 42697 40023 42706 40057
rect 42654 40014 42706 40023
rect 42814 40057 42866 40066
rect 42814 40023 42823 40057
rect 42823 40023 42857 40057
rect 42857 40023 42866 40057
rect 42814 40014 42866 40023
rect 42974 40057 43026 40066
rect 42974 40023 42983 40057
rect 42983 40023 43017 40057
rect 43017 40023 43026 40057
rect 42974 40014 43026 40023
rect 43134 40057 43186 40066
rect 43134 40023 43143 40057
rect 43143 40023 43177 40057
rect 43177 40023 43186 40057
rect 43134 40014 43186 40023
rect 41054 39737 41106 39746
rect 41054 39703 41063 39737
rect 41063 39703 41097 39737
rect 41097 39703 41106 39737
rect 41054 39694 41106 39703
rect 41214 39737 41266 39746
rect 41214 39703 41223 39737
rect 41223 39703 41257 39737
rect 41257 39703 41266 39737
rect 41214 39694 41266 39703
rect 41374 39737 41426 39746
rect 41374 39703 41383 39737
rect 41383 39703 41417 39737
rect 41417 39703 41426 39737
rect 41374 39694 41426 39703
rect 41534 39737 41586 39746
rect 41534 39703 41543 39737
rect 41543 39703 41577 39737
rect 41577 39703 41586 39737
rect 41534 39694 41586 39703
rect 41694 39737 41746 39746
rect 41694 39703 41703 39737
rect 41703 39703 41737 39737
rect 41737 39703 41746 39737
rect 41694 39694 41746 39703
rect 41854 39737 41906 39746
rect 41854 39703 41863 39737
rect 41863 39703 41897 39737
rect 41897 39703 41906 39737
rect 41854 39694 41906 39703
rect 42014 39737 42066 39746
rect 42014 39703 42023 39737
rect 42023 39703 42057 39737
rect 42057 39703 42066 39737
rect 42014 39694 42066 39703
rect 42174 39737 42226 39746
rect 42174 39703 42183 39737
rect 42183 39703 42217 39737
rect 42217 39703 42226 39737
rect 42174 39694 42226 39703
rect 42334 39737 42386 39746
rect 42334 39703 42343 39737
rect 42343 39703 42377 39737
rect 42377 39703 42386 39737
rect 42334 39694 42386 39703
rect 42494 39737 42546 39746
rect 42494 39703 42503 39737
rect 42503 39703 42537 39737
rect 42537 39703 42546 39737
rect 42494 39694 42546 39703
rect 42654 39737 42706 39746
rect 42654 39703 42663 39737
rect 42663 39703 42697 39737
rect 42697 39703 42706 39737
rect 42654 39694 42706 39703
rect 42814 39737 42866 39746
rect 42814 39703 42823 39737
rect 42823 39703 42857 39737
rect 42857 39703 42866 39737
rect 42814 39694 42866 39703
rect 42974 39737 43026 39746
rect 42974 39703 42983 39737
rect 42983 39703 43017 39737
rect 43017 39703 43026 39737
rect 42974 39694 43026 39703
rect 43134 39737 43186 39746
rect 43134 39703 43143 39737
rect 43143 39703 43177 39737
rect 43177 39703 43186 39737
rect 43134 39694 43186 39703
rect -33106 37737 -33054 37746
rect -33106 37703 -33097 37737
rect -33097 37703 -33063 37737
rect -33063 37703 -33054 37737
rect -33106 37694 -33054 37703
rect -32946 37737 -32894 37746
rect -32946 37703 -32937 37737
rect -32937 37703 -32903 37737
rect -32903 37703 -32894 37737
rect -32946 37694 -32894 37703
rect -32786 37737 -32734 37746
rect -32786 37703 -32777 37737
rect -32777 37703 -32743 37737
rect -32743 37703 -32734 37737
rect -32786 37694 -32734 37703
rect -32626 37737 -32574 37746
rect -32626 37703 -32617 37737
rect -32617 37703 -32583 37737
rect -32583 37703 -32574 37737
rect -32626 37694 -32574 37703
rect -32466 37737 -32414 37746
rect -32466 37703 -32457 37737
rect -32457 37703 -32423 37737
rect -32423 37703 -32414 37737
rect -32466 37694 -32414 37703
rect -32306 37737 -32254 37746
rect -32306 37703 -32297 37737
rect -32297 37703 -32263 37737
rect -32263 37703 -32254 37737
rect -32306 37694 -32254 37703
rect -32146 37737 -32094 37746
rect -32146 37703 -32137 37737
rect -32137 37703 -32103 37737
rect -32103 37703 -32094 37737
rect -32146 37694 -32094 37703
rect -31986 37737 -31934 37746
rect -31986 37703 -31977 37737
rect -31977 37703 -31943 37737
rect -31943 37703 -31934 37737
rect -31986 37694 -31934 37703
rect -31826 37737 -31774 37746
rect -31826 37703 -31817 37737
rect -31817 37703 -31783 37737
rect -31783 37703 -31774 37737
rect -31826 37694 -31774 37703
rect -31666 37737 -31614 37746
rect -31666 37703 -31657 37737
rect -31657 37703 -31623 37737
rect -31623 37703 -31614 37737
rect -31666 37694 -31614 37703
rect -31506 37737 -31454 37746
rect -31506 37703 -31497 37737
rect -31497 37703 -31463 37737
rect -31463 37703 -31454 37737
rect -31506 37694 -31454 37703
rect -31346 37737 -31294 37746
rect -31346 37703 -31337 37737
rect -31337 37703 -31303 37737
rect -31303 37703 -31294 37737
rect -31346 37694 -31294 37703
rect -31186 37737 -31134 37746
rect -31186 37703 -31177 37737
rect -31177 37703 -31143 37737
rect -31143 37703 -31134 37737
rect -31186 37694 -31134 37703
rect -33106 37417 -33054 37426
rect -33106 37383 -33097 37417
rect -33097 37383 -33063 37417
rect -33063 37383 -33054 37417
rect -33106 37374 -33054 37383
rect -32946 37417 -32894 37426
rect -32946 37383 -32937 37417
rect -32937 37383 -32903 37417
rect -32903 37383 -32894 37417
rect -32946 37374 -32894 37383
rect -32786 37417 -32734 37426
rect -32786 37383 -32777 37417
rect -32777 37383 -32743 37417
rect -32743 37383 -32734 37417
rect -32786 37374 -32734 37383
rect -32626 37417 -32574 37426
rect -32626 37383 -32617 37417
rect -32617 37383 -32583 37417
rect -32583 37383 -32574 37417
rect -32626 37374 -32574 37383
rect -32466 37417 -32414 37426
rect -32466 37383 -32457 37417
rect -32457 37383 -32423 37417
rect -32423 37383 -32414 37417
rect -32466 37374 -32414 37383
rect -32306 37417 -32254 37426
rect -32306 37383 -32297 37417
rect -32297 37383 -32263 37417
rect -32263 37383 -32254 37417
rect -32306 37374 -32254 37383
rect -32146 37417 -32094 37426
rect -32146 37383 -32137 37417
rect -32137 37383 -32103 37417
rect -32103 37383 -32094 37417
rect -32146 37374 -32094 37383
rect -31986 37417 -31934 37426
rect -31986 37383 -31977 37417
rect -31977 37383 -31943 37417
rect -31943 37383 -31934 37417
rect -31986 37374 -31934 37383
rect -31826 37417 -31774 37426
rect -31826 37383 -31817 37417
rect -31817 37383 -31783 37417
rect -31783 37383 -31774 37417
rect -31826 37374 -31774 37383
rect -31666 37417 -31614 37426
rect -31666 37383 -31657 37417
rect -31657 37383 -31623 37417
rect -31623 37383 -31614 37417
rect -31666 37374 -31614 37383
rect -31506 37417 -31454 37426
rect -31506 37383 -31497 37417
rect -31497 37383 -31463 37417
rect -31463 37383 -31454 37417
rect -31506 37374 -31454 37383
rect -31346 37417 -31294 37426
rect -31346 37383 -31337 37417
rect -31337 37383 -31303 37417
rect -31303 37383 -31294 37417
rect -31346 37374 -31294 37383
rect -31186 37417 -31134 37426
rect -31186 37383 -31177 37417
rect -31177 37383 -31143 37417
rect -31143 37383 -31134 37417
rect -31186 37374 -31134 37383
rect -33106 37097 -33054 37106
rect -33106 37063 -33097 37097
rect -33097 37063 -33063 37097
rect -33063 37063 -33054 37097
rect -33106 37054 -33054 37063
rect -32946 37097 -32894 37106
rect -32946 37063 -32937 37097
rect -32937 37063 -32903 37097
rect -32903 37063 -32894 37097
rect -32946 37054 -32894 37063
rect -32786 37097 -32734 37106
rect -32786 37063 -32777 37097
rect -32777 37063 -32743 37097
rect -32743 37063 -32734 37097
rect -32786 37054 -32734 37063
rect -32626 37097 -32574 37106
rect -32626 37063 -32617 37097
rect -32617 37063 -32583 37097
rect -32583 37063 -32574 37097
rect -32626 37054 -32574 37063
rect -32466 37097 -32414 37106
rect -32466 37063 -32457 37097
rect -32457 37063 -32423 37097
rect -32423 37063 -32414 37097
rect -32466 37054 -32414 37063
rect -32306 37097 -32254 37106
rect -32306 37063 -32297 37097
rect -32297 37063 -32263 37097
rect -32263 37063 -32254 37097
rect -32306 37054 -32254 37063
rect -32146 37097 -32094 37106
rect -32146 37063 -32137 37097
rect -32137 37063 -32103 37097
rect -32103 37063 -32094 37097
rect -32146 37054 -32094 37063
rect -31986 37097 -31934 37106
rect -31986 37063 -31977 37097
rect -31977 37063 -31943 37097
rect -31943 37063 -31934 37097
rect -31986 37054 -31934 37063
rect -31826 37097 -31774 37106
rect -31826 37063 -31817 37097
rect -31817 37063 -31783 37097
rect -31783 37063 -31774 37097
rect -31826 37054 -31774 37063
rect -31666 37097 -31614 37106
rect -31666 37063 -31657 37097
rect -31657 37063 -31623 37097
rect -31623 37063 -31614 37097
rect -31666 37054 -31614 37063
rect -31506 37097 -31454 37106
rect -31506 37063 -31497 37097
rect -31497 37063 -31463 37097
rect -31463 37063 -31454 37097
rect -31506 37054 -31454 37063
rect -31346 37097 -31294 37106
rect -31346 37063 -31337 37097
rect -31337 37063 -31303 37097
rect -31303 37063 -31294 37097
rect -31346 37054 -31294 37063
rect -31186 37097 -31134 37106
rect -31186 37063 -31177 37097
rect -31177 37063 -31143 37097
rect -31143 37063 -31134 37097
rect -31186 37054 -31134 37063
rect 41054 36057 41106 36066
rect 41054 36023 41063 36057
rect 41063 36023 41097 36057
rect 41097 36023 41106 36057
rect 41054 36014 41106 36023
rect 41214 36057 41266 36066
rect 41214 36023 41223 36057
rect 41223 36023 41257 36057
rect 41257 36023 41266 36057
rect 41214 36014 41266 36023
rect 41374 36057 41426 36066
rect 41374 36023 41383 36057
rect 41383 36023 41417 36057
rect 41417 36023 41426 36057
rect 41374 36014 41426 36023
rect 41534 36057 41586 36066
rect 41534 36023 41543 36057
rect 41543 36023 41577 36057
rect 41577 36023 41586 36057
rect 41534 36014 41586 36023
rect 41694 36057 41746 36066
rect 41694 36023 41703 36057
rect 41703 36023 41737 36057
rect 41737 36023 41746 36057
rect 41694 36014 41746 36023
rect 41854 36057 41906 36066
rect 41854 36023 41863 36057
rect 41863 36023 41897 36057
rect 41897 36023 41906 36057
rect 41854 36014 41906 36023
rect 42014 36057 42066 36066
rect 42014 36023 42023 36057
rect 42023 36023 42057 36057
rect 42057 36023 42066 36057
rect 42014 36014 42066 36023
rect 42174 36057 42226 36066
rect 42174 36023 42183 36057
rect 42183 36023 42217 36057
rect 42217 36023 42226 36057
rect 42174 36014 42226 36023
rect 42334 36057 42386 36066
rect 42334 36023 42343 36057
rect 42343 36023 42377 36057
rect 42377 36023 42386 36057
rect 42334 36014 42386 36023
rect 42494 36057 42546 36066
rect 42494 36023 42503 36057
rect 42503 36023 42537 36057
rect 42537 36023 42546 36057
rect 42494 36014 42546 36023
rect 42654 36057 42706 36066
rect 42654 36023 42663 36057
rect 42663 36023 42697 36057
rect 42697 36023 42706 36057
rect 42654 36014 42706 36023
rect 42814 36057 42866 36066
rect 42814 36023 42823 36057
rect 42823 36023 42857 36057
rect 42857 36023 42866 36057
rect 42814 36014 42866 36023
rect 42974 36057 43026 36066
rect 42974 36023 42983 36057
rect 42983 36023 43017 36057
rect 43017 36023 43026 36057
rect 42974 36014 43026 36023
rect 43134 36057 43186 36066
rect 43134 36023 43143 36057
rect 43143 36023 43177 36057
rect 43177 36023 43186 36057
rect 43134 36014 43186 36023
rect 41054 35737 41106 35746
rect 41054 35703 41063 35737
rect 41063 35703 41097 35737
rect 41097 35703 41106 35737
rect 41054 35694 41106 35703
rect 41214 35737 41266 35746
rect 41214 35703 41223 35737
rect 41223 35703 41257 35737
rect 41257 35703 41266 35737
rect 41214 35694 41266 35703
rect 41374 35737 41426 35746
rect 41374 35703 41383 35737
rect 41383 35703 41417 35737
rect 41417 35703 41426 35737
rect 41374 35694 41426 35703
rect 41534 35737 41586 35746
rect 41534 35703 41543 35737
rect 41543 35703 41577 35737
rect 41577 35703 41586 35737
rect 41534 35694 41586 35703
rect 41694 35737 41746 35746
rect 41694 35703 41703 35737
rect 41703 35703 41737 35737
rect 41737 35703 41746 35737
rect 41694 35694 41746 35703
rect 41854 35737 41906 35746
rect 41854 35703 41863 35737
rect 41863 35703 41897 35737
rect 41897 35703 41906 35737
rect 41854 35694 41906 35703
rect 42014 35737 42066 35746
rect 42014 35703 42023 35737
rect 42023 35703 42057 35737
rect 42057 35703 42066 35737
rect 42014 35694 42066 35703
rect 42174 35737 42226 35746
rect 42174 35703 42183 35737
rect 42183 35703 42217 35737
rect 42217 35703 42226 35737
rect 42174 35694 42226 35703
rect 42334 35737 42386 35746
rect 42334 35703 42343 35737
rect 42343 35703 42377 35737
rect 42377 35703 42386 35737
rect 42334 35694 42386 35703
rect 42494 35737 42546 35746
rect 42494 35703 42503 35737
rect 42503 35703 42537 35737
rect 42537 35703 42546 35737
rect 42494 35694 42546 35703
rect 42654 35737 42706 35746
rect 42654 35703 42663 35737
rect 42663 35703 42697 35737
rect 42697 35703 42706 35737
rect 42654 35694 42706 35703
rect 42814 35737 42866 35746
rect 42814 35703 42823 35737
rect 42823 35703 42857 35737
rect 42857 35703 42866 35737
rect 42814 35694 42866 35703
rect 42974 35737 43026 35746
rect 42974 35703 42983 35737
rect 42983 35703 43017 35737
rect 43017 35703 43026 35737
rect 42974 35694 43026 35703
rect 43134 35737 43186 35746
rect 43134 35703 43143 35737
rect 43143 35703 43177 35737
rect 43177 35703 43186 35737
rect 43134 35694 43186 35703
rect -33106 34697 -33054 34706
rect -33106 34663 -33097 34697
rect -33097 34663 -33063 34697
rect -33063 34663 -33054 34697
rect -33106 34654 -33054 34663
rect -32946 34697 -32894 34706
rect -32946 34663 -32937 34697
rect -32937 34663 -32903 34697
rect -32903 34663 -32894 34697
rect -32946 34654 -32894 34663
rect -32786 34697 -32734 34706
rect -32786 34663 -32777 34697
rect -32777 34663 -32743 34697
rect -32743 34663 -32734 34697
rect -32786 34654 -32734 34663
rect -32626 34697 -32574 34706
rect -32626 34663 -32617 34697
rect -32617 34663 -32583 34697
rect -32583 34663 -32574 34697
rect -32626 34654 -32574 34663
rect -32466 34697 -32414 34706
rect -32466 34663 -32457 34697
rect -32457 34663 -32423 34697
rect -32423 34663 -32414 34697
rect -32466 34654 -32414 34663
rect -32306 34697 -32254 34706
rect -32306 34663 -32297 34697
rect -32297 34663 -32263 34697
rect -32263 34663 -32254 34697
rect -32306 34654 -32254 34663
rect -32146 34697 -32094 34706
rect -32146 34663 -32137 34697
rect -32137 34663 -32103 34697
rect -32103 34663 -32094 34697
rect -32146 34654 -32094 34663
rect -31986 34697 -31934 34706
rect -31986 34663 -31977 34697
rect -31977 34663 -31943 34697
rect -31943 34663 -31934 34697
rect -31986 34654 -31934 34663
rect -31826 34697 -31774 34706
rect -31826 34663 -31817 34697
rect -31817 34663 -31783 34697
rect -31783 34663 -31774 34697
rect -31826 34654 -31774 34663
rect -31666 34697 -31614 34706
rect -31666 34663 -31657 34697
rect -31657 34663 -31623 34697
rect -31623 34663 -31614 34697
rect -31666 34654 -31614 34663
rect -31506 34697 -31454 34706
rect -31506 34663 -31497 34697
rect -31497 34663 -31463 34697
rect -31463 34663 -31454 34697
rect -31506 34654 -31454 34663
rect -31346 34697 -31294 34706
rect -31346 34663 -31337 34697
rect -31337 34663 -31303 34697
rect -31303 34663 -31294 34697
rect -31346 34654 -31294 34663
rect -31186 34697 -31134 34706
rect -31186 34663 -31177 34697
rect -31177 34663 -31143 34697
rect -31143 34663 -31134 34697
rect -31186 34654 -31134 34663
rect -29906 34697 -29854 34706
rect -29906 34663 -29897 34697
rect -29897 34663 -29863 34697
rect -29863 34663 -29854 34697
rect -29906 34654 -29854 34663
rect -29746 34697 -29694 34706
rect -29746 34663 -29737 34697
rect -29737 34663 -29703 34697
rect -29703 34663 -29694 34697
rect -29746 34654 -29694 34663
rect -29586 34697 -29534 34706
rect -29586 34663 -29577 34697
rect -29577 34663 -29543 34697
rect -29543 34663 -29534 34697
rect -29586 34654 -29534 34663
rect -29426 34697 -29374 34706
rect -29426 34663 -29417 34697
rect -29417 34663 -29383 34697
rect -29383 34663 -29374 34697
rect -29426 34654 -29374 34663
rect -29266 34697 -29214 34706
rect -29266 34663 -29257 34697
rect -29257 34663 -29223 34697
rect -29223 34663 -29214 34697
rect -29266 34654 -29214 34663
rect -29106 34697 -29054 34706
rect -29106 34663 -29097 34697
rect -29097 34663 -29063 34697
rect -29063 34663 -29054 34697
rect -29106 34654 -29054 34663
rect -28946 34697 -28894 34706
rect -28946 34663 -28937 34697
rect -28937 34663 -28903 34697
rect -28903 34663 -28894 34697
rect -28946 34654 -28894 34663
rect -28786 34697 -28734 34706
rect -28786 34663 -28777 34697
rect -28777 34663 -28743 34697
rect -28743 34663 -28734 34697
rect -28786 34654 -28734 34663
rect -28626 34697 -28574 34706
rect -28626 34663 -28617 34697
rect -28617 34663 -28583 34697
rect -28583 34663 -28574 34697
rect -28626 34654 -28574 34663
rect -28466 34697 -28414 34706
rect -28466 34663 -28457 34697
rect -28457 34663 -28423 34697
rect -28423 34663 -28414 34697
rect -28466 34654 -28414 34663
rect -28306 34697 -28254 34706
rect -28306 34663 -28297 34697
rect -28297 34663 -28263 34697
rect -28263 34663 -28254 34697
rect -28306 34654 -28254 34663
rect -28146 34697 -28094 34706
rect -28146 34663 -28137 34697
rect -28137 34663 -28103 34697
rect -28103 34663 -28094 34697
rect -28146 34654 -28094 34663
rect -27986 34697 -27934 34706
rect -27986 34663 -27977 34697
rect -27977 34663 -27943 34697
rect -27943 34663 -27934 34697
rect -27986 34654 -27934 34663
rect -27826 34697 -27774 34706
rect -27826 34663 -27817 34697
rect -27817 34663 -27783 34697
rect -27783 34663 -27774 34697
rect -27826 34654 -27774 34663
rect -27666 34697 -27614 34706
rect -27666 34663 -27657 34697
rect -27657 34663 -27623 34697
rect -27623 34663 -27614 34697
rect -27666 34654 -27614 34663
rect -27506 34697 -27454 34706
rect -27506 34663 -27497 34697
rect -27497 34663 -27463 34697
rect -27463 34663 -27454 34697
rect -27506 34654 -27454 34663
rect -27346 34697 -27294 34706
rect -27346 34663 -27337 34697
rect -27337 34663 -27303 34697
rect -27303 34663 -27294 34697
rect -27346 34654 -27294 34663
rect -27186 34697 -27134 34706
rect -27186 34663 -27177 34697
rect -27177 34663 -27143 34697
rect -27143 34663 -27134 34697
rect -27186 34654 -27134 34663
rect -27026 34697 -26974 34706
rect -27026 34663 -27017 34697
rect -27017 34663 -26983 34697
rect -26983 34663 -26974 34697
rect -27026 34654 -26974 34663
rect -26866 34697 -26814 34706
rect -26866 34663 -26857 34697
rect -26857 34663 -26823 34697
rect -26823 34663 -26814 34697
rect -26866 34654 -26814 34663
rect -26706 34697 -26654 34706
rect -26706 34663 -26697 34697
rect -26697 34663 -26663 34697
rect -26663 34663 -26654 34697
rect -26706 34654 -26654 34663
rect -26546 34697 -26494 34706
rect -26546 34663 -26537 34697
rect -26537 34663 -26503 34697
rect -26503 34663 -26494 34697
rect -26546 34654 -26494 34663
rect -26386 34697 -26334 34706
rect -26386 34663 -26377 34697
rect -26377 34663 -26343 34697
rect -26343 34663 -26334 34697
rect -26386 34654 -26334 34663
rect -26226 34697 -26174 34706
rect -26226 34663 -26217 34697
rect -26217 34663 -26183 34697
rect -26183 34663 -26174 34697
rect -26226 34654 -26174 34663
rect -26066 34697 -26014 34706
rect -26066 34663 -26057 34697
rect -26057 34663 -26023 34697
rect -26023 34663 -26014 34697
rect -26066 34654 -26014 34663
rect -25906 34697 -25854 34706
rect -25906 34663 -25897 34697
rect -25897 34663 -25863 34697
rect -25863 34663 -25854 34697
rect -25906 34654 -25854 34663
rect -25746 34697 -25694 34706
rect -25746 34663 -25737 34697
rect -25737 34663 -25703 34697
rect -25703 34663 -25694 34697
rect -25746 34654 -25694 34663
rect -25586 34697 -25534 34706
rect -25586 34663 -25577 34697
rect -25577 34663 -25543 34697
rect -25543 34663 -25534 34697
rect -25586 34654 -25534 34663
rect -25426 34697 -25374 34706
rect -25426 34663 -25417 34697
rect -25417 34663 -25383 34697
rect -25383 34663 -25374 34697
rect -25426 34654 -25374 34663
rect -25266 34697 -25214 34706
rect -25266 34663 -25257 34697
rect -25257 34663 -25223 34697
rect -25223 34663 -25214 34697
rect -25266 34654 -25214 34663
rect -25106 34697 -25054 34706
rect -25106 34663 -25097 34697
rect -25097 34663 -25063 34697
rect -25063 34663 -25054 34697
rect -25106 34654 -25054 34663
rect -24946 34697 -24894 34706
rect -24946 34663 -24937 34697
rect -24937 34663 -24903 34697
rect -24903 34663 -24894 34697
rect -24946 34654 -24894 34663
rect -24786 34697 -24734 34706
rect -24786 34663 -24777 34697
rect -24777 34663 -24743 34697
rect -24743 34663 -24734 34697
rect -24786 34654 -24734 34663
rect -24626 34697 -24574 34706
rect -24626 34663 -24617 34697
rect -24617 34663 -24583 34697
rect -24583 34663 -24574 34697
rect -24626 34654 -24574 34663
rect -24466 34697 -24414 34706
rect -24466 34663 -24457 34697
rect -24457 34663 -24423 34697
rect -24423 34663 -24414 34697
rect -24466 34654 -24414 34663
rect -24306 34697 -24254 34706
rect -24306 34663 -24297 34697
rect -24297 34663 -24263 34697
rect -24263 34663 -24254 34697
rect -24306 34654 -24254 34663
rect -24146 34697 -24094 34706
rect -24146 34663 -24137 34697
rect -24137 34663 -24103 34697
rect -24103 34663 -24094 34697
rect -24146 34654 -24094 34663
rect -23986 34697 -23934 34706
rect -23986 34663 -23977 34697
rect -23977 34663 -23943 34697
rect -23943 34663 -23934 34697
rect -23986 34654 -23934 34663
rect -23826 34697 -23774 34706
rect -23826 34663 -23817 34697
rect -23817 34663 -23783 34697
rect -23783 34663 -23774 34697
rect -23826 34654 -23774 34663
rect -23666 34697 -23614 34706
rect -23666 34663 -23657 34697
rect -23657 34663 -23623 34697
rect -23623 34663 -23614 34697
rect -23666 34654 -23614 34663
rect -23506 34697 -23454 34706
rect -23506 34663 -23497 34697
rect -23497 34663 -23463 34697
rect -23463 34663 -23454 34697
rect -23506 34654 -23454 34663
rect -23346 34697 -23294 34706
rect -23346 34663 -23337 34697
rect -23337 34663 -23303 34697
rect -23303 34663 -23294 34697
rect -23346 34654 -23294 34663
rect -23186 34697 -23134 34706
rect -23186 34663 -23177 34697
rect -23177 34663 -23143 34697
rect -23143 34663 -23134 34697
rect -23186 34654 -23134 34663
rect -23026 34697 -22974 34706
rect -23026 34663 -23017 34697
rect -23017 34663 -22983 34697
rect -22983 34663 -22974 34697
rect -23026 34654 -22974 34663
rect -22866 34697 -22814 34706
rect -22866 34663 -22857 34697
rect -22857 34663 -22823 34697
rect -22823 34663 -22814 34697
rect -22866 34654 -22814 34663
rect -22706 34697 -22654 34706
rect -22706 34663 -22697 34697
rect -22697 34663 -22663 34697
rect -22663 34663 -22654 34697
rect -22706 34654 -22654 34663
rect -22546 34697 -22494 34706
rect -22546 34663 -22537 34697
rect -22537 34663 -22503 34697
rect -22503 34663 -22494 34697
rect -22546 34654 -22494 34663
rect -22386 34697 -22334 34706
rect -22386 34663 -22377 34697
rect -22377 34663 -22343 34697
rect -22343 34663 -22334 34697
rect -22386 34654 -22334 34663
rect -22226 34697 -22174 34706
rect -22226 34663 -22217 34697
rect -22217 34663 -22183 34697
rect -22183 34663 -22174 34697
rect -22226 34654 -22174 34663
rect -22066 34697 -22014 34706
rect -22066 34663 -22057 34697
rect -22057 34663 -22023 34697
rect -22023 34663 -22014 34697
rect -22066 34654 -22014 34663
rect -21906 34697 -21854 34706
rect -21906 34663 -21897 34697
rect -21897 34663 -21863 34697
rect -21863 34663 -21854 34697
rect -21906 34654 -21854 34663
rect -21746 34697 -21694 34706
rect -21746 34663 -21737 34697
rect -21737 34663 -21703 34697
rect -21703 34663 -21694 34697
rect -21746 34654 -21694 34663
rect -21586 34697 -21534 34706
rect -21586 34663 -21577 34697
rect -21577 34663 -21543 34697
rect -21543 34663 -21534 34697
rect -21586 34654 -21534 34663
rect -21426 34697 -21374 34706
rect -21426 34663 -21417 34697
rect -21417 34663 -21383 34697
rect -21383 34663 -21374 34697
rect -21426 34654 -21374 34663
rect -21266 34697 -21214 34706
rect -21266 34663 -21257 34697
rect -21257 34663 -21223 34697
rect -21223 34663 -21214 34697
rect -21266 34654 -21214 34663
rect -21106 34697 -21054 34706
rect -21106 34663 -21097 34697
rect -21097 34663 -21063 34697
rect -21063 34663 -21054 34697
rect -21106 34654 -21054 34663
rect -20946 34697 -20894 34706
rect -20946 34663 -20937 34697
rect -20937 34663 -20903 34697
rect -20903 34663 -20894 34697
rect -20946 34654 -20894 34663
rect -20786 34697 -20734 34706
rect -20786 34663 -20777 34697
rect -20777 34663 -20743 34697
rect -20743 34663 -20734 34697
rect -20786 34654 -20734 34663
rect -20626 34697 -20574 34706
rect -20626 34663 -20617 34697
rect -20617 34663 -20583 34697
rect -20583 34663 -20574 34697
rect -20626 34654 -20574 34663
rect -20466 34697 -20414 34706
rect -20466 34663 -20457 34697
rect -20457 34663 -20423 34697
rect -20423 34663 -20414 34697
rect -20466 34654 -20414 34663
rect -20306 34697 -20254 34706
rect -20306 34663 -20297 34697
rect -20297 34663 -20263 34697
rect -20263 34663 -20254 34697
rect -20306 34654 -20254 34663
rect -20146 34697 -20094 34706
rect -20146 34663 -20137 34697
rect -20137 34663 -20103 34697
rect -20103 34663 -20094 34697
rect -20146 34654 -20094 34663
rect -19986 34697 -19934 34706
rect -19986 34663 -19977 34697
rect -19977 34663 -19943 34697
rect -19943 34663 -19934 34697
rect -19986 34654 -19934 34663
rect -19826 34697 -19774 34706
rect -19826 34663 -19817 34697
rect -19817 34663 -19783 34697
rect -19783 34663 -19774 34697
rect -19826 34654 -19774 34663
rect -19666 34697 -19614 34706
rect -19666 34663 -19657 34697
rect -19657 34663 -19623 34697
rect -19623 34663 -19614 34697
rect -19666 34654 -19614 34663
rect -19506 34697 -19454 34706
rect -19506 34663 -19497 34697
rect -19497 34663 -19463 34697
rect -19463 34663 -19454 34697
rect -19506 34654 -19454 34663
rect -19346 34697 -19294 34706
rect -19346 34663 -19337 34697
rect -19337 34663 -19303 34697
rect -19303 34663 -19294 34697
rect -19346 34654 -19294 34663
rect -19186 34697 -19134 34706
rect -19186 34663 -19177 34697
rect -19177 34663 -19143 34697
rect -19143 34663 -19134 34697
rect -19186 34654 -19134 34663
rect -19026 34697 -18974 34706
rect -19026 34663 -19017 34697
rect -19017 34663 -18983 34697
rect -18983 34663 -18974 34697
rect -19026 34654 -18974 34663
rect -18866 34697 -18814 34706
rect -18866 34663 -18857 34697
rect -18857 34663 -18823 34697
rect -18823 34663 -18814 34697
rect -18866 34654 -18814 34663
rect -18706 34697 -18654 34706
rect -18706 34663 -18697 34697
rect -18697 34663 -18663 34697
rect -18663 34663 -18654 34697
rect -18706 34654 -18654 34663
rect -18546 34697 -18494 34706
rect -18546 34663 -18537 34697
rect -18537 34663 -18503 34697
rect -18503 34663 -18494 34697
rect -18546 34654 -18494 34663
rect -18386 34697 -18334 34706
rect -18386 34663 -18377 34697
rect -18377 34663 -18343 34697
rect -18343 34663 -18334 34697
rect -18386 34654 -18334 34663
rect -18226 34697 -18174 34706
rect -18226 34663 -18217 34697
rect -18217 34663 -18183 34697
rect -18183 34663 -18174 34697
rect -18226 34654 -18174 34663
rect -18066 34697 -18014 34706
rect -18066 34663 -18057 34697
rect -18057 34663 -18023 34697
rect -18023 34663 -18014 34697
rect -18066 34654 -18014 34663
rect -17906 34697 -17854 34706
rect -17906 34663 -17897 34697
rect -17897 34663 -17863 34697
rect -17863 34663 -17854 34697
rect -17906 34654 -17854 34663
rect -17746 34697 -17694 34706
rect -17746 34663 -17737 34697
rect -17737 34663 -17703 34697
rect -17703 34663 -17694 34697
rect -17746 34654 -17694 34663
rect -17586 34697 -17534 34706
rect -17586 34663 -17577 34697
rect -17577 34663 -17543 34697
rect -17543 34663 -17534 34697
rect -17586 34654 -17534 34663
rect -17426 34697 -17374 34706
rect -17426 34663 -17417 34697
rect -17417 34663 -17383 34697
rect -17383 34663 -17374 34697
rect -17426 34654 -17374 34663
rect -17266 34697 -17214 34706
rect -17266 34663 -17257 34697
rect -17257 34663 -17223 34697
rect -17223 34663 -17214 34697
rect -17266 34654 -17214 34663
rect -17106 34697 -17054 34706
rect -17106 34663 -17097 34697
rect -17097 34663 -17063 34697
rect -17063 34663 -17054 34697
rect -17106 34654 -17054 34663
rect -16946 34697 -16894 34706
rect -16946 34663 -16937 34697
rect -16937 34663 -16903 34697
rect -16903 34663 -16894 34697
rect -16946 34654 -16894 34663
rect -16786 34697 -16734 34706
rect -16786 34663 -16777 34697
rect -16777 34663 -16743 34697
rect -16743 34663 -16734 34697
rect -16786 34654 -16734 34663
rect -16626 34697 -16574 34706
rect -16626 34663 -16617 34697
rect -16617 34663 -16583 34697
rect -16583 34663 -16574 34697
rect -16626 34654 -16574 34663
rect -16466 34697 -16414 34706
rect -16466 34663 -16457 34697
rect -16457 34663 -16423 34697
rect -16423 34663 -16414 34697
rect -16466 34654 -16414 34663
rect -16306 34697 -16254 34706
rect -16306 34663 -16297 34697
rect -16297 34663 -16263 34697
rect -16263 34663 -16254 34697
rect -16306 34654 -16254 34663
rect -16146 34697 -16094 34706
rect -16146 34663 -16137 34697
rect -16137 34663 -16103 34697
rect -16103 34663 -16094 34697
rect -16146 34654 -16094 34663
rect -15986 34697 -15934 34706
rect -15986 34663 -15977 34697
rect -15977 34663 -15943 34697
rect -15943 34663 -15934 34697
rect -15986 34654 -15934 34663
rect -15826 34697 -15774 34706
rect -15826 34663 -15817 34697
rect -15817 34663 -15783 34697
rect -15783 34663 -15774 34697
rect -15826 34654 -15774 34663
rect -15666 34697 -15614 34706
rect -15666 34663 -15657 34697
rect -15657 34663 -15623 34697
rect -15623 34663 -15614 34697
rect -15666 34654 -15614 34663
rect -15506 34697 -15454 34706
rect -15506 34663 -15497 34697
rect -15497 34663 -15463 34697
rect -15463 34663 -15454 34697
rect -15506 34654 -15454 34663
rect -15346 34697 -15294 34706
rect -15346 34663 -15337 34697
rect -15337 34663 -15303 34697
rect -15303 34663 -15294 34697
rect -15346 34654 -15294 34663
rect -15186 34697 -15134 34706
rect -15186 34663 -15177 34697
rect -15177 34663 -15143 34697
rect -15143 34663 -15134 34697
rect -15186 34654 -15134 34663
rect -15026 34697 -14974 34706
rect -15026 34663 -15017 34697
rect -15017 34663 -14983 34697
rect -14983 34663 -14974 34697
rect -15026 34654 -14974 34663
rect -14866 34697 -14814 34706
rect -14866 34663 -14857 34697
rect -14857 34663 -14823 34697
rect -14823 34663 -14814 34697
rect -14866 34654 -14814 34663
rect -14706 34697 -14654 34706
rect -14706 34663 -14697 34697
rect -14697 34663 -14663 34697
rect -14663 34663 -14654 34697
rect -14706 34654 -14654 34663
rect -14546 34697 -14494 34706
rect -14546 34663 -14537 34697
rect -14537 34663 -14503 34697
rect -14503 34663 -14494 34697
rect -14546 34654 -14494 34663
rect -14386 34697 -14334 34706
rect -14386 34663 -14377 34697
rect -14377 34663 -14343 34697
rect -14343 34663 -14334 34697
rect -14386 34654 -14334 34663
rect -14226 34697 -14174 34706
rect -14226 34663 -14217 34697
rect -14217 34663 -14183 34697
rect -14183 34663 -14174 34697
rect -14226 34654 -14174 34663
rect -14066 34697 -14014 34706
rect -14066 34663 -14057 34697
rect -14057 34663 -14023 34697
rect -14023 34663 -14014 34697
rect -14066 34654 -14014 34663
rect -13906 34697 -13854 34706
rect -13906 34663 -13897 34697
rect -13897 34663 -13863 34697
rect -13863 34663 -13854 34697
rect -13906 34654 -13854 34663
rect -13746 34697 -13694 34706
rect -13746 34663 -13737 34697
rect -13737 34663 -13703 34697
rect -13703 34663 -13694 34697
rect -13746 34654 -13694 34663
rect -13586 34697 -13534 34706
rect -13586 34663 -13577 34697
rect -13577 34663 -13543 34697
rect -13543 34663 -13534 34697
rect -13586 34654 -13534 34663
rect -13426 34697 -13374 34706
rect -13426 34663 -13417 34697
rect -13417 34663 -13383 34697
rect -13383 34663 -13374 34697
rect -13426 34654 -13374 34663
rect -13266 34697 -13214 34706
rect -13266 34663 -13257 34697
rect -13257 34663 -13223 34697
rect -13223 34663 -13214 34697
rect -13266 34654 -13214 34663
rect -13106 34697 -13054 34706
rect -13106 34663 -13097 34697
rect -13097 34663 -13063 34697
rect -13063 34663 -13054 34697
rect -13106 34654 -13054 34663
rect -12946 34697 -12894 34706
rect -12946 34663 -12937 34697
rect -12937 34663 -12903 34697
rect -12903 34663 -12894 34697
rect -12946 34654 -12894 34663
rect -12786 34697 -12734 34706
rect -12786 34663 -12777 34697
rect -12777 34663 -12743 34697
rect -12743 34663 -12734 34697
rect -12786 34654 -12734 34663
rect -12626 34697 -12574 34706
rect -12626 34663 -12617 34697
rect -12617 34663 -12583 34697
rect -12583 34663 -12574 34697
rect -12626 34654 -12574 34663
rect -12466 34697 -12414 34706
rect -12466 34663 -12457 34697
rect -12457 34663 -12423 34697
rect -12423 34663 -12414 34697
rect -12466 34654 -12414 34663
rect -12306 34697 -12254 34706
rect -12306 34663 -12297 34697
rect -12297 34663 -12263 34697
rect -12263 34663 -12254 34697
rect -12306 34654 -12254 34663
rect -12146 34697 -12094 34706
rect -12146 34663 -12137 34697
rect -12137 34663 -12103 34697
rect -12103 34663 -12094 34697
rect -12146 34654 -12094 34663
rect -11986 34697 -11934 34706
rect -11986 34663 -11977 34697
rect -11977 34663 -11943 34697
rect -11943 34663 -11934 34697
rect -11986 34654 -11934 34663
rect -11826 34697 -11774 34706
rect -11826 34663 -11817 34697
rect -11817 34663 -11783 34697
rect -11783 34663 -11774 34697
rect -11826 34654 -11774 34663
rect -11666 34697 -11614 34706
rect -11666 34663 -11657 34697
rect -11657 34663 -11623 34697
rect -11623 34663 -11614 34697
rect -11666 34654 -11614 34663
rect -11506 34697 -11454 34706
rect -11506 34663 -11497 34697
rect -11497 34663 -11463 34697
rect -11463 34663 -11454 34697
rect -11506 34654 -11454 34663
rect -10866 34697 -10814 34706
rect -10866 34663 -10857 34697
rect -10857 34663 -10823 34697
rect -10823 34663 -10814 34697
rect -10866 34654 -10814 34663
rect -10546 34697 -10494 34706
rect -10546 34663 -10537 34697
rect -10537 34663 -10503 34697
rect -10503 34663 -10494 34697
rect -10546 34654 -10494 34663
rect -33106 34377 -33054 34386
rect -33106 34343 -33097 34377
rect -33097 34343 -33063 34377
rect -33063 34343 -33054 34377
rect -33106 34334 -33054 34343
rect -32946 34377 -32894 34386
rect -32946 34343 -32937 34377
rect -32937 34343 -32903 34377
rect -32903 34343 -32894 34377
rect -32946 34334 -32894 34343
rect -32786 34377 -32734 34386
rect -32786 34343 -32777 34377
rect -32777 34343 -32743 34377
rect -32743 34343 -32734 34377
rect -32786 34334 -32734 34343
rect -32626 34377 -32574 34386
rect -32626 34343 -32617 34377
rect -32617 34343 -32583 34377
rect -32583 34343 -32574 34377
rect -32626 34334 -32574 34343
rect -32466 34377 -32414 34386
rect -32466 34343 -32457 34377
rect -32457 34343 -32423 34377
rect -32423 34343 -32414 34377
rect -32466 34334 -32414 34343
rect -32306 34377 -32254 34386
rect -32306 34343 -32297 34377
rect -32297 34343 -32263 34377
rect -32263 34343 -32254 34377
rect -32306 34334 -32254 34343
rect -32146 34377 -32094 34386
rect -32146 34343 -32137 34377
rect -32137 34343 -32103 34377
rect -32103 34343 -32094 34377
rect -32146 34334 -32094 34343
rect -31986 34377 -31934 34386
rect -31986 34343 -31977 34377
rect -31977 34343 -31943 34377
rect -31943 34343 -31934 34377
rect -31986 34334 -31934 34343
rect -31826 34377 -31774 34386
rect -31826 34343 -31817 34377
rect -31817 34343 -31783 34377
rect -31783 34343 -31774 34377
rect -31826 34334 -31774 34343
rect -31666 34377 -31614 34386
rect -31666 34343 -31657 34377
rect -31657 34343 -31623 34377
rect -31623 34343 -31614 34377
rect -31666 34334 -31614 34343
rect -31506 34377 -31454 34386
rect -31506 34343 -31497 34377
rect -31497 34343 -31463 34377
rect -31463 34343 -31454 34377
rect -31506 34334 -31454 34343
rect -31346 34377 -31294 34386
rect -31346 34343 -31337 34377
rect -31337 34343 -31303 34377
rect -31303 34343 -31294 34377
rect -31346 34334 -31294 34343
rect -31186 34377 -31134 34386
rect -31186 34343 -31177 34377
rect -31177 34343 -31143 34377
rect -31143 34343 -31134 34377
rect -31186 34334 -31134 34343
rect -29906 34377 -29854 34386
rect -29906 34343 -29897 34377
rect -29897 34343 -29863 34377
rect -29863 34343 -29854 34377
rect -29906 34334 -29854 34343
rect -29746 34377 -29694 34386
rect -29746 34343 -29737 34377
rect -29737 34343 -29703 34377
rect -29703 34343 -29694 34377
rect -29746 34334 -29694 34343
rect -29586 34377 -29534 34386
rect -29586 34343 -29577 34377
rect -29577 34343 -29543 34377
rect -29543 34343 -29534 34377
rect -29586 34334 -29534 34343
rect -29426 34377 -29374 34386
rect -29426 34343 -29417 34377
rect -29417 34343 -29383 34377
rect -29383 34343 -29374 34377
rect -29426 34334 -29374 34343
rect -29266 34377 -29214 34386
rect -29266 34343 -29257 34377
rect -29257 34343 -29223 34377
rect -29223 34343 -29214 34377
rect -29266 34334 -29214 34343
rect -29106 34377 -29054 34386
rect -29106 34343 -29097 34377
rect -29097 34343 -29063 34377
rect -29063 34343 -29054 34377
rect -29106 34334 -29054 34343
rect -28946 34377 -28894 34386
rect -28946 34343 -28937 34377
rect -28937 34343 -28903 34377
rect -28903 34343 -28894 34377
rect -28946 34334 -28894 34343
rect -28786 34377 -28734 34386
rect -28786 34343 -28777 34377
rect -28777 34343 -28743 34377
rect -28743 34343 -28734 34377
rect -28786 34334 -28734 34343
rect -28626 34377 -28574 34386
rect -28626 34343 -28617 34377
rect -28617 34343 -28583 34377
rect -28583 34343 -28574 34377
rect -28626 34334 -28574 34343
rect -28466 34377 -28414 34386
rect -28466 34343 -28457 34377
rect -28457 34343 -28423 34377
rect -28423 34343 -28414 34377
rect -28466 34334 -28414 34343
rect -28306 34377 -28254 34386
rect -28306 34343 -28297 34377
rect -28297 34343 -28263 34377
rect -28263 34343 -28254 34377
rect -28306 34334 -28254 34343
rect -28146 34377 -28094 34386
rect -28146 34343 -28137 34377
rect -28137 34343 -28103 34377
rect -28103 34343 -28094 34377
rect -28146 34334 -28094 34343
rect -27986 34377 -27934 34386
rect -27986 34343 -27977 34377
rect -27977 34343 -27943 34377
rect -27943 34343 -27934 34377
rect -27986 34334 -27934 34343
rect -27826 34377 -27774 34386
rect -27826 34343 -27817 34377
rect -27817 34343 -27783 34377
rect -27783 34343 -27774 34377
rect -27826 34334 -27774 34343
rect -27666 34377 -27614 34386
rect -27666 34343 -27657 34377
rect -27657 34343 -27623 34377
rect -27623 34343 -27614 34377
rect -27666 34334 -27614 34343
rect -27506 34377 -27454 34386
rect -27506 34343 -27497 34377
rect -27497 34343 -27463 34377
rect -27463 34343 -27454 34377
rect -27506 34334 -27454 34343
rect -27346 34377 -27294 34386
rect -27346 34343 -27337 34377
rect -27337 34343 -27303 34377
rect -27303 34343 -27294 34377
rect -27346 34334 -27294 34343
rect -27186 34377 -27134 34386
rect -27186 34343 -27177 34377
rect -27177 34343 -27143 34377
rect -27143 34343 -27134 34377
rect -27186 34334 -27134 34343
rect -27026 34377 -26974 34386
rect -27026 34343 -27017 34377
rect -27017 34343 -26983 34377
rect -26983 34343 -26974 34377
rect -27026 34334 -26974 34343
rect -26866 34377 -26814 34386
rect -26866 34343 -26857 34377
rect -26857 34343 -26823 34377
rect -26823 34343 -26814 34377
rect -26866 34334 -26814 34343
rect -26706 34377 -26654 34386
rect -26706 34343 -26697 34377
rect -26697 34343 -26663 34377
rect -26663 34343 -26654 34377
rect -26706 34334 -26654 34343
rect -26546 34377 -26494 34386
rect -26546 34343 -26537 34377
rect -26537 34343 -26503 34377
rect -26503 34343 -26494 34377
rect -26546 34334 -26494 34343
rect -26386 34377 -26334 34386
rect -26386 34343 -26377 34377
rect -26377 34343 -26343 34377
rect -26343 34343 -26334 34377
rect -26386 34334 -26334 34343
rect -26226 34377 -26174 34386
rect -26226 34343 -26217 34377
rect -26217 34343 -26183 34377
rect -26183 34343 -26174 34377
rect -26226 34334 -26174 34343
rect -26066 34377 -26014 34386
rect -26066 34343 -26057 34377
rect -26057 34343 -26023 34377
rect -26023 34343 -26014 34377
rect -26066 34334 -26014 34343
rect -25906 34377 -25854 34386
rect -25906 34343 -25897 34377
rect -25897 34343 -25863 34377
rect -25863 34343 -25854 34377
rect -25906 34334 -25854 34343
rect -25746 34377 -25694 34386
rect -25746 34343 -25737 34377
rect -25737 34343 -25703 34377
rect -25703 34343 -25694 34377
rect -25746 34334 -25694 34343
rect -25586 34377 -25534 34386
rect -25586 34343 -25577 34377
rect -25577 34343 -25543 34377
rect -25543 34343 -25534 34377
rect -25586 34334 -25534 34343
rect -25426 34377 -25374 34386
rect -25426 34343 -25417 34377
rect -25417 34343 -25383 34377
rect -25383 34343 -25374 34377
rect -25426 34334 -25374 34343
rect -25266 34377 -25214 34386
rect -25266 34343 -25257 34377
rect -25257 34343 -25223 34377
rect -25223 34343 -25214 34377
rect -25266 34334 -25214 34343
rect -25106 34377 -25054 34386
rect -25106 34343 -25097 34377
rect -25097 34343 -25063 34377
rect -25063 34343 -25054 34377
rect -25106 34334 -25054 34343
rect -24946 34377 -24894 34386
rect -24946 34343 -24937 34377
rect -24937 34343 -24903 34377
rect -24903 34343 -24894 34377
rect -24946 34334 -24894 34343
rect -24786 34377 -24734 34386
rect -24786 34343 -24777 34377
rect -24777 34343 -24743 34377
rect -24743 34343 -24734 34377
rect -24786 34334 -24734 34343
rect -24626 34377 -24574 34386
rect -24626 34343 -24617 34377
rect -24617 34343 -24583 34377
rect -24583 34343 -24574 34377
rect -24626 34334 -24574 34343
rect -24466 34377 -24414 34386
rect -24466 34343 -24457 34377
rect -24457 34343 -24423 34377
rect -24423 34343 -24414 34377
rect -24466 34334 -24414 34343
rect -24306 34377 -24254 34386
rect -24306 34343 -24297 34377
rect -24297 34343 -24263 34377
rect -24263 34343 -24254 34377
rect -24306 34334 -24254 34343
rect -24146 34377 -24094 34386
rect -24146 34343 -24137 34377
rect -24137 34343 -24103 34377
rect -24103 34343 -24094 34377
rect -24146 34334 -24094 34343
rect -23986 34377 -23934 34386
rect -23986 34343 -23977 34377
rect -23977 34343 -23943 34377
rect -23943 34343 -23934 34377
rect -23986 34334 -23934 34343
rect -23826 34377 -23774 34386
rect -23826 34343 -23817 34377
rect -23817 34343 -23783 34377
rect -23783 34343 -23774 34377
rect -23826 34334 -23774 34343
rect -23666 34377 -23614 34386
rect -23666 34343 -23657 34377
rect -23657 34343 -23623 34377
rect -23623 34343 -23614 34377
rect -23666 34334 -23614 34343
rect -23506 34377 -23454 34386
rect -23506 34343 -23497 34377
rect -23497 34343 -23463 34377
rect -23463 34343 -23454 34377
rect -23506 34334 -23454 34343
rect -23346 34377 -23294 34386
rect -23346 34343 -23337 34377
rect -23337 34343 -23303 34377
rect -23303 34343 -23294 34377
rect -23346 34334 -23294 34343
rect -23186 34377 -23134 34386
rect -23186 34343 -23177 34377
rect -23177 34343 -23143 34377
rect -23143 34343 -23134 34377
rect -23186 34334 -23134 34343
rect -23026 34377 -22974 34386
rect -23026 34343 -23017 34377
rect -23017 34343 -22983 34377
rect -22983 34343 -22974 34377
rect -23026 34334 -22974 34343
rect -22866 34377 -22814 34386
rect -22866 34343 -22857 34377
rect -22857 34343 -22823 34377
rect -22823 34343 -22814 34377
rect -22866 34334 -22814 34343
rect -22706 34377 -22654 34386
rect -22706 34343 -22697 34377
rect -22697 34343 -22663 34377
rect -22663 34343 -22654 34377
rect -22706 34334 -22654 34343
rect -22546 34377 -22494 34386
rect -22546 34343 -22537 34377
rect -22537 34343 -22503 34377
rect -22503 34343 -22494 34377
rect -22546 34334 -22494 34343
rect -22386 34377 -22334 34386
rect -22386 34343 -22377 34377
rect -22377 34343 -22343 34377
rect -22343 34343 -22334 34377
rect -22386 34334 -22334 34343
rect -22226 34377 -22174 34386
rect -22226 34343 -22217 34377
rect -22217 34343 -22183 34377
rect -22183 34343 -22174 34377
rect -22226 34334 -22174 34343
rect -22066 34377 -22014 34386
rect -22066 34343 -22057 34377
rect -22057 34343 -22023 34377
rect -22023 34343 -22014 34377
rect -22066 34334 -22014 34343
rect -21906 34377 -21854 34386
rect -21906 34343 -21897 34377
rect -21897 34343 -21863 34377
rect -21863 34343 -21854 34377
rect -21906 34334 -21854 34343
rect -21746 34377 -21694 34386
rect -21746 34343 -21737 34377
rect -21737 34343 -21703 34377
rect -21703 34343 -21694 34377
rect -21746 34334 -21694 34343
rect -21586 34377 -21534 34386
rect -21586 34343 -21577 34377
rect -21577 34343 -21543 34377
rect -21543 34343 -21534 34377
rect -21586 34334 -21534 34343
rect -21426 34377 -21374 34386
rect -21426 34343 -21417 34377
rect -21417 34343 -21383 34377
rect -21383 34343 -21374 34377
rect -21426 34334 -21374 34343
rect -21266 34377 -21214 34386
rect -21266 34343 -21257 34377
rect -21257 34343 -21223 34377
rect -21223 34343 -21214 34377
rect -21266 34334 -21214 34343
rect -21106 34377 -21054 34386
rect -21106 34343 -21097 34377
rect -21097 34343 -21063 34377
rect -21063 34343 -21054 34377
rect -21106 34334 -21054 34343
rect -20946 34377 -20894 34386
rect -20946 34343 -20937 34377
rect -20937 34343 -20903 34377
rect -20903 34343 -20894 34377
rect -20946 34334 -20894 34343
rect -20786 34377 -20734 34386
rect -20786 34343 -20777 34377
rect -20777 34343 -20743 34377
rect -20743 34343 -20734 34377
rect -20786 34334 -20734 34343
rect -20626 34377 -20574 34386
rect -20626 34343 -20617 34377
rect -20617 34343 -20583 34377
rect -20583 34343 -20574 34377
rect -20626 34334 -20574 34343
rect -20466 34377 -20414 34386
rect -20466 34343 -20457 34377
rect -20457 34343 -20423 34377
rect -20423 34343 -20414 34377
rect -20466 34334 -20414 34343
rect -20306 34377 -20254 34386
rect -20306 34343 -20297 34377
rect -20297 34343 -20263 34377
rect -20263 34343 -20254 34377
rect -20306 34334 -20254 34343
rect -20146 34377 -20094 34386
rect -20146 34343 -20137 34377
rect -20137 34343 -20103 34377
rect -20103 34343 -20094 34377
rect -20146 34334 -20094 34343
rect -19986 34377 -19934 34386
rect -19986 34343 -19977 34377
rect -19977 34343 -19943 34377
rect -19943 34343 -19934 34377
rect -19986 34334 -19934 34343
rect -19826 34377 -19774 34386
rect -19826 34343 -19817 34377
rect -19817 34343 -19783 34377
rect -19783 34343 -19774 34377
rect -19826 34334 -19774 34343
rect -19666 34377 -19614 34386
rect -19666 34343 -19657 34377
rect -19657 34343 -19623 34377
rect -19623 34343 -19614 34377
rect -19666 34334 -19614 34343
rect -19506 34377 -19454 34386
rect -19506 34343 -19497 34377
rect -19497 34343 -19463 34377
rect -19463 34343 -19454 34377
rect -19506 34334 -19454 34343
rect -19346 34377 -19294 34386
rect -19346 34343 -19337 34377
rect -19337 34343 -19303 34377
rect -19303 34343 -19294 34377
rect -19346 34334 -19294 34343
rect -19186 34377 -19134 34386
rect -19186 34343 -19177 34377
rect -19177 34343 -19143 34377
rect -19143 34343 -19134 34377
rect -19186 34334 -19134 34343
rect -19026 34377 -18974 34386
rect -19026 34343 -19017 34377
rect -19017 34343 -18983 34377
rect -18983 34343 -18974 34377
rect -19026 34334 -18974 34343
rect -18866 34377 -18814 34386
rect -18866 34343 -18857 34377
rect -18857 34343 -18823 34377
rect -18823 34343 -18814 34377
rect -18866 34334 -18814 34343
rect -18706 34377 -18654 34386
rect -18706 34343 -18697 34377
rect -18697 34343 -18663 34377
rect -18663 34343 -18654 34377
rect -18706 34334 -18654 34343
rect -18546 34377 -18494 34386
rect -18546 34343 -18537 34377
rect -18537 34343 -18503 34377
rect -18503 34343 -18494 34377
rect -18546 34334 -18494 34343
rect -18386 34377 -18334 34386
rect -18386 34343 -18377 34377
rect -18377 34343 -18343 34377
rect -18343 34343 -18334 34377
rect -18386 34334 -18334 34343
rect -18226 34377 -18174 34386
rect -18226 34343 -18217 34377
rect -18217 34343 -18183 34377
rect -18183 34343 -18174 34377
rect -18226 34334 -18174 34343
rect -18066 34377 -18014 34386
rect -18066 34343 -18057 34377
rect -18057 34343 -18023 34377
rect -18023 34343 -18014 34377
rect -18066 34334 -18014 34343
rect -17906 34377 -17854 34386
rect -17906 34343 -17897 34377
rect -17897 34343 -17863 34377
rect -17863 34343 -17854 34377
rect -17906 34334 -17854 34343
rect -17746 34377 -17694 34386
rect -17746 34343 -17737 34377
rect -17737 34343 -17703 34377
rect -17703 34343 -17694 34377
rect -17746 34334 -17694 34343
rect -17586 34377 -17534 34386
rect -17586 34343 -17577 34377
rect -17577 34343 -17543 34377
rect -17543 34343 -17534 34377
rect -17586 34334 -17534 34343
rect -17426 34377 -17374 34386
rect -17426 34343 -17417 34377
rect -17417 34343 -17383 34377
rect -17383 34343 -17374 34377
rect -17426 34334 -17374 34343
rect -17266 34377 -17214 34386
rect -17266 34343 -17257 34377
rect -17257 34343 -17223 34377
rect -17223 34343 -17214 34377
rect -17266 34334 -17214 34343
rect -17106 34377 -17054 34386
rect -17106 34343 -17097 34377
rect -17097 34343 -17063 34377
rect -17063 34343 -17054 34377
rect -17106 34334 -17054 34343
rect -16946 34377 -16894 34386
rect -16946 34343 -16937 34377
rect -16937 34343 -16903 34377
rect -16903 34343 -16894 34377
rect -16946 34334 -16894 34343
rect -16786 34377 -16734 34386
rect -16786 34343 -16777 34377
rect -16777 34343 -16743 34377
rect -16743 34343 -16734 34377
rect -16786 34334 -16734 34343
rect -16626 34377 -16574 34386
rect -16626 34343 -16617 34377
rect -16617 34343 -16583 34377
rect -16583 34343 -16574 34377
rect -16626 34334 -16574 34343
rect -16466 34377 -16414 34386
rect -16466 34343 -16457 34377
rect -16457 34343 -16423 34377
rect -16423 34343 -16414 34377
rect -16466 34334 -16414 34343
rect -16306 34377 -16254 34386
rect -16306 34343 -16297 34377
rect -16297 34343 -16263 34377
rect -16263 34343 -16254 34377
rect -16306 34334 -16254 34343
rect -16146 34377 -16094 34386
rect -16146 34343 -16137 34377
rect -16137 34343 -16103 34377
rect -16103 34343 -16094 34377
rect -16146 34334 -16094 34343
rect -15986 34377 -15934 34386
rect -15986 34343 -15977 34377
rect -15977 34343 -15943 34377
rect -15943 34343 -15934 34377
rect -15986 34334 -15934 34343
rect -15826 34377 -15774 34386
rect -15826 34343 -15817 34377
rect -15817 34343 -15783 34377
rect -15783 34343 -15774 34377
rect -15826 34334 -15774 34343
rect -15666 34377 -15614 34386
rect -15666 34343 -15657 34377
rect -15657 34343 -15623 34377
rect -15623 34343 -15614 34377
rect -15666 34334 -15614 34343
rect -15506 34377 -15454 34386
rect -15506 34343 -15497 34377
rect -15497 34343 -15463 34377
rect -15463 34343 -15454 34377
rect -15506 34334 -15454 34343
rect -15346 34377 -15294 34386
rect -15346 34343 -15337 34377
rect -15337 34343 -15303 34377
rect -15303 34343 -15294 34377
rect -15346 34334 -15294 34343
rect -15186 34377 -15134 34386
rect -15186 34343 -15177 34377
rect -15177 34343 -15143 34377
rect -15143 34343 -15134 34377
rect -15186 34334 -15134 34343
rect -15026 34377 -14974 34386
rect -15026 34343 -15017 34377
rect -15017 34343 -14983 34377
rect -14983 34343 -14974 34377
rect -15026 34334 -14974 34343
rect -14866 34377 -14814 34386
rect -14866 34343 -14857 34377
rect -14857 34343 -14823 34377
rect -14823 34343 -14814 34377
rect -14866 34334 -14814 34343
rect -14706 34377 -14654 34386
rect -14706 34343 -14697 34377
rect -14697 34343 -14663 34377
rect -14663 34343 -14654 34377
rect -14706 34334 -14654 34343
rect -14546 34377 -14494 34386
rect -14546 34343 -14537 34377
rect -14537 34343 -14503 34377
rect -14503 34343 -14494 34377
rect -14546 34334 -14494 34343
rect -14386 34377 -14334 34386
rect -14386 34343 -14377 34377
rect -14377 34343 -14343 34377
rect -14343 34343 -14334 34377
rect -14386 34334 -14334 34343
rect -14226 34377 -14174 34386
rect -14226 34343 -14217 34377
rect -14217 34343 -14183 34377
rect -14183 34343 -14174 34377
rect -14226 34334 -14174 34343
rect -14066 34377 -14014 34386
rect -14066 34343 -14057 34377
rect -14057 34343 -14023 34377
rect -14023 34343 -14014 34377
rect -14066 34334 -14014 34343
rect -13906 34377 -13854 34386
rect -13906 34343 -13897 34377
rect -13897 34343 -13863 34377
rect -13863 34343 -13854 34377
rect -13906 34334 -13854 34343
rect -13746 34377 -13694 34386
rect -13746 34343 -13737 34377
rect -13737 34343 -13703 34377
rect -13703 34343 -13694 34377
rect -13746 34334 -13694 34343
rect -13586 34377 -13534 34386
rect -13586 34343 -13577 34377
rect -13577 34343 -13543 34377
rect -13543 34343 -13534 34377
rect -13586 34334 -13534 34343
rect -13426 34377 -13374 34386
rect -13426 34343 -13417 34377
rect -13417 34343 -13383 34377
rect -13383 34343 -13374 34377
rect -13426 34334 -13374 34343
rect -13266 34377 -13214 34386
rect -13266 34343 -13257 34377
rect -13257 34343 -13223 34377
rect -13223 34343 -13214 34377
rect -13266 34334 -13214 34343
rect -13106 34377 -13054 34386
rect -13106 34343 -13097 34377
rect -13097 34343 -13063 34377
rect -13063 34343 -13054 34377
rect -13106 34334 -13054 34343
rect -12946 34377 -12894 34386
rect -12946 34343 -12937 34377
rect -12937 34343 -12903 34377
rect -12903 34343 -12894 34377
rect -12946 34334 -12894 34343
rect -12786 34377 -12734 34386
rect -12786 34343 -12777 34377
rect -12777 34343 -12743 34377
rect -12743 34343 -12734 34377
rect -12786 34334 -12734 34343
rect -12626 34377 -12574 34386
rect -12626 34343 -12617 34377
rect -12617 34343 -12583 34377
rect -12583 34343 -12574 34377
rect -12626 34334 -12574 34343
rect -12466 34377 -12414 34386
rect -12466 34343 -12457 34377
rect -12457 34343 -12423 34377
rect -12423 34343 -12414 34377
rect -12466 34334 -12414 34343
rect -12306 34377 -12254 34386
rect -12306 34343 -12297 34377
rect -12297 34343 -12263 34377
rect -12263 34343 -12254 34377
rect -12306 34334 -12254 34343
rect -12146 34377 -12094 34386
rect -12146 34343 -12137 34377
rect -12137 34343 -12103 34377
rect -12103 34343 -12094 34377
rect -12146 34334 -12094 34343
rect -11986 34377 -11934 34386
rect -11986 34343 -11977 34377
rect -11977 34343 -11943 34377
rect -11943 34343 -11934 34377
rect -11986 34334 -11934 34343
rect -11826 34377 -11774 34386
rect -11826 34343 -11817 34377
rect -11817 34343 -11783 34377
rect -11783 34343 -11774 34377
rect -11826 34334 -11774 34343
rect -11666 34377 -11614 34386
rect -11666 34343 -11657 34377
rect -11657 34343 -11623 34377
rect -11623 34343 -11614 34377
rect -11666 34334 -11614 34343
rect -11506 34377 -11454 34386
rect -11506 34343 -11497 34377
rect -11497 34343 -11463 34377
rect -11463 34343 -11454 34377
rect -11506 34334 -11454 34343
rect -10866 34377 -10814 34386
rect -10866 34343 -10857 34377
rect -10857 34343 -10823 34377
rect -10823 34343 -10814 34377
rect -10866 34334 -10814 34343
rect -10546 34377 -10494 34386
rect -10546 34343 -10537 34377
rect -10537 34343 -10503 34377
rect -10503 34343 -10494 34377
rect -10546 34334 -10494 34343
rect -29906 32937 -29854 32946
rect -29906 32903 -29897 32937
rect -29897 32903 -29863 32937
rect -29863 32903 -29854 32937
rect -29906 32894 -29854 32903
rect -29746 32937 -29694 32946
rect -29746 32903 -29737 32937
rect -29737 32903 -29703 32937
rect -29703 32903 -29694 32937
rect -29746 32894 -29694 32903
rect -29586 32937 -29534 32946
rect -29586 32903 -29577 32937
rect -29577 32903 -29543 32937
rect -29543 32903 -29534 32937
rect -29586 32894 -29534 32903
rect -29426 32937 -29374 32946
rect -29426 32903 -29417 32937
rect -29417 32903 -29383 32937
rect -29383 32903 -29374 32937
rect -29426 32894 -29374 32903
rect -29266 32937 -29214 32946
rect -29266 32903 -29257 32937
rect -29257 32903 -29223 32937
rect -29223 32903 -29214 32937
rect -29266 32894 -29214 32903
rect -29106 32937 -29054 32946
rect -29106 32903 -29097 32937
rect -29097 32903 -29063 32937
rect -29063 32903 -29054 32937
rect -29106 32894 -29054 32903
rect -28946 32937 -28894 32946
rect -28946 32903 -28937 32937
rect -28937 32903 -28903 32937
rect -28903 32903 -28894 32937
rect -28946 32894 -28894 32903
rect -28786 32937 -28734 32946
rect -28786 32903 -28777 32937
rect -28777 32903 -28743 32937
rect -28743 32903 -28734 32937
rect -28786 32894 -28734 32903
rect -28626 32937 -28574 32946
rect -28626 32903 -28617 32937
rect -28617 32903 -28583 32937
rect -28583 32903 -28574 32937
rect -28626 32894 -28574 32903
rect -28466 32937 -28414 32946
rect -28466 32903 -28457 32937
rect -28457 32903 -28423 32937
rect -28423 32903 -28414 32937
rect -28466 32894 -28414 32903
rect -28306 32937 -28254 32946
rect -28306 32903 -28297 32937
rect -28297 32903 -28263 32937
rect -28263 32903 -28254 32937
rect -28306 32894 -28254 32903
rect -28146 32937 -28094 32946
rect -28146 32903 -28137 32937
rect -28137 32903 -28103 32937
rect -28103 32903 -28094 32937
rect -28146 32894 -28094 32903
rect -27986 32937 -27934 32946
rect -27986 32903 -27977 32937
rect -27977 32903 -27943 32937
rect -27943 32903 -27934 32937
rect -27986 32894 -27934 32903
rect -27826 32937 -27774 32946
rect -27826 32903 -27817 32937
rect -27817 32903 -27783 32937
rect -27783 32903 -27774 32937
rect -27826 32894 -27774 32903
rect -27666 32937 -27614 32946
rect -27666 32903 -27657 32937
rect -27657 32903 -27623 32937
rect -27623 32903 -27614 32937
rect -27666 32894 -27614 32903
rect -27506 32937 -27454 32946
rect -27506 32903 -27497 32937
rect -27497 32903 -27463 32937
rect -27463 32903 -27454 32937
rect -27506 32894 -27454 32903
rect -27346 32937 -27294 32946
rect -27346 32903 -27337 32937
rect -27337 32903 -27303 32937
rect -27303 32903 -27294 32937
rect -27346 32894 -27294 32903
rect -27186 32937 -27134 32946
rect -27186 32903 -27177 32937
rect -27177 32903 -27143 32937
rect -27143 32903 -27134 32937
rect -27186 32894 -27134 32903
rect -27026 32937 -26974 32946
rect -27026 32903 -27017 32937
rect -27017 32903 -26983 32937
rect -26983 32903 -26974 32937
rect -27026 32894 -26974 32903
rect -26866 32937 -26814 32946
rect -26866 32903 -26857 32937
rect -26857 32903 -26823 32937
rect -26823 32903 -26814 32937
rect -26866 32894 -26814 32903
rect -26706 32937 -26654 32946
rect -26706 32903 -26697 32937
rect -26697 32903 -26663 32937
rect -26663 32903 -26654 32937
rect -26706 32894 -26654 32903
rect -26546 32937 -26494 32946
rect -26546 32903 -26537 32937
rect -26537 32903 -26503 32937
rect -26503 32903 -26494 32937
rect -26546 32894 -26494 32903
rect -26386 32937 -26334 32946
rect -26386 32903 -26377 32937
rect -26377 32903 -26343 32937
rect -26343 32903 -26334 32937
rect -26386 32894 -26334 32903
rect -26226 32937 -26174 32946
rect -26226 32903 -26217 32937
rect -26217 32903 -26183 32937
rect -26183 32903 -26174 32937
rect -26226 32894 -26174 32903
rect -26066 32937 -26014 32946
rect -26066 32903 -26057 32937
rect -26057 32903 -26023 32937
rect -26023 32903 -26014 32937
rect -26066 32894 -26014 32903
rect -25906 32937 -25854 32946
rect -25906 32903 -25897 32937
rect -25897 32903 -25863 32937
rect -25863 32903 -25854 32937
rect -25906 32894 -25854 32903
rect -25746 32937 -25694 32946
rect -25746 32903 -25737 32937
rect -25737 32903 -25703 32937
rect -25703 32903 -25694 32937
rect -25746 32894 -25694 32903
rect -25586 32937 -25534 32946
rect -25586 32903 -25577 32937
rect -25577 32903 -25543 32937
rect -25543 32903 -25534 32937
rect -25586 32894 -25534 32903
rect -25426 32937 -25374 32946
rect -25426 32903 -25417 32937
rect -25417 32903 -25383 32937
rect -25383 32903 -25374 32937
rect -25426 32894 -25374 32903
rect -25266 32937 -25214 32946
rect -25266 32903 -25257 32937
rect -25257 32903 -25223 32937
rect -25223 32903 -25214 32937
rect -25266 32894 -25214 32903
rect -25106 32937 -25054 32946
rect -25106 32903 -25097 32937
rect -25097 32903 -25063 32937
rect -25063 32903 -25054 32937
rect -25106 32894 -25054 32903
rect -24946 32937 -24894 32946
rect -24946 32903 -24937 32937
rect -24937 32903 -24903 32937
rect -24903 32903 -24894 32937
rect -24946 32894 -24894 32903
rect -24786 32937 -24734 32946
rect -24786 32903 -24777 32937
rect -24777 32903 -24743 32937
rect -24743 32903 -24734 32937
rect -24786 32894 -24734 32903
rect -24626 32937 -24574 32946
rect -24626 32903 -24617 32937
rect -24617 32903 -24583 32937
rect -24583 32903 -24574 32937
rect -24626 32894 -24574 32903
rect -24466 32937 -24414 32946
rect -24466 32903 -24457 32937
rect -24457 32903 -24423 32937
rect -24423 32903 -24414 32937
rect -24466 32894 -24414 32903
rect -24306 32937 -24254 32946
rect -24306 32903 -24297 32937
rect -24297 32903 -24263 32937
rect -24263 32903 -24254 32937
rect -24306 32894 -24254 32903
rect -24146 32937 -24094 32946
rect -24146 32903 -24137 32937
rect -24137 32903 -24103 32937
rect -24103 32903 -24094 32937
rect -24146 32894 -24094 32903
rect -23986 32937 -23934 32946
rect -23986 32903 -23977 32937
rect -23977 32903 -23943 32937
rect -23943 32903 -23934 32937
rect -23986 32894 -23934 32903
rect -23826 32937 -23774 32946
rect -23826 32903 -23817 32937
rect -23817 32903 -23783 32937
rect -23783 32903 -23774 32937
rect -23826 32894 -23774 32903
rect -23666 32937 -23614 32946
rect -23666 32903 -23657 32937
rect -23657 32903 -23623 32937
rect -23623 32903 -23614 32937
rect -23666 32894 -23614 32903
rect -23506 32937 -23454 32946
rect -23506 32903 -23497 32937
rect -23497 32903 -23463 32937
rect -23463 32903 -23454 32937
rect -23506 32894 -23454 32903
rect -23346 32937 -23294 32946
rect -23346 32903 -23337 32937
rect -23337 32903 -23303 32937
rect -23303 32903 -23294 32937
rect -23346 32894 -23294 32903
rect -23186 32937 -23134 32946
rect -23186 32903 -23177 32937
rect -23177 32903 -23143 32937
rect -23143 32903 -23134 32937
rect -23186 32894 -23134 32903
rect -23026 32937 -22974 32946
rect -23026 32903 -23017 32937
rect -23017 32903 -22983 32937
rect -22983 32903 -22974 32937
rect -23026 32894 -22974 32903
rect -22866 32937 -22814 32946
rect -22866 32903 -22857 32937
rect -22857 32903 -22823 32937
rect -22823 32903 -22814 32937
rect -22866 32894 -22814 32903
rect -22706 32937 -22654 32946
rect -22706 32903 -22697 32937
rect -22697 32903 -22663 32937
rect -22663 32903 -22654 32937
rect -22706 32894 -22654 32903
rect -22546 32937 -22494 32946
rect -22546 32903 -22537 32937
rect -22537 32903 -22503 32937
rect -22503 32903 -22494 32937
rect -22546 32894 -22494 32903
rect -22386 32937 -22334 32946
rect -22386 32903 -22377 32937
rect -22377 32903 -22343 32937
rect -22343 32903 -22334 32937
rect -22386 32894 -22334 32903
rect -22226 32937 -22174 32946
rect -22226 32903 -22217 32937
rect -22217 32903 -22183 32937
rect -22183 32903 -22174 32937
rect -22226 32894 -22174 32903
rect -22066 32937 -22014 32946
rect -22066 32903 -22057 32937
rect -22057 32903 -22023 32937
rect -22023 32903 -22014 32937
rect -22066 32894 -22014 32903
rect -21906 32937 -21854 32946
rect -21906 32903 -21897 32937
rect -21897 32903 -21863 32937
rect -21863 32903 -21854 32937
rect -21906 32894 -21854 32903
rect -21746 32937 -21694 32946
rect -21746 32903 -21737 32937
rect -21737 32903 -21703 32937
rect -21703 32903 -21694 32937
rect -21746 32894 -21694 32903
rect -21586 32937 -21534 32946
rect -21586 32903 -21577 32937
rect -21577 32903 -21543 32937
rect -21543 32903 -21534 32937
rect -21586 32894 -21534 32903
rect -21426 32937 -21374 32946
rect -21426 32903 -21417 32937
rect -21417 32903 -21383 32937
rect -21383 32903 -21374 32937
rect -21426 32894 -21374 32903
rect -21266 32937 -21214 32946
rect -21266 32903 -21257 32937
rect -21257 32903 -21223 32937
rect -21223 32903 -21214 32937
rect -21266 32894 -21214 32903
rect -21106 32937 -21054 32946
rect -21106 32903 -21097 32937
rect -21097 32903 -21063 32937
rect -21063 32903 -21054 32937
rect -21106 32894 -21054 32903
rect -20946 32937 -20894 32946
rect -20946 32903 -20937 32937
rect -20937 32903 -20903 32937
rect -20903 32903 -20894 32937
rect -20946 32894 -20894 32903
rect -20786 32937 -20734 32946
rect -20786 32903 -20777 32937
rect -20777 32903 -20743 32937
rect -20743 32903 -20734 32937
rect -20786 32894 -20734 32903
rect -20626 32937 -20574 32946
rect -20626 32903 -20617 32937
rect -20617 32903 -20583 32937
rect -20583 32903 -20574 32937
rect -20626 32894 -20574 32903
rect -20466 32937 -20414 32946
rect -20466 32903 -20457 32937
rect -20457 32903 -20423 32937
rect -20423 32903 -20414 32937
rect -20466 32894 -20414 32903
rect -20306 32937 -20254 32946
rect -20306 32903 -20297 32937
rect -20297 32903 -20263 32937
rect -20263 32903 -20254 32937
rect -20306 32894 -20254 32903
rect -20146 32937 -20094 32946
rect -20146 32903 -20137 32937
rect -20137 32903 -20103 32937
rect -20103 32903 -20094 32937
rect -20146 32894 -20094 32903
rect -19986 32937 -19934 32946
rect -19986 32903 -19977 32937
rect -19977 32903 -19943 32937
rect -19943 32903 -19934 32937
rect -19986 32894 -19934 32903
rect -19826 32937 -19774 32946
rect -19826 32903 -19817 32937
rect -19817 32903 -19783 32937
rect -19783 32903 -19774 32937
rect -19826 32894 -19774 32903
rect -19666 32937 -19614 32946
rect -19666 32903 -19657 32937
rect -19657 32903 -19623 32937
rect -19623 32903 -19614 32937
rect -19666 32894 -19614 32903
rect -19506 32937 -19454 32946
rect -19506 32903 -19497 32937
rect -19497 32903 -19463 32937
rect -19463 32903 -19454 32937
rect -19506 32894 -19454 32903
rect -19346 32937 -19294 32946
rect -19346 32903 -19337 32937
rect -19337 32903 -19303 32937
rect -19303 32903 -19294 32937
rect -19346 32894 -19294 32903
rect -19186 32937 -19134 32946
rect -19186 32903 -19177 32937
rect -19177 32903 -19143 32937
rect -19143 32903 -19134 32937
rect -19186 32894 -19134 32903
rect -19026 32937 -18974 32946
rect -19026 32903 -19017 32937
rect -19017 32903 -18983 32937
rect -18983 32903 -18974 32937
rect -19026 32894 -18974 32903
rect -18866 32937 -18814 32946
rect -18866 32903 -18857 32937
rect -18857 32903 -18823 32937
rect -18823 32903 -18814 32937
rect -18866 32894 -18814 32903
rect -18706 32937 -18654 32946
rect -18706 32903 -18697 32937
rect -18697 32903 -18663 32937
rect -18663 32903 -18654 32937
rect -18706 32894 -18654 32903
rect -18546 32937 -18494 32946
rect -18546 32903 -18537 32937
rect -18537 32903 -18503 32937
rect -18503 32903 -18494 32937
rect -18546 32894 -18494 32903
rect -18386 32937 -18334 32946
rect -18386 32903 -18377 32937
rect -18377 32903 -18343 32937
rect -18343 32903 -18334 32937
rect -18386 32894 -18334 32903
rect -18226 32937 -18174 32946
rect -18226 32903 -18217 32937
rect -18217 32903 -18183 32937
rect -18183 32903 -18174 32937
rect -18226 32894 -18174 32903
rect -18066 32937 -18014 32946
rect -18066 32903 -18057 32937
rect -18057 32903 -18023 32937
rect -18023 32903 -18014 32937
rect -18066 32894 -18014 32903
rect -17906 32937 -17854 32946
rect -17906 32903 -17897 32937
rect -17897 32903 -17863 32937
rect -17863 32903 -17854 32937
rect -17906 32894 -17854 32903
rect -17746 32937 -17694 32946
rect -17746 32903 -17737 32937
rect -17737 32903 -17703 32937
rect -17703 32903 -17694 32937
rect -17746 32894 -17694 32903
rect -17586 32937 -17534 32946
rect -17586 32903 -17577 32937
rect -17577 32903 -17543 32937
rect -17543 32903 -17534 32937
rect -17586 32894 -17534 32903
rect -17426 32937 -17374 32946
rect -17426 32903 -17417 32937
rect -17417 32903 -17383 32937
rect -17383 32903 -17374 32937
rect -17426 32894 -17374 32903
rect -17266 32937 -17214 32946
rect -17266 32903 -17257 32937
rect -17257 32903 -17223 32937
rect -17223 32903 -17214 32937
rect -17266 32894 -17214 32903
rect -17106 32937 -17054 32946
rect -17106 32903 -17097 32937
rect -17097 32903 -17063 32937
rect -17063 32903 -17054 32937
rect -17106 32894 -17054 32903
rect -16946 32937 -16894 32946
rect -16946 32903 -16937 32937
rect -16937 32903 -16903 32937
rect -16903 32903 -16894 32937
rect -16946 32894 -16894 32903
rect -16786 32937 -16734 32946
rect -16786 32903 -16777 32937
rect -16777 32903 -16743 32937
rect -16743 32903 -16734 32937
rect -16786 32894 -16734 32903
rect -16626 32937 -16574 32946
rect -16626 32903 -16617 32937
rect -16617 32903 -16583 32937
rect -16583 32903 -16574 32937
rect -16626 32894 -16574 32903
rect -16466 32937 -16414 32946
rect -16466 32903 -16457 32937
rect -16457 32903 -16423 32937
rect -16423 32903 -16414 32937
rect -16466 32894 -16414 32903
rect -16306 32937 -16254 32946
rect -16306 32903 -16297 32937
rect -16297 32903 -16263 32937
rect -16263 32903 -16254 32937
rect -16306 32894 -16254 32903
rect -16146 32937 -16094 32946
rect -16146 32903 -16137 32937
rect -16137 32903 -16103 32937
rect -16103 32903 -16094 32937
rect -16146 32894 -16094 32903
rect -15986 32937 -15934 32946
rect -15986 32903 -15977 32937
rect -15977 32903 -15943 32937
rect -15943 32903 -15934 32937
rect -15986 32894 -15934 32903
rect -15826 32937 -15774 32946
rect -15826 32903 -15817 32937
rect -15817 32903 -15783 32937
rect -15783 32903 -15774 32937
rect -15826 32894 -15774 32903
rect -15666 32937 -15614 32946
rect -15666 32903 -15657 32937
rect -15657 32903 -15623 32937
rect -15623 32903 -15614 32937
rect -15666 32894 -15614 32903
rect -15506 32937 -15454 32946
rect -15506 32903 -15497 32937
rect -15497 32903 -15463 32937
rect -15463 32903 -15454 32937
rect -15506 32894 -15454 32903
rect -15346 32937 -15294 32946
rect -15346 32903 -15337 32937
rect -15337 32903 -15303 32937
rect -15303 32903 -15294 32937
rect -15346 32894 -15294 32903
rect -15186 32937 -15134 32946
rect -15186 32903 -15177 32937
rect -15177 32903 -15143 32937
rect -15143 32903 -15134 32937
rect -15186 32894 -15134 32903
rect -15026 32937 -14974 32946
rect -15026 32903 -15017 32937
rect -15017 32903 -14983 32937
rect -14983 32903 -14974 32937
rect -15026 32894 -14974 32903
rect -14866 32937 -14814 32946
rect -14866 32903 -14857 32937
rect -14857 32903 -14823 32937
rect -14823 32903 -14814 32937
rect -14866 32894 -14814 32903
rect -14706 32937 -14654 32946
rect -14706 32903 -14697 32937
rect -14697 32903 -14663 32937
rect -14663 32903 -14654 32937
rect -14706 32894 -14654 32903
rect -14546 32937 -14494 32946
rect -14546 32903 -14537 32937
rect -14537 32903 -14503 32937
rect -14503 32903 -14494 32937
rect -14546 32894 -14494 32903
rect -14386 32937 -14334 32946
rect -14386 32903 -14377 32937
rect -14377 32903 -14343 32937
rect -14343 32903 -14334 32937
rect -14386 32894 -14334 32903
rect -14226 32937 -14174 32946
rect -14226 32903 -14217 32937
rect -14217 32903 -14183 32937
rect -14183 32903 -14174 32937
rect -14226 32894 -14174 32903
rect -14066 32937 -14014 32946
rect -14066 32903 -14057 32937
rect -14057 32903 -14023 32937
rect -14023 32903 -14014 32937
rect -14066 32894 -14014 32903
rect -13906 32937 -13854 32946
rect -13906 32903 -13897 32937
rect -13897 32903 -13863 32937
rect -13863 32903 -13854 32937
rect -13906 32894 -13854 32903
rect -13746 32937 -13694 32946
rect -13746 32903 -13737 32937
rect -13737 32903 -13703 32937
rect -13703 32903 -13694 32937
rect -13746 32894 -13694 32903
rect -13586 32937 -13534 32946
rect -13586 32903 -13577 32937
rect -13577 32903 -13543 32937
rect -13543 32903 -13534 32937
rect -13586 32894 -13534 32903
rect -13426 32937 -13374 32946
rect -13426 32903 -13417 32937
rect -13417 32903 -13383 32937
rect -13383 32903 -13374 32937
rect -13426 32894 -13374 32903
rect -13266 32937 -13214 32946
rect -13266 32903 -13257 32937
rect -13257 32903 -13223 32937
rect -13223 32903 -13214 32937
rect -13266 32894 -13214 32903
rect -13106 32937 -13054 32946
rect -13106 32903 -13097 32937
rect -13097 32903 -13063 32937
rect -13063 32903 -13054 32937
rect -13106 32894 -13054 32903
rect -12946 32937 -12894 32946
rect -12946 32903 -12937 32937
rect -12937 32903 -12903 32937
rect -12903 32903 -12894 32937
rect -12946 32894 -12894 32903
rect -12786 32937 -12734 32946
rect -12786 32903 -12777 32937
rect -12777 32903 -12743 32937
rect -12743 32903 -12734 32937
rect -12786 32894 -12734 32903
rect -12626 32937 -12574 32946
rect -12626 32903 -12617 32937
rect -12617 32903 -12583 32937
rect -12583 32903 -12574 32937
rect -12626 32894 -12574 32903
rect -12466 32937 -12414 32946
rect -12466 32903 -12457 32937
rect -12457 32903 -12423 32937
rect -12423 32903 -12414 32937
rect -12466 32894 -12414 32903
rect -12306 32937 -12254 32946
rect -12306 32903 -12297 32937
rect -12297 32903 -12263 32937
rect -12263 32903 -12254 32937
rect -12306 32894 -12254 32903
rect -12146 32937 -12094 32946
rect -12146 32903 -12137 32937
rect -12137 32903 -12103 32937
rect -12103 32903 -12094 32937
rect -12146 32894 -12094 32903
rect -11986 32937 -11934 32946
rect -11986 32903 -11977 32937
rect -11977 32903 -11943 32937
rect -11943 32903 -11934 32937
rect -11986 32894 -11934 32903
rect -11826 32937 -11774 32946
rect -11826 32903 -11817 32937
rect -11817 32903 -11783 32937
rect -11783 32903 -11774 32937
rect -11826 32894 -11774 32903
rect -11666 32937 -11614 32946
rect -11666 32903 -11657 32937
rect -11657 32903 -11623 32937
rect -11623 32903 -11614 32937
rect -11666 32894 -11614 32903
rect -11506 32937 -11454 32946
rect -11506 32903 -11497 32937
rect -11497 32903 -11463 32937
rect -11463 32903 -11454 32937
rect -11506 32894 -11454 32903
rect -11186 32937 -11134 32946
rect -11186 32903 -11177 32937
rect -11177 32903 -11143 32937
rect -11143 32903 -11134 32937
rect -11186 32894 -11134 32903
rect -10866 32937 -10814 32946
rect -10866 32903 -10857 32937
rect -10857 32903 -10823 32937
rect -10823 32903 -10814 32937
rect -10866 32894 -10814 32903
rect -10706 32937 -10654 32946
rect -10706 32903 -10697 32937
rect -10697 32903 -10663 32937
rect -10663 32903 -10654 32937
rect -10706 32894 -10654 32903
rect -10546 32937 -10494 32946
rect -10546 32903 -10537 32937
rect -10537 32903 -10503 32937
rect -10503 32903 -10494 32937
rect -10546 32894 -10494 32903
rect -10386 32937 -10334 32946
rect -10386 32903 -10377 32937
rect -10377 32903 -10343 32937
rect -10343 32903 -10334 32937
rect -10386 32894 -10334 32903
rect -10226 32937 -10174 32946
rect -10226 32903 -10217 32937
rect -10217 32903 -10183 32937
rect -10183 32903 -10174 32937
rect -10226 32894 -10174 32903
rect -10066 32937 -10014 32946
rect -10066 32903 -10057 32937
rect -10057 32903 -10023 32937
rect -10023 32903 -10014 32937
rect -10066 32894 -10014 32903
rect -9906 32937 -9854 32946
rect -9906 32903 -9897 32937
rect -9897 32903 -9863 32937
rect -9863 32903 -9854 32937
rect -9906 32894 -9854 32903
rect -9746 32937 -9694 32946
rect -9746 32903 -9737 32937
rect -9737 32903 -9703 32937
rect -9703 32903 -9694 32937
rect -9746 32894 -9694 32903
rect -9586 32937 -9534 32946
rect -9586 32903 -9577 32937
rect -9577 32903 -9543 32937
rect -9543 32903 -9534 32937
rect -9586 32894 -9534 32903
rect -9426 32937 -9374 32946
rect -9426 32903 -9417 32937
rect -9417 32903 -9383 32937
rect -9383 32903 -9374 32937
rect -9426 32894 -9374 32903
rect -9266 32937 -9214 32946
rect -9266 32903 -9257 32937
rect -9257 32903 -9223 32937
rect -9223 32903 -9214 32937
rect -9266 32894 -9214 32903
rect -9106 32937 -9054 32946
rect -9106 32903 -9097 32937
rect -9097 32903 -9063 32937
rect -9063 32903 -9054 32937
rect -9106 32894 -9054 32903
rect -8946 32937 -8894 32946
rect -8946 32903 -8937 32937
rect -8937 32903 -8903 32937
rect -8903 32903 -8894 32937
rect -8946 32894 -8894 32903
rect -8786 32937 -8734 32946
rect -8786 32903 -8777 32937
rect -8777 32903 -8743 32937
rect -8743 32903 -8734 32937
rect -8786 32894 -8734 32903
rect -8626 32937 -8574 32946
rect -8626 32903 -8617 32937
rect -8617 32903 -8583 32937
rect -8583 32903 -8574 32937
rect -8626 32894 -8574 32903
rect -8466 32937 -8414 32946
rect -8466 32903 -8457 32937
rect -8457 32903 -8423 32937
rect -8423 32903 -8414 32937
rect -8466 32894 -8414 32903
rect -8306 32937 -8254 32946
rect -8306 32903 -8297 32937
rect -8297 32903 -8263 32937
rect -8263 32903 -8254 32937
rect -8306 32894 -8254 32903
rect -8146 32937 -8094 32946
rect -8146 32903 -8137 32937
rect -8137 32903 -8103 32937
rect -8103 32903 -8094 32937
rect -8146 32894 -8094 32903
rect -7986 32937 -7934 32946
rect -7986 32903 -7977 32937
rect -7977 32903 -7943 32937
rect -7943 32903 -7934 32937
rect -7986 32894 -7934 32903
rect -7826 32937 -7774 32946
rect -7826 32903 -7817 32937
rect -7817 32903 -7783 32937
rect -7783 32903 -7774 32937
rect -7826 32894 -7774 32903
rect -7666 32937 -7614 32946
rect -7666 32903 -7657 32937
rect -7657 32903 -7623 32937
rect -7623 32903 -7614 32937
rect -7666 32894 -7614 32903
rect -7506 32937 -7454 32946
rect -7506 32903 -7497 32937
rect -7497 32903 -7463 32937
rect -7463 32903 -7454 32937
rect -7506 32894 -7454 32903
rect -7346 32937 -7294 32946
rect -7346 32903 -7337 32937
rect -7337 32903 -7303 32937
rect -7303 32903 -7294 32937
rect -7346 32894 -7294 32903
rect -7186 32937 -7134 32946
rect -7186 32903 -7177 32937
rect -7177 32903 -7143 32937
rect -7143 32903 -7134 32937
rect -7186 32894 -7134 32903
rect -7026 32937 -6974 32946
rect -7026 32903 -7017 32937
rect -7017 32903 -6983 32937
rect -6983 32903 -6974 32937
rect -7026 32894 -6974 32903
rect -6866 32937 -6814 32946
rect -6866 32903 -6857 32937
rect -6857 32903 -6823 32937
rect -6823 32903 -6814 32937
rect -6866 32894 -6814 32903
rect -6706 32937 -6654 32946
rect -6706 32903 -6697 32937
rect -6697 32903 -6663 32937
rect -6663 32903 -6654 32937
rect -6706 32894 -6654 32903
rect -6546 32937 -6494 32946
rect -6546 32903 -6537 32937
rect -6537 32903 -6503 32937
rect -6503 32903 -6494 32937
rect -6546 32894 -6494 32903
rect -6386 32937 -6334 32946
rect -6386 32903 -6377 32937
rect -6377 32903 -6343 32937
rect -6343 32903 -6334 32937
rect -6386 32894 -6334 32903
rect -6226 32937 -6174 32946
rect -6226 32903 -6217 32937
rect -6217 32903 -6183 32937
rect -6183 32903 -6174 32937
rect -6226 32894 -6174 32903
rect -6066 32937 -6014 32946
rect -6066 32903 -6057 32937
rect -6057 32903 -6023 32937
rect -6023 32903 -6014 32937
rect -6066 32894 -6014 32903
rect -5906 32937 -5854 32946
rect -5906 32903 -5897 32937
rect -5897 32903 -5863 32937
rect -5863 32903 -5854 32937
rect -5906 32894 -5854 32903
rect -5746 32937 -5694 32946
rect -5746 32903 -5737 32937
rect -5737 32903 -5703 32937
rect -5703 32903 -5694 32937
rect -5746 32894 -5694 32903
rect -5586 32937 -5534 32946
rect -5586 32903 -5577 32937
rect -5577 32903 -5543 32937
rect -5543 32903 -5534 32937
rect -5586 32894 -5534 32903
rect -5426 32937 -5374 32946
rect -5426 32903 -5417 32937
rect -5417 32903 -5383 32937
rect -5383 32903 -5374 32937
rect -5426 32894 -5374 32903
rect -5266 32937 -5214 32946
rect -5266 32903 -5257 32937
rect -5257 32903 -5223 32937
rect -5223 32903 -5214 32937
rect -5266 32894 -5214 32903
rect -5106 32937 -5054 32946
rect -5106 32903 -5097 32937
rect -5097 32903 -5063 32937
rect -5063 32903 -5054 32937
rect -5106 32894 -5054 32903
rect -4946 32937 -4894 32946
rect -4946 32903 -4937 32937
rect -4937 32903 -4903 32937
rect -4903 32903 -4894 32937
rect -4946 32894 -4894 32903
rect -4786 32937 -4734 32946
rect -4786 32903 -4777 32937
rect -4777 32903 -4743 32937
rect -4743 32903 -4734 32937
rect -4786 32894 -4734 32903
rect -4626 32937 -4574 32946
rect -4626 32903 -4617 32937
rect -4617 32903 -4583 32937
rect -4583 32903 -4574 32937
rect -4626 32894 -4574 32903
rect -4466 32937 -4414 32946
rect -4466 32903 -4457 32937
rect -4457 32903 -4423 32937
rect -4423 32903 -4414 32937
rect -4466 32894 -4414 32903
rect -4306 32937 -4254 32946
rect -4306 32903 -4297 32937
rect -4297 32903 -4263 32937
rect -4263 32903 -4254 32937
rect -4306 32894 -4254 32903
rect -4146 32937 -4094 32946
rect -4146 32903 -4137 32937
rect -4137 32903 -4103 32937
rect -4103 32903 -4094 32937
rect -4146 32894 -4094 32903
rect -3986 32937 -3934 32946
rect -3986 32903 -3977 32937
rect -3977 32903 -3943 32937
rect -3943 32903 -3934 32937
rect -3986 32894 -3934 32903
rect -3666 32937 -3614 32946
rect -3666 32903 -3657 32937
rect -3657 32903 -3623 32937
rect -3623 32903 -3614 32937
rect -3666 32894 -3614 32903
rect -3506 32937 -3454 32946
rect -3506 32903 -3497 32937
rect -3497 32903 -3463 32937
rect -3463 32903 -3454 32937
rect -3506 32894 -3454 32903
rect -3346 32937 -3294 32946
rect -3346 32903 -3337 32937
rect -3337 32903 -3303 32937
rect -3303 32903 -3294 32937
rect -3346 32894 -3294 32903
rect -3186 32937 -3134 32946
rect -3186 32903 -3177 32937
rect -3177 32903 -3143 32937
rect -3143 32903 -3134 32937
rect -3186 32894 -3134 32903
rect -3026 32937 -2974 32946
rect -3026 32903 -3017 32937
rect -3017 32903 -2983 32937
rect -2983 32903 -2974 32937
rect -3026 32894 -2974 32903
rect -2866 32937 -2814 32946
rect -2866 32903 -2857 32937
rect -2857 32903 -2823 32937
rect -2823 32903 -2814 32937
rect -2866 32894 -2814 32903
rect -2706 32937 -2654 32946
rect -2706 32903 -2697 32937
rect -2697 32903 -2663 32937
rect -2663 32903 -2654 32937
rect -2706 32894 -2654 32903
rect -2386 32937 -2334 32946
rect -2386 32903 -2377 32937
rect -2377 32903 -2343 32937
rect -2343 32903 -2334 32937
rect -2386 32894 -2334 32903
rect -2066 32937 -2014 32946
rect -2066 32903 -2057 32937
rect -2057 32903 -2023 32937
rect -2023 32903 -2014 32937
rect -2066 32894 -2014 32903
rect -1746 32937 -1694 32946
rect -1746 32903 -1737 32937
rect -1737 32903 -1703 32937
rect -1703 32903 -1694 32937
rect -1746 32894 -1694 32903
rect -1426 32937 -1374 32946
rect -1426 32903 -1417 32937
rect -1417 32903 -1383 32937
rect -1383 32903 -1374 32937
rect -1426 32894 -1374 32903
rect -1106 32937 -1054 32946
rect -1106 32903 -1097 32937
rect -1097 32903 -1063 32937
rect -1063 32903 -1054 32937
rect -1106 32894 -1054 32903
rect -29906 32617 -29854 32626
rect -29906 32583 -29897 32617
rect -29897 32583 -29863 32617
rect -29863 32583 -29854 32617
rect -29906 32574 -29854 32583
rect -29746 32617 -29694 32626
rect -29746 32583 -29737 32617
rect -29737 32583 -29703 32617
rect -29703 32583 -29694 32617
rect -29746 32574 -29694 32583
rect -29586 32617 -29534 32626
rect -29586 32583 -29577 32617
rect -29577 32583 -29543 32617
rect -29543 32583 -29534 32617
rect -29586 32574 -29534 32583
rect -29426 32617 -29374 32626
rect -29426 32583 -29417 32617
rect -29417 32583 -29383 32617
rect -29383 32583 -29374 32617
rect -29426 32574 -29374 32583
rect -29266 32617 -29214 32626
rect -29266 32583 -29257 32617
rect -29257 32583 -29223 32617
rect -29223 32583 -29214 32617
rect -29266 32574 -29214 32583
rect -29106 32617 -29054 32626
rect -29106 32583 -29097 32617
rect -29097 32583 -29063 32617
rect -29063 32583 -29054 32617
rect -29106 32574 -29054 32583
rect -28946 32617 -28894 32626
rect -28946 32583 -28937 32617
rect -28937 32583 -28903 32617
rect -28903 32583 -28894 32617
rect -28946 32574 -28894 32583
rect -28786 32617 -28734 32626
rect -28786 32583 -28777 32617
rect -28777 32583 -28743 32617
rect -28743 32583 -28734 32617
rect -28786 32574 -28734 32583
rect -28626 32617 -28574 32626
rect -28626 32583 -28617 32617
rect -28617 32583 -28583 32617
rect -28583 32583 -28574 32617
rect -28626 32574 -28574 32583
rect -28466 32617 -28414 32626
rect -28466 32583 -28457 32617
rect -28457 32583 -28423 32617
rect -28423 32583 -28414 32617
rect -28466 32574 -28414 32583
rect -28306 32617 -28254 32626
rect -28306 32583 -28297 32617
rect -28297 32583 -28263 32617
rect -28263 32583 -28254 32617
rect -28306 32574 -28254 32583
rect -28146 32617 -28094 32626
rect -28146 32583 -28137 32617
rect -28137 32583 -28103 32617
rect -28103 32583 -28094 32617
rect -28146 32574 -28094 32583
rect -27986 32617 -27934 32626
rect -27986 32583 -27977 32617
rect -27977 32583 -27943 32617
rect -27943 32583 -27934 32617
rect -27986 32574 -27934 32583
rect -27826 32617 -27774 32626
rect -27826 32583 -27817 32617
rect -27817 32583 -27783 32617
rect -27783 32583 -27774 32617
rect -27826 32574 -27774 32583
rect -27666 32617 -27614 32626
rect -27666 32583 -27657 32617
rect -27657 32583 -27623 32617
rect -27623 32583 -27614 32617
rect -27666 32574 -27614 32583
rect -27506 32617 -27454 32626
rect -27506 32583 -27497 32617
rect -27497 32583 -27463 32617
rect -27463 32583 -27454 32617
rect -27506 32574 -27454 32583
rect -27346 32617 -27294 32626
rect -27346 32583 -27337 32617
rect -27337 32583 -27303 32617
rect -27303 32583 -27294 32617
rect -27346 32574 -27294 32583
rect -27186 32617 -27134 32626
rect -27186 32583 -27177 32617
rect -27177 32583 -27143 32617
rect -27143 32583 -27134 32617
rect -27186 32574 -27134 32583
rect -27026 32617 -26974 32626
rect -27026 32583 -27017 32617
rect -27017 32583 -26983 32617
rect -26983 32583 -26974 32617
rect -27026 32574 -26974 32583
rect -26866 32617 -26814 32626
rect -26866 32583 -26857 32617
rect -26857 32583 -26823 32617
rect -26823 32583 -26814 32617
rect -26866 32574 -26814 32583
rect -26706 32617 -26654 32626
rect -26706 32583 -26697 32617
rect -26697 32583 -26663 32617
rect -26663 32583 -26654 32617
rect -26706 32574 -26654 32583
rect -26546 32617 -26494 32626
rect -26546 32583 -26537 32617
rect -26537 32583 -26503 32617
rect -26503 32583 -26494 32617
rect -26546 32574 -26494 32583
rect -26386 32617 -26334 32626
rect -26386 32583 -26377 32617
rect -26377 32583 -26343 32617
rect -26343 32583 -26334 32617
rect -26386 32574 -26334 32583
rect -26226 32617 -26174 32626
rect -26226 32583 -26217 32617
rect -26217 32583 -26183 32617
rect -26183 32583 -26174 32617
rect -26226 32574 -26174 32583
rect -26066 32617 -26014 32626
rect -26066 32583 -26057 32617
rect -26057 32583 -26023 32617
rect -26023 32583 -26014 32617
rect -26066 32574 -26014 32583
rect -25906 32617 -25854 32626
rect -25906 32583 -25897 32617
rect -25897 32583 -25863 32617
rect -25863 32583 -25854 32617
rect -25906 32574 -25854 32583
rect -25746 32617 -25694 32626
rect -25746 32583 -25737 32617
rect -25737 32583 -25703 32617
rect -25703 32583 -25694 32617
rect -25746 32574 -25694 32583
rect -25586 32617 -25534 32626
rect -25586 32583 -25577 32617
rect -25577 32583 -25543 32617
rect -25543 32583 -25534 32617
rect -25586 32574 -25534 32583
rect -25426 32617 -25374 32626
rect -25426 32583 -25417 32617
rect -25417 32583 -25383 32617
rect -25383 32583 -25374 32617
rect -25426 32574 -25374 32583
rect -25266 32617 -25214 32626
rect -25266 32583 -25257 32617
rect -25257 32583 -25223 32617
rect -25223 32583 -25214 32617
rect -25266 32574 -25214 32583
rect -25106 32617 -25054 32626
rect -25106 32583 -25097 32617
rect -25097 32583 -25063 32617
rect -25063 32583 -25054 32617
rect -25106 32574 -25054 32583
rect -24946 32617 -24894 32626
rect -24946 32583 -24937 32617
rect -24937 32583 -24903 32617
rect -24903 32583 -24894 32617
rect -24946 32574 -24894 32583
rect -24786 32617 -24734 32626
rect -24786 32583 -24777 32617
rect -24777 32583 -24743 32617
rect -24743 32583 -24734 32617
rect -24786 32574 -24734 32583
rect -24626 32617 -24574 32626
rect -24626 32583 -24617 32617
rect -24617 32583 -24583 32617
rect -24583 32583 -24574 32617
rect -24626 32574 -24574 32583
rect -24466 32617 -24414 32626
rect -24466 32583 -24457 32617
rect -24457 32583 -24423 32617
rect -24423 32583 -24414 32617
rect -24466 32574 -24414 32583
rect -24306 32617 -24254 32626
rect -24306 32583 -24297 32617
rect -24297 32583 -24263 32617
rect -24263 32583 -24254 32617
rect -24306 32574 -24254 32583
rect -24146 32617 -24094 32626
rect -24146 32583 -24137 32617
rect -24137 32583 -24103 32617
rect -24103 32583 -24094 32617
rect -24146 32574 -24094 32583
rect -23986 32617 -23934 32626
rect -23986 32583 -23977 32617
rect -23977 32583 -23943 32617
rect -23943 32583 -23934 32617
rect -23986 32574 -23934 32583
rect -23826 32617 -23774 32626
rect -23826 32583 -23817 32617
rect -23817 32583 -23783 32617
rect -23783 32583 -23774 32617
rect -23826 32574 -23774 32583
rect -23666 32617 -23614 32626
rect -23666 32583 -23657 32617
rect -23657 32583 -23623 32617
rect -23623 32583 -23614 32617
rect -23666 32574 -23614 32583
rect -23506 32617 -23454 32626
rect -23506 32583 -23497 32617
rect -23497 32583 -23463 32617
rect -23463 32583 -23454 32617
rect -23506 32574 -23454 32583
rect -23346 32617 -23294 32626
rect -23346 32583 -23337 32617
rect -23337 32583 -23303 32617
rect -23303 32583 -23294 32617
rect -23346 32574 -23294 32583
rect -23186 32617 -23134 32626
rect -23186 32583 -23177 32617
rect -23177 32583 -23143 32617
rect -23143 32583 -23134 32617
rect -23186 32574 -23134 32583
rect -23026 32617 -22974 32626
rect -23026 32583 -23017 32617
rect -23017 32583 -22983 32617
rect -22983 32583 -22974 32617
rect -23026 32574 -22974 32583
rect -22866 32617 -22814 32626
rect -22866 32583 -22857 32617
rect -22857 32583 -22823 32617
rect -22823 32583 -22814 32617
rect -22866 32574 -22814 32583
rect -22706 32617 -22654 32626
rect -22706 32583 -22697 32617
rect -22697 32583 -22663 32617
rect -22663 32583 -22654 32617
rect -22706 32574 -22654 32583
rect -22546 32617 -22494 32626
rect -22546 32583 -22537 32617
rect -22537 32583 -22503 32617
rect -22503 32583 -22494 32617
rect -22546 32574 -22494 32583
rect -22386 32617 -22334 32626
rect -22386 32583 -22377 32617
rect -22377 32583 -22343 32617
rect -22343 32583 -22334 32617
rect -22386 32574 -22334 32583
rect -22226 32617 -22174 32626
rect -22226 32583 -22217 32617
rect -22217 32583 -22183 32617
rect -22183 32583 -22174 32617
rect -22226 32574 -22174 32583
rect -22066 32617 -22014 32626
rect -22066 32583 -22057 32617
rect -22057 32583 -22023 32617
rect -22023 32583 -22014 32617
rect -22066 32574 -22014 32583
rect -21906 32617 -21854 32626
rect -21906 32583 -21897 32617
rect -21897 32583 -21863 32617
rect -21863 32583 -21854 32617
rect -21906 32574 -21854 32583
rect -21746 32617 -21694 32626
rect -21746 32583 -21737 32617
rect -21737 32583 -21703 32617
rect -21703 32583 -21694 32617
rect -21746 32574 -21694 32583
rect -21586 32617 -21534 32626
rect -21586 32583 -21577 32617
rect -21577 32583 -21543 32617
rect -21543 32583 -21534 32617
rect -21586 32574 -21534 32583
rect -21426 32617 -21374 32626
rect -21426 32583 -21417 32617
rect -21417 32583 -21383 32617
rect -21383 32583 -21374 32617
rect -21426 32574 -21374 32583
rect -21266 32617 -21214 32626
rect -21266 32583 -21257 32617
rect -21257 32583 -21223 32617
rect -21223 32583 -21214 32617
rect -21266 32574 -21214 32583
rect -21106 32617 -21054 32626
rect -21106 32583 -21097 32617
rect -21097 32583 -21063 32617
rect -21063 32583 -21054 32617
rect -21106 32574 -21054 32583
rect -20946 32617 -20894 32626
rect -20946 32583 -20937 32617
rect -20937 32583 -20903 32617
rect -20903 32583 -20894 32617
rect -20946 32574 -20894 32583
rect -20786 32617 -20734 32626
rect -20786 32583 -20777 32617
rect -20777 32583 -20743 32617
rect -20743 32583 -20734 32617
rect -20786 32574 -20734 32583
rect -20626 32617 -20574 32626
rect -20626 32583 -20617 32617
rect -20617 32583 -20583 32617
rect -20583 32583 -20574 32617
rect -20626 32574 -20574 32583
rect -20466 32617 -20414 32626
rect -20466 32583 -20457 32617
rect -20457 32583 -20423 32617
rect -20423 32583 -20414 32617
rect -20466 32574 -20414 32583
rect -20306 32617 -20254 32626
rect -20306 32583 -20297 32617
rect -20297 32583 -20263 32617
rect -20263 32583 -20254 32617
rect -20306 32574 -20254 32583
rect -20146 32617 -20094 32626
rect -20146 32583 -20137 32617
rect -20137 32583 -20103 32617
rect -20103 32583 -20094 32617
rect -20146 32574 -20094 32583
rect -19986 32617 -19934 32626
rect -19986 32583 -19977 32617
rect -19977 32583 -19943 32617
rect -19943 32583 -19934 32617
rect -19986 32574 -19934 32583
rect -19826 32617 -19774 32626
rect -19826 32583 -19817 32617
rect -19817 32583 -19783 32617
rect -19783 32583 -19774 32617
rect -19826 32574 -19774 32583
rect -19666 32617 -19614 32626
rect -19666 32583 -19657 32617
rect -19657 32583 -19623 32617
rect -19623 32583 -19614 32617
rect -19666 32574 -19614 32583
rect -19506 32617 -19454 32626
rect -19506 32583 -19497 32617
rect -19497 32583 -19463 32617
rect -19463 32583 -19454 32617
rect -19506 32574 -19454 32583
rect -19346 32617 -19294 32626
rect -19346 32583 -19337 32617
rect -19337 32583 -19303 32617
rect -19303 32583 -19294 32617
rect -19346 32574 -19294 32583
rect -19186 32617 -19134 32626
rect -19186 32583 -19177 32617
rect -19177 32583 -19143 32617
rect -19143 32583 -19134 32617
rect -19186 32574 -19134 32583
rect -19026 32617 -18974 32626
rect -19026 32583 -19017 32617
rect -19017 32583 -18983 32617
rect -18983 32583 -18974 32617
rect -19026 32574 -18974 32583
rect -18866 32617 -18814 32626
rect -18866 32583 -18857 32617
rect -18857 32583 -18823 32617
rect -18823 32583 -18814 32617
rect -18866 32574 -18814 32583
rect -18706 32617 -18654 32626
rect -18706 32583 -18697 32617
rect -18697 32583 -18663 32617
rect -18663 32583 -18654 32617
rect -18706 32574 -18654 32583
rect -18546 32617 -18494 32626
rect -18546 32583 -18537 32617
rect -18537 32583 -18503 32617
rect -18503 32583 -18494 32617
rect -18546 32574 -18494 32583
rect -18386 32617 -18334 32626
rect -18386 32583 -18377 32617
rect -18377 32583 -18343 32617
rect -18343 32583 -18334 32617
rect -18386 32574 -18334 32583
rect -18226 32617 -18174 32626
rect -18226 32583 -18217 32617
rect -18217 32583 -18183 32617
rect -18183 32583 -18174 32617
rect -18226 32574 -18174 32583
rect -18066 32617 -18014 32626
rect -18066 32583 -18057 32617
rect -18057 32583 -18023 32617
rect -18023 32583 -18014 32617
rect -18066 32574 -18014 32583
rect -17906 32617 -17854 32626
rect -17906 32583 -17897 32617
rect -17897 32583 -17863 32617
rect -17863 32583 -17854 32617
rect -17906 32574 -17854 32583
rect -17746 32617 -17694 32626
rect -17746 32583 -17737 32617
rect -17737 32583 -17703 32617
rect -17703 32583 -17694 32617
rect -17746 32574 -17694 32583
rect -17586 32617 -17534 32626
rect -17586 32583 -17577 32617
rect -17577 32583 -17543 32617
rect -17543 32583 -17534 32617
rect -17586 32574 -17534 32583
rect -17426 32617 -17374 32626
rect -17426 32583 -17417 32617
rect -17417 32583 -17383 32617
rect -17383 32583 -17374 32617
rect -17426 32574 -17374 32583
rect -17266 32617 -17214 32626
rect -17266 32583 -17257 32617
rect -17257 32583 -17223 32617
rect -17223 32583 -17214 32617
rect -17266 32574 -17214 32583
rect -17106 32617 -17054 32626
rect -17106 32583 -17097 32617
rect -17097 32583 -17063 32617
rect -17063 32583 -17054 32617
rect -17106 32574 -17054 32583
rect -16946 32617 -16894 32626
rect -16946 32583 -16937 32617
rect -16937 32583 -16903 32617
rect -16903 32583 -16894 32617
rect -16946 32574 -16894 32583
rect -16786 32617 -16734 32626
rect -16786 32583 -16777 32617
rect -16777 32583 -16743 32617
rect -16743 32583 -16734 32617
rect -16786 32574 -16734 32583
rect -16626 32617 -16574 32626
rect -16626 32583 -16617 32617
rect -16617 32583 -16583 32617
rect -16583 32583 -16574 32617
rect -16626 32574 -16574 32583
rect -16466 32617 -16414 32626
rect -16466 32583 -16457 32617
rect -16457 32583 -16423 32617
rect -16423 32583 -16414 32617
rect -16466 32574 -16414 32583
rect -16306 32617 -16254 32626
rect -16306 32583 -16297 32617
rect -16297 32583 -16263 32617
rect -16263 32583 -16254 32617
rect -16306 32574 -16254 32583
rect -16146 32617 -16094 32626
rect -16146 32583 -16137 32617
rect -16137 32583 -16103 32617
rect -16103 32583 -16094 32617
rect -16146 32574 -16094 32583
rect -15986 32617 -15934 32626
rect -15986 32583 -15977 32617
rect -15977 32583 -15943 32617
rect -15943 32583 -15934 32617
rect -15986 32574 -15934 32583
rect -15826 32617 -15774 32626
rect -15826 32583 -15817 32617
rect -15817 32583 -15783 32617
rect -15783 32583 -15774 32617
rect -15826 32574 -15774 32583
rect -15666 32617 -15614 32626
rect -15666 32583 -15657 32617
rect -15657 32583 -15623 32617
rect -15623 32583 -15614 32617
rect -15666 32574 -15614 32583
rect -15506 32617 -15454 32626
rect -15506 32583 -15497 32617
rect -15497 32583 -15463 32617
rect -15463 32583 -15454 32617
rect -15506 32574 -15454 32583
rect -15346 32617 -15294 32626
rect -15346 32583 -15337 32617
rect -15337 32583 -15303 32617
rect -15303 32583 -15294 32617
rect -15346 32574 -15294 32583
rect -15186 32617 -15134 32626
rect -15186 32583 -15177 32617
rect -15177 32583 -15143 32617
rect -15143 32583 -15134 32617
rect -15186 32574 -15134 32583
rect -15026 32617 -14974 32626
rect -15026 32583 -15017 32617
rect -15017 32583 -14983 32617
rect -14983 32583 -14974 32617
rect -15026 32574 -14974 32583
rect -14866 32617 -14814 32626
rect -14866 32583 -14857 32617
rect -14857 32583 -14823 32617
rect -14823 32583 -14814 32617
rect -14866 32574 -14814 32583
rect -14706 32617 -14654 32626
rect -14706 32583 -14697 32617
rect -14697 32583 -14663 32617
rect -14663 32583 -14654 32617
rect -14706 32574 -14654 32583
rect -14546 32617 -14494 32626
rect -14546 32583 -14537 32617
rect -14537 32583 -14503 32617
rect -14503 32583 -14494 32617
rect -14546 32574 -14494 32583
rect -14386 32617 -14334 32626
rect -14386 32583 -14377 32617
rect -14377 32583 -14343 32617
rect -14343 32583 -14334 32617
rect -14386 32574 -14334 32583
rect -14226 32617 -14174 32626
rect -14226 32583 -14217 32617
rect -14217 32583 -14183 32617
rect -14183 32583 -14174 32617
rect -14226 32574 -14174 32583
rect -14066 32617 -14014 32626
rect -14066 32583 -14057 32617
rect -14057 32583 -14023 32617
rect -14023 32583 -14014 32617
rect -14066 32574 -14014 32583
rect -13906 32617 -13854 32626
rect -13906 32583 -13897 32617
rect -13897 32583 -13863 32617
rect -13863 32583 -13854 32617
rect -13906 32574 -13854 32583
rect -13746 32617 -13694 32626
rect -13746 32583 -13737 32617
rect -13737 32583 -13703 32617
rect -13703 32583 -13694 32617
rect -13746 32574 -13694 32583
rect -13586 32617 -13534 32626
rect -13586 32583 -13577 32617
rect -13577 32583 -13543 32617
rect -13543 32583 -13534 32617
rect -13586 32574 -13534 32583
rect -13426 32617 -13374 32626
rect -13426 32583 -13417 32617
rect -13417 32583 -13383 32617
rect -13383 32583 -13374 32617
rect -13426 32574 -13374 32583
rect -13266 32617 -13214 32626
rect -13266 32583 -13257 32617
rect -13257 32583 -13223 32617
rect -13223 32583 -13214 32617
rect -13266 32574 -13214 32583
rect -13106 32617 -13054 32626
rect -13106 32583 -13097 32617
rect -13097 32583 -13063 32617
rect -13063 32583 -13054 32617
rect -13106 32574 -13054 32583
rect -12946 32617 -12894 32626
rect -12946 32583 -12937 32617
rect -12937 32583 -12903 32617
rect -12903 32583 -12894 32617
rect -12946 32574 -12894 32583
rect -12786 32617 -12734 32626
rect -12786 32583 -12777 32617
rect -12777 32583 -12743 32617
rect -12743 32583 -12734 32617
rect -12786 32574 -12734 32583
rect -12626 32617 -12574 32626
rect -12626 32583 -12617 32617
rect -12617 32583 -12583 32617
rect -12583 32583 -12574 32617
rect -12626 32574 -12574 32583
rect -12466 32617 -12414 32626
rect -12466 32583 -12457 32617
rect -12457 32583 -12423 32617
rect -12423 32583 -12414 32617
rect -12466 32574 -12414 32583
rect -12306 32617 -12254 32626
rect -12306 32583 -12297 32617
rect -12297 32583 -12263 32617
rect -12263 32583 -12254 32617
rect -12306 32574 -12254 32583
rect -12146 32617 -12094 32626
rect -12146 32583 -12137 32617
rect -12137 32583 -12103 32617
rect -12103 32583 -12094 32617
rect -12146 32574 -12094 32583
rect -11986 32617 -11934 32626
rect -11986 32583 -11977 32617
rect -11977 32583 -11943 32617
rect -11943 32583 -11934 32617
rect -11986 32574 -11934 32583
rect -11826 32617 -11774 32626
rect -11826 32583 -11817 32617
rect -11817 32583 -11783 32617
rect -11783 32583 -11774 32617
rect -11826 32574 -11774 32583
rect -11666 32617 -11614 32626
rect -11666 32583 -11657 32617
rect -11657 32583 -11623 32617
rect -11623 32583 -11614 32617
rect -11666 32574 -11614 32583
rect -11506 32617 -11454 32626
rect -11506 32583 -11497 32617
rect -11497 32583 -11463 32617
rect -11463 32583 -11454 32617
rect -11506 32574 -11454 32583
rect -11186 32617 -11134 32626
rect -11186 32583 -11177 32617
rect -11177 32583 -11143 32617
rect -11143 32583 -11134 32617
rect -11186 32574 -11134 32583
rect -10866 32617 -10814 32626
rect -10866 32583 -10857 32617
rect -10857 32583 -10823 32617
rect -10823 32583 -10814 32617
rect -10866 32574 -10814 32583
rect -10706 32617 -10654 32626
rect -10706 32583 -10697 32617
rect -10697 32583 -10663 32617
rect -10663 32583 -10654 32617
rect -10706 32574 -10654 32583
rect -10546 32617 -10494 32626
rect -10546 32583 -10537 32617
rect -10537 32583 -10503 32617
rect -10503 32583 -10494 32617
rect -10546 32574 -10494 32583
rect -10386 32617 -10334 32626
rect -10386 32583 -10377 32617
rect -10377 32583 -10343 32617
rect -10343 32583 -10334 32617
rect -10386 32574 -10334 32583
rect -10226 32617 -10174 32626
rect -10226 32583 -10217 32617
rect -10217 32583 -10183 32617
rect -10183 32583 -10174 32617
rect -10226 32574 -10174 32583
rect -10066 32617 -10014 32626
rect -10066 32583 -10057 32617
rect -10057 32583 -10023 32617
rect -10023 32583 -10014 32617
rect -10066 32574 -10014 32583
rect -9906 32617 -9854 32626
rect -9906 32583 -9897 32617
rect -9897 32583 -9863 32617
rect -9863 32583 -9854 32617
rect -9906 32574 -9854 32583
rect -9746 32617 -9694 32626
rect -9746 32583 -9737 32617
rect -9737 32583 -9703 32617
rect -9703 32583 -9694 32617
rect -9746 32574 -9694 32583
rect -9586 32617 -9534 32626
rect -9586 32583 -9577 32617
rect -9577 32583 -9543 32617
rect -9543 32583 -9534 32617
rect -9586 32574 -9534 32583
rect -9426 32617 -9374 32626
rect -9426 32583 -9417 32617
rect -9417 32583 -9383 32617
rect -9383 32583 -9374 32617
rect -9426 32574 -9374 32583
rect -9266 32617 -9214 32626
rect -9266 32583 -9257 32617
rect -9257 32583 -9223 32617
rect -9223 32583 -9214 32617
rect -9266 32574 -9214 32583
rect -9106 32617 -9054 32626
rect -9106 32583 -9097 32617
rect -9097 32583 -9063 32617
rect -9063 32583 -9054 32617
rect -9106 32574 -9054 32583
rect -8946 32617 -8894 32626
rect -8946 32583 -8937 32617
rect -8937 32583 -8903 32617
rect -8903 32583 -8894 32617
rect -8946 32574 -8894 32583
rect -8786 32617 -8734 32626
rect -8786 32583 -8777 32617
rect -8777 32583 -8743 32617
rect -8743 32583 -8734 32617
rect -8786 32574 -8734 32583
rect -8626 32617 -8574 32626
rect -8626 32583 -8617 32617
rect -8617 32583 -8583 32617
rect -8583 32583 -8574 32617
rect -8626 32574 -8574 32583
rect -8466 32617 -8414 32626
rect -8466 32583 -8457 32617
rect -8457 32583 -8423 32617
rect -8423 32583 -8414 32617
rect -8466 32574 -8414 32583
rect -8306 32617 -8254 32626
rect -8306 32583 -8297 32617
rect -8297 32583 -8263 32617
rect -8263 32583 -8254 32617
rect -8306 32574 -8254 32583
rect -8146 32617 -8094 32626
rect -8146 32583 -8137 32617
rect -8137 32583 -8103 32617
rect -8103 32583 -8094 32617
rect -8146 32574 -8094 32583
rect -7986 32617 -7934 32626
rect -7986 32583 -7977 32617
rect -7977 32583 -7943 32617
rect -7943 32583 -7934 32617
rect -7986 32574 -7934 32583
rect -7826 32617 -7774 32626
rect -7826 32583 -7817 32617
rect -7817 32583 -7783 32617
rect -7783 32583 -7774 32617
rect -7826 32574 -7774 32583
rect -7666 32617 -7614 32626
rect -7666 32583 -7657 32617
rect -7657 32583 -7623 32617
rect -7623 32583 -7614 32617
rect -7666 32574 -7614 32583
rect -7506 32617 -7454 32626
rect -7506 32583 -7497 32617
rect -7497 32583 -7463 32617
rect -7463 32583 -7454 32617
rect -7506 32574 -7454 32583
rect -7346 32617 -7294 32626
rect -7346 32583 -7337 32617
rect -7337 32583 -7303 32617
rect -7303 32583 -7294 32617
rect -7346 32574 -7294 32583
rect -7186 32617 -7134 32626
rect -7186 32583 -7177 32617
rect -7177 32583 -7143 32617
rect -7143 32583 -7134 32617
rect -7186 32574 -7134 32583
rect -7026 32617 -6974 32626
rect -7026 32583 -7017 32617
rect -7017 32583 -6983 32617
rect -6983 32583 -6974 32617
rect -7026 32574 -6974 32583
rect -6866 32617 -6814 32626
rect -6866 32583 -6857 32617
rect -6857 32583 -6823 32617
rect -6823 32583 -6814 32617
rect -6866 32574 -6814 32583
rect -6706 32617 -6654 32626
rect -6706 32583 -6697 32617
rect -6697 32583 -6663 32617
rect -6663 32583 -6654 32617
rect -6706 32574 -6654 32583
rect -6546 32617 -6494 32626
rect -6546 32583 -6537 32617
rect -6537 32583 -6503 32617
rect -6503 32583 -6494 32617
rect -6546 32574 -6494 32583
rect -6386 32617 -6334 32626
rect -6386 32583 -6377 32617
rect -6377 32583 -6343 32617
rect -6343 32583 -6334 32617
rect -6386 32574 -6334 32583
rect -6226 32617 -6174 32626
rect -6226 32583 -6217 32617
rect -6217 32583 -6183 32617
rect -6183 32583 -6174 32617
rect -6226 32574 -6174 32583
rect -6066 32617 -6014 32626
rect -6066 32583 -6057 32617
rect -6057 32583 -6023 32617
rect -6023 32583 -6014 32617
rect -6066 32574 -6014 32583
rect -5906 32617 -5854 32626
rect -5906 32583 -5897 32617
rect -5897 32583 -5863 32617
rect -5863 32583 -5854 32617
rect -5906 32574 -5854 32583
rect -5746 32617 -5694 32626
rect -5746 32583 -5737 32617
rect -5737 32583 -5703 32617
rect -5703 32583 -5694 32617
rect -5746 32574 -5694 32583
rect -5586 32617 -5534 32626
rect -5586 32583 -5577 32617
rect -5577 32583 -5543 32617
rect -5543 32583 -5534 32617
rect -5586 32574 -5534 32583
rect -5426 32617 -5374 32626
rect -5426 32583 -5417 32617
rect -5417 32583 -5383 32617
rect -5383 32583 -5374 32617
rect -5426 32574 -5374 32583
rect -5266 32617 -5214 32626
rect -5266 32583 -5257 32617
rect -5257 32583 -5223 32617
rect -5223 32583 -5214 32617
rect -5266 32574 -5214 32583
rect -5106 32617 -5054 32626
rect -5106 32583 -5097 32617
rect -5097 32583 -5063 32617
rect -5063 32583 -5054 32617
rect -5106 32574 -5054 32583
rect -4946 32617 -4894 32626
rect -4946 32583 -4937 32617
rect -4937 32583 -4903 32617
rect -4903 32583 -4894 32617
rect -4946 32574 -4894 32583
rect -4786 32617 -4734 32626
rect -4786 32583 -4777 32617
rect -4777 32583 -4743 32617
rect -4743 32583 -4734 32617
rect -4786 32574 -4734 32583
rect -4626 32617 -4574 32626
rect -4626 32583 -4617 32617
rect -4617 32583 -4583 32617
rect -4583 32583 -4574 32617
rect -4626 32574 -4574 32583
rect -4466 32617 -4414 32626
rect -4466 32583 -4457 32617
rect -4457 32583 -4423 32617
rect -4423 32583 -4414 32617
rect -4466 32574 -4414 32583
rect -4306 32617 -4254 32626
rect -4306 32583 -4297 32617
rect -4297 32583 -4263 32617
rect -4263 32583 -4254 32617
rect -4306 32574 -4254 32583
rect -4146 32617 -4094 32626
rect -4146 32583 -4137 32617
rect -4137 32583 -4103 32617
rect -4103 32583 -4094 32617
rect -4146 32574 -4094 32583
rect -3986 32617 -3934 32626
rect -3986 32583 -3977 32617
rect -3977 32583 -3943 32617
rect -3943 32583 -3934 32617
rect -3986 32574 -3934 32583
rect -3666 32617 -3614 32626
rect -3666 32583 -3657 32617
rect -3657 32583 -3623 32617
rect -3623 32583 -3614 32617
rect -3666 32574 -3614 32583
rect -3506 32617 -3454 32626
rect -3506 32583 -3497 32617
rect -3497 32583 -3463 32617
rect -3463 32583 -3454 32617
rect -3506 32574 -3454 32583
rect -3346 32617 -3294 32626
rect -3346 32583 -3337 32617
rect -3337 32583 -3303 32617
rect -3303 32583 -3294 32617
rect -3346 32574 -3294 32583
rect -3186 32617 -3134 32626
rect -3186 32583 -3177 32617
rect -3177 32583 -3143 32617
rect -3143 32583 -3134 32617
rect -3186 32574 -3134 32583
rect -3026 32617 -2974 32626
rect -3026 32583 -3017 32617
rect -3017 32583 -2983 32617
rect -2983 32583 -2974 32617
rect -3026 32574 -2974 32583
rect -2866 32617 -2814 32626
rect -2866 32583 -2857 32617
rect -2857 32583 -2823 32617
rect -2823 32583 -2814 32617
rect -2866 32574 -2814 32583
rect -2706 32617 -2654 32626
rect -2706 32583 -2697 32617
rect -2697 32583 -2663 32617
rect -2663 32583 -2654 32617
rect -2706 32574 -2654 32583
rect -2386 32617 -2334 32626
rect -2386 32583 -2377 32617
rect -2377 32583 -2343 32617
rect -2343 32583 -2334 32617
rect -2386 32574 -2334 32583
rect -2066 32617 -2014 32626
rect -2066 32583 -2057 32617
rect -2057 32583 -2023 32617
rect -2023 32583 -2014 32617
rect -2066 32574 -2014 32583
rect -1746 32617 -1694 32626
rect -1746 32583 -1737 32617
rect -1737 32583 -1703 32617
rect -1703 32583 -1694 32617
rect -1746 32574 -1694 32583
rect -1426 32617 -1374 32626
rect -1426 32583 -1417 32617
rect -1417 32583 -1383 32617
rect -1383 32583 -1374 32617
rect -1426 32574 -1374 32583
rect -1106 32617 -1054 32626
rect -1106 32583 -1097 32617
rect -1097 32583 -1063 32617
rect -1063 32583 -1054 32617
rect -1106 32574 -1054 32583
rect -29906 32297 -29854 32306
rect -29906 32263 -29897 32297
rect -29897 32263 -29863 32297
rect -29863 32263 -29854 32297
rect -29906 32254 -29854 32263
rect -29746 32297 -29694 32306
rect -29746 32263 -29737 32297
rect -29737 32263 -29703 32297
rect -29703 32263 -29694 32297
rect -29746 32254 -29694 32263
rect -29586 32297 -29534 32306
rect -29586 32263 -29577 32297
rect -29577 32263 -29543 32297
rect -29543 32263 -29534 32297
rect -29586 32254 -29534 32263
rect -29426 32297 -29374 32306
rect -29426 32263 -29417 32297
rect -29417 32263 -29383 32297
rect -29383 32263 -29374 32297
rect -29426 32254 -29374 32263
rect -29266 32297 -29214 32306
rect -29266 32263 -29257 32297
rect -29257 32263 -29223 32297
rect -29223 32263 -29214 32297
rect -29266 32254 -29214 32263
rect -29106 32297 -29054 32306
rect -29106 32263 -29097 32297
rect -29097 32263 -29063 32297
rect -29063 32263 -29054 32297
rect -29106 32254 -29054 32263
rect -28946 32297 -28894 32306
rect -28946 32263 -28937 32297
rect -28937 32263 -28903 32297
rect -28903 32263 -28894 32297
rect -28946 32254 -28894 32263
rect -28786 32297 -28734 32306
rect -28786 32263 -28777 32297
rect -28777 32263 -28743 32297
rect -28743 32263 -28734 32297
rect -28786 32254 -28734 32263
rect -28626 32297 -28574 32306
rect -28626 32263 -28617 32297
rect -28617 32263 -28583 32297
rect -28583 32263 -28574 32297
rect -28626 32254 -28574 32263
rect -28466 32297 -28414 32306
rect -28466 32263 -28457 32297
rect -28457 32263 -28423 32297
rect -28423 32263 -28414 32297
rect -28466 32254 -28414 32263
rect -28306 32297 -28254 32306
rect -28306 32263 -28297 32297
rect -28297 32263 -28263 32297
rect -28263 32263 -28254 32297
rect -28306 32254 -28254 32263
rect -28146 32297 -28094 32306
rect -28146 32263 -28137 32297
rect -28137 32263 -28103 32297
rect -28103 32263 -28094 32297
rect -28146 32254 -28094 32263
rect -27986 32297 -27934 32306
rect -27986 32263 -27977 32297
rect -27977 32263 -27943 32297
rect -27943 32263 -27934 32297
rect -27986 32254 -27934 32263
rect -27826 32297 -27774 32306
rect -27826 32263 -27817 32297
rect -27817 32263 -27783 32297
rect -27783 32263 -27774 32297
rect -27826 32254 -27774 32263
rect -27666 32297 -27614 32306
rect -27666 32263 -27657 32297
rect -27657 32263 -27623 32297
rect -27623 32263 -27614 32297
rect -27666 32254 -27614 32263
rect -27506 32297 -27454 32306
rect -27506 32263 -27497 32297
rect -27497 32263 -27463 32297
rect -27463 32263 -27454 32297
rect -27506 32254 -27454 32263
rect -27346 32297 -27294 32306
rect -27346 32263 -27337 32297
rect -27337 32263 -27303 32297
rect -27303 32263 -27294 32297
rect -27346 32254 -27294 32263
rect -27186 32297 -27134 32306
rect -27186 32263 -27177 32297
rect -27177 32263 -27143 32297
rect -27143 32263 -27134 32297
rect -27186 32254 -27134 32263
rect -27026 32297 -26974 32306
rect -27026 32263 -27017 32297
rect -27017 32263 -26983 32297
rect -26983 32263 -26974 32297
rect -27026 32254 -26974 32263
rect -26866 32297 -26814 32306
rect -26866 32263 -26857 32297
rect -26857 32263 -26823 32297
rect -26823 32263 -26814 32297
rect -26866 32254 -26814 32263
rect -26706 32297 -26654 32306
rect -26706 32263 -26697 32297
rect -26697 32263 -26663 32297
rect -26663 32263 -26654 32297
rect -26706 32254 -26654 32263
rect -26546 32297 -26494 32306
rect -26546 32263 -26537 32297
rect -26537 32263 -26503 32297
rect -26503 32263 -26494 32297
rect -26546 32254 -26494 32263
rect -26386 32297 -26334 32306
rect -26386 32263 -26377 32297
rect -26377 32263 -26343 32297
rect -26343 32263 -26334 32297
rect -26386 32254 -26334 32263
rect -26226 32297 -26174 32306
rect -26226 32263 -26217 32297
rect -26217 32263 -26183 32297
rect -26183 32263 -26174 32297
rect -26226 32254 -26174 32263
rect -26066 32297 -26014 32306
rect -26066 32263 -26057 32297
rect -26057 32263 -26023 32297
rect -26023 32263 -26014 32297
rect -26066 32254 -26014 32263
rect -25906 32297 -25854 32306
rect -25906 32263 -25897 32297
rect -25897 32263 -25863 32297
rect -25863 32263 -25854 32297
rect -25906 32254 -25854 32263
rect -25746 32297 -25694 32306
rect -25746 32263 -25737 32297
rect -25737 32263 -25703 32297
rect -25703 32263 -25694 32297
rect -25746 32254 -25694 32263
rect -25586 32297 -25534 32306
rect -25586 32263 -25577 32297
rect -25577 32263 -25543 32297
rect -25543 32263 -25534 32297
rect -25586 32254 -25534 32263
rect -25426 32297 -25374 32306
rect -25426 32263 -25417 32297
rect -25417 32263 -25383 32297
rect -25383 32263 -25374 32297
rect -25426 32254 -25374 32263
rect -25266 32297 -25214 32306
rect -25266 32263 -25257 32297
rect -25257 32263 -25223 32297
rect -25223 32263 -25214 32297
rect -25266 32254 -25214 32263
rect -25106 32297 -25054 32306
rect -25106 32263 -25097 32297
rect -25097 32263 -25063 32297
rect -25063 32263 -25054 32297
rect -25106 32254 -25054 32263
rect -24946 32297 -24894 32306
rect -24946 32263 -24937 32297
rect -24937 32263 -24903 32297
rect -24903 32263 -24894 32297
rect -24946 32254 -24894 32263
rect -24786 32297 -24734 32306
rect -24786 32263 -24777 32297
rect -24777 32263 -24743 32297
rect -24743 32263 -24734 32297
rect -24786 32254 -24734 32263
rect -24626 32297 -24574 32306
rect -24626 32263 -24617 32297
rect -24617 32263 -24583 32297
rect -24583 32263 -24574 32297
rect -24626 32254 -24574 32263
rect -24466 32297 -24414 32306
rect -24466 32263 -24457 32297
rect -24457 32263 -24423 32297
rect -24423 32263 -24414 32297
rect -24466 32254 -24414 32263
rect -24306 32297 -24254 32306
rect -24306 32263 -24297 32297
rect -24297 32263 -24263 32297
rect -24263 32263 -24254 32297
rect -24306 32254 -24254 32263
rect -24146 32297 -24094 32306
rect -24146 32263 -24137 32297
rect -24137 32263 -24103 32297
rect -24103 32263 -24094 32297
rect -24146 32254 -24094 32263
rect -23986 32297 -23934 32306
rect -23986 32263 -23977 32297
rect -23977 32263 -23943 32297
rect -23943 32263 -23934 32297
rect -23986 32254 -23934 32263
rect -23826 32297 -23774 32306
rect -23826 32263 -23817 32297
rect -23817 32263 -23783 32297
rect -23783 32263 -23774 32297
rect -23826 32254 -23774 32263
rect -23666 32297 -23614 32306
rect -23666 32263 -23657 32297
rect -23657 32263 -23623 32297
rect -23623 32263 -23614 32297
rect -23666 32254 -23614 32263
rect -23506 32297 -23454 32306
rect -23506 32263 -23497 32297
rect -23497 32263 -23463 32297
rect -23463 32263 -23454 32297
rect -23506 32254 -23454 32263
rect -23346 32297 -23294 32306
rect -23346 32263 -23337 32297
rect -23337 32263 -23303 32297
rect -23303 32263 -23294 32297
rect -23346 32254 -23294 32263
rect -23186 32297 -23134 32306
rect -23186 32263 -23177 32297
rect -23177 32263 -23143 32297
rect -23143 32263 -23134 32297
rect -23186 32254 -23134 32263
rect -23026 32297 -22974 32306
rect -23026 32263 -23017 32297
rect -23017 32263 -22983 32297
rect -22983 32263 -22974 32297
rect -23026 32254 -22974 32263
rect -22866 32297 -22814 32306
rect -22866 32263 -22857 32297
rect -22857 32263 -22823 32297
rect -22823 32263 -22814 32297
rect -22866 32254 -22814 32263
rect -22706 32297 -22654 32306
rect -22706 32263 -22697 32297
rect -22697 32263 -22663 32297
rect -22663 32263 -22654 32297
rect -22706 32254 -22654 32263
rect -22546 32297 -22494 32306
rect -22546 32263 -22537 32297
rect -22537 32263 -22503 32297
rect -22503 32263 -22494 32297
rect -22546 32254 -22494 32263
rect -22386 32297 -22334 32306
rect -22386 32263 -22377 32297
rect -22377 32263 -22343 32297
rect -22343 32263 -22334 32297
rect -22386 32254 -22334 32263
rect -22226 32297 -22174 32306
rect -22226 32263 -22217 32297
rect -22217 32263 -22183 32297
rect -22183 32263 -22174 32297
rect -22226 32254 -22174 32263
rect -22066 32297 -22014 32306
rect -22066 32263 -22057 32297
rect -22057 32263 -22023 32297
rect -22023 32263 -22014 32297
rect -22066 32254 -22014 32263
rect -21906 32297 -21854 32306
rect -21906 32263 -21897 32297
rect -21897 32263 -21863 32297
rect -21863 32263 -21854 32297
rect -21906 32254 -21854 32263
rect -21746 32297 -21694 32306
rect -21746 32263 -21737 32297
rect -21737 32263 -21703 32297
rect -21703 32263 -21694 32297
rect -21746 32254 -21694 32263
rect -21586 32297 -21534 32306
rect -21586 32263 -21577 32297
rect -21577 32263 -21543 32297
rect -21543 32263 -21534 32297
rect -21586 32254 -21534 32263
rect -21426 32297 -21374 32306
rect -21426 32263 -21417 32297
rect -21417 32263 -21383 32297
rect -21383 32263 -21374 32297
rect -21426 32254 -21374 32263
rect -21266 32297 -21214 32306
rect -21266 32263 -21257 32297
rect -21257 32263 -21223 32297
rect -21223 32263 -21214 32297
rect -21266 32254 -21214 32263
rect -21106 32297 -21054 32306
rect -21106 32263 -21097 32297
rect -21097 32263 -21063 32297
rect -21063 32263 -21054 32297
rect -21106 32254 -21054 32263
rect -20946 32297 -20894 32306
rect -20946 32263 -20937 32297
rect -20937 32263 -20903 32297
rect -20903 32263 -20894 32297
rect -20946 32254 -20894 32263
rect -20786 32297 -20734 32306
rect -20786 32263 -20777 32297
rect -20777 32263 -20743 32297
rect -20743 32263 -20734 32297
rect -20786 32254 -20734 32263
rect -20626 32297 -20574 32306
rect -20626 32263 -20617 32297
rect -20617 32263 -20583 32297
rect -20583 32263 -20574 32297
rect -20626 32254 -20574 32263
rect -20466 32297 -20414 32306
rect -20466 32263 -20457 32297
rect -20457 32263 -20423 32297
rect -20423 32263 -20414 32297
rect -20466 32254 -20414 32263
rect -20306 32297 -20254 32306
rect -20306 32263 -20297 32297
rect -20297 32263 -20263 32297
rect -20263 32263 -20254 32297
rect -20306 32254 -20254 32263
rect -20146 32297 -20094 32306
rect -20146 32263 -20137 32297
rect -20137 32263 -20103 32297
rect -20103 32263 -20094 32297
rect -20146 32254 -20094 32263
rect -19986 32297 -19934 32306
rect -19986 32263 -19977 32297
rect -19977 32263 -19943 32297
rect -19943 32263 -19934 32297
rect -19986 32254 -19934 32263
rect -19826 32297 -19774 32306
rect -19826 32263 -19817 32297
rect -19817 32263 -19783 32297
rect -19783 32263 -19774 32297
rect -19826 32254 -19774 32263
rect -19666 32297 -19614 32306
rect -19666 32263 -19657 32297
rect -19657 32263 -19623 32297
rect -19623 32263 -19614 32297
rect -19666 32254 -19614 32263
rect -19506 32297 -19454 32306
rect -19506 32263 -19497 32297
rect -19497 32263 -19463 32297
rect -19463 32263 -19454 32297
rect -19506 32254 -19454 32263
rect -19346 32297 -19294 32306
rect -19346 32263 -19337 32297
rect -19337 32263 -19303 32297
rect -19303 32263 -19294 32297
rect -19346 32254 -19294 32263
rect -19186 32297 -19134 32306
rect -19186 32263 -19177 32297
rect -19177 32263 -19143 32297
rect -19143 32263 -19134 32297
rect -19186 32254 -19134 32263
rect -19026 32297 -18974 32306
rect -19026 32263 -19017 32297
rect -19017 32263 -18983 32297
rect -18983 32263 -18974 32297
rect -19026 32254 -18974 32263
rect -18866 32297 -18814 32306
rect -18866 32263 -18857 32297
rect -18857 32263 -18823 32297
rect -18823 32263 -18814 32297
rect -18866 32254 -18814 32263
rect -18706 32297 -18654 32306
rect -18706 32263 -18697 32297
rect -18697 32263 -18663 32297
rect -18663 32263 -18654 32297
rect -18706 32254 -18654 32263
rect -18546 32297 -18494 32306
rect -18546 32263 -18537 32297
rect -18537 32263 -18503 32297
rect -18503 32263 -18494 32297
rect -18546 32254 -18494 32263
rect -18386 32297 -18334 32306
rect -18386 32263 -18377 32297
rect -18377 32263 -18343 32297
rect -18343 32263 -18334 32297
rect -18386 32254 -18334 32263
rect -18226 32297 -18174 32306
rect -18226 32263 -18217 32297
rect -18217 32263 -18183 32297
rect -18183 32263 -18174 32297
rect -18226 32254 -18174 32263
rect -18066 32297 -18014 32306
rect -18066 32263 -18057 32297
rect -18057 32263 -18023 32297
rect -18023 32263 -18014 32297
rect -18066 32254 -18014 32263
rect -17906 32297 -17854 32306
rect -17906 32263 -17897 32297
rect -17897 32263 -17863 32297
rect -17863 32263 -17854 32297
rect -17906 32254 -17854 32263
rect -17746 32297 -17694 32306
rect -17746 32263 -17737 32297
rect -17737 32263 -17703 32297
rect -17703 32263 -17694 32297
rect -17746 32254 -17694 32263
rect -17586 32297 -17534 32306
rect -17586 32263 -17577 32297
rect -17577 32263 -17543 32297
rect -17543 32263 -17534 32297
rect -17586 32254 -17534 32263
rect -17426 32297 -17374 32306
rect -17426 32263 -17417 32297
rect -17417 32263 -17383 32297
rect -17383 32263 -17374 32297
rect -17426 32254 -17374 32263
rect -17266 32297 -17214 32306
rect -17266 32263 -17257 32297
rect -17257 32263 -17223 32297
rect -17223 32263 -17214 32297
rect -17266 32254 -17214 32263
rect -17106 32297 -17054 32306
rect -17106 32263 -17097 32297
rect -17097 32263 -17063 32297
rect -17063 32263 -17054 32297
rect -17106 32254 -17054 32263
rect -16946 32297 -16894 32306
rect -16946 32263 -16937 32297
rect -16937 32263 -16903 32297
rect -16903 32263 -16894 32297
rect -16946 32254 -16894 32263
rect -16786 32297 -16734 32306
rect -16786 32263 -16777 32297
rect -16777 32263 -16743 32297
rect -16743 32263 -16734 32297
rect -16786 32254 -16734 32263
rect -16626 32297 -16574 32306
rect -16626 32263 -16617 32297
rect -16617 32263 -16583 32297
rect -16583 32263 -16574 32297
rect -16626 32254 -16574 32263
rect -16466 32297 -16414 32306
rect -16466 32263 -16457 32297
rect -16457 32263 -16423 32297
rect -16423 32263 -16414 32297
rect -16466 32254 -16414 32263
rect -16306 32297 -16254 32306
rect -16306 32263 -16297 32297
rect -16297 32263 -16263 32297
rect -16263 32263 -16254 32297
rect -16306 32254 -16254 32263
rect -16146 32297 -16094 32306
rect -16146 32263 -16137 32297
rect -16137 32263 -16103 32297
rect -16103 32263 -16094 32297
rect -16146 32254 -16094 32263
rect -15986 32297 -15934 32306
rect -15986 32263 -15977 32297
rect -15977 32263 -15943 32297
rect -15943 32263 -15934 32297
rect -15986 32254 -15934 32263
rect -15826 32297 -15774 32306
rect -15826 32263 -15817 32297
rect -15817 32263 -15783 32297
rect -15783 32263 -15774 32297
rect -15826 32254 -15774 32263
rect -15666 32297 -15614 32306
rect -15666 32263 -15657 32297
rect -15657 32263 -15623 32297
rect -15623 32263 -15614 32297
rect -15666 32254 -15614 32263
rect -15506 32297 -15454 32306
rect -15506 32263 -15497 32297
rect -15497 32263 -15463 32297
rect -15463 32263 -15454 32297
rect -15506 32254 -15454 32263
rect -15346 32297 -15294 32306
rect -15346 32263 -15337 32297
rect -15337 32263 -15303 32297
rect -15303 32263 -15294 32297
rect -15346 32254 -15294 32263
rect -15186 32297 -15134 32306
rect -15186 32263 -15177 32297
rect -15177 32263 -15143 32297
rect -15143 32263 -15134 32297
rect -15186 32254 -15134 32263
rect -15026 32297 -14974 32306
rect -15026 32263 -15017 32297
rect -15017 32263 -14983 32297
rect -14983 32263 -14974 32297
rect -15026 32254 -14974 32263
rect -14866 32297 -14814 32306
rect -14866 32263 -14857 32297
rect -14857 32263 -14823 32297
rect -14823 32263 -14814 32297
rect -14866 32254 -14814 32263
rect -14706 32297 -14654 32306
rect -14706 32263 -14697 32297
rect -14697 32263 -14663 32297
rect -14663 32263 -14654 32297
rect -14706 32254 -14654 32263
rect -14546 32297 -14494 32306
rect -14546 32263 -14537 32297
rect -14537 32263 -14503 32297
rect -14503 32263 -14494 32297
rect -14546 32254 -14494 32263
rect -14386 32297 -14334 32306
rect -14386 32263 -14377 32297
rect -14377 32263 -14343 32297
rect -14343 32263 -14334 32297
rect -14386 32254 -14334 32263
rect -14226 32297 -14174 32306
rect -14226 32263 -14217 32297
rect -14217 32263 -14183 32297
rect -14183 32263 -14174 32297
rect -14226 32254 -14174 32263
rect -14066 32297 -14014 32306
rect -14066 32263 -14057 32297
rect -14057 32263 -14023 32297
rect -14023 32263 -14014 32297
rect -14066 32254 -14014 32263
rect -13906 32297 -13854 32306
rect -13906 32263 -13897 32297
rect -13897 32263 -13863 32297
rect -13863 32263 -13854 32297
rect -13906 32254 -13854 32263
rect -13746 32297 -13694 32306
rect -13746 32263 -13737 32297
rect -13737 32263 -13703 32297
rect -13703 32263 -13694 32297
rect -13746 32254 -13694 32263
rect -13586 32297 -13534 32306
rect -13586 32263 -13577 32297
rect -13577 32263 -13543 32297
rect -13543 32263 -13534 32297
rect -13586 32254 -13534 32263
rect -13426 32297 -13374 32306
rect -13426 32263 -13417 32297
rect -13417 32263 -13383 32297
rect -13383 32263 -13374 32297
rect -13426 32254 -13374 32263
rect -13266 32297 -13214 32306
rect -13266 32263 -13257 32297
rect -13257 32263 -13223 32297
rect -13223 32263 -13214 32297
rect -13266 32254 -13214 32263
rect -13106 32297 -13054 32306
rect -13106 32263 -13097 32297
rect -13097 32263 -13063 32297
rect -13063 32263 -13054 32297
rect -13106 32254 -13054 32263
rect -12946 32297 -12894 32306
rect -12946 32263 -12937 32297
rect -12937 32263 -12903 32297
rect -12903 32263 -12894 32297
rect -12946 32254 -12894 32263
rect -12786 32297 -12734 32306
rect -12786 32263 -12777 32297
rect -12777 32263 -12743 32297
rect -12743 32263 -12734 32297
rect -12786 32254 -12734 32263
rect -12626 32297 -12574 32306
rect -12626 32263 -12617 32297
rect -12617 32263 -12583 32297
rect -12583 32263 -12574 32297
rect -12626 32254 -12574 32263
rect -12466 32297 -12414 32306
rect -12466 32263 -12457 32297
rect -12457 32263 -12423 32297
rect -12423 32263 -12414 32297
rect -12466 32254 -12414 32263
rect -12306 32297 -12254 32306
rect -12306 32263 -12297 32297
rect -12297 32263 -12263 32297
rect -12263 32263 -12254 32297
rect -12306 32254 -12254 32263
rect -12146 32297 -12094 32306
rect -12146 32263 -12137 32297
rect -12137 32263 -12103 32297
rect -12103 32263 -12094 32297
rect -12146 32254 -12094 32263
rect -11986 32297 -11934 32306
rect -11986 32263 -11977 32297
rect -11977 32263 -11943 32297
rect -11943 32263 -11934 32297
rect -11986 32254 -11934 32263
rect -11826 32297 -11774 32306
rect -11826 32263 -11817 32297
rect -11817 32263 -11783 32297
rect -11783 32263 -11774 32297
rect -11826 32254 -11774 32263
rect -11666 32297 -11614 32306
rect -11666 32263 -11657 32297
rect -11657 32263 -11623 32297
rect -11623 32263 -11614 32297
rect -11666 32254 -11614 32263
rect -11506 32297 -11454 32306
rect -11506 32263 -11497 32297
rect -11497 32263 -11463 32297
rect -11463 32263 -11454 32297
rect -11506 32254 -11454 32263
rect -11346 32297 -11294 32306
rect -11346 32263 -11337 32297
rect -11337 32263 -11303 32297
rect -11303 32263 -11294 32297
rect -11346 32254 -11294 32263
rect -11186 32297 -11134 32306
rect -11186 32263 -11177 32297
rect -11177 32263 -11143 32297
rect -11143 32263 -11134 32297
rect -11186 32254 -11134 32263
rect -10866 32297 -10814 32306
rect -10866 32263 -10857 32297
rect -10857 32263 -10823 32297
rect -10823 32263 -10814 32297
rect -10866 32254 -10814 32263
rect -10706 32297 -10654 32306
rect -10706 32263 -10697 32297
rect -10697 32263 -10663 32297
rect -10663 32263 -10654 32297
rect -10706 32254 -10654 32263
rect -10546 32297 -10494 32306
rect -10546 32263 -10537 32297
rect -10537 32263 -10503 32297
rect -10503 32263 -10494 32297
rect -10546 32254 -10494 32263
rect -10386 32297 -10334 32306
rect -10386 32263 -10377 32297
rect -10377 32263 -10343 32297
rect -10343 32263 -10334 32297
rect -10386 32254 -10334 32263
rect -10226 32297 -10174 32306
rect -10226 32263 -10217 32297
rect -10217 32263 -10183 32297
rect -10183 32263 -10174 32297
rect -10226 32254 -10174 32263
rect -10066 32297 -10014 32306
rect -10066 32263 -10057 32297
rect -10057 32263 -10023 32297
rect -10023 32263 -10014 32297
rect -10066 32254 -10014 32263
rect -9906 32297 -9854 32306
rect -9906 32263 -9897 32297
rect -9897 32263 -9863 32297
rect -9863 32263 -9854 32297
rect -9906 32254 -9854 32263
rect -9746 32297 -9694 32306
rect -9746 32263 -9737 32297
rect -9737 32263 -9703 32297
rect -9703 32263 -9694 32297
rect -9746 32254 -9694 32263
rect -9586 32297 -9534 32306
rect -9586 32263 -9577 32297
rect -9577 32263 -9543 32297
rect -9543 32263 -9534 32297
rect -9586 32254 -9534 32263
rect -9426 32297 -9374 32306
rect -9426 32263 -9417 32297
rect -9417 32263 -9383 32297
rect -9383 32263 -9374 32297
rect -9426 32254 -9374 32263
rect -9266 32297 -9214 32306
rect -9266 32263 -9257 32297
rect -9257 32263 -9223 32297
rect -9223 32263 -9214 32297
rect -9266 32254 -9214 32263
rect -9106 32297 -9054 32306
rect -9106 32263 -9097 32297
rect -9097 32263 -9063 32297
rect -9063 32263 -9054 32297
rect -9106 32254 -9054 32263
rect -8946 32297 -8894 32306
rect -8946 32263 -8937 32297
rect -8937 32263 -8903 32297
rect -8903 32263 -8894 32297
rect -8946 32254 -8894 32263
rect -8786 32297 -8734 32306
rect -8786 32263 -8777 32297
rect -8777 32263 -8743 32297
rect -8743 32263 -8734 32297
rect -8786 32254 -8734 32263
rect -8626 32297 -8574 32306
rect -8626 32263 -8617 32297
rect -8617 32263 -8583 32297
rect -8583 32263 -8574 32297
rect -8626 32254 -8574 32263
rect -8466 32297 -8414 32306
rect -8466 32263 -8457 32297
rect -8457 32263 -8423 32297
rect -8423 32263 -8414 32297
rect -8466 32254 -8414 32263
rect -8306 32297 -8254 32306
rect -8306 32263 -8297 32297
rect -8297 32263 -8263 32297
rect -8263 32263 -8254 32297
rect -8306 32254 -8254 32263
rect -8146 32297 -8094 32306
rect -8146 32263 -8137 32297
rect -8137 32263 -8103 32297
rect -8103 32263 -8094 32297
rect -8146 32254 -8094 32263
rect -7986 32297 -7934 32306
rect -7986 32263 -7977 32297
rect -7977 32263 -7943 32297
rect -7943 32263 -7934 32297
rect -7986 32254 -7934 32263
rect -7826 32297 -7774 32306
rect -7826 32263 -7817 32297
rect -7817 32263 -7783 32297
rect -7783 32263 -7774 32297
rect -7826 32254 -7774 32263
rect -7666 32297 -7614 32306
rect -7666 32263 -7657 32297
rect -7657 32263 -7623 32297
rect -7623 32263 -7614 32297
rect -7666 32254 -7614 32263
rect -7506 32297 -7454 32306
rect -7506 32263 -7497 32297
rect -7497 32263 -7463 32297
rect -7463 32263 -7454 32297
rect -7506 32254 -7454 32263
rect -7346 32297 -7294 32306
rect -7346 32263 -7337 32297
rect -7337 32263 -7303 32297
rect -7303 32263 -7294 32297
rect -7346 32254 -7294 32263
rect -7186 32297 -7134 32306
rect -7186 32263 -7177 32297
rect -7177 32263 -7143 32297
rect -7143 32263 -7134 32297
rect -7186 32254 -7134 32263
rect -7026 32297 -6974 32306
rect -7026 32263 -7017 32297
rect -7017 32263 -6983 32297
rect -6983 32263 -6974 32297
rect -7026 32254 -6974 32263
rect -6866 32297 -6814 32306
rect -6866 32263 -6857 32297
rect -6857 32263 -6823 32297
rect -6823 32263 -6814 32297
rect -6866 32254 -6814 32263
rect -6706 32297 -6654 32306
rect -6706 32263 -6697 32297
rect -6697 32263 -6663 32297
rect -6663 32263 -6654 32297
rect -6706 32254 -6654 32263
rect -6546 32297 -6494 32306
rect -6546 32263 -6537 32297
rect -6537 32263 -6503 32297
rect -6503 32263 -6494 32297
rect -6546 32254 -6494 32263
rect -6386 32297 -6334 32306
rect -6386 32263 -6377 32297
rect -6377 32263 -6343 32297
rect -6343 32263 -6334 32297
rect -6386 32254 -6334 32263
rect -6226 32297 -6174 32306
rect -6226 32263 -6217 32297
rect -6217 32263 -6183 32297
rect -6183 32263 -6174 32297
rect -6226 32254 -6174 32263
rect -6066 32297 -6014 32306
rect -6066 32263 -6057 32297
rect -6057 32263 -6023 32297
rect -6023 32263 -6014 32297
rect -6066 32254 -6014 32263
rect -5906 32297 -5854 32306
rect -5906 32263 -5897 32297
rect -5897 32263 -5863 32297
rect -5863 32263 -5854 32297
rect -5906 32254 -5854 32263
rect -5746 32297 -5694 32306
rect -5746 32263 -5737 32297
rect -5737 32263 -5703 32297
rect -5703 32263 -5694 32297
rect -5746 32254 -5694 32263
rect -5586 32297 -5534 32306
rect -5586 32263 -5577 32297
rect -5577 32263 -5543 32297
rect -5543 32263 -5534 32297
rect -5586 32254 -5534 32263
rect -5426 32297 -5374 32306
rect -5426 32263 -5417 32297
rect -5417 32263 -5383 32297
rect -5383 32263 -5374 32297
rect -5426 32254 -5374 32263
rect -5266 32297 -5214 32306
rect -5266 32263 -5257 32297
rect -5257 32263 -5223 32297
rect -5223 32263 -5214 32297
rect -5266 32254 -5214 32263
rect -5106 32297 -5054 32306
rect -5106 32263 -5097 32297
rect -5097 32263 -5063 32297
rect -5063 32263 -5054 32297
rect -5106 32254 -5054 32263
rect -4946 32297 -4894 32306
rect -4946 32263 -4937 32297
rect -4937 32263 -4903 32297
rect -4903 32263 -4894 32297
rect -4946 32254 -4894 32263
rect -4786 32297 -4734 32306
rect -4786 32263 -4777 32297
rect -4777 32263 -4743 32297
rect -4743 32263 -4734 32297
rect -4786 32254 -4734 32263
rect -4626 32297 -4574 32306
rect -4626 32263 -4617 32297
rect -4617 32263 -4583 32297
rect -4583 32263 -4574 32297
rect -4626 32254 -4574 32263
rect -4466 32297 -4414 32306
rect -4466 32263 -4457 32297
rect -4457 32263 -4423 32297
rect -4423 32263 -4414 32297
rect -4466 32254 -4414 32263
rect -4306 32297 -4254 32306
rect -4306 32263 -4297 32297
rect -4297 32263 -4263 32297
rect -4263 32263 -4254 32297
rect -4306 32254 -4254 32263
rect -4146 32297 -4094 32306
rect -4146 32263 -4137 32297
rect -4137 32263 -4103 32297
rect -4103 32263 -4094 32297
rect -4146 32254 -4094 32263
rect -3986 32297 -3934 32306
rect -3986 32263 -3977 32297
rect -3977 32263 -3943 32297
rect -3943 32263 -3934 32297
rect -3986 32254 -3934 32263
rect -3666 32297 -3614 32306
rect -3666 32263 -3657 32297
rect -3657 32263 -3623 32297
rect -3623 32263 -3614 32297
rect -3666 32254 -3614 32263
rect -3506 32297 -3454 32306
rect -3506 32263 -3497 32297
rect -3497 32263 -3463 32297
rect -3463 32263 -3454 32297
rect -3506 32254 -3454 32263
rect -3346 32297 -3294 32306
rect -3346 32263 -3337 32297
rect -3337 32263 -3303 32297
rect -3303 32263 -3294 32297
rect -3346 32254 -3294 32263
rect -3186 32297 -3134 32306
rect -3186 32263 -3177 32297
rect -3177 32263 -3143 32297
rect -3143 32263 -3134 32297
rect -3186 32254 -3134 32263
rect -3026 32297 -2974 32306
rect -3026 32263 -3017 32297
rect -3017 32263 -2983 32297
rect -2983 32263 -2974 32297
rect -3026 32254 -2974 32263
rect -2866 32297 -2814 32306
rect -2866 32263 -2857 32297
rect -2857 32263 -2823 32297
rect -2823 32263 -2814 32297
rect -2866 32254 -2814 32263
rect -2706 32297 -2654 32306
rect -2706 32263 -2697 32297
rect -2697 32263 -2663 32297
rect -2663 32263 -2654 32297
rect -2706 32254 -2654 32263
rect -2386 32297 -2334 32306
rect -2386 32263 -2377 32297
rect -2377 32263 -2343 32297
rect -2343 32263 -2334 32297
rect -2386 32254 -2334 32263
rect -2066 32297 -2014 32306
rect -2066 32263 -2057 32297
rect -2057 32263 -2023 32297
rect -2023 32263 -2014 32297
rect -2066 32254 -2014 32263
rect -1746 32297 -1694 32306
rect -1746 32263 -1737 32297
rect -1737 32263 -1703 32297
rect -1703 32263 -1694 32297
rect -1746 32254 -1694 32263
rect -1426 32297 -1374 32306
rect -1426 32263 -1417 32297
rect -1417 32263 -1383 32297
rect -1383 32263 -1374 32297
rect -1426 32254 -1374 32263
rect -1106 32297 -1054 32306
rect -1106 32263 -1097 32297
rect -1097 32263 -1063 32297
rect -1063 32263 -1054 32297
rect -1106 32254 -1054 32263
rect -29906 31977 -29854 31986
rect -29906 31943 -29897 31977
rect -29897 31943 -29863 31977
rect -29863 31943 -29854 31977
rect -29906 31934 -29854 31943
rect -29746 31977 -29694 31986
rect -29746 31943 -29737 31977
rect -29737 31943 -29703 31977
rect -29703 31943 -29694 31977
rect -29746 31934 -29694 31943
rect -29586 31977 -29534 31986
rect -29586 31943 -29577 31977
rect -29577 31943 -29543 31977
rect -29543 31943 -29534 31977
rect -29586 31934 -29534 31943
rect -29426 31977 -29374 31986
rect -29426 31943 -29417 31977
rect -29417 31943 -29383 31977
rect -29383 31943 -29374 31977
rect -29426 31934 -29374 31943
rect -29266 31977 -29214 31986
rect -29266 31943 -29257 31977
rect -29257 31943 -29223 31977
rect -29223 31943 -29214 31977
rect -29266 31934 -29214 31943
rect -29106 31977 -29054 31986
rect -29106 31943 -29097 31977
rect -29097 31943 -29063 31977
rect -29063 31943 -29054 31977
rect -29106 31934 -29054 31943
rect -28946 31977 -28894 31986
rect -28946 31943 -28937 31977
rect -28937 31943 -28903 31977
rect -28903 31943 -28894 31977
rect -28946 31934 -28894 31943
rect -28786 31977 -28734 31986
rect -28786 31943 -28777 31977
rect -28777 31943 -28743 31977
rect -28743 31943 -28734 31977
rect -28786 31934 -28734 31943
rect -28626 31977 -28574 31986
rect -28626 31943 -28617 31977
rect -28617 31943 -28583 31977
rect -28583 31943 -28574 31977
rect -28626 31934 -28574 31943
rect -28466 31977 -28414 31986
rect -28466 31943 -28457 31977
rect -28457 31943 -28423 31977
rect -28423 31943 -28414 31977
rect -28466 31934 -28414 31943
rect -28306 31977 -28254 31986
rect -28306 31943 -28297 31977
rect -28297 31943 -28263 31977
rect -28263 31943 -28254 31977
rect -28306 31934 -28254 31943
rect -28146 31977 -28094 31986
rect -28146 31943 -28137 31977
rect -28137 31943 -28103 31977
rect -28103 31943 -28094 31977
rect -28146 31934 -28094 31943
rect -27986 31977 -27934 31986
rect -27986 31943 -27977 31977
rect -27977 31943 -27943 31977
rect -27943 31943 -27934 31977
rect -27986 31934 -27934 31943
rect -27826 31977 -27774 31986
rect -27826 31943 -27817 31977
rect -27817 31943 -27783 31977
rect -27783 31943 -27774 31977
rect -27826 31934 -27774 31943
rect -27666 31977 -27614 31986
rect -27666 31943 -27657 31977
rect -27657 31943 -27623 31977
rect -27623 31943 -27614 31977
rect -27666 31934 -27614 31943
rect -27506 31977 -27454 31986
rect -27506 31943 -27497 31977
rect -27497 31943 -27463 31977
rect -27463 31943 -27454 31977
rect -27506 31934 -27454 31943
rect -27346 31977 -27294 31986
rect -27346 31943 -27337 31977
rect -27337 31943 -27303 31977
rect -27303 31943 -27294 31977
rect -27346 31934 -27294 31943
rect -27186 31977 -27134 31986
rect -27186 31943 -27177 31977
rect -27177 31943 -27143 31977
rect -27143 31943 -27134 31977
rect -27186 31934 -27134 31943
rect -27026 31977 -26974 31986
rect -27026 31943 -27017 31977
rect -27017 31943 -26983 31977
rect -26983 31943 -26974 31977
rect -27026 31934 -26974 31943
rect -26866 31977 -26814 31986
rect -26866 31943 -26857 31977
rect -26857 31943 -26823 31977
rect -26823 31943 -26814 31977
rect -26866 31934 -26814 31943
rect -26706 31977 -26654 31986
rect -26706 31943 -26697 31977
rect -26697 31943 -26663 31977
rect -26663 31943 -26654 31977
rect -26706 31934 -26654 31943
rect -26546 31977 -26494 31986
rect -26546 31943 -26537 31977
rect -26537 31943 -26503 31977
rect -26503 31943 -26494 31977
rect -26546 31934 -26494 31943
rect -26386 31977 -26334 31986
rect -26386 31943 -26377 31977
rect -26377 31943 -26343 31977
rect -26343 31943 -26334 31977
rect -26386 31934 -26334 31943
rect -26226 31977 -26174 31986
rect -26226 31943 -26217 31977
rect -26217 31943 -26183 31977
rect -26183 31943 -26174 31977
rect -26226 31934 -26174 31943
rect -26066 31977 -26014 31986
rect -26066 31943 -26057 31977
rect -26057 31943 -26023 31977
rect -26023 31943 -26014 31977
rect -26066 31934 -26014 31943
rect -25906 31977 -25854 31986
rect -25906 31943 -25897 31977
rect -25897 31943 -25863 31977
rect -25863 31943 -25854 31977
rect -25906 31934 -25854 31943
rect -25746 31977 -25694 31986
rect -25746 31943 -25737 31977
rect -25737 31943 -25703 31977
rect -25703 31943 -25694 31977
rect -25746 31934 -25694 31943
rect -25586 31977 -25534 31986
rect -25586 31943 -25577 31977
rect -25577 31943 -25543 31977
rect -25543 31943 -25534 31977
rect -25586 31934 -25534 31943
rect -25426 31977 -25374 31986
rect -25426 31943 -25417 31977
rect -25417 31943 -25383 31977
rect -25383 31943 -25374 31977
rect -25426 31934 -25374 31943
rect -25266 31977 -25214 31986
rect -25266 31943 -25257 31977
rect -25257 31943 -25223 31977
rect -25223 31943 -25214 31977
rect -25266 31934 -25214 31943
rect -25106 31977 -25054 31986
rect -25106 31943 -25097 31977
rect -25097 31943 -25063 31977
rect -25063 31943 -25054 31977
rect -25106 31934 -25054 31943
rect -24946 31977 -24894 31986
rect -24946 31943 -24937 31977
rect -24937 31943 -24903 31977
rect -24903 31943 -24894 31977
rect -24946 31934 -24894 31943
rect -24786 31977 -24734 31986
rect -24786 31943 -24777 31977
rect -24777 31943 -24743 31977
rect -24743 31943 -24734 31977
rect -24786 31934 -24734 31943
rect -24626 31977 -24574 31986
rect -24626 31943 -24617 31977
rect -24617 31943 -24583 31977
rect -24583 31943 -24574 31977
rect -24626 31934 -24574 31943
rect -24466 31977 -24414 31986
rect -24466 31943 -24457 31977
rect -24457 31943 -24423 31977
rect -24423 31943 -24414 31977
rect -24466 31934 -24414 31943
rect -24306 31977 -24254 31986
rect -24306 31943 -24297 31977
rect -24297 31943 -24263 31977
rect -24263 31943 -24254 31977
rect -24306 31934 -24254 31943
rect -24146 31977 -24094 31986
rect -24146 31943 -24137 31977
rect -24137 31943 -24103 31977
rect -24103 31943 -24094 31977
rect -24146 31934 -24094 31943
rect -23986 31977 -23934 31986
rect -23986 31943 -23977 31977
rect -23977 31943 -23943 31977
rect -23943 31943 -23934 31977
rect -23986 31934 -23934 31943
rect -23826 31977 -23774 31986
rect -23826 31943 -23817 31977
rect -23817 31943 -23783 31977
rect -23783 31943 -23774 31977
rect -23826 31934 -23774 31943
rect -23666 31977 -23614 31986
rect -23666 31943 -23657 31977
rect -23657 31943 -23623 31977
rect -23623 31943 -23614 31977
rect -23666 31934 -23614 31943
rect -23506 31977 -23454 31986
rect -23506 31943 -23497 31977
rect -23497 31943 -23463 31977
rect -23463 31943 -23454 31977
rect -23506 31934 -23454 31943
rect -23346 31977 -23294 31986
rect -23346 31943 -23337 31977
rect -23337 31943 -23303 31977
rect -23303 31943 -23294 31977
rect -23346 31934 -23294 31943
rect -23186 31977 -23134 31986
rect -23186 31943 -23177 31977
rect -23177 31943 -23143 31977
rect -23143 31943 -23134 31977
rect -23186 31934 -23134 31943
rect -23026 31977 -22974 31986
rect -23026 31943 -23017 31977
rect -23017 31943 -22983 31977
rect -22983 31943 -22974 31977
rect -23026 31934 -22974 31943
rect -22866 31977 -22814 31986
rect -22866 31943 -22857 31977
rect -22857 31943 -22823 31977
rect -22823 31943 -22814 31977
rect -22866 31934 -22814 31943
rect -22706 31977 -22654 31986
rect -22706 31943 -22697 31977
rect -22697 31943 -22663 31977
rect -22663 31943 -22654 31977
rect -22706 31934 -22654 31943
rect -22546 31977 -22494 31986
rect -22546 31943 -22537 31977
rect -22537 31943 -22503 31977
rect -22503 31943 -22494 31977
rect -22546 31934 -22494 31943
rect -22386 31977 -22334 31986
rect -22386 31943 -22377 31977
rect -22377 31943 -22343 31977
rect -22343 31943 -22334 31977
rect -22386 31934 -22334 31943
rect -22226 31977 -22174 31986
rect -22226 31943 -22217 31977
rect -22217 31943 -22183 31977
rect -22183 31943 -22174 31977
rect -22226 31934 -22174 31943
rect -22066 31977 -22014 31986
rect -22066 31943 -22057 31977
rect -22057 31943 -22023 31977
rect -22023 31943 -22014 31977
rect -22066 31934 -22014 31943
rect -21906 31977 -21854 31986
rect -21906 31943 -21897 31977
rect -21897 31943 -21863 31977
rect -21863 31943 -21854 31977
rect -21906 31934 -21854 31943
rect -21746 31977 -21694 31986
rect -21746 31943 -21737 31977
rect -21737 31943 -21703 31977
rect -21703 31943 -21694 31977
rect -21746 31934 -21694 31943
rect -21586 31977 -21534 31986
rect -21586 31943 -21577 31977
rect -21577 31943 -21543 31977
rect -21543 31943 -21534 31977
rect -21586 31934 -21534 31943
rect -21426 31977 -21374 31986
rect -21426 31943 -21417 31977
rect -21417 31943 -21383 31977
rect -21383 31943 -21374 31977
rect -21426 31934 -21374 31943
rect -21266 31977 -21214 31986
rect -21266 31943 -21257 31977
rect -21257 31943 -21223 31977
rect -21223 31943 -21214 31977
rect -21266 31934 -21214 31943
rect -21106 31977 -21054 31986
rect -21106 31943 -21097 31977
rect -21097 31943 -21063 31977
rect -21063 31943 -21054 31977
rect -21106 31934 -21054 31943
rect -20946 31977 -20894 31986
rect -20946 31943 -20937 31977
rect -20937 31943 -20903 31977
rect -20903 31943 -20894 31977
rect -20946 31934 -20894 31943
rect -20786 31977 -20734 31986
rect -20786 31943 -20777 31977
rect -20777 31943 -20743 31977
rect -20743 31943 -20734 31977
rect -20786 31934 -20734 31943
rect -20626 31977 -20574 31986
rect -20626 31943 -20617 31977
rect -20617 31943 -20583 31977
rect -20583 31943 -20574 31977
rect -20626 31934 -20574 31943
rect -20466 31977 -20414 31986
rect -20466 31943 -20457 31977
rect -20457 31943 -20423 31977
rect -20423 31943 -20414 31977
rect -20466 31934 -20414 31943
rect -20306 31977 -20254 31986
rect -20306 31943 -20297 31977
rect -20297 31943 -20263 31977
rect -20263 31943 -20254 31977
rect -20306 31934 -20254 31943
rect -20146 31977 -20094 31986
rect -20146 31943 -20137 31977
rect -20137 31943 -20103 31977
rect -20103 31943 -20094 31977
rect -20146 31934 -20094 31943
rect -19986 31977 -19934 31986
rect -19986 31943 -19977 31977
rect -19977 31943 -19943 31977
rect -19943 31943 -19934 31977
rect -19986 31934 -19934 31943
rect -19826 31977 -19774 31986
rect -19826 31943 -19817 31977
rect -19817 31943 -19783 31977
rect -19783 31943 -19774 31977
rect -19826 31934 -19774 31943
rect -19666 31977 -19614 31986
rect -19666 31943 -19657 31977
rect -19657 31943 -19623 31977
rect -19623 31943 -19614 31977
rect -19666 31934 -19614 31943
rect -19506 31977 -19454 31986
rect -19506 31943 -19497 31977
rect -19497 31943 -19463 31977
rect -19463 31943 -19454 31977
rect -19506 31934 -19454 31943
rect -19346 31977 -19294 31986
rect -19346 31943 -19337 31977
rect -19337 31943 -19303 31977
rect -19303 31943 -19294 31977
rect -19346 31934 -19294 31943
rect -19186 31977 -19134 31986
rect -19186 31943 -19177 31977
rect -19177 31943 -19143 31977
rect -19143 31943 -19134 31977
rect -19186 31934 -19134 31943
rect -19026 31977 -18974 31986
rect -19026 31943 -19017 31977
rect -19017 31943 -18983 31977
rect -18983 31943 -18974 31977
rect -19026 31934 -18974 31943
rect -18866 31977 -18814 31986
rect -18866 31943 -18857 31977
rect -18857 31943 -18823 31977
rect -18823 31943 -18814 31977
rect -18866 31934 -18814 31943
rect -18706 31977 -18654 31986
rect -18706 31943 -18697 31977
rect -18697 31943 -18663 31977
rect -18663 31943 -18654 31977
rect -18706 31934 -18654 31943
rect -18546 31977 -18494 31986
rect -18546 31943 -18537 31977
rect -18537 31943 -18503 31977
rect -18503 31943 -18494 31977
rect -18546 31934 -18494 31943
rect -18386 31977 -18334 31986
rect -18386 31943 -18377 31977
rect -18377 31943 -18343 31977
rect -18343 31943 -18334 31977
rect -18386 31934 -18334 31943
rect -18226 31977 -18174 31986
rect -18226 31943 -18217 31977
rect -18217 31943 -18183 31977
rect -18183 31943 -18174 31977
rect -18226 31934 -18174 31943
rect -18066 31977 -18014 31986
rect -18066 31943 -18057 31977
rect -18057 31943 -18023 31977
rect -18023 31943 -18014 31977
rect -18066 31934 -18014 31943
rect -17906 31977 -17854 31986
rect -17906 31943 -17897 31977
rect -17897 31943 -17863 31977
rect -17863 31943 -17854 31977
rect -17906 31934 -17854 31943
rect -17746 31977 -17694 31986
rect -17746 31943 -17737 31977
rect -17737 31943 -17703 31977
rect -17703 31943 -17694 31977
rect -17746 31934 -17694 31943
rect -17586 31977 -17534 31986
rect -17586 31943 -17577 31977
rect -17577 31943 -17543 31977
rect -17543 31943 -17534 31977
rect -17586 31934 -17534 31943
rect -17426 31977 -17374 31986
rect -17426 31943 -17417 31977
rect -17417 31943 -17383 31977
rect -17383 31943 -17374 31977
rect -17426 31934 -17374 31943
rect -17266 31977 -17214 31986
rect -17266 31943 -17257 31977
rect -17257 31943 -17223 31977
rect -17223 31943 -17214 31977
rect -17266 31934 -17214 31943
rect -17106 31977 -17054 31986
rect -17106 31943 -17097 31977
rect -17097 31943 -17063 31977
rect -17063 31943 -17054 31977
rect -17106 31934 -17054 31943
rect -16946 31977 -16894 31986
rect -16946 31943 -16937 31977
rect -16937 31943 -16903 31977
rect -16903 31943 -16894 31977
rect -16946 31934 -16894 31943
rect -16786 31977 -16734 31986
rect -16786 31943 -16777 31977
rect -16777 31943 -16743 31977
rect -16743 31943 -16734 31977
rect -16786 31934 -16734 31943
rect -16626 31977 -16574 31986
rect -16626 31943 -16617 31977
rect -16617 31943 -16583 31977
rect -16583 31943 -16574 31977
rect -16626 31934 -16574 31943
rect -16466 31977 -16414 31986
rect -16466 31943 -16457 31977
rect -16457 31943 -16423 31977
rect -16423 31943 -16414 31977
rect -16466 31934 -16414 31943
rect -16306 31977 -16254 31986
rect -16306 31943 -16297 31977
rect -16297 31943 -16263 31977
rect -16263 31943 -16254 31977
rect -16306 31934 -16254 31943
rect -16146 31977 -16094 31986
rect -16146 31943 -16137 31977
rect -16137 31943 -16103 31977
rect -16103 31943 -16094 31977
rect -16146 31934 -16094 31943
rect -15986 31977 -15934 31986
rect -15986 31943 -15977 31977
rect -15977 31943 -15943 31977
rect -15943 31943 -15934 31977
rect -15986 31934 -15934 31943
rect -15826 31977 -15774 31986
rect -15826 31943 -15817 31977
rect -15817 31943 -15783 31977
rect -15783 31943 -15774 31977
rect -15826 31934 -15774 31943
rect -15666 31977 -15614 31986
rect -15666 31943 -15657 31977
rect -15657 31943 -15623 31977
rect -15623 31943 -15614 31977
rect -15666 31934 -15614 31943
rect -15506 31977 -15454 31986
rect -15506 31943 -15497 31977
rect -15497 31943 -15463 31977
rect -15463 31943 -15454 31977
rect -15506 31934 -15454 31943
rect -15346 31977 -15294 31986
rect -15346 31943 -15337 31977
rect -15337 31943 -15303 31977
rect -15303 31943 -15294 31977
rect -15346 31934 -15294 31943
rect -15186 31977 -15134 31986
rect -15186 31943 -15177 31977
rect -15177 31943 -15143 31977
rect -15143 31943 -15134 31977
rect -15186 31934 -15134 31943
rect -15026 31977 -14974 31986
rect -15026 31943 -15017 31977
rect -15017 31943 -14983 31977
rect -14983 31943 -14974 31977
rect -15026 31934 -14974 31943
rect -14866 31977 -14814 31986
rect -14866 31943 -14857 31977
rect -14857 31943 -14823 31977
rect -14823 31943 -14814 31977
rect -14866 31934 -14814 31943
rect -14706 31977 -14654 31986
rect -14706 31943 -14697 31977
rect -14697 31943 -14663 31977
rect -14663 31943 -14654 31977
rect -14706 31934 -14654 31943
rect -14546 31977 -14494 31986
rect -14546 31943 -14537 31977
rect -14537 31943 -14503 31977
rect -14503 31943 -14494 31977
rect -14546 31934 -14494 31943
rect -14386 31977 -14334 31986
rect -14386 31943 -14377 31977
rect -14377 31943 -14343 31977
rect -14343 31943 -14334 31977
rect -14386 31934 -14334 31943
rect -14226 31977 -14174 31986
rect -14226 31943 -14217 31977
rect -14217 31943 -14183 31977
rect -14183 31943 -14174 31977
rect -14226 31934 -14174 31943
rect -14066 31977 -14014 31986
rect -14066 31943 -14057 31977
rect -14057 31943 -14023 31977
rect -14023 31943 -14014 31977
rect -14066 31934 -14014 31943
rect -13906 31977 -13854 31986
rect -13906 31943 -13897 31977
rect -13897 31943 -13863 31977
rect -13863 31943 -13854 31977
rect -13906 31934 -13854 31943
rect -13746 31977 -13694 31986
rect -13746 31943 -13737 31977
rect -13737 31943 -13703 31977
rect -13703 31943 -13694 31977
rect -13746 31934 -13694 31943
rect -13586 31977 -13534 31986
rect -13586 31943 -13577 31977
rect -13577 31943 -13543 31977
rect -13543 31943 -13534 31977
rect -13586 31934 -13534 31943
rect -13426 31977 -13374 31986
rect -13426 31943 -13417 31977
rect -13417 31943 -13383 31977
rect -13383 31943 -13374 31977
rect -13426 31934 -13374 31943
rect -13266 31977 -13214 31986
rect -13266 31943 -13257 31977
rect -13257 31943 -13223 31977
rect -13223 31943 -13214 31977
rect -13266 31934 -13214 31943
rect -13106 31977 -13054 31986
rect -13106 31943 -13097 31977
rect -13097 31943 -13063 31977
rect -13063 31943 -13054 31977
rect -13106 31934 -13054 31943
rect -12946 31977 -12894 31986
rect -12946 31943 -12937 31977
rect -12937 31943 -12903 31977
rect -12903 31943 -12894 31977
rect -12946 31934 -12894 31943
rect -12786 31977 -12734 31986
rect -12786 31943 -12777 31977
rect -12777 31943 -12743 31977
rect -12743 31943 -12734 31977
rect -12786 31934 -12734 31943
rect -12626 31977 -12574 31986
rect -12626 31943 -12617 31977
rect -12617 31943 -12583 31977
rect -12583 31943 -12574 31977
rect -12626 31934 -12574 31943
rect -12466 31977 -12414 31986
rect -12466 31943 -12457 31977
rect -12457 31943 -12423 31977
rect -12423 31943 -12414 31977
rect -12466 31934 -12414 31943
rect -12306 31977 -12254 31986
rect -12306 31943 -12297 31977
rect -12297 31943 -12263 31977
rect -12263 31943 -12254 31977
rect -12306 31934 -12254 31943
rect -12146 31977 -12094 31986
rect -12146 31943 -12137 31977
rect -12137 31943 -12103 31977
rect -12103 31943 -12094 31977
rect -12146 31934 -12094 31943
rect -11986 31977 -11934 31986
rect -11986 31943 -11977 31977
rect -11977 31943 -11943 31977
rect -11943 31943 -11934 31977
rect -11986 31934 -11934 31943
rect -11826 31977 -11774 31986
rect -11826 31943 -11817 31977
rect -11817 31943 -11783 31977
rect -11783 31943 -11774 31977
rect -11826 31934 -11774 31943
rect -11666 31977 -11614 31986
rect -11666 31943 -11657 31977
rect -11657 31943 -11623 31977
rect -11623 31943 -11614 31977
rect -11666 31934 -11614 31943
rect -11506 31977 -11454 31986
rect -11506 31943 -11497 31977
rect -11497 31943 -11463 31977
rect -11463 31943 -11454 31977
rect -11506 31934 -11454 31943
rect -11346 31977 -11294 31986
rect -11346 31943 -11337 31977
rect -11337 31943 -11303 31977
rect -11303 31943 -11294 31977
rect -11346 31934 -11294 31943
rect -11186 31977 -11134 31986
rect -11186 31943 -11177 31977
rect -11177 31943 -11143 31977
rect -11143 31943 -11134 31977
rect -11186 31934 -11134 31943
rect -10866 31977 -10814 31986
rect -10866 31943 -10857 31977
rect -10857 31943 -10823 31977
rect -10823 31943 -10814 31977
rect -10866 31934 -10814 31943
rect -10706 31977 -10654 31986
rect -10706 31943 -10697 31977
rect -10697 31943 -10663 31977
rect -10663 31943 -10654 31977
rect -10706 31934 -10654 31943
rect -10546 31977 -10494 31986
rect -10546 31943 -10537 31977
rect -10537 31943 -10503 31977
rect -10503 31943 -10494 31977
rect -10546 31934 -10494 31943
rect -10386 31977 -10334 31986
rect -10386 31943 -10377 31977
rect -10377 31943 -10343 31977
rect -10343 31943 -10334 31977
rect -10386 31934 -10334 31943
rect -10226 31977 -10174 31986
rect -10226 31943 -10217 31977
rect -10217 31943 -10183 31977
rect -10183 31943 -10174 31977
rect -10226 31934 -10174 31943
rect -10066 31977 -10014 31986
rect -10066 31943 -10057 31977
rect -10057 31943 -10023 31977
rect -10023 31943 -10014 31977
rect -10066 31934 -10014 31943
rect -9906 31977 -9854 31986
rect -9906 31943 -9897 31977
rect -9897 31943 -9863 31977
rect -9863 31943 -9854 31977
rect -9906 31934 -9854 31943
rect -9746 31977 -9694 31986
rect -9746 31943 -9737 31977
rect -9737 31943 -9703 31977
rect -9703 31943 -9694 31977
rect -9746 31934 -9694 31943
rect -9586 31977 -9534 31986
rect -9586 31943 -9577 31977
rect -9577 31943 -9543 31977
rect -9543 31943 -9534 31977
rect -9586 31934 -9534 31943
rect -9426 31977 -9374 31986
rect -9426 31943 -9417 31977
rect -9417 31943 -9383 31977
rect -9383 31943 -9374 31977
rect -9426 31934 -9374 31943
rect -9266 31977 -9214 31986
rect -9266 31943 -9257 31977
rect -9257 31943 -9223 31977
rect -9223 31943 -9214 31977
rect -9266 31934 -9214 31943
rect -9106 31977 -9054 31986
rect -9106 31943 -9097 31977
rect -9097 31943 -9063 31977
rect -9063 31943 -9054 31977
rect -9106 31934 -9054 31943
rect -8946 31977 -8894 31986
rect -8946 31943 -8937 31977
rect -8937 31943 -8903 31977
rect -8903 31943 -8894 31977
rect -8946 31934 -8894 31943
rect -8786 31977 -8734 31986
rect -8786 31943 -8777 31977
rect -8777 31943 -8743 31977
rect -8743 31943 -8734 31977
rect -8786 31934 -8734 31943
rect -8626 31977 -8574 31986
rect -8626 31943 -8617 31977
rect -8617 31943 -8583 31977
rect -8583 31943 -8574 31977
rect -8626 31934 -8574 31943
rect -8466 31977 -8414 31986
rect -8466 31943 -8457 31977
rect -8457 31943 -8423 31977
rect -8423 31943 -8414 31977
rect -8466 31934 -8414 31943
rect -8306 31977 -8254 31986
rect -8306 31943 -8297 31977
rect -8297 31943 -8263 31977
rect -8263 31943 -8254 31977
rect -8306 31934 -8254 31943
rect -8146 31977 -8094 31986
rect -8146 31943 -8137 31977
rect -8137 31943 -8103 31977
rect -8103 31943 -8094 31977
rect -8146 31934 -8094 31943
rect -7986 31977 -7934 31986
rect -7986 31943 -7977 31977
rect -7977 31943 -7943 31977
rect -7943 31943 -7934 31977
rect -7986 31934 -7934 31943
rect -7826 31977 -7774 31986
rect -7826 31943 -7817 31977
rect -7817 31943 -7783 31977
rect -7783 31943 -7774 31977
rect -7826 31934 -7774 31943
rect -7666 31977 -7614 31986
rect -7666 31943 -7657 31977
rect -7657 31943 -7623 31977
rect -7623 31943 -7614 31977
rect -7666 31934 -7614 31943
rect -7506 31977 -7454 31986
rect -7506 31943 -7497 31977
rect -7497 31943 -7463 31977
rect -7463 31943 -7454 31977
rect -7506 31934 -7454 31943
rect -7346 31977 -7294 31986
rect -7346 31943 -7337 31977
rect -7337 31943 -7303 31977
rect -7303 31943 -7294 31977
rect -7346 31934 -7294 31943
rect -7186 31977 -7134 31986
rect -7186 31943 -7177 31977
rect -7177 31943 -7143 31977
rect -7143 31943 -7134 31977
rect -7186 31934 -7134 31943
rect -7026 31977 -6974 31986
rect -7026 31943 -7017 31977
rect -7017 31943 -6983 31977
rect -6983 31943 -6974 31977
rect -7026 31934 -6974 31943
rect -6866 31977 -6814 31986
rect -6866 31943 -6857 31977
rect -6857 31943 -6823 31977
rect -6823 31943 -6814 31977
rect -6866 31934 -6814 31943
rect -6706 31977 -6654 31986
rect -6706 31943 -6697 31977
rect -6697 31943 -6663 31977
rect -6663 31943 -6654 31977
rect -6706 31934 -6654 31943
rect -6546 31977 -6494 31986
rect -6546 31943 -6537 31977
rect -6537 31943 -6503 31977
rect -6503 31943 -6494 31977
rect -6546 31934 -6494 31943
rect -6386 31977 -6334 31986
rect -6386 31943 -6377 31977
rect -6377 31943 -6343 31977
rect -6343 31943 -6334 31977
rect -6386 31934 -6334 31943
rect -6226 31977 -6174 31986
rect -6226 31943 -6217 31977
rect -6217 31943 -6183 31977
rect -6183 31943 -6174 31977
rect -6226 31934 -6174 31943
rect -6066 31977 -6014 31986
rect -6066 31943 -6057 31977
rect -6057 31943 -6023 31977
rect -6023 31943 -6014 31977
rect -6066 31934 -6014 31943
rect -5906 31977 -5854 31986
rect -5906 31943 -5897 31977
rect -5897 31943 -5863 31977
rect -5863 31943 -5854 31977
rect -5906 31934 -5854 31943
rect -5746 31977 -5694 31986
rect -5746 31943 -5737 31977
rect -5737 31943 -5703 31977
rect -5703 31943 -5694 31977
rect -5746 31934 -5694 31943
rect -5586 31977 -5534 31986
rect -5586 31943 -5577 31977
rect -5577 31943 -5543 31977
rect -5543 31943 -5534 31977
rect -5586 31934 -5534 31943
rect -5426 31977 -5374 31986
rect -5426 31943 -5417 31977
rect -5417 31943 -5383 31977
rect -5383 31943 -5374 31977
rect -5426 31934 -5374 31943
rect -5266 31977 -5214 31986
rect -5266 31943 -5257 31977
rect -5257 31943 -5223 31977
rect -5223 31943 -5214 31977
rect -5266 31934 -5214 31943
rect -5106 31977 -5054 31986
rect -5106 31943 -5097 31977
rect -5097 31943 -5063 31977
rect -5063 31943 -5054 31977
rect -5106 31934 -5054 31943
rect -4946 31977 -4894 31986
rect -4946 31943 -4937 31977
rect -4937 31943 -4903 31977
rect -4903 31943 -4894 31977
rect -4946 31934 -4894 31943
rect -4786 31977 -4734 31986
rect -4786 31943 -4777 31977
rect -4777 31943 -4743 31977
rect -4743 31943 -4734 31977
rect -4786 31934 -4734 31943
rect -4626 31977 -4574 31986
rect -4626 31943 -4617 31977
rect -4617 31943 -4583 31977
rect -4583 31943 -4574 31977
rect -4626 31934 -4574 31943
rect -4466 31977 -4414 31986
rect -4466 31943 -4457 31977
rect -4457 31943 -4423 31977
rect -4423 31943 -4414 31977
rect -4466 31934 -4414 31943
rect -4306 31977 -4254 31986
rect -4306 31943 -4297 31977
rect -4297 31943 -4263 31977
rect -4263 31943 -4254 31977
rect -4306 31934 -4254 31943
rect -4146 31977 -4094 31986
rect -4146 31943 -4137 31977
rect -4137 31943 -4103 31977
rect -4103 31943 -4094 31977
rect -4146 31934 -4094 31943
rect -3986 31977 -3934 31986
rect -3986 31943 -3977 31977
rect -3977 31943 -3943 31977
rect -3943 31943 -3934 31977
rect -3986 31934 -3934 31943
rect -3666 31977 -3614 31986
rect -3666 31943 -3657 31977
rect -3657 31943 -3623 31977
rect -3623 31943 -3614 31977
rect -3666 31934 -3614 31943
rect -3506 31977 -3454 31986
rect -3506 31943 -3497 31977
rect -3497 31943 -3463 31977
rect -3463 31943 -3454 31977
rect -3506 31934 -3454 31943
rect -3346 31977 -3294 31986
rect -3346 31943 -3337 31977
rect -3337 31943 -3303 31977
rect -3303 31943 -3294 31977
rect -3346 31934 -3294 31943
rect -3186 31977 -3134 31986
rect -3186 31943 -3177 31977
rect -3177 31943 -3143 31977
rect -3143 31943 -3134 31977
rect -3186 31934 -3134 31943
rect -3026 31977 -2974 31986
rect -3026 31943 -3017 31977
rect -3017 31943 -2983 31977
rect -2983 31943 -2974 31977
rect -3026 31934 -2974 31943
rect -2866 31977 -2814 31986
rect -2866 31943 -2857 31977
rect -2857 31943 -2823 31977
rect -2823 31943 -2814 31977
rect -2866 31934 -2814 31943
rect -2706 31977 -2654 31986
rect -2706 31943 -2697 31977
rect -2697 31943 -2663 31977
rect -2663 31943 -2654 31977
rect -2706 31934 -2654 31943
rect -2386 31977 -2334 31986
rect -2386 31943 -2377 31977
rect -2377 31943 -2343 31977
rect -2343 31943 -2334 31977
rect -2386 31934 -2334 31943
rect -2066 31977 -2014 31986
rect -2066 31943 -2057 31977
rect -2057 31943 -2023 31977
rect -2023 31943 -2014 31977
rect -2066 31934 -2014 31943
rect -1746 31977 -1694 31986
rect -1746 31943 -1737 31977
rect -1737 31943 -1703 31977
rect -1703 31943 -1694 31977
rect -1746 31934 -1694 31943
rect -1426 31977 -1374 31986
rect -1426 31943 -1417 31977
rect -1417 31943 -1383 31977
rect -1383 31943 -1374 31977
rect -1426 31934 -1374 31943
rect -1106 31977 -1054 31986
rect -1106 31943 -1097 31977
rect -1097 31943 -1063 31977
rect -1063 31943 -1054 31977
rect -1106 31934 -1054 31943
<< metal2 >>
rect -31040 42868 -1040 42880
rect -31040 42812 -31028 42868
rect -30972 42812 -30708 42868
rect -30652 42812 -30388 42868
rect -30332 42812 -30068 42868
rect -30012 42812 -29908 42868
rect -29852 42812 -29748 42868
rect -29692 42812 -29588 42868
rect -29532 42812 -29428 42868
rect -29372 42812 -29268 42868
rect -29212 42812 -29108 42868
rect -29052 42812 -28948 42868
rect -28892 42812 -28788 42868
rect -28732 42812 -28628 42868
rect -28572 42812 -28468 42868
rect -28412 42812 -28308 42868
rect -28252 42812 -28148 42868
rect -28092 42812 -27988 42868
rect -27932 42812 -27828 42868
rect -27772 42812 -27668 42868
rect -27612 42812 -27508 42868
rect -27452 42812 -27348 42868
rect -27292 42812 -27188 42868
rect -27132 42812 -27028 42868
rect -26972 42812 -26868 42868
rect -26812 42812 -26708 42868
rect -26652 42812 -26548 42868
rect -26492 42812 -26388 42868
rect -26332 42812 -26228 42868
rect -26172 42812 -26068 42868
rect -26012 42812 -25908 42868
rect -25852 42812 -25748 42868
rect -25692 42812 -25588 42868
rect -25532 42812 -25428 42868
rect -25372 42812 -25268 42868
rect -25212 42812 -25108 42868
rect -25052 42812 -24948 42868
rect -24892 42812 -24788 42868
rect -24732 42812 -24628 42868
rect -24572 42812 -24468 42868
rect -24412 42812 -24308 42868
rect -24252 42812 -24148 42868
rect -24092 42812 -23988 42868
rect -23932 42812 -23828 42868
rect -23772 42812 -23668 42868
rect -23612 42812 -23508 42868
rect -23452 42812 -23348 42868
rect -23292 42812 -23188 42868
rect -23132 42812 -23028 42868
rect -22972 42812 -22868 42868
rect -22812 42812 -22708 42868
rect -22652 42812 -22548 42868
rect -22492 42812 -22388 42868
rect -22332 42812 -22228 42868
rect -22172 42812 -22068 42868
rect -22012 42812 -21908 42868
rect -21852 42812 -21748 42868
rect -21692 42812 -21588 42868
rect -21532 42812 -21428 42868
rect -21372 42812 -21268 42868
rect -21212 42812 -21108 42868
rect -21052 42812 -20948 42868
rect -20892 42812 -20788 42868
rect -20732 42812 -20628 42868
rect -20572 42812 -20468 42868
rect -20412 42812 -20308 42868
rect -20252 42812 -20148 42868
rect -20092 42812 -19988 42868
rect -19932 42812 -19828 42868
rect -19772 42812 -19668 42868
rect -19612 42812 -19508 42868
rect -19452 42812 -19348 42868
rect -19292 42812 -19188 42868
rect -19132 42812 -19028 42868
rect -18972 42812 -18868 42868
rect -18812 42812 -18708 42868
rect -18652 42812 -18548 42868
rect -18492 42812 -18388 42868
rect -18332 42812 -18228 42868
rect -18172 42812 -18068 42868
rect -18012 42812 -17908 42868
rect -17852 42812 -17748 42868
rect -17692 42812 -17588 42868
rect -17532 42812 -17428 42868
rect -17372 42812 -17268 42868
rect -17212 42812 -17108 42868
rect -17052 42812 -16948 42868
rect -16892 42812 -16788 42868
rect -16732 42812 -16628 42868
rect -16572 42812 -16468 42868
rect -16412 42812 -16308 42868
rect -16252 42812 -16148 42868
rect -16092 42812 -15988 42868
rect -15932 42812 -15828 42868
rect -15772 42812 -15668 42868
rect -15612 42812 -15508 42868
rect -15452 42812 -15348 42868
rect -15292 42812 -15188 42868
rect -15132 42812 -15028 42868
rect -14972 42812 -14868 42868
rect -14812 42812 -14708 42868
rect -14652 42812 -14548 42868
rect -14492 42812 -14388 42868
rect -14332 42812 -14228 42868
rect -14172 42812 -14068 42868
rect -14012 42812 -13908 42868
rect -13852 42812 -13748 42868
rect -13692 42812 -13588 42868
rect -13532 42812 -13428 42868
rect -13372 42812 -13268 42868
rect -13212 42812 -13108 42868
rect -13052 42812 -12948 42868
rect -12892 42812 -12788 42868
rect -12732 42812 -12628 42868
rect -12572 42812 -12468 42868
rect -12412 42812 -12308 42868
rect -12252 42812 -12148 42868
rect -12092 42812 -11828 42868
rect -11772 42812 -11508 42868
rect -11452 42812 -11348 42868
rect -11292 42812 -11188 42868
rect -11132 42812 -11028 42868
rect -10972 42812 -10868 42868
rect -10812 42812 -10708 42868
rect -10652 42812 -10548 42868
rect -10492 42812 -10388 42868
rect -10332 42812 -10228 42868
rect -10172 42812 -10068 42868
rect -10012 42812 -9908 42868
rect -9852 42812 -9748 42868
rect -9692 42812 -9588 42868
rect -9532 42812 -9428 42868
rect -9372 42812 -9268 42868
rect -9212 42812 -9108 42868
rect -9052 42812 -8948 42868
rect -8892 42812 -8788 42868
rect -8732 42812 -8628 42868
rect -8572 42812 -8468 42868
rect -8412 42812 -8308 42868
rect -8252 42812 -8148 42868
rect -8092 42812 -7988 42868
rect -7932 42812 -7828 42868
rect -7772 42812 -7668 42868
rect -7612 42812 -7508 42868
rect -7452 42812 -7348 42868
rect -7292 42812 -7188 42868
rect -7132 42812 -7028 42868
rect -6972 42812 -6868 42868
rect -6812 42812 -6708 42868
rect -6652 42812 -6548 42868
rect -6492 42812 -6388 42868
rect -6332 42812 -6228 42868
rect -6172 42812 -6068 42868
rect -6012 42812 -5908 42868
rect -5852 42812 -5748 42868
rect -5692 42812 -5588 42868
rect -5532 42812 -5428 42868
rect -5372 42812 -5268 42868
rect -5212 42812 -5108 42868
rect -5052 42812 -4948 42868
rect -4892 42812 -4788 42868
rect -4732 42812 -4628 42868
rect -4572 42812 -4468 42868
rect -4412 42812 -4308 42868
rect -4252 42812 -4148 42868
rect -4092 42812 -3988 42868
rect -3932 42812 -3668 42868
rect -3612 42812 -3508 42868
rect -3452 42812 -3348 42868
rect -3292 42812 -3188 42868
rect -3132 42812 -3028 42868
rect -2972 42812 -2708 42868
rect -2652 42812 -2548 42868
rect -2492 42812 -2388 42868
rect -2332 42812 -2228 42868
rect -2172 42812 -2068 42868
rect -2012 42812 -1748 42868
rect -1692 42812 -1428 42868
rect -1372 42812 -1108 42868
rect -1052 42812 -1040 42868
rect -31040 42800 -1040 42812
rect -31040 42708 -30320 42720
rect -31040 42652 -31028 42708
rect -30972 42652 -30708 42708
rect -30652 42652 -30388 42708
rect -30332 42652 -30320 42708
rect -31040 42640 -30320 42652
rect -30240 42708 -2800 42720
rect -30240 42652 -30228 42708
rect -30172 42652 -11988 42708
rect -11932 42652 -2868 42708
rect -2812 42652 -2800 42708
rect -30240 42640 -2800 42652
rect -2720 42640 -2640 42720
rect -2560 42640 -2480 42720
rect -2400 42640 -2320 42720
rect -2240 42640 -2160 42720
rect -2080 42640 -2000 42720
rect -1760 42640 -1680 42720
rect -1440 42640 -1360 42720
rect -1120 42640 -1040 42720
rect -31040 42548 -1040 42560
rect -31040 42492 -31028 42548
rect -30972 42492 -30708 42548
rect -30652 42492 -30388 42548
rect -30332 42492 -30068 42548
rect -30012 42492 -29908 42548
rect -29852 42492 -29748 42548
rect -29692 42492 -29588 42548
rect -29532 42492 -29428 42548
rect -29372 42492 -29268 42548
rect -29212 42492 -29108 42548
rect -29052 42492 -28948 42548
rect -28892 42492 -28788 42548
rect -28732 42492 -28628 42548
rect -28572 42492 -28468 42548
rect -28412 42492 -28308 42548
rect -28252 42492 -28148 42548
rect -28092 42492 -27988 42548
rect -27932 42492 -27828 42548
rect -27772 42492 -27668 42548
rect -27612 42492 -27508 42548
rect -27452 42492 -27348 42548
rect -27292 42492 -27188 42548
rect -27132 42492 -27028 42548
rect -26972 42492 -26868 42548
rect -26812 42492 -26708 42548
rect -26652 42492 -26548 42548
rect -26492 42492 -26388 42548
rect -26332 42492 -26228 42548
rect -26172 42492 -26068 42548
rect -26012 42492 -25908 42548
rect -25852 42492 -25748 42548
rect -25692 42492 -25588 42548
rect -25532 42492 -25428 42548
rect -25372 42492 -25268 42548
rect -25212 42492 -25108 42548
rect -25052 42492 -24948 42548
rect -24892 42492 -24788 42548
rect -24732 42492 -24628 42548
rect -24572 42492 -24468 42548
rect -24412 42492 -24308 42548
rect -24252 42492 -24148 42548
rect -24092 42492 -23988 42548
rect -23932 42492 -23828 42548
rect -23772 42492 -23668 42548
rect -23612 42492 -23508 42548
rect -23452 42492 -23348 42548
rect -23292 42492 -23188 42548
rect -23132 42492 -23028 42548
rect -22972 42492 -22868 42548
rect -22812 42492 -22708 42548
rect -22652 42492 -22548 42548
rect -22492 42492 -22388 42548
rect -22332 42492 -22228 42548
rect -22172 42492 -22068 42548
rect -22012 42492 -21908 42548
rect -21852 42492 -21748 42548
rect -21692 42492 -21588 42548
rect -21532 42492 -21428 42548
rect -21372 42492 -21268 42548
rect -21212 42492 -21108 42548
rect -21052 42492 -20948 42548
rect -20892 42492 -20788 42548
rect -20732 42492 -20628 42548
rect -20572 42492 -20468 42548
rect -20412 42492 -20308 42548
rect -20252 42492 -20148 42548
rect -20092 42492 -19988 42548
rect -19932 42492 -19828 42548
rect -19772 42492 -19668 42548
rect -19612 42492 -19508 42548
rect -19452 42492 -19348 42548
rect -19292 42492 -19188 42548
rect -19132 42492 -19028 42548
rect -18972 42492 -18868 42548
rect -18812 42492 -18708 42548
rect -18652 42492 -18548 42548
rect -18492 42492 -18388 42548
rect -18332 42492 -18228 42548
rect -18172 42492 -18068 42548
rect -18012 42492 -17908 42548
rect -17852 42492 -17748 42548
rect -17692 42492 -17588 42548
rect -17532 42492 -17428 42548
rect -17372 42492 -17268 42548
rect -17212 42492 -17108 42548
rect -17052 42492 -16948 42548
rect -16892 42492 -16788 42548
rect -16732 42492 -16628 42548
rect -16572 42492 -16468 42548
rect -16412 42492 -16308 42548
rect -16252 42492 -16148 42548
rect -16092 42492 -15988 42548
rect -15932 42492 -15828 42548
rect -15772 42492 -15668 42548
rect -15612 42492 -15508 42548
rect -15452 42492 -15348 42548
rect -15292 42492 -15188 42548
rect -15132 42492 -15028 42548
rect -14972 42492 -14868 42548
rect -14812 42492 -14708 42548
rect -14652 42492 -14548 42548
rect -14492 42492 -14388 42548
rect -14332 42492 -14228 42548
rect -14172 42492 -14068 42548
rect -14012 42492 -13908 42548
rect -13852 42492 -13748 42548
rect -13692 42492 -13588 42548
rect -13532 42492 -13428 42548
rect -13372 42492 -13268 42548
rect -13212 42492 -13108 42548
rect -13052 42492 -12948 42548
rect -12892 42492 -12788 42548
rect -12732 42492 -12628 42548
rect -12572 42492 -12468 42548
rect -12412 42492 -12308 42548
rect -12252 42492 -12148 42548
rect -12092 42492 -11828 42548
rect -11772 42492 -11508 42548
rect -11452 42492 -11348 42548
rect -11292 42492 -11188 42548
rect -11132 42492 -11028 42548
rect -10972 42492 -10868 42548
rect -10812 42492 -10708 42548
rect -10652 42492 -10548 42548
rect -10492 42492 -10388 42548
rect -10332 42492 -10228 42548
rect -10172 42492 -10068 42548
rect -10012 42492 -9908 42548
rect -9852 42492 -9748 42548
rect -9692 42492 -9588 42548
rect -9532 42492 -9428 42548
rect -9372 42492 -9268 42548
rect -9212 42492 -9108 42548
rect -9052 42492 -8948 42548
rect -8892 42492 -8788 42548
rect -8732 42492 -8628 42548
rect -8572 42492 -8468 42548
rect -8412 42492 -8308 42548
rect -8252 42492 -8148 42548
rect -8092 42492 -7988 42548
rect -7932 42492 -7828 42548
rect -7772 42492 -7668 42548
rect -7612 42492 -7508 42548
rect -7452 42492 -7348 42548
rect -7292 42492 -7188 42548
rect -7132 42492 -7028 42548
rect -6972 42492 -6868 42548
rect -6812 42492 -6708 42548
rect -6652 42492 -6548 42548
rect -6492 42492 -6388 42548
rect -6332 42492 -6228 42548
rect -6172 42492 -6068 42548
rect -6012 42492 -5908 42548
rect -5852 42492 -5748 42548
rect -5692 42492 -5588 42548
rect -5532 42492 -5428 42548
rect -5372 42492 -5268 42548
rect -5212 42492 -5108 42548
rect -5052 42492 -4948 42548
rect -4892 42492 -4788 42548
rect -4732 42492 -4628 42548
rect -4572 42492 -4468 42548
rect -4412 42492 -4308 42548
rect -4252 42492 -4148 42548
rect -4092 42492 -3988 42548
rect -3932 42492 -3668 42548
rect -3612 42492 -3508 42548
rect -3452 42492 -3348 42548
rect -3292 42492 -3188 42548
rect -3132 42492 -3028 42548
rect -2972 42492 -2708 42548
rect -2652 42492 -2548 42548
rect -2492 42492 -2388 42548
rect -2332 42492 -2228 42548
rect -2172 42492 -2068 42548
rect -2012 42492 -1748 42548
rect -1692 42492 -1428 42548
rect -1372 42492 -1108 42548
rect -1052 42492 -1040 42548
rect -31040 42480 -1040 42492
rect -31040 42388 -30640 42400
rect -31040 42332 -31028 42388
rect -30972 42332 -30708 42388
rect -30652 42332 -30640 42388
rect -31040 42320 -30640 42332
rect -30560 42388 -3120 42400
rect -30560 42332 -30548 42388
rect -30492 42332 -11668 42388
rect -11612 42332 -3188 42388
rect -3132 42332 -3120 42388
rect -30560 42320 -3120 42332
rect -3040 42320 -2960 42400
rect -2720 42320 -2640 42400
rect -2560 42320 -2480 42400
rect -2400 42320 -2320 42400
rect -2240 42320 -2160 42400
rect -2080 42320 -2000 42400
rect -1760 42320 -1680 42400
rect -1440 42320 -1360 42400
rect -1120 42320 -1040 42400
rect -31040 42228 -1040 42240
rect -31040 42172 -31028 42228
rect -30972 42172 -30708 42228
rect -30652 42172 -30388 42228
rect -30332 42172 -30068 42228
rect -30012 42172 -29908 42228
rect -29852 42172 -29748 42228
rect -29692 42172 -29588 42228
rect -29532 42172 -29428 42228
rect -29372 42172 -29268 42228
rect -29212 42172 -29108 42228
rect -29052 42172 -28948 42228
rect -28892 42172 -28788 42228
rect -28732 42172 -28628 42228
rect -28572 42172 -28468 42228
rect -28412 42172 -28308 42228
rect -28252 42172 -28148 42228
rect -28092 42172 -27988 42228
rect -27932 42172 -27828 42228
rect -27772 42172 -27668 42228
rect -27612 42172 -27508 42228
rect -27452 42172 -27348 42228
rect -27292 42172 -27188 42228
rect -27132 42172 -27028 42228
rect -26972 42172 -26868 42228
rect -26812 42172 -26708 42228
rect -26652 42172 -26548 42228
rect -26492 42172 -26388 42228
rect -26332 42172 -26228 42228
rect -26172 42172 -26068 42228
rect -26012 42172 -25908 42228
rect -25852 42172 -25748 42228
rect -25692 42172 -25588 42228
rect -25532 42172 -25428 42228
rect -25372 42172 -25268 42228
rect -25212 42172 -25108 42228
rect -25052 42172 -24948 42228
rect -24892 42172 -24788 42228
rect -24732 42172 -24628 42228
rect -24572 42172 -24468 42228
rect -24412 42172 -24308 42228
rect -24252 42172 -24148 42228
rect -24092 42172 -23988 42228
rect -23932 42172 -23828 42228
rect -23772 42172 -23668 42228
rect -23612 42172 -23508 42228
rect -23452 42172 -23348 42228
rect -23292 42172 -23188 42228
rect -23132 42172 -23028 42228
rect -22972 42172 -22868 42228
rect -22812 42172 -22708 42228
rect -22652 42172 -22548 42228
rect -22492 42172 -22388 42228
rect -22332 42172 -22228 42228
rect -22172 42172 -22068 42228
rect -22012 42172 -21908 42228
rect -21852 42172 -21748 42228
rect -21692 42172 -21588 42228
rect -21532 42172 -21428 42228
rect -21372 42172 -21268 42228
rect -21212 42172 -21108 42228
rect -21052 42172 -20948 42228
rect -20892 42172 -20788 42228
rect -20732 42172 -20628 42228
rect -20572 42172 -20468 42228
rect -20412 42172 -20308 42228
rect -20252 42172 -20148 42228
rect -20092 42172 -19988 42228
rect -19932 42172 -19828 42228
rect -19772 42172 -19668 42228
rect -19612 42172 -19508 42228
rect -19452 42172 -19348 42228
rect -19292 42172 -19188 42228
rect -19132 42172 -19028 42228
rect -18972 42172 -18868 42228
rect -18812 42172 -18708 42228
rect -18652 42172 -18548 42228
rect -18492 42172 -18388 42228
rect -18332 42172 -18228 42228
rect -18172 42172 -18068 42228
rect -18012 42172 -17908 42228
rect -17852 42172 -17748 42228
rect -17692 42172 -17588 42228
rect -17532 42172 -17428 42228
rect -17372 42172 -17268 42228
rect -17212 42172 -17108 42228
rect -17052 42172 -16948 42228
rect -16892 42172 -16788 42228
rect -16732 42172 -16628 42228
rect -16572 42172 -16468 42228
rect -16412 42172 -16308 42228
rect -16252 42172 -16148 42228
rect -16092 42172 -15988 42228
rect -15932 42172 -15828 42228
rect -15772 42172 -15668 42228
rect -15612 42172 -15508 42228
rect -15452 42172 -15348 42228
rect -15292 42172 -15188 42228
rect -15132 42172 -15028 42228
rect -14972 42172 -14868 42228
rect -14812 42172 -14708 42228
rect -14652 42172 -14548 42228
rect -14492 42172 -14388 42228
rect -14332 42172 -14228 42228
rect -14172 42172 -14068 42228
rect -14012 42172 -13908 42228
rect -13852 42172 -13748 42228
rect -13692 42172 -13588 42228
rect -13532 42172 -13428 42228
rect -13372 42172 -13268 42228
rect -13212 42172 -13108 42228
rect -13052 42172 -12948 42228
rect -12892 42172 -12788 42228
rect -12732 42172 -12628 42228
rect -12572 42172 -12468 42228
rect -12412 42172 -12308 42228
rect -12252 42172 -12148 42228
rect -12092 42172 -11828 42228
rect -11772 42172 -11508 42228
rect -11452 42172 -11348 42228
rect -11292 42172 -11188 42228
rect -11132 42172 -11028 42228
rect -10972 42172 -10868 42228
rect -10812 42172 -10708 42228
rect -10652 42172 -10548 42228
rect -10492 42172 -10388 42228
rect -10332 42172 -10228 42228
rect -10172 42172 -10068 42228
rect -10012 42172 -9908 42228
rect -9852 42172 -9748 42228
rect -9692 42172 -9588 42228
rect -9532 42172 -9428 42228
rect -9372 42172 -9268 42228
rect -9212 42172 -9108 42228
rect -9052 42172 -8948 42228
rect -8892 42172 -8788 42228
rect -8732 42172 -8628 42228
rect -8572 42172 -8468 42228
rect -8412 42172 -8308 42228
rect -8252 42172 -8148 42228
rect -8092 42172 -7988 42228
rect -7932 42172 -7828 42228
rect -7772 42172 -7668 42228
rect -7612 42172 -7508 42228
rect -7452 42172 -7348 42228
rect -7292 42172 -7188 42228
rect -7132 42172 -7028 42228
rect -6972 42172 -6868 42228
rect -6812 42172 -6708 42228
rect -6652 42172 -6548 42228
rect -6492 42172 -6388 42228
rect -6332 42172 -6228 42228
rect -6172 42172 -6068 42228
rect -6012 42172 -5908 42228
rect -5852 42172 -5748 42228
rect -5692 42172 -5588 42228
rect -5532 42172 -5428 42228
rect -5372 42172 -5268 42228
rect -5212 42172 -5108 42228
rect -5052 42172 -4948 42228
rect -4892 42172 -4788 42228
rect -4732 42172 -4628 42228
rect -4572 42172 -4468 42228
rect -4412 42172 -4308 42228
rect -4252 42172 -4148 42228
rect -4092 42172 -3988 42228
rect -3932 42172 -3668 42228
rect -3612 42172 -3508 42228
rect -3452 42172 -3348 42228
rect -3292 42172 -3028 42228
rect -2972 42172 -2708 42228
rect -2652 42172 -2548 42228
rect -2492 42172 -2388 42228
rect -2332 42172 -2228 42228
rect -2172 42172 -2068 42228
rect -2012 42172 -1748 42228
rect -1692 42172 -1428 42228
rect -1372 42172 -1108 42228
rect -1052 42172 -1040 42228
rect -31040 42160 -1040 42172
rect -31040 42068 -30320 42080
rect -31040 42012 -31028 42068
rect -30972 42012 -30708 42068
rect -30652 42012 -30388 42068
rect -30332 42012 -30320 42068
rect -31040 42000 -30320 42012
rect -30240 42068 -1200 42080
rect -30240 42012 -30228 42068
rect -30172 42012 -1268 42068
rect -1212 42012 -1200 42068
rect -30240 42000 -1200 42012
rect -1120 42000 -1040 42080
rect -31040 41908 -1040 41920
rect -31040 41852 -31028 41908
rect -30972 41852 -30708 41908
rect -30652 41852 -30388 41908
rect -30332 41852 -30068 41908
rect -30012 41852 -29908 41908
rect -29852 41852 -29748 41908
rect -29692 41852 -29588 41908
rect -29532 41852 -29428 41908
rect -29372 41852 -29268 41908
rect -29212 41852 -29108 41908
rect -29052 41852 -28948 41908
rect -28892 41852 -28788 41908
rect -28732 41852 -28628 41908
rect -28572 41852 -28468 41908
rect -28412 41852 -28308 41908
rect -28252 41852 -28148 41908
rect -28092 41852 -27988 41908
rect -27932 41852 -27828 41908
rect -27772 41852 -27668 41908
rect -27612 41852 -27508 41908
rect -27452 41852 -27348 41908
rect -27292 41852 -27188 41908
rect -27132 41852 -27028 41908
rect -26972 41852 -26868 41908
rect -26812 41852 -26708 41908
rect -26652 41852 -26548 41908
rect -26492 41852 -26388 41908
rect -26332 41852 -26228 41908
rect -26172 41852 -26068 41908
rect -26012 41852 -25908 41908
rect -25852 41852 -25748 41908
rect -25692 41852 -25588 41908
rect -25532 41852 -25428 41908
rect -25372 41852 -25268 41908
rect -25212 41852 -25108 41908
rect -25052 41852 -24948 41908
rect -24892 41852 -24788 41908
rect -24732 41852 -24628 41908
rect -24572 41852 -24468 41908
rect -24412 41852 -24308 41908
rect -24252 41852 -24148 41908
rect -24092 41852 -23988 41908
rect -23932 41852 -23828 41908
rect -23772 41852 -23668 41908
rect -23612 41852 -23508 41908
rect -23452 41852 -23348 41908
rect -23292 41852 -23188 41908
rect -23132 41852 -23028 41908
rect -22972 41852 -22868 41908
rect -22812 41852 -22708 41908
rect -22652 41852 -22548 41908
rect -22492 41852 -22388 41908
rect -22332 41852 -22228 41908
rect -22172 41852 -22068 41908
rect -22012 41852 -21908 41908
rect -21852 41852 -21748 41908
rect -21692 41852 -21588 41908
rect -21532 41852 -21428 41908
rect -21372 41852 -21268 41908
rect -21212 41852 -21108 41908
rect -21052 41852 -20948 41908
rect -20892 41852 -20788 41908
rect -20732 41852 -20628 41908
rect -20572 41852 -20468 41908
rect -20412 41852 -20308 41908
rect -20252 41852 -20148 41908
rect -20092 41852 -19988 41908
rect -19932 41852 -19828 41908
rect -19772 41852 -19668 41908
rect -19612 41852 -19508 41908
rect -19452 41852 -19348 41908
rect -19292 41852 -19188 41908
rect -19132 41852 -19028 41908
rect -18972 41852 -18868 41908
rect -18812 41852 -18708 41908
rect -18652 41852 -18548 41908
rect -18492 41852 -18388 41908
rect -18332 41852 -18228 41908
rect -18172 41852 -18068 41908
rect -18012 41852 -17908 41908
rect -17852 41852 -17748 41908
rect -17692 41852 -17588 41908
rect -17532 41852 -17428 41908
rect -17372 41852 -17268 41908
rect -17212 41852 -17108 41908
rect -17052 41852 -16948 41908
rect -16892 41852 -16788 41908
rect -16732 41852 -16628 41908
rect -16572 41852 -16468 41908
rect -16412 41852 -16308 41908
rect -16252 41852 -16148 41908
rect -16092 41852 -15988 41908
rect -15932 41852 -15828 41908
rect -15772 41852 -15668 41908
rect -15612 41852 -15508 41908
rect -15452 41852 -15348 41908
rect -15292 41852 -15188 41908
rect -15132 41852 -15028 41908
rect -14972 41852 -14868 41908
rect -14812 41852 -14708 41908
rect -14652 41852 -14548 41908
rect -14492 41852 -14388 41908
rect -14332 41852 -14228 41908
rect -14172 41852 -14068 41908
rect -14012 41852 -13908 41908
rect -13852 41852 -13748 41908
rect -13692 41852 -13588 41908
rect -13532 41852 -13428 41908
rect -13372 41852 -13268 41908
rect -13212 41852 -13108 41908
rect -13052 41852 -12948 41908
rect -12892 41852 -12788 41908
rect -12732 41852 -12628 41908
rect -12572 41852 -12468 41908
rect -12412 41852 -12308 41908
rect -12252 41852 -12148 41908
rect -12092 41852 -11828 41908
rect -11772 41852 -11508 41908
rect -11452 41852 -11348 41908
rect -11292 41852 -11188 41908
rect -11132 41852 -11028 41908
rect -10972 41852 -10868 41908
rect -10812 41852 -10708 41908
rect -10652 41852 -10548 41908
rect -10492 41852 -10388 41908
rect -10332 41852 -10228 41908
rect -10172 41852 -10068 41908
rect -10012 41852 -9908 41908
rect -9852 41852 -9748 41908
rect -9692 41852 -9588 41908
rect -9532 41852 -9428 41908
rect -9372 41852 -9268 41908
rect -9212 41852 -9108 41908
rect -9052 41852 -8948 41908
rect -8892 41852 -8788 41908
rect -8732 41852 -8628 41908
rect -8572 41852 -8468 41908
rect -8412 41852 -8308 41908
rect -8252 41852 -8148 41908
rect -8092 41852 -7988 41908
rect -7932 41852 -7828 41908
rect -7772 41852 -7668 41908
rect -7612 41852 -7508 41908
rect -7452 41852 -7348 41908
rect -7292 41852 -7188 41908
rect -7132 41852 -7028 41908
rect -6972 41852 -6868 41908
rect -6812 41852 -6708 41908
rect -6652 41852 -6548 41908
rect -6492 41852 -6388 41908
rect -6332 41852 -6228 41908
rect -6172 41852 -6068 41908
rect -6012 41852 -5908 41908
rect -5852 41852 -5748 41908
rect -5692 41852 -5588 41908
rect -5532 41852 -5428 41908
rect -5372 41852 -5268 41908
rect -5212 41852 -5108 41908
rect -5052 41852 -4948 41908
rect -4892 41852 -4788 41908
rect -4732 41852 -4628 41908
rect -4572 41852 -4468 41908
rect -4412 41852 -4308 41908
rect -4252 41852 -4148 41908
rect -4092 41852 -3988 41908
rect -3932 41852 -3668 41908
rect -3612 41852 -3508 41908
rect -3452 41852 -3348 41908
rect -3292 41852 -3028 41908
rect -2972 41852 -2708 41908
rect -2652 41852 -2548 41908
rect -2492 41852 -2388 41908
rect -2332 41852 -2228 41908
rect -2172 41852 -2068 41908
rect -2012 41852 -1748 41908
rect -1692 41852 -1428 41908
rect -1372 41852 -1108 41908
rect -1052 41852 -1040 41908
rect -31040 41840 -1040 41852
rect -31040 41748 -30000 41760
rect -31040 41692 -31028 41748
rect -30972 41692 -30708 41748
rect -30652 41692 -30388 41748
rect -30332 41692 -30068 41748
rect -30012 41692 -30000 41748
rect -31040 41680 -30000 41692
rect -12160 41748 -11440 41760
rect -12160 41692 -12148 41748
rect -12092 41692 -11828 41748
rect -11772 41692 -11508 41748
rect -11452 41692 -11440 41748
rect -12160 41680 -11440 41692
rect -3360 41748 -1040 41760
rect -3360 41692 -3348 41748
rect -3292 41692 -3028 41748
rect -2972 41692 -2708 41748
rect -2652 41692 -2388 41748
rect -2332 41692 -2068 41748
rect -2012 41692 -1748 41748
rect -1692 41692 -1428 41748
rect -1372 41692 -1108 41748
rect -1052 41692 -1040 41748
rect -3360 41680 -1040 41692
rect -31040 41588 -30000 41600
rect -31040 41532 -31028 41588
rect -30972 41532 -30708 41588
rect -30652 41532 -30388 41588
rect -30332 41532 -30068 41588
rect -30012 41532 -30000 41588
rect -31040 41520 -30000 41532
rect -12160 41588 -11440 41600
rect -12160 41532 -12148 41588
rect -12092 41532 -11828 41588
rect -11772 41532 -11508 41588
rect -11452 41532 -11440 41588
rect -12160 41520 -11440 41532
rect -3360 41588 -1040 41600
rect -3360 41532 -3348 41588
rect -3292 41532 -3028 41588
rect -2972 41532 -2708 41588
rect -2652 41532 -2388 41588
rect -2332 41532 -2068 41588
rect -2012 41532 -1748 41588
rect -1692 41532 -1428 41588
rect -1372 41532 -1108 41588
rect -1052 41532 -1040 41588
rect -3360 41520 -1040 41532
rect -33120 41348 -960 41360
rect -33120 41292 -33108 41348
rect -33052 41292 -32948 41348
rect -32892 41292 -32788 41348
rect -32732 41292 -32628 41348
rect -32572 41292 -32468 41348
rect -32412 41292 -32308 41348
rect -32252 41292 -32148 41348
rect -32092 41292 -31988 41348
rect -31932 41292 -31828 41348
rect -31772 41292 -31668 41348
rect -31612 41292 -31508 41348
rect -31452 41292 -31348 41348
rect -31292 41292 -31188 41348
rect -31132 41292 -29908 41348
rect -29852 41292 -29748 41348
rect -29692 41292 -29588 41348
rect -29532 41292 -29428 41348
rect -29372 41292 -29268 41348
rect -29212 41292 -29108 41348
rect -29052 41292 -28948 41348
rect -28892 41292 -28788 41348
rect -28732 41292 -28628 41348
rect -28572 41292 -28468 41348
rect -28412 41292 -28308 41348
rect -28252 41292 -28148 41348
rect -28092 41292 -27988 41348
rect -27932 41292 -27828 41348
rect -27772 41292 -27668 41348
rect -27612 41292 -27508 41348
rect -27452 41292 -27348 41348
rect -27292 41292 -27188 41348
rect -27132 41292 -27028 41348
rect -26972 41292 -26868 41348
rect -26812 41292 -26708 41348
rect -26652 41292 -26548 41348
rect -26492 41292 -26388 41348
rect -26332 41292 -26228 41348
rect -26172 41292 -26068 41348
rect -26012 41292 -25908 41348
rect -25852 41292 -25748 41348
rect -25692 41292 -25588 41348
rect -25532 41292 -25428 41348
rect -25372 41292 -25268 41348
rect -25212 41292 -25108 41348
rect -25052 41292 -24948 41348
rect -24892 41292 -24788 41348
rect -24732 41292 -24628 41348
rect -24572 41292 -24468 41348
rect -24412 41292 -24308 41348
rect -24252 41292 -24148 41348
rect -24092 41292 -23988 41348
rect -23932 41292 -23828 41348
rect -23772 41292 -23668 41348
rect -23612 41292 -23508 41348
rect -23452 41292 -23348 41348
rect -23292 41292 -23188 41348
rect -23132 41292 -23028 41348
rect -22972 41292 -22868 41348
rect -22812 41292 -22708 41348
rect -22652 41292 -22548 41348
rect -22492 41292 -22388 41348
rect -22332 41292 -22228 41348
rect -22172 41292 -22068 41348
rect -22012 41292 -21908 41348
rect -21852 41292 -21748 41348
rect -21692 41292 -21588 41348
rect -21532 41292 -21428 41348
rect -21372 41292 -21268 41348
rect -21212 41292 -21108 41348
rect -21052 41292 -20948 41348
rect -20892 41292 -20788 41348
rect -20732 41292 -20628 41348
rect -20572 41292 -20468 41348
rect -20412 41292 -20308 41348
rect -20252 41292 -20148 41348
rect -20092 41292 -19988 41348
rect -19932 41292 -19828 41348
rect -19772 41292 -19668 41348
rect -19612 41292 -19508 41348
rect -19452 41292 -19348 41348
rect -19292 41292 -19188 41348
rect -19132 41292 -19028 41348
rect -18972 41292 -18868 41348
rect -18812 41292 -18708 41348
rect -18652 41292 -18548 41348
rect -18492 41292 -18388 41348
rect -18332 41292 -18228 41348
rect -18172 41292 -18068 41348
rect -18012 41292 -17908 41348
rect -17852 41292 -17748 41348
rect -17692 41292 -17588 41348
rect -17532 41292 -17428 41348
rect -17372 41292 -17268 41348
rect -17212 41292 -17108 41348
rect -17052 41292 -16948 41348
rect -16892 41292 -16788 41348
rect -16732 41292 -16628 41348
rect -16572 41292 -16468 41348
rect -16412 41292 -16308 41348
rect -16252 41292 -16148 41348
rect -16092 41292 -15988 41348
rect -15932 41292 -15828 41348
rect -15772 41292 -15668 41348
rect -15612 41292 -15508 41348
rect -15452 41292 -15348 41348
rect -15292 41292 -15188 41348
rect -15132 41292 -15028 41348
rect -14972 41292 -14868 41348
rect -14812 41292 -14708 41348
rect -14652 41292 -14548 41348
rect -14492 41292 -14388 41348
rect -14332 41292 -14228 41348
rect -14172 41292 -14068 41348
rect -14012 41292 -13908 41348
rect -13852 41292 -13748 41348
rect -13692 41292 -13588 41348
rect -13532 41292 -13428 41348
rect -13372 41292 -13268 41348
rect -13212 41292 -13108 41348
rect -13052 41292 -12948 41348
rect -12892 41292 -12788 41348
rect -12732 41292 -12628 41348
rect -12572 41292 -12468 41348
rect -12412 41292 -12308 41348
rect -12252 41292 -11348 41348
rect -11292 41292 -11188 41348
rect -11132 41292 -11028 41348
rect -10972 41292 -10868 41348
rect -10812 41292 -10708 41348
rect -10652 41292 -10548 41348
rect -10492 41292 -10388 41348
rect -10332 41292 -10228 41348
rect -10172 41292 -10068 41348
rect -10012 41292 -9908 41348
rect -9852 41292 -9748 41348
rect -9692 41292 -9588 41348
rect -9532 41292 -9428 41348
rect -9372 41292 -9268 41348
rect -9212 41292 -9108 41348
rect -9052 41292 -8948 41348
rect -8892 41292 -8788 41348
rect -8732 41292 -8628 41348
rect -8572 41292 -8468 41348
rect -8412 41292 -8308 41348
rect -8252 41292 -8148 41348
rect -8092 41292 -7988 41348
rect -7932 41292 -7828 41348
rect -7772 41292 -7668 41348
rect -7612 41292 -7508 41348
rect -7452 41292 -7348 41348
rect -7292 41292 -7188 41348
rect -7132 41292 -7028 41348
rect -6972 41292 -6868 41348
rect -6812 41292 -6708 41348
rect -6652 41292 -6548 41348
rect -6492 41292 -6388 41348
rect -6332 41292 -6228 41348
rect -6172 41292 -6068 41348
rect -6012 41292 -5908 41348
rect -5852 41292 -5748 41348
rect -5692 41292 -5588 41348
rect -5532 41292 -5428 41348
rect -5372 41292 -5268 41348
rect -5212 41292 -5108 41348
rect -5052 41292 -4948 41348
rect -4892 41292 -4788 41348
rect -4732 41292 -4628 41348
rect -4572 41292 -4468 41348
rect -4412 41292 -4308 41348
rect -4252 41292 -4148 41348
rect -4092 41292 -3988 41348
rect -3932 41292 -3828 41348
rect -3772 41292 -3668 41348
rect -3612 41292 -3508 41348
rect -3452 41292 -960 41348
rect -33120 41280 -960 41292
rect 40960 41348 43200 41360
rect 40960 41292 41052 41348
rect 41108 41292 41212 41348
rect 41268 41292 41372 41348
rect 41428 41292 41532 41348
rect 41588 41292 41692 41348
rect 41748 41292 41852 41348
rect 41908 41292 42012 41348
rect 42068 41292 42172 41348
rect 42228 41292 42332 41348
rect 42388 41292 42492 41348
rect 42548 41292 42652 41348
rect 42708 41292 42812 41348
rect 42868 41292 42972 41348
rect 43028 41292 43132 41348
rect 43188 41292 43200 41348
rect 40960 41280 43200 41292
rect -33280 41120 43360 41200
rect -33120 41028 -960 41040
rect -33120 40972 -33108 41028
rect -33052 40972 -32948 41028
rect -32892 40972 -32788 41028
rect -32732 40972 -32628 41028
rect -32572 40972 -32468 41028
rect -32412 40972 -32308 41028
rect -32252 40972 -32148 41028
rect -32092 40972 -31988 41028
rect -31932 40972 -31828 41028
rect -31772 40972 -31668 41028
rect -31612 40972 -31508 41028
rect -31452 40972 -31348 41028
rect -31292 40972 -31188 41028
rect -31132 40972 -29908 41028
rect -29852 40972 -29748 41028
rect -29692 40972 -29588 41028
rect -29532 40972 -29428 41028
rect -29372 40972 -29268 41028
rect -29212 40972 -29108 41028
rect -29052 40972 -28948 41028
rect -28892 40972 -28788 41028
rect -28732 40972 -28628 41028
rect -28572 40972 -28468 41028
rect -28412 40972 -28308 41028
rect -28252 40972 -28148 41028
rect -28092 40972 -27988 41028
rect -27932 40972 -27828 41028
rect -27772 40972 -27668 41028
rect -27612 40972 -27508 41028
rect -27452 40972 -27348 41028
rect -27292 40972 -27188 41028
rect -27132 40972 -27028 41028
rect -26972 40972 -26868 41028
rect -26812 40972 -26708 41028
rect -26652 40972 -26548 41028
rect -26492 40972 -26388 41028
rect -26332 40972 -26228 41028
rect -26172 40972 -26068 41028
rect -26012 40972 -25908 41028
rect -25852 40972 -25748 41028
rect -25692 40972 -25588 41028
rect -25532 40972 -25428 41028
rect -25372 40972 -25268 41028
rect -25212 40972 -25108 41028
rect -25052 40972 -24948 41028
rect -24892 40972 -24788 41028
rect -24732 40972 -24628 41028
rect -24572 40972 -24468 41028
rect -24412 40972 -24308 41028
rect -24252 40972 -24148 41028
rect -24092 40972 -23988 41028
rect -23932 40972 -23828 41028
rect -23772 40972 -23668 41028
rect -23612 40972 -23508 41028
rect -23452 40972 -23348 41028
rect -23292 40972 -23188 41028
rect -23132 40972 -23028 41028
rect -22972 40972 -22868 41028
rect -22812 40972 -22708 41028
rect -22652 40972 -22548 41028
rect -22492 40972 -22388 41028
rect -22332 40972 -22228 41028
rect -22172 40972 -22068 41028
rect -22012 40972 -21908 41028
rect -21852 40972 -21748 41028
rect -21692 40972 -21588 41028
rect -21532 40972 -21428 41028
rect -21372 40972 -21268 41028
rect -21212 40972 -21108 41028
rect -21052 40972 -20948 41028
rect -20892 40972 -20788 41028
rect -20732 40972 -20628 41028
rect -20572 40972 -20468 41028
rect -20412 40972 -20308 41028
rect -20252 40972 -20148 41028
rect -20092 40972 -19988 41028
rect -19932 40972 -19828 41028
rect -19772 40972 -19668 41028
rect -19612 40972 -19508 41028
rect -19452 40972 -19348 41028
rect -19292 40972 -19188 41028
rect -19132 40972 -19028 41028
rect -18972 40972 -18868 41028
rect -18812 40972 -18708 41028
rect -18652 40972 -18548 41028
rect -18492 40972 -18388 41028
rect -18332 40972 -18228 41028
rect -18172 40972 -18068 41028
rect -18012 40972 -17908 41028
rect -17852 40972 -17748 41028
rect -17692 40972 -17588 41028
rect -17532 40972 -17428 41028
rect -17372 40972 -17268 41028
rect -17212 40972 -17108 41028
rect -17052 40972 -16948 41028
rect -16892 40972 -16788 41028
rect -16732 40972 -16628 41028
rect -16572 40972 -16468 41028
rect -16412 40972 -16308 41028
rect -16252 40972 -16148 41028
rect -16092 40972 -15988 41028
rect -15932 40972 -15828 41028
rect -15772 40972 -15668 41028
rect -15612 40972 -15508 41028
rect -15452 40972 -15348 41028
rect -15292 40972 -15188 41028
rect -15132 40972 -15028 41028
rect -14972 40972 -14868 41028
rect -14812 40972 -14708 41028
rect -14652 40972 -14548 41028
rect -14492 40972 -14388 41028
rect -14332 40972 -14228 41028
rect -14172 40972 -14068 41028
rect -14012 40972 -13908 41028
rect -13852 40972 -13748 41028
rect -13692 40972 -13588 41028
rect -13532 40972 -13428 41028
rect -13372 40972 -13268 41028
rect -13212 40972 -13108 41028
rect -13052 40972 -12948 41028
rect -12892 40972 -12788 41028
rect -12732 40972 -12628 41028
rect -12572 40972 -12468 41028
rect -12412 40972 -12308 41028
rect -12252 40972 -11348 41028
rect -11292 40972 -11188 41028
rect -11132 40972 -11028 41028
rect -10972 40972 -10868 41028
rect -10812 40972 -10708 41028
rect -10652 40972 -10548 41028
rect -10492 40972 -10388 41028
rect -10332 40972 -10228 41028
rect -10172 40972 -10068 41028
rect -10012 40972 -9908 41028
rect -9852 40972 -9748 41028
rect -9692 40972 -9588 41028
rect -9532 40972 -9428 41028
rect -9372 40972 -9268 41028
rect -9212 40972 -9108 41028
rect -9052 40972 -8948 41028
rect -8892 40972 -8788 41028
rect -8732 40972 -8628 41028
rect -8572 40972 -8468 41028
rect -8412 40972 -8308 41028
rect -8252 40972 -8148 41028
rect -8092 40972 -7988 41028
rect -7932 40972 -7828 41028
rect -7772 40972 -7668 41028
rect -7612 40972 -7508 41028
rect -7452 40972 -7348 41028
rect -7292 40972 -7188 41028
rect -7132 40972 -7028 41028
rect -6972 40972 -6868 41028
rect -6812 40972 -6708 41028
rect -6652 40972 -6548 41028
rect -6492 40972 -6388 41028
rect -6332 40972 -6228 41028
rect -6172 40972 -6068 41028
rect -6012 40972 -5908 41028
rect -5852 40972 -5748 41028
rect -5692 40972 -5588 41028
rect -5532 40972 -5428 41028
rect -5372 40972 -5268 41028
rect -5212 40972 -5108 41028
rect -5052 40972 -4948 41028
rect -4892 40972 -4788 41028
rect -4732 40972 -4628 41028
rect -4572 40972 -4468 41028
rect -4412 40972 -4308 41028
rect -4252 40972 -4148 41028
rect -4092 40972 -3988 41028
rect -3932 40972 -3828 41028
rect -3772 40972 -3668 41028
rect -3612 40972 -3508 41028
rect -3452 40972 -960 41028
rect -33120 40960 -960 40972
rect 40960 41028 43200 41040
rect 40960 40972 41052 41028
rect 41108 40972 41212 41028
rect 41268 40972 41372 41028
rect 41428 40972 41532 41028
rect 41588 40972 41692 41028
rect 41748 40972 41852 41028
rect 41908 40972 42012 41028
rect 42068 40972 42172 41028
rect 42228 40972 42332 41028
rect 42388 40972 42492 41028
rect 42548 40972 42652 41028
rect 42708 40972 42812 41028
rect 42868 40972 42972 41028
rect 43028 40972 43132 41028
rect 43188 40972 43200 41028
rect 40960 40960 43200 40972
rect -12160 40868 -11440 40880
rect -12160 40812 -12148 40868
rect -12092 40812 -11828 40868
rect -11772 40812 -11508 40868
rect -11452 40812 -11440 40868
rect -12160 40800 -11440 40812
rect -3360 40868 -1040 40880
rect -3360 40812 -3348 40868
rect -3292 40812 -3028 40868
rect -2972 40812 -2708 40868
rect -2652 40812 -2388 40868
rect -2332 40812 -2068 40868
rect -2012 40812 -1748 40868
rect -1692 40812 -1428 40868
rect -1372 40812 -1108 40868
rect -1052 40812 -1040 40868
rect -3360 40800 -1040 40812
rect -31040 40788 -30000 40800
rect -31040 40732 -31028 40788
rect -30972 40732 -30708 40788
rect -30652 40732 -30388 40788
rect -30332 40732 -30068 40788
rect -30012 40732 -30000 40788
rect -31040 40720 -30000 40732
rect -12160 40708 -11440 40720
rect -12160 40652 -12148 40708
rect -12092 40652 -11828 40708
rect -11772 40652 -11508 40708
rect -11452 40652 -11440 40708
rect -12160 40640 -11440 40652
rect -10560 40708 -1040 40720
rect -10560 40652 -10548 40708
rect -10492 40652 -10228 40708
rect -10172 40652 -10068 40708
rect -10012 40652 -9908 40708
rect -9852 40652 -9748 40708
rect -9692 40652 -9588 40708
rect -9532 40652 -9428 40708
rect -9372 40652 -9268 40708
rect -9212 40652 -9108 40708
rect -9052 40652 -8948 40708
rect -8892 40652 -8788 40708
rect -8732 40652 -8628 40708
rect -8572 40652 -8468 40708
rect -8412 40652 -8308 40708
rect -8252 40652 -8148 40708
rect -8092 40652 -7988 40708
rect -7932 40652 -7828 40708
rect -7772 40652 -7668 40708
rect -7612 40652 -7508 40708
rect -7452 40652 -7348 40708
rect -7292 40652 -7188 40708
rect -7132 40652 -7028 40708
rect -6972 40652 -6868 40708
rect -6812 40652 -6708 40708
rect -6652 40652 -6548 40708
rect -6492 40652 -6388 40708
rect -6332 40652 -6228 40708
rect -6172 40652 -6068 40708
rect -6012 40652 -5908 40708
rect -5852 40652 -5748 40708
rect -5692 40652 -5588 40708
rect -5532 40652 -5428 40708
rect -5372 40652 -5268 40708
rect -5212 40652 -5108 40708
rect -5052 40652 -4948 40708
rect -4892 40652 -4788 40708
rect -4732 40652 -4628 40708
rect -4572 40652 -4468 40708
rect -4412 40652 -4308 40708
rect -4252 40652 -4148 40708
rect -4092 40652 -3988 40708
rect -3932 40652 -3668 40708
rect -3612 40652 -3508 40708
rect -3452 40652 -3348 40708
rect -3292 40652 -3028 40708
rect -2972 40652 -2708 40708
rect -2652 40652 -2388 40708
rect -2332 40652 -2068 40708
rect -2012 40652 -1748 40708
rect -1692 40652 -1428 40708
rect -1372 40652 -1108 40708
rect -1052 40652 -1040 40708
rect -10560 40640 -1040 40652
rect -31040 40628 -30000 40640
rect -31040 40572 -31028 40628
rect -30972 40572 -30708 40628
rect -30652 40572 -30388 40628
rect -30332 40572 -30068 40628
rect -30012 40572 -30000 40628
rect -31040 40560 -30000 40572
rect -10400 40548 -1200 40560
rect -10400 40492 -10388 40548
rect -10332 40492 -1268 40548
rect -1212 40492 -1200 40548
rect -10400 40480 -1200 40492
rect -31040 40468 -30000 40480
rect -31040 40412 -31028 40468
rect -30972 40412 -30708 40468
rect -30652 40412 -30388 40468
rect -30332 40412 -30068 40468
rect -30012 40412 -30000 40468
rect -31040 40400 -30000 40412
rect -12160 40388 -11440 40400
rect -12160 40332 -12148 40388
rect -12092 40332 -11828 40388
rect -11772 40332 -11508 40388
rect -11452 40332 -11440 40388
rect -12160 40320 -11440 40332
rect -10560 40388 -1040 40400
rect -10560 40332 -10548 40388
rect -10492 40332 -10228 40388
rect -10172 40332 -10068 40388
rect -10012 40332 -9908 40388
rect -9852 40332 -9748 40388
rect -9692 40332 -9588 40388
rect -9532 40332 -9428 40388
rect -9372 40332 -9268 40388
rect -9212 40332 -9108 40388
rect -9052 40332 -8948 40388
rect -8892 40332 -8788 40388
rect -8732 40332 -8628 40388
rect -8572 40332 -8468 40388
rect -8412 40332 -8308 40388
rect -8252 40332 -8148 40388
rect -8092 40332 -7988 40388
rect -7932 40332 -7828 40388
rect -7772 40332 -7668 40388
rect -7612 40332 -7508 40388
rect -7452 40332 -7348 40388
rect -7292 40332 -7188 40388
rect -7132 40332 -7028 40388
rect -6972 40332 -6868 40388
rect -6812 40332 -6708 40388
rect -6652 40332 -6548 40388
rect -6492 40332 -6388 40388
rect -6332 40332 -6228 40388
rect -6172 40332 -6068 40388
rect -6012 40332 -5908 40388
rect -5852 40332 -5748 40388
rect -5692 40332 -5588 40388
rect -5532 40332 -5428 40388
rect -5372 40332 -5268 40388
rect -5212 40332 -5108 40388
rect -5052 40332 -4948 40388
rect -4892 40332 -4788 40388
rect -4732 40332 -4628 40388
rect -4572 40332 -4468 40388
rect -4412 40332 -4308 40388
rect -4252 40332 -4148 40388
rect -4092 40332 -3988 40388
rect -3932 40332 -3668 40388
rect -3612 40332 -3508 40388
rect -3452 40332 -3348 40388
rect -3292 40332 -3028 40388
rect -2972 40332 -2708 40388
rect -2652 40332 -2388 40388
rect -2332 40332 -2068 40388
rect -2012 40332 -1748 40388
rect -1692 40332 -1428 40388
rect -1372 40332 -1108 40388
rect -1052 40332 -1040 40388
rect -10560 40320 -1040 40332
rect -31040 40308 -30000 40320
rect -31040 40252 -31028 40308
rect -30972 40252 -30708 40308
rect -30652 40252 -30388 40308
rect -30332 40252 -30068 40308
rect -30012 40252 -30000 40308
rect -31040 40240 -30000 40252
rect -3360 40228 -2640 40240
rect -3360 40172 -3348 40228
rect -3292 40172 -3028 40228
rect -2972 40172 -2708 40228
rect -2652 40172 -2640 40228
rect -3360 40160 -2640 40172
rect -2560 40228 -960 40240
rect -2560 40172 -2548 40228
rect -2492 40172 -1908 40228
rect -1852 40172 -960 40228
rect -2560 40160 -960 40172
rect -31040 40148 -30000 40160
rect -31040 40092 -31028 40148
rect -30972 40092 -30708 40148
rect -30652 40092 -30388 40148
rect -30332 40092 -30068 40148
rect -30012 40092 -30000 40148
rect -31040 40080 -30000 40092
rect -3360 40068 -1040 40080
rect -3360 40012 -3348 40068
rect -3292 40012 -3028 40068
rect -2972 40012 -2708 40068
rect -2652 40012 -2388 40068
rect -2332 40012 -2068 40068
rect -2012 40012 -1748 40068
rect -1692 40012 -1428 40068
rect -1372 40012 -1108 40068
rect -1052 40012 -1040 40068
rect -3360 40000 -1040 40012
rect 40960 40068 43200 40080
rect 40960 40012 41052 40068
rect 41108 40012 41212 40068
rect 41268 40012 41372 40068
rect 41428 40012 41532 40068
rect 41588 40012 41692 40068
rect 41748 40012 41852 40068
rect 41908 40012 42012 40068
rect 42068 40012 42172 40068
rect 42228 40012 42332 40068
rect 42388 40012 42492 40068
rect 42548 40012 42652 40068
rect 42708 40012 42812 40068
rect 42868 40012 42972 40068
rect 43028 40012 43132 40068
rect 43188 40012 43200 40068
rect 40960 40000 43200 40012
rect -31040 39988 -30000 40000
rect -31040 39932 -31028 39988
rect -30972 39932 -30708 39988
rect -30652 39932 -30388 39988
rect -30332 39932 -30068 39988
rect -30012 39932 -30000 39988
rect -31040 39920 -30000 39932
rect -3360 39908 -2320 39920
rect -3360 39852 -3348 39908
rect -3292 39852 -3028 39908
rect -2972 39852 -2708 39908
rect -2652 39852 -2388 39908
rect -2332 39852 -2320 39908
rect -3360 39840 -2320 39852
rect -2240 39908 43360 39920
rect -2240 39852 -2228 39908
rect -2172 39852 -1588 39908
rect -1532 39852 43360 39908
rect -2240 39840 43360 39852
rect -31040 39828 -30000 39840
rect -31040 39772 -31028 39828
rect -30972 39772 -30708 39828
rect -30652 39772 -30388 39828
rect -30332 39772 -30068 39828
rect -30012 39772 -30000 39828
rect -31040 39760 -30000 39772
rect -3360 39748 -1040 39760
rect -3360 39692 -3348 39748
rect -3292 39692 -3028 39748
rect -2972 39692 -2708 39748
rect -2652 39692 -2388 39748
rect -2332 39692 -2068 39748
rect -2012 39692 -1748 39748
rect -1692 39692 -1428 39748
rect -1372 39692 -1108 39748
rect -1052 39692 -1040 39748
rect -3360 39680 -1040 39692
rect 40960 39748 43200 39760
rect 40960 39692 41052 39748
rect 41108 39692 41212 39748
rect 41268 39692 41372 39748
rect 41428 39692 41532 39748
rect 41588 39692 41692 39748
rect 41748 39692 41852 39748
rect 41908 39692 42012 39748
rect 42068 39692 42172 39748
rect 42228 39692 42332 39748
rect 42388 39692 42492 39748
rect 42548 39692 42652 39748
rect 42708 39692 42812 39748
rect 42868 39692 42972 39748
rect 43028 39692 43132 39748
rect 43188 39692 43200 39748
rect 40960 39680 43200 39692
rect -31040 39668 -30000 39680
rect -31040 39612 -31028 39668
rect -30972 39612 -30708 39668
rect -30652 39612 -30388 39668
rect -30332 39612 -30068 39668
rect -30012 39612 -30000 39668
rect -31040 39600 -30000 39612
rect -3360 39588 -1040 39600
rect -3360 39532 -3348 39588
rect -3292 39532 -3028 39588
rect -2972 39532 -2708 39588
rect -2652 39532 -2388 39588
rect -2332 39532 -2068 39588
rect -2012 39532 -1748 39588
rect -1692 39532 -1428 39588
rect -1372 39532 -1108 39588
rect -1052 39532 -1040 39588
rect -3360 39520 -1040 39532
rect -31040 39508 -30000 39520
rect -31040 39452 -31028 39508
rect -30972 39452 -30708 39508
rect -30652 39452 -30388 39508
rect -30332 39452 -30068 39508
rect -30012 39452 -30000 39508
rect -31040 39440 -30000 39452
rect -3360 39428 -1040 39440
rect -3360 39372 -3348 39428
rect -3292 39372 -3028 39428
rect -2972 39372 -2708 39428
rect -2652 39372 -2388 39428
rect -2332 39372 -2068 39428
rect -2012 39372 -1748 39428
rect -1692 39372 -1428 39428
rect -1372 39372 -1108 39428
rect -1052 39372 -1040 39428
rect -3360 39360 -1040 39372
rect -31040 39348 -30000 39360
rect -31040 39292 -31028 39348
rect -30972 39292 -30708 39348
rect -30652 39292 -30388 39348
rect -30332 39292 -30068 39348
rect -30012 39292 -30000 39348
rect -31040 39280 -30000 39292
rect -3360 39268 -1040 39280
rect -3360 39212 -3348 39268
rect -3292 39212 -3028 39268
rect -2972 39212 -2708 39268
rect -2652 39212 -2388 39268
rect -2332 39212 -2068 39268
rect -2012 39212 -1748 39268
rect -1692 39212 -1428 39268
rect -1372 39212 -1108 39268
rect -1052 39212 -1040 39268
rect -3360 39200 -1040 39212
rect -31040 39188 -30000 39200
rect -31040 39132 -31028 39188
rect -30972 39132 -30708 39188
rect -30652 39132 -30388 39188
rect -30332 39132 -30068 39188
rect -30012 39132 -30000 39188
rect -31040 39120 -30000 39132
rect -3360 39108 -1040 39120
rect -3360 39052 -3348 39108
rect -3292 39052 -3028 39108
rect -2972 39052 -2708 39108
rect -2652 39052 -2388 39108
rect -2332 39052 -2068 39108
rect -2012 39052 -1748 39108
rect -1692 39052 -1428 39108
rect -1372 39052 -1108 39108
rect -1052 39052 -1040 39108
rect -3360 39040 -1040 39052
rect -31040 39028 -30000 39040
rect -31040 38972 -31028 39028
rect -30972 38972 -30708 39028
rect -30652 38972 -30388 39028
rect -30332 38972 -30068 39028
rect -30012 38972 -30000 39028
rect -31040 38960 -30000 38972
rect -3360 38948 -1040 38960
rect -3360 38892 -3348 38948
rect -3292 38892 -3028 38948
rect -2972 38892 -2708 38948
rect -2652 38892 -2388 38948
rect -2332 38892 -2068 38948
rect -2012 38892 -1748 38948
rect -1692 38892 -1428 38948
rect -1372 38892 -1108 38948
rect -1052 38892 -1040 38948
rect -3360 38880 -1040 38892
rect -31040 38868 -30000 38880
rect -31040 38812 -31028 38868
rect -30972 38812 -30708 38868
rect -30652 38812 -30388 38868
rect -30332 38812 -30068 38868
rect -30012 38812 -30000 38868
rect -31040 38800 -30000 38812
rect -3360 38788 -1040 38800
rect -3360 38732 -3348 38788
rect -3292 38732 -3028 38788
rect -2972 38732 -2708 38788
rect -2652 38732 -2388 38788
rect -2332 38732 -2068 38788
rect -2012 38732 -1748 38788
rect -1692 38732 -1428 38788
rect -1372 38732 -1108 38788
rect -1052 38732 -1040 38788
rect -3360 38720 -1040 38732
rect -31040 38708 -30000 38720
rect -31040 38652 -31028 38708
rect -30972 38652 -30708 38708
rect -30652 38652 -30388 38708
rect -30332 38652 -30068 38708
rect -30012 38652 -30000 38708
rect -31040 38640 -30000 38652
rect -3360 38628 -1040 38640
rect -3360 38572 -3348 38628
rect -3292 38572 -3028 38628
rect -2972 38572 -2708 38628
rect -2652 38572 -2388 38628
rect -2332 38572 -2068 38628
rect -2012 38572 -1748 38628
rect -1692 38572 -1428 38628
rect -1372 38572 -1108 38628
rect -1052 38572 -1040 38628
rect -3360 38560 -1040 38572
rect -31040 38548 -30000 38560
rect -31040 38492 -31028 38548
rect -30972 38492 -30708 38548
rect -30652 38492 -30388 38548
rect -30332 38492 -30068 38548
rect -30012 38492 -30000 38548
rect -31040 38480 -30000 38492
rect -3360 38468 -1040 38480
rect -3360 38412 -3348 38468
rect -3292 38412 -3028 38468
rect -2972 38412 -2708 38468
rect -2652 38412 -2388 38468
rect -2332 38412 -2068 38468
rect -2012 38412 -1748 38468
rect -1692 38412 -1428 38468
rect -1372 38412 -1108 38468
rect -1052 38412 -1040 38468
rect -3360 38400 -1040 38412
rect -31040 38388 -30000 38400
rect -31040 38332 -31028 38388
rect -30972 38332 -30708 38388
rect -30652 38332 -30388 38388
rect -30332 38332 -30068 38388
rect -30012 38332 -30000 38388
rect -31040 38320 -30000 38332
rect -3360 38308 -1040 38320
rect -3360 38252 -3348 38308
rect -3292 38252 -3028 38308
rect -2972 38252 -2708 38308
rect -2652 38252 -2388 38308
rect -2332 38252 -2068 38308
rect -2012 38252 -1748 38308
rect -1692 38252 -1428 38308
rect -1372 38252 -1108 38308
rect -1052 38252 -1040 38308
rect -3360 38240 -1040 38252
rect -31040 38228 -30000 38240
rect -31040 38172 -31028 38228
rect -30972 38172 -30708 38228
rect -30652 38172 -30388 38228
rect -30332 38172 -30068 38228
rect -30012 38172 -30000 38228
rect -31040 38160 -30000 38172
rect -3360 38148 -1040 38160
rect -3360 38092 -3348 38148
rect -3292 38092 -3028 38148
rect -2972 38092 -2708 38148
rect -2652 38092 -2388 38148
rect -2332 38092 -2068 38148
rect -2012 38092 -1748 38148
rect -1692 38092 -1428 38148
rect -1372 38092 -1108 38148
rect -1052 38092 -1040 38148
rect -3360 38080 -1040 38092
rect -31040 38068 -30000 38080
rect -31040 38012 -31028 38068
rect -30972 38012 -30708 38068
rect -30652 38012 -30388 38068
rect -30332 38012 -30068 38068
rect -30012 38012 -30000 38068
rect -31040 38000 -30000 38012
rect -3360 37988 -1040 38000
rect -3360 37932 -3348 37988
rect -3292 37932 -3028 37988
rect -2972 37932 -2708 37988
rect -2652 37932 -2388 37988
rect -2332 37932 -2068 37988
rect -2012 37932 -1748 37988
rect -1692 37932 -1428 37988
rect -1372 37932 -1108 37988
rect -1052 37932 -1040 37988
rect -3360 37920 -1040 37932
rect -31040 37908 -30000 37920
rect -31040 37852 -31028 37908
rect -30972 37852 -30708 37908
rect -30652 37852 -30388 37908
rect -30332 37852 -30068 37908
rect -30012 37852 -30000 37908
rect -31040 37840 -30000 37852
rect -3360 37828 -1040 37840
rect -3360 37772 -3348 37828
rect -3292 37772 -3028 37828
rect -2972 37772 -2708 37828
rect -2652 37772 -2388 37828
rect -2332 37772 -2068 37828
rect -2012 37772 -1748 37828
rect -1692 37772 -1428 37828
rect -1372 37772 -1108 37828
rect -1052 37772 -1040 37828
rect -3360 37760 -1040 37772
rect -33120 37748 -30000 37760
rect -33120 37692 -33108 37748
rect -33052 37692 -32948 37748
rect -32892 37692 -32788 37748
rect -32732 37692 -32628 37748
rect -32572 37692 -32468 37748
rect -32412 37692 -32308 37748
rect -32252 37692 -32148 37748
rect -32092 37692 -31988 37748
rect -31932 37692 -31828 37748
rect -31772 37692 -31668 37748
rect -31612 37692 -31508 37748
rect -31452 37692 -31348 37748
rect -31292 37692 -31188 37748
rect -31132 37692 -31028 37748
rect -30972 37692 -30708 37748
rect -30652 37692 -30388 37748
rect -30332 37692 -30068 37748
rect -30012 37692 -30000 37748
rect -33120 37680 -30000 37692
rect -3360 37668 -1360 37680
rect -3360 37612 -3348 37668
rect -3292 37612 -3028 37668
rect -2972 37612 -2708 37668
rect -2652 37612 -2388 37668
rect -2332 37612 -2068 37668
rect -2012 37612 -1748 37668
rect -1692 37612 -1428 37668
rect -1372 37612 -1360 37668
rect -3360 37600 -1360 37612
rect -1280 37668 40960 37680
rect -1280 37612 -1268 37668
rect -1212 37612 40960 37668
rect -1280 37600 40960 37612
rect -33280 37588 -30480 37600
rect -33280 37532 -30868 37588
rect -30812 37532 -30548 37588
rect -30492 37532 -30480 37588
rect -33280 37520 -30480 37532
rect -3360 37508 -1040 37520
rect -3360 37452 -3348 37508
rect -3292 37452 -3028 37508
rect -2972 37452 -2708 37508
rect -2652 37452 -2388 37508
rect -2332 37452 -2068 37508
rect -2012 37452 -1748 37508
rect -1692 37452 -1428 37508
rect -1372 37452 -1108 37508
rect -1052 37452 -1040 37508
rect -3360 37440 -1040 37452
rect -33120 37428 -30000 37440
rect -33120 37372 -33108 37428
rect -33052 37372 -32948 37428
rect -32892 37372 -32788 37428
rect -32732 37372 -32628 37428
rect -32572 37372 -32468 37428
rect -32412 37372 -32308 37428
rect -32252 37372 -32148 37428
rect -32092 37372 -31988 37428
rect -31932 37372 -31828 37428
rect -31772 37372 -31668 37428
rect -31612 37372 -31508 37428
rect -31452 37372 -31348 37428
rect -31292 37372 -31188 37428
rect -31132 37372 -31028 37428
rect -30972 37372 -30708 37428
rect -30652 37372 -30388 37428
rect -30332 37372 -30068 37428
rect -30012 37372 -30000 37428
rect -33120 37360 -30000 37372
rect -3360 37348 -1040 37360
rect -3360 37292 -3348 37348
rect -3292 37292 -3028 37348
rect -2972 37292 -2708 37348
rect -2652 37292 -2388 37348
rect -2332 37292 -2068 37348
rect -2012 37292 -1748 37348
rect -1692 37292 -1428 37348
rect -1372 37292 -1108 37348
rect -1052 37292 -1040 37348
rect -3360 37280 -1040 37292
rect -33280 37268 -30160 37280
rect -33280 37212 -30868 37268
rect -30812 37212 -30228 37268
rect -30172 37212 -30160 37268
rect -33280 37200 -30160 37212
rect -3360 37188 -1040 37200
rect -3360 37132 -3348 37188
rect -3292 37132 -3028 37188
rect -2972 37132 -2708 37188
rect -2652 37132 -2388 37188
rect -2332 37132 -2068 37188
rect -2012 37132 -1748 37188
rect -1692 37132 -1428 37188
rect -1372 37132 -1108 37188
rect -1052 37132 -1040 37188
rect -3360 37120 -1040 37132
rect -33120 37108 -30000 37120
rect -33120 37052 -33108 37108
rect -33052 37052 -32948 37108
rect -32892 37052 -32788 37108
rect -32732 37052 -32628 37108
rect -32572 37052 -32468 37108
rect -32412 37052 -32308 37108
rect -32252 37052 -32148 37108
rect -32092 37052 -31988 37108
rect -31932 37052 -31828 37108
rect -31772 37052 -31668 37108
rect -31612 37052 -31508 37108
rect -31452 37052 -31348 37108
rect -31292 37052 -31188 37108
rect -31132 37052 -31028 37108
rect -30972 37052 -30708 37108
rect -30652 37052 -30388 37108
rect -30332 37052 -30068 37108
rect -30012 37052 -30000 37108
rect -33120 37040 -30000 37052
rect -3360 37028 -1040 37040
rect -3360 36972 -3348 37028
rect -3292 36972 -3028 37028
rect -2972 36972 -2708 37028
rect -2652 36972 -2388 37028
rect -2332 36972 -2068 37028
rect -2012 36972 -1748 37028
rect -1692 36972 -1428 37028
rect -1372 36972 -1108 37028
rect -1052 36972 -1040 37028
rect -3360 36960 -1040 36972
rect -31040 36948 -30000 36960
rect -31040 36892 -31028 36948
rect -30972 36892 -30708 36948
rect -30652 36892 -30388 36948
rect -30332 36892 -30068 36948
rect -30012 36892 -30000 36948
rect -31040 36880 -30000 36892
rect -3360 36868 -1040 36880
rect -3360 36812 -3348 36868
rect -3292 36812 -3028 36868
rect -2972 36812 -2708 36868
rect -2652 36812 -2388 36868
rect -2332 36812 -2068 36868
rect -2012 36812 -1748 36868
rect -1692 36812 -1428 36868
rect -1372 36812 -1108 36868
rect -1052 36812 -1040 36868
rect -3360 36800 -1040 36812
rect -31040 36788 -30000 36800
rect -31040 36732 -31028 36788
rect -30972 36732 -30708 36788
rect -30652 36732 -30388 36788
rect -30332 36732 -30068 36788
rect -30012 36732 -30000 36788
rect -31040 36720 -30000 36732
rect -3360 36708 -1040 36720
rect -3360 36652 -3348 36708
rect -3292 36652 -3028 36708
rect -2972 36652 -2708 36708
rect -2652 36652 -2388 36708
rect -2332 36652 -2068 36708
rect -2012 36652 -1748 36708
rect -1692 36652 -1428 36708
rect -1372 36652 -1108 36708
rect -1052 36652 -1040 36708
rect -3360 36640 -1040 36652
rect -31040 36628 -30000 36640
rect -31040 36572 -31028 36628
rect -30972 36572 -30708 36628
rect -30652 36572 -30388 36628
rect -30332 36572 -30068 36628
rect -30012 36572 -30000 36628
rect -31040 36560 -30000 36572
rect -3360 36548 -1040 36560
rect -3360 36492 -3348 36548
rect -3292 36492 -3028 36548
rect -2972 36492 -2708 36548
rect -2652 36492 -2388 36548
rect -2332 36492 -2068 36548
rect -2012 36492 -1748 36548
rect -1692 36492 -1428 36548
rect -1372 36492 -1108 36548
rect -1052 36492 -1040 36548
rect -3360 36480 -1040 36492
rect -31040 36468 -30000 36480
rect -31040 36412 -31028 36468
rect -30972 36412 -30708 36468
rect -30652 36412 -30388 36468
rect -30332 36412 -30068 36468
rect -30012 36412 -30000 36468
rect -31040 36400 -30000 36412
rect -3360 36388 -1040 36400
rect -3360 36332 -3348 36388
rect -3292 36332 -3028 36388
rect -2972 36332 -2708 36388
rect -2652 36332 -2388 36388
rect -2332 36332 -2068 36388
rect -2012 36332 -1748 36388
rect -1692 36332 -1428 36388
rect -1372 36332 -1108 36388
rect -1052 36332 -1040 36388
rect -3360 36320 -1040 36332
rect -31040 36308 -30000 36320
rect -31040 36252 -31028 36308
rect -30972 36252 -30708 36308
rect -30652 36252 -30388 36308
rect -30332 36252 -30068 36308
rect -30012 36252 -30000 36308
rect -31040 36240 -30000 36252
rect -3360 36228 -2960 36240
rect -3360 36172 -3348 36228
rect -3292 36172 -3028 36228
rect -2972 36172 -2960 36228
rect -3360 36160 -2960 36172
rect -2880 36228 -960 36240
rect -2880 36172 -2868 36228
rect -2812 36172 -1908 36228
rect -1852 36172 -960 36228
rect -2880 36160 -960 36172
rect -31040 36148 -30000 36160
rect -31040 36092 -31028 36148
rect -30972 36092 -30708 36148
rect -30652 36092 -30388 36148
rect -30332 36092 -30068 36148
rect -30012 36092 -30000 36148
rect -31040 36080 -30000 36092
rect -3360 36068 -1040 36080
rect -3360 36012 -3348 36068
rect -3292 36012 -3028 36068
rect -2972 36012 -2708 36068
rect -2652 36012 -2388 36068
rect -2332 36012 -2068 36068
rect -2012 36012 -1748 36068
rect -1692 36012 -1428 36068
rect -1372 36012 -1108 36068
rect -1052 36012 -1040 36068
rect -3360 36000 -1040 36012
rect 40960 36068 43200 36080
rect 40960 36012 41052 36068
rect 41108 36012 41212 36068
rect 41268 36012 41372 36068
rect 41428 36012 41532 36068
rect 41588 36012 41692 36068
rect 41748 36012 41852 36068
rect 41908 36012 42012 36068
rect 42068 36012 42172 36068
rect 42228 36012 42332 36068
rect 42388 36012 42492 36068
rect 42548 36012 42652 36068
rect 42708 36012 42812 36068
rect 42868 36012 42972 36068
rect 43028 36012 43132 36068
rect 43188 36012 43200 36068
rect 40960 36000 43200 36012
rect -31040 35988 -30000 36000
rect -31040 35932 -31028 35988
rect -30972 35932 -30708 35988
rect -30652 35932 -30388 35988
rect -30332 35932 -30068 35988
rect -30012 35932 -30000 35988
rect -31040 35920 -30000 35932
rect -3200 35908 43360 35920
rect -3200 35852 -3188 35908
rect -3132 35852 -1588 35908
rect -1532 35852 43360 35908
rect -3200 35840 43360 35852
rect -31040 35828 -30000 35840
rect -31040 35772 -31028 35828
rect -30972 35772 -30708 35828
rect -30652 35772 -30388 35828
rect -30332 35772 -30068 35828
rect -30012 35772 -30000 35828
rect -31040 35760 -30000 35772
rect -3360 35748 -1040 35760
rect -3360 35692 -3348 35748
rect -3292 35692 -3028 35748
rect -2972 35692 -2708 35748
rect -2652 35692 -2388 35748
rect -2332 35692 -2068 35748
rect -2012 35692 -1748 35748
rect -1692 35692 -1428 35748
rect -1372 35692 -1108 35748
rect -1052 35692 -1040 35748
rect -3360 35680 -1040 35692
rect 40960 35748 43200 35760
rect 40960 35692 41052 35748
rect 41108 35692 41212 35748
rect 41268 35692 41372 35748
rect 41428 35692 41532 35748
rect 41588 35692 41692 35748
rect 41748 35692 41852 35748
rect 41908 35692 42012 35748
rect 42068 35692 42172 35748
rect 42228 35692 42332 35748
rect 42388 35692 42492 35748
rect 42548 35692 42652 35748
rect 42708 35692 42812 35748
rect 42868 35692 42972 35748
rect 43028 35692 43132 35748
rect 43188 35692 43200 35748
rect 40960 35680 43200 35692
rect -31040 35668 -30000 35680
rect -31040 35612 -31028 35668
rect -30972 35612 -30708 35668
rect -30652 35612 -30388 35668
rect -30332 35612 -30068 35668
rect -30012 35612 -30000 35668
rect -31040 35600 -30000 35612
rect -3360 35588 -1040 35600
rect -3360 35532 -3348 35588
rect -3292 35532 -3028 35588
rect -2972 35532 -2708 35588
rect -2652 35532 -2388 35588
rect -2332 35532 -2068 35588
rect -2012 35532 -1748 35588
rect -1692 35532 -1428 35588
rect -1372 35532 -1108 35588
rect -1052 35532 -1040 35588
rect -3360 35520 -1040 35532
rect -31040 35508 -30000 35520
rect -31040 35452 -31028 35508
rect -30972 35452 -30708 35508
rect -30652 35452 -30388 35508
rect -30332 35452 -30068 35508
rect -30012 35452 -30000 35508
rect -31040 35440 -30000 35452
rect -3360 35428 -1040 35440
rect -3360 35372 -3348 35428
rect -3292 35372 -3028 35428
rect -2972 35372 -2708 35428
rect -2652 35372 -2388 35428
rect -2332 35372 -2068 35428
rect -2012 35372 -1748 35428
rect -1692 35372 -1428 35428
rect -1372 35372 -1108 35428
rect -1052 35372 -1040 35428
rect -3360 35360 -1040 35372
rect -31040 35348 -30000 35360
rect -31040 35292 -31028 35348
rect -30972 35292 -30708 35348
rect -30652 35292 -30388 35348
rect -30332 35292 -30068 35348
rect -30012 35292 -30000 35348
rect -31040 35280 -30000 35292
rect -3360 35268 -1040 35280
rect -3360 35212 -3348 35268
rect -3292 35212 -3028 35268
rect -2972 35212 -2708 35268
rect -2652 35212 -2388 35268
rect -2332 35212 -2068 35268
rect -2012 35212 -1748 35268
rect -1692 35212 -1428 35268
rect -1372 35212 -1108 35268
rect -1052 35212 -1040 35268
rect -3360 35200 -1040 35212
rect -31040 35188 -30000 35200
rect -31040 35132 -31028 35188
rect -30972 35132 -30708 35188
rect -30652 35132 -30388 35188
rect -30332 35132 -30068 35188
rect -30012 35132 -30000 35188
rect -31040 35120 -30000 35132
rect -3360 35108 -1040 35120
rect -3360 35052 -3348 35108
rect -3292 35052 -3028 35108
rect -2972 35052 -2708 35108
rect -2652 35052 -2388 35108
rect -2332 35052 -2068 35108
rect -2012 35052 -1748 35108
rect -1692 35052 -1428 35108
rect -1372 35052 -1108 35108
rect -1052 35052 -1040 35108
rect -3360 35040 -1040 35052
rect -31040 35028 -30000 35040
rect -31040 34972 -31028 35028
rect -30972 34972 -30708 35028
rect -30652 34972 -30388 35028
rect -30332 34972 -30068 35028
rect -30012 34972 -30000 35028
rect -31040 34960 -30000 34972
rect -3360 34948 -1040 34960
rect -3360 34892 -3348 34948
rect -3292 34892 -3028 34948
rect -2972 34892 -2708 34948
rect -2652 34892 -2388 34948
rect -2332 34892 -2068 34948
rect -2012 34892 -1748 34948
rect -1692 34892 -1428 34948
rect -1372 34892 -1108 34948
rect -1052 34892 -1040 34948
rect -3360 34880 -1040 34892
rect -31040 34868 -30000 34880
rect -31040 34812 -31028 34868
rect -30972 34812 -30708 34868
rect -30652 34812 -30388 34868
rect -30332 34812 -30068 34868
rect -30012 34812 -30000 34868
rect -31040 34800 -30000 34812
rect -3360 34788 -1040 34800
rect -3360 34732 -3348 34788
rect -3292 34732 -3028 34788
rect -2972 34732 -2708 34788
rect -2652 34732 -2388 34788
rect -2332 34732 -2068 34788
rect -2012 34732 -1748 34788
rect -1692 34732 -1428 34788
rect -1372 34732 -1108 34788
rect -1052 34732 -1040 34788
rect -3360 34720 -1040 34732
rect -33120 34708 -10480 34720
rect -33120 34652 -33108 34708
rect -33052 34652 -32948 34708
rect -32892 34652 -32788 34708
rect -32732 34652 -32628 34708
rect -32572 34652 -32468 34708
rect -32412 34652 -32308 34708
rect -32252 34652 -32148 34708
rect -32092 34652 -31988 34708
rect -31932 34652 -31828 34708
rect -31772 34652 -31668 34708
rect -31612 34652 -31508 34708
rect -31452 34652 -31348 34708
rect -31292 34652 -31188 34708
rect -31132 34652 -31028 34708
rect -30972 34652 -30708 34708
rect -30652 34652 -30388 34708
rect -30332 34652 -30068 34708
rect -30012 34652 -29908 34708
rect -29852 34652 -29748 34708
rect -29692 34652 -29588 34708
rect -29532 34652 -29428 34708
rect -29372 34652 -29268 34708
rect -29212 34652 -29108 34708
rect -29052 34652 -28948 34708
rect -28892 34652 -28788 34708
rect -28732 34652 -28628 34708
rect -28572 34652 -28468 34708
rect -28412 34652 -28308 34708
rect -28252 34652 -28148 34708
rect -28092 34652 -27988 34708
rect -27932 34652 -27828 34708
rect -27772 34652 -27668 34708
rect -27612 34652 -27508 34708
rect -27452 34652 -27348 34708
rect -27292 34652 -27188 34708
rect -27132 34652 -27028 34708
rect -26972 34652 -26868 34708
rect -26812 34652 -26708 34708
rect -26652 34652 -26548 34708
rect -26492 34652 -26388 34708
rect -26332 34652 -26228 34708
rect -26172 34652 -26068 34708
rect -26012 34652 -25908 34708
rect -25852 34652 -25748 34708
rect -25692 34652 -25588 34708
rect -25532 34652 -25428 34708
rect -25372 34652 -25268 34708
rect -25212 34652 -25108 34708
rect -25052 34652 -24948 34708
rect -24892 34652 -24788 34708
rect -24732 34652 -24628 34708
rect -24572 34652 -24468 34708
rect -24412 34652 -24308 34708
rect -24252 34652 -24148 34708
rect -24092 34652 -23988 34708
rect -23932 34652 -23828 34708
rect -23772 34652 -23668 34708
rect -23612 34652 -23508 34708
rect -23452 34652 -23348 34708
rect -23292 34652 -23188 34708
rect -23132 34652 -23028 34708
rect -22972 34652 -22868 34708
rect -22812 34652 -22708 34708
rect -22652 34652 -22548 34708
rect -22492 34652 -22388 34708
rect -22332 34652 -22228 34708
rect -22172 34652 -22068 34708
rect -22012 34652 -21908 34708
rect -21852 34652 -21748 34708
rect -21692 34652 -21588 34708
rect -21532 34652 -21428 34708
rect -21372 34652 -21268 34708
rect -21212 34652 -21108 34708
rect -21052 34652 -20948 34708
rect -20892 34652 -20788 34708
rect -20732 34652 -20628 34708
rect -20572 34652 -20468 34708
rect -20412 34652 -20308 34708
rect -20252 34652 -20148 34708
rect -20092 34652 -19988 34708
rect -19932 34652 -19828 34708
rect -19772 34652 -19668 34708
rect -19612 34652 -19508 34708
rect -19452 34652 -19348 34708
rect -19292 34652 -19188 34708
rect -19132 34652 -19028 34708
rect -18972 34652 -18868 34708
rect -18812 34652 -18708 34708
rect -18652 34652 -18548 34708
rect -18492 34652 -18388 34708
rect -18332 34652 -18228 34708
rect -18172 34652 -18068 34708
rect -18012 34652 -17908 34708
rect -17852 34652 -17748 34708
rect -17692 34652 -17588 34708
rect -17532 34652 -17428 34708
rect -17372 34652 -17268 34708
rect -17212 34652 -17108 34708
rect -17052 34652 -16948 34708
rect -16892 34652 -16788 34708
rect -16732 34652 -16628 34708
rect -16572 34652 -16468 34708
rect -16412 34652 -16308 34708
rect -16252 34652 -16148 34708
rect -16092 34652 -15988 34708
rect -15932 34652 -15828 34708
rect -15772 34652 -15668 34708
rect -15612 34652 -15508 34708
rect -15452 34652 -15348 34708
rect -15292 34652 -15188 34708
rect -15132 34652 -15028 34708
rect -14972 34652 -14868 34708
rect -14812 34652 -14708 34708
rect -14652 34652 -14548 34708
rect -14492 34652 -14388 34708
rect -14332 34652 -14228 34708
rect -14172 34652 -14068 34708
rect -14012 34652 -13908 34708
rect -13852 34652 -13748 34708
rect -13692 34652 -13588 34708
rect -13532 34652 -13428 34708
rect -13372 34652 -13268 34708
rect -13212 34652 -13108 34708
rect -13052 34652 -12948 34708
rect -12892 34652 -12788 34708
rect -12732 34652 -12628 34708
rect -12572 34652 -12468 34708
rect -12412 34652 -12308 34708
rect -12252 34652 -12148 34708
rect -12092 34652 -11988 34708
rect -11932 34652 -11828 34708
rect -11772 34652 -11668 34708
rect -11612 34652 -11508 34708
rect -11452 34652 -11188 34708
rect -11132 34652 -10868 34708
rect -10812 34652 -10548 34708
rect -10492 34652 -10480 34708
rect -33120 34640 -10480 34652
rect -3360 34628 -1040 34640
rect -3360 34572 -3348 34628
rect -3292 34572 -3028 34628
rect -2972 34572 -2708 34628
rect -2652 34572 -2388 34628
rect -2332 34572 -2068 34628
rect -2012 34572 -1748 34628
rect -1692 34572 -1428 34628
rect -1372 34572 -1108 34628
rect -1052 34572 -1040 34628
rect -3360 34560 -1040 34572
rect -33280 34548 -10640 34560
rect -33280 34492 -10708 34548
rect -10652 34492 -10640 34548
rect -33280 34480 -10640 34492
rect -10560 34480 -10480 34560
rect -3360 34468 -1040 34480
rect -3360 34412 -3348 34468
rect -3292 34412 -3028 34468
rect -2972 34412 -2708 34468
rect -2652 34412 -2388 34468
rect -2332 34412 -2068 34468
rect -2012 34412 -1748 34468
rect -1692 34412 -1428 34468
rect -1372 34412 -1108 34468
rect -1052 34412 -1040 34468
rect -3360 34400 -1040 34412
rect -33120 34388 -10480 34400
rect -33120 34332 -33108 34388
rect -33052 34332 -32948 34388
rect -32892 34332 -32788 34388
rect -32732 34332 -32628 34388
rect -32572 34332 -32468 34388
rect -32412 34332 -32308 34388
rect -32252 34332 -32148 34388
rect -32092 34332 -31988 34388
rect -31932 34332 -31828 34388
rect -31772 34332 -31668 34388
rect -31612 34332 -31508 34388
rect -31452 34332 -31348 34388
rect -31292 34332 -31188 34388
rect -31132 34332 -31028 34388
rect -30972 34332 -30708 34388
rect -30652 34332 -30388 34388
rect -30332 34332 -30068 34388
rect -30012 34332 -29908 34388
rect -29852 34332 -29748 34388
rect -29692 34332 -29588 34388
rect -29532 34332 -29428 34388
rect -29372 34332 -29268 34388
rect -29212 34332 -29108 34388
rect -29052 34332 -28948 34388
rect -28892 34332 -28788 34388
rect -28732 34332 -28628 34388
rect -28572 34332 -28468 34388
rect -28412 34332 -28308 34388
rect -28252 34332 -28148 34388
rect -28092 34332 -27988 34388
rect -27932 34332 -27828 34388
rect -27772 34332 -27668 34388
rect -27612 34332 -27508 34388
rect -27452 34332 -27348 34388
rect -27292 34332 -27188 34388
rect -27132 34332 -27028 34388
rect -26972 34332 -26868 34388
rect -26812 34332 -26708 34388
rect -26652 34332 -26548 34388
rect -26492 34332 -26388 34388
rect -26332 34332 -26228 34388
rect -26172 34332 -26068 34388
rect -26012 34332 -25908 34388
rect -25852 34332 -25748 34388
rect -25692 34332 -25588 34388
rect -25532 34332 -25428 34388
rect -25372 34332 -25268 34388
rect -25212 34332 -25108 34388
rect -25052 34332 -24948 34388
rect -24892 34332 -24788 34388
rect -24732 34332 -24628 34388
rect -24572 34332 -24468 34388
rect -24412 34332 -24308 34388
rect -24252 34332 -24148 34388
rect -24092 34332 -23988 34388
rect -23932 34332 -23828 34388
rect -23772 34332 -23668 34388
rect -23612 34332 -23508 34388
rect -23452 34332 -23348 34388
rect -23292 34332 -23188 34388
rect -23132 34332 -23028 34388
rect -22972 34332 -22868 34388
rect -22812 34332 -22708 34388
rect -22652 34332 -22548 34388
rect -22492 34332 -22388 34388
rect -22332 34332 -22228 34388
rect -22172 34332 -22068 34388
rect -22012 34332 -21908 34388
rect -21852 34332 -21748 34388
rect -21692 34332 -21588 34388
rect -21532 34332 -21428 34388
rect -21372 34332 -21268 34388
rect -21212 34332 -21108 34388
rect -21052 34332 -20948 34388
rect -20892 34332 -20788 34388
rect -20732 34332 -20628 34388
rect -20572 34332 -20468 34388
rect -20412 34332 -20308 34388
rect -20252 34332 -20148 34388
rect -20092 34332 -19988 34388
rect -19932 34332 -19828 34388
rect -19772 34332 -19668 34388
rect -19612 34332 -19508 34388
rect -19452 34332 -19348 34388
rect -19292 34332 -19188 34388
rect -19132 34332 -19028 34388
rect -18972 34332 -18868 34388
rect -18812 34332 -18708 34388
rect -18652 34332 -18548 34388
rect -18492 34332 -18388 34388
rect -18332 34332 -18228 34388
rect -18172 34332 -18068 34388
rect -18012 34332 -17908 34388
rect -17852 34332 -17748 34388
rect -17692 34332 -17588 34388
rect -17532 34332 -17428 34388
rect -17372 34332 -17268 34388
rect -17212 34332 -17108 34388
rect -17052 34332 -16948 34388
rect -16892 34332 -16788 34388
rect -16732 34332 -16628 34388
rect -16572 34332 -16468 34388
rect -16412 34332 -16308 34388
rect -16252 34332 -16148 34388
rect -16092 34332 -15988 34388
rect -15932 34332 -15828 34388
rect -15772 34332 -15668 34388
rect -15612 34332 -15508 34388
rect -15452 34332 -15348 34388
rect -15292 34332 -15188 34388
rect -15132 34332 -15028 34388
rect -14972 34332 -14868 34388
rect -14812 34332 -14708 34388
rect -14652 34332 -14548 34388
rect -14492 34332 -14388 34388
rect -14332 34332 -14228 34388
rect -14172 34332 -14068 34388
rect -14012 34332 -13908 34388
rect -13852 34332 -13748 34388
rect -13692 34332 -13588 34388
rect -13532 34332 -13428 34388
rect -13372 34332 -13268 34388
rect -13212 34332 -13108 34388
rect -13052 34332 -12948 34388
rect -12892 34332 -12788 34388
rect -12732 34332 -12628 34388
rect -12572 34332 -12468 34388
rect -12412 34332 -12308 34388
rect -12252 34332 -12148 34388
rect -12092 34332 -11988 34388
rect -11932 34332 -11828 34388
rect -11772 34332 -11668 34388
rect -11612 34332 -11508 34388
rect -11452 34332 -11188 34388
rect -11132 34332 -10868 34388
rect -10812 34332 -10548 34388
rect -10492 34332 -10480 34388
rect -33120 34320 -10480 34332
rect -3360 34308 -1040 34320
rect -3360 34252 -3348 34308
rect -3292 34252 -3028 34308
rect -2972 34252 -2708 34308
rect -2652 34252 -2388 34308
rect -2332 34252 -2068 34308
rect -2012 34252 -1748 34308
rect -1692 34252 -1428 34308
rect -1372 34252 -1108 34308
rect -1052 34252 -1040 34308
rect -3360 34240 -1040 34252
rect -31040 34228 -30000 34240
rect -31040 34172 -31028 34228
rect -30972 34172 -30708 34228
rect -30652 34172 -30388 34228
rect -30332 34172 -30068 34228
rect -30012 34172 -30000 34228
rect -31040 34160 -30000 34172
rect -3360 34148 -1040 34160
rect -3360 34092 -3348 34148
rect -3292 34092 -3028 34148
rect -2972 34092 -2708 34148
rect -2652 34092 -2388 34148
rect -2332 34092 -2068 34148
rect -2012 34092 -1748 34148
rect -1692 34092 -1428 34148
rect -1372 34092 -1108 34148
rect -1052 34092 -1040 34148
rect -3360 34080 -1040 34092
rect -31040 34068 -30000 34080
rect -31040 34012 -31028 34068
rect -30972 34012 -30708 34068
rect -30652 34012 -30388 34068
rect -30332 34012 -30068 34068
rect -30012 34012 -30000 34068
rect -31040 34000 -30000 34012
rect -3360 33988 -1040 34000
rect -3360 33932 -3348 33988
rect -3292 33932 -3028 33988
rect -2972 33932 -2708 33988
rect -2652 33932 -2388 33988
rect -2332 33932 -2068 33988
rect -2012 33932 -1748 33988
rect -1692 33932 -1428 33988
rect -1372 33932 -1108 33988
rect -1052 33932 -1040 33988
rect -3360 33920 -1040 33932
rect -31040 33908 -30000 33920
rect -31040 33852 -31028 33908
rect -30972 33852 -30708 33908
rect -30652 33852 -30388 33908
rect -30332 33852 -30068 33908
rect -30012 33852 -30000 33908
rect -31040 33840 -30000 33852
rect -3360 33828 -1040 33840
rect -3360 33772 -3348 33828
rect -3292 33772 -3028 33828
rect -2972 33772 -2708 33828
rect -2652 33772 -2388 33828
rect -2332 33772 -2068 33828
rect -2012 33772 -1748 33828
rect -1692 33772 -1428 33828
rect -1372 33772 -1108 33828
rect -1052 33772 -1040 33828
rect -3360 33760 -1040 33772
rect -31040 33748 -30000 33760
rect -31040 33692 -31028 33748
rect -30972 33692 -30708 33748
rect -30652 33692 -30388 33748
rect -30332 33692 -30068 33748
rect -30012 33692 -30000 33748
rect -31040 33680 -30000 33692
rect -3360 33668 -1040 33680
rect -3360 33612 -3348 33668
rect -3292 33612 -3028 33668
rect -2972 33612 -2708 33668
rect -2652 33612 -2388 33668
rect -2332 33612 -2068 33668
rect -2012 33612 -1748 33668
rect -1692 33612 -1428 33668
rect -1372 33612 -1108 33668
rect -1052 33612 -1040 33668
rect -3360 33600 -1040 33612
rect -31040 33588 -30000 33600
rect -31040 33532 -31028 33588
rect -30972 33532 -30708 33588
rect -30652 33532 -30388 33588
rect -30332 33532 -30068 33588
rect -30012 33532 -30000 33588
rect -31040 33520 -30000 33532
rect -3360 33508 -1040 33520
rect -3360 33452 -3348 33508
rect -3292 33452 -3028 33508
rect -2972 33452 -2708 33508
rect -2652 33452 -2388 33508
rect -2332 33452 -2068 33508
rect -2012 33452 -1748 33508
rect -1692 33452 -1428 33508
rect -1372 33452 -1108 33508
rect -1052 33452 -1040 33508
rect -3360 33440 -1040 33452
rect -31040 33428 -30000 33440
rect -31040 33372 -31028 33428
rect -30972 33372 -30708 33428
rect -30652 33372 -30388 33428
rect -30332 33372 -30068 33428
rect -30012 33372 -30000 33428
rect -31040 33360 -30000 33372
rect -31040 33268 -30000 33280
rect -31040 33212 -31028 33268
rect -30972 33212 -30708 33268
rect -30652 33212 -30388 33268
rect -30332 33212 -30068 33268
rect -30012 33212 -30000 33268
rect -31040 33200 -30000 33212
rect -3360 33268 -1040 33280
rect -3360 33212 -3348 33268
rect -3292 33212 -3028 33268
rect -2972 33212 -2708 33268
rect -2652 33212 -2388 33268
rect -2332 33212 -2068 33268
rect -2012 33212 -1748 33268
rect -1692 33212 -1428 33268
rect -1372 33212 -1108 33268
rect -1052 33212 -1040 33268
rect -3360 33200 -1040 33212
rect -31040 33108 -30000 33120
rect -31040 33052 -31028 33108
rect -30972 33052 -30708 33108
rect -30652 33052 -30388 33108
rect -30332 33052 -30068 33108
rect -30012 33052 -30000 33108
rect -31040 33040 -30000 33052
rect -3360 33108 -1040 33120
rect -3360 33052 -3348 33108
rect -3292 33052 -3028 33108
rect -2972 33052 -2708 33108
rect -2652 33052 -2388 33108
rect -2332 33052 -2068 33108
rect -2012 33052 -1748 33108
rect -1692 33052 -1428 33108
rect -1372 33052 -1108 33108
rect -1052 33052 -1040 33108
rect -3360 33040 -1040 33052
rect -31040 32948 -1040 32960
rect -31040 32892 -31028 32948
rect -30972 32892 -30708 32948
rect -30652 32892 -30388 32948
rect -30332 32892 -30068 32948
rect -30012 32892 -29908 32948
rect -29852 32892 -29748 32948
rect -29692 32892 -29588 32948
rect -29532 32892 -29428 32948
rect -29372 32892 -29268 32948
rect -29212 32892 -29108 32948
rect -29052 32892 -28948 32948
rect -28892 32892 -28788 32948
rect -28732 32892 -28628 32948
rect -28572 32892 -28468 32948
rect -28412 32892 -28308 32948
rect -28252 32892 -28148 32948
rect -28092 32892 -27988 32948
rect -27932 32892 -27828 32948
rect -27772 32892 -27668 32948
rect -27612 32892 -27508 32948
rect -27452 32892 -27348 32948
rect -27292 32892 -27188 32948
rect -27132 32892 -27028 32948
rect -26972 32892 -26868 32948
rect -26812 32892 -26708 32948
rect -26652 32892 -26548 32948
rect -26492 32892 -26388 32948
rect -26332 32892 -26228 32948
rect -26172 32892 -26068 32948
rect -26012 32892 -25908 32948
rect -25852 32892 -25748 32948
rect -25692 32892 -25588 32948
rect -25532 32892 -25428 32948
rect -25372 32892 -25268 32948
rect -25212 32892 -25108 32948
rect -25052 32892 -24948 32948
rect -24892 32892 -24788 32948
rect -24732 32892 -24628 32948
rect -24572 32892 -24468 32948
rect -24412 32892 -24308 32948
rect -24252 32892 -24148 32948
rect -24092 32892 -23988 32948
rect -23932 32892 -23828 32948
rect -23772 32892 -23668 32948
rect -23612 32892 -23508 32948
rect -23452 32892 -23348 32948
rect -23292 32892 -23188 32948
rect -23132 32892 -23028 32948
rect -22972 32892 -22868 32948
rect -22812 32892 -22708 32948
rect -22652 32892 -22548 32948
rect -22492 32892 -22388 32948
rect -22332 32892 -22228 32948
rect -22172 32892 -22068 32948
rect -22012 32892 -21908 32948
rect -21852 32892 -21748 32948
rect -21692 32892 -21588 32948
rect -21532 32892 -21428 32948
rect -21372 32892 -21268 32948
rect -21212 32892 -21108 32948
rect -21052 32892 -20948 32948
rect -20892 32892 -20788 32948
rect -20732 32892 -20628 32948
rect -20572 32892 -20468 32948
rect -20412 32892 -20308 32948
rect -20252 32892 -20148 32948
rect -20092 32892 -19988 32948
rect -19932 32892 -19828 32948
rect -19772 32892 -19668 32948
rect -19612 32892 -19508 32948
rect -19452 32892 -19348 32948
rect -19292 32892 -19188 32948
rect -19132 32892 -19028 32948
rect -18972 32892 -18868 32948
rect -18812 32892 -18708 32948
rect -18652 32892 -18548 32948
rect -18492 32892 -18388 32948
rect -18332 32892 -18228 32948
rect -18172 32892 -18068 32948
rect -18012 32892 -17908 32948
rect -17852 32892 -17748 32948
rect -17692 32892 -17588 32948
rect -17532 32892 -17428 32948
rect -17372 32892 -17268 32948
rect -17212 32892 -17108 32948
rect -17052 32892 -16948 32948
rect -16892 32892 -16788 32948
rect -16732 32892 -16628 32948
rect -16572 32892 -16468 32948
rect -16412 32892 -16308 32948
rect -16252 32892 -16148 32948
rect -16092 32892 -15988 32948
rect -15932 32892 -15828 32948
rect -15772 32892 -15668 32948
rect -15612 32892 -15508 32948
rect -15452 32892 -15348 32948
rect -15292 32892 -15188 32948
rect -15132 32892 -15028 32948
rect -14972 32892 -14868 32948
rect -14812 32892 -14708 32948
rect -14652 32892 -14548 32948
rect -14492 32892 -14388 32948
rect -14332 32892 -14228 32948
rect -14172 32892 -14068 32948
rect -14012 32892 -13908 32948
rect -13852 32892 -13748 32948
rect -13692 32892 -13588 32948
rect -13532 32892 -13428 32948
rect -13372 32892 -13268 32948
rect -13212 32892 -13108 32948
rect -13052 32892 -12948 32948
rect -12892 32892 -12788 32948
rect -12732 32892 -12628 32948
rect -12572 32892 -12468 32948
rect -12412 32892 -12308 32948
rect -12252 32892 -12148 32948
rect -12092 32892 -11988 32948
rect -11932 32892 -11828 32948
rect -11772 32892 -11668 32948
rect -11612 32892 -11508 32948
rect -11452 32892 -11188 32948
rect -11132 32892 -10868 32948
rect -10812 32892 -10708 32948
rect -10652 32892 -10548 32948
rect -10492 32892 -10388 32948
rect -10332 32892 -10228 32948
rect -10172 32892 -10068 32948
rect -10012 32892 -9908 32948
rect -9852 32892 -9748 32948
rect -9692 32892 -9588 32948
rect -9532 32892 -9428 32948
rect -9372 32892 -9268 32948
rect -9212 32892 -9108 32948
rect -9052 32892 -8948 32948
rect -8892 32892 -8788 32948
rect -8732 32892 -8628 32948
rect -8572 32892 -8468 32948
rect -8412 32892 -8308 32948
rect -8252 32892 -8148 32948
rect -8092 32892 -7988 32948
rect -7932 32892 -7828 32948
rect -7772 32892 -7668 32948
rect -7612 32892 -7508 32948
rect -7452 32892 -7348 32948
rect -7292 32892 -7188 32948
rect -7132 32892 -7028 32948
rect -6972 32892 -6868 32948
rect -6812 32892 -6708 32948
rect -6652 32892 -6548 32948
rect -6492 32892 -6388 32948
rect -6332 32892 -6228 32948
rect -6172 32892 -6068 32948
rect -6012 32892 -5908 32948
rect -5852 32892 -5748 32948
rect -5692 32892 -5588 32948
rect -5532 32892 -5428 32948
rect -5372 32892 -5268 32948
rect -5212 32892 -5108 32948
rect -5052 32892 -4948 32948
rect -4892 32892 -4788 32948
rect -4732 32892 -4628 32948
rect -4572 32892 -4468 32948
rect -4412 32892 -4308 32948
rect -4252 32892 -4148 32948
rect -4092 32892 -3988 32948
rect -3932 32892 -3668 32948
rect -3612 32892 -3508 32948
rect -3452 32892 -3348 32948
rect -3292 32892 -3188 32948
rect -3132 32892 -3028 32948
rect -2972 32892 -2868 32948
rect -2812 32892 -2708 32948
rect -2652 32892 -2388 32948
rect -2332 32892 -2068 32948
rect -2012 32892 -1748 32948
rect -1692 32892 -1428 32948
rect -1372 32892 -1108 32948
rect -1052 32892 -1040 32948
rect -31040 32880 -1040 32892
rect -31040 32788 -30640 32800
rect -31040 32732 -31028 32788
rect -30972 32732 -30708 32788
rect -30652 32732 -30640 32788
rect -31040 32720 -30640 32732
rect -30560 32788 -1200 32800
rect -30560 32732 -30548 32788
rect -30492 32732 -1268 32788
rect -1212 32732 -1200 32788
rect -30560 32720 -1200 32732
rect -1120 32720 -1040 32800
rect -31040 32628 -1040 32640
rect -31040 32572 -31028 32628
rect -30972 32572 -30708 32628
rect -30652 32572 -30388 32628
rect -30332 32572 -30068 32628
rect -30012 32572 -29908 32628
rect -29852 32572 -29748 32628
rect -29692 32572 -29588 32628
rect -29532 32572 -29428 32628
rect -29372 32572 -29268 32628
rect -29212 32572 -29108 32628
rect -29052 32572 -28948 32628
rect -28892 32572 -28788 32628
rect -28732 32572 -28628 32628
rect -28572 32572 -28468 32628
rect -28412 32572 -28308 32628
rect -28252 32572 -28148 32628
rect -28092 32572 -27988 32628
rect -27932 32572 -27828 32628
rect -27772 32572 -27668 32628
rect -27612 32572 -27508 32628
rect -27452 32572 -27348 32628
rect -27292 32572 -27188 32628
rect -27132 32572 -27028 32628
rect -26972 32572 -26868 32628
rect -26812 32572 -26708 32628
rect -26652 32572 -26548 32628
rect -26492 32572 -26388 32628
rect -26332 32572 -26228 32628
rect -26172 32572 -26068 32628
rect -26012 32572 -25908 32628
rect -25852 32572 -25748 32628
rect -25692 32572 -25588 32628
rect -25532 32572 -25428 32628
rect -25372 32572 -25268 32628
rect -25212 32572 -25108 32628
rect -25052 32572 -24948 32628
rect -24892 32572 -24788 32628
rect -24732 32572 -24628 32628
rect -24572 32572 -24468 32628
rect -24412 32572 -24308 32628
rect -24252 32572 -24148 32628
rect -24092 32572 -23988 32628
rect -23932 32572 -23828 32628
rect -23772 32572 -23668 32628
rect -23612 32572 -23508 32628
rect -23452 32572 -23348 32628
rect -23292 32572 -23188 32628
rect -23132 32572 -23028 32628
rect -22972 32572 -22868 32628
rect -22812 32572 -22708 32628
rect -22652 32572 -22548 32628
rect -22492 32572 -22388 32628
rect -22332 32572 -22228 32628
rect -22172 32572 -22068 32628
rect -22012 32572 -21908 32628
rect -21852 32572 -21748 32628
rect -21692 32572 -21588 32628
rect -21532 32572 -21428 32628
rect -21372 32572 -21268 32628
rect -21212 32572 -21108 32628
rect -21052 32572 -20948 32628
rect -20892 32572 -20788 32628
rect -20732 32572 -20628 32628
rect -20572 32572 -20468 32628
rect -20412 32572 -20308 32628
rect -20252 32572 -20148 32628
rect -20092 32572 -19988 32628
rect -19932 32572 -19828 32628
rect -19772 32572 -19668 32628
rect -19612 32572 -19508 32628
rect -19452 32572 -19348 32628
rect -19292 32572 -19188 32628
rect -19132 32572 -19028 32628
rect -18972 32572 -18868 32628
rect -18812 32572 -18708 32628
rect -18652 32572 -18548 32628
rect -18492 32572 -18388 32628
rect -18332 32572 -18228 32628
rect -18172 32572 -18068 32628
rect -18012 32572 -17908 32628
rect -17852 32572 -17748 32628
rect -17692 32572 -17588 32628
rect -17532 32572 -17428 32628
rect -17372 32572 -17268 32628
rect -17212 32572 -17108 32628
rect -17052 32572 -16948 32628
rect -16892 32572 -16788 32628
rect -16732 32572 -16628 32628
rect -16572 32572 -16468 32628
rect -16412 32572 -16308 32628
rect -16252 32572 -16148 32628
rect -16092 32572 -15988 32628
rect -15932 32572 -15828 32628
rect -15772 32572 -15668 32628
rect -15612 32572 -15508 32628
rect -15452 32572 -15348 32628
rect -15292 32572 -15188 32628
rect -15132 32572 -15028 32628
rect -14972 32572 -14868 32628
rect -14812 32572 -14708 32628
rect -14652 32572 -14548 32628
rect -14492 32572 -14388 32628
rect -14332 32572 -14228 32628
rect -14172 32572 -14068 32628
rect -14012 32572 -13908 32628
rect -13852 32572 -13748 32628
rect -13692 32572 -13588 32628
rect -13532 32572 -13428 32628
rect -13372 32572 -13268 32628
rect -13212 32572 -13108 32628
rect -13052 32572 -12948 32628
rect -12892 32572 -12788 32628
rect -12732 32572 -12628 32628
rect -12572 32572 -12468 32628
rect -12412 32572 -12308 32628
rect -12252 32572 -12148 32628
rect -12092 32572 -11988 32628
rect -11932 32572 -11828 32628
rect -11772 32572 -11668 32628
rect -11612 32572 -11508 32628
rect -11452 32572 -11188 32628
rect -11132 32572 -10868 32628
rect -10812 32572 -10708 32628
rect -10652 32572 -10548 32628
rect -10492 32572 -10388 32628
rect -10332 32572 -10228 32628
rect -10172 32572 -10068 32628
rect -10012 32572 -9908 32628
rect -9852 32572 -9748 32628
rect -9692 32572 -9588 32628
rect -9532 32572 -9428 32628
rect -9372 32572 -9268 32628
rect -9212 32572 -9108 32628
rect -9052 32572 -8948 32628
rect -8892 32572 -8788 32628
rect -8732 32572 -8628 32628
rect -8572 32572 -8468 32628
rect -8412 32572 -8308 32628
rect -8252 32572 -8148 32628
rect -8092 32572 -7988 32628
rect -7932 32572 -7828 32628
rect -7772 32572 -7668 32628
rect -7612 32572 -7508 32628
rect -7452 32572 -7348 32628
rect -7292 32572 -7188 32628
rect -7132 32572 -7028 32628
rect -6972 32572 -6868 32628
rect -6812 32572 -6708 32628
rect -6652 32572 -6548 32628
rect -6492 32572 -6388 32628
rect -6332 32572 -6228 32628
rect -6172 32572 -6068 32628
rect -6012 32572 -5908 32628
rect -5852 32572 -5748 32628
rect -5692 32572 -5588 32628
rect -5532 32572 -5428 32628
rect -5372 32572 -5268 32628
rect -5212 32572 -5108 32628
rect -5052 32572 -4948 32628
rect -4892 32572 -4788 32628
rect -4732 32572 -4628 32628
rect -4572 32572 -4468 32628
rect -4412 32572 -4308 32628
rect -4252 32572 -4148 32628
rect -4092 32572 -3988 32628
rect -3932 32572 -3668 32628
rect -3612 32572 -3508 32628
rect -3452 32572 -3348 32628
rect -3292 32572 -3188 32628
rect -3132 32572 -3028 32628
rect -2972 32572 -2868 32628
rect -2812 32572 -2708 32628
rect -2652 32572 -2388 32628
rect -2332 32572 -2068 32628
rect -2012 32572 -1748 32628
rect -1692 32572 -1428 32628
rect -1372 32572 -1108 32628
rect -1052 32572 -1040 32628
rect -31040 32560 -1040 32572
rect -31040 32468 -30320 32480
rect -31040 32412 -31028 32468
rect -30972 32412 -30708 32468
rect -30652 32412 -30320 32468
rect -31040 32400 -30320 32412
rect -30240 32468 -2480 32480
rect -30240 32412 -30228 32468
rect -30172 32412 -11348 32468
rect -11292 32412 -2548 32468
rect -2492 32412 -2480 32468
rect -30240 32400 -2480 32412
rect -2400 32400 -2320 32480
rect -2080 32400 -2000 32480
rect -1760 32400 -1680 32480
rect -1440 32400 -1360 32480
rect -1120 32400 -1040 32480
rect -31040 32308 -1040 32320
rect -31040 32252 -31028 32308
rect -30972 32252 -30708 32308
rect -30652 32252 -30388 32308
rect -30332 32252 -30068 32308
rect -30012 32252 -29908 32308
rect -29852 32252 -29748 32308
rect -29692 32252 -29588 32308
rect -29532 32252 -29428 32308
rect -29372 32252 -29268 32308
rect -29212 32252 -29108 32308
rect -29052 32252 -28948 32308
rect -28892 32252 -28788 32308
rect -28732 32252 -28628 32308
rect -28572 32252 -28468 32308
rect -28412 32252 -28308 32308
rect -28252 32252 -28148 32308
rect -28092 32252 -27988 32308
rect -27932 32252 -27828 32308
rect -27772 32252 -27668 32308
rect -27612 32252 -27508 32308
rect -27452 32252 -27348 32308
rect -27292 32252 -27188 32308
rect -27132 32252 -27028 32308
rect -26972 32252 -26868 32308
rect -26812 32252 -26708 32308
rect -26652 32252 -26548 32308
rect -26492 32252 -26388 32308
rect -26332 32252 -26228 32308
rect -26172 32252 -26068 32308
rect -26012 32252 -25908 32308
rect -25852 32252 -25748 32308
rect -25692 32252 -25588 32308
rect -25532 32252 -25428 32308
rect -25372 32252 -25268 32308
rect -25212 32252 -25108 32308
rect -25052 32252 -24948 32308
rect -24892 32252 -24788 32308
rect -24732 32252 -24628 32308
rect -24572 32252 -24468 32308
rect -24412 32252 -24308 32308
rect -24252 32252 -24148 32308
rect -24092 32252 -23988 32308
rect -23932 32252 -23828 32308
rect -23772 32252 -23668 32308
rect -23612 32252 -23508 32308
rect -23452 32252 -23348 32308
rect -23292 32252 -23188 32308
rect -23132 32252 -23028 32308
rect -22972 32252 -22868 32308
rect -22812 32252 -22708 32308
rect -22652 32252 -22548 32308
rect -22492 32252 -22388 32308
rect -22332 32252 -22228 32308
rect -22172 32252 -22068 32308
rect -22012 32252 -21908 32308
rect -21852 32252 -21748 32308
rect -21692 32252 -21588 32308
rect -21532 32252 -21428 32308
rect -21372 32252 -21268 32308
rect -21212 32252 -21108 32308
rect -21052 32252 -20948 32308
rect -20892 32252 -20788 32308
rect -20732 32252 -20628 32308
rect -20572 32252 -20468 32308
rect -20412 32252 -20308 32308
rect -20252 32252 -20148 32308
rect -20092 32252 -19988 32308
rect -19932 32252 -19828 32308
rect -19772 32252 -19668 32308
rect -19612 32252 -19508 32308
rect -19452 32252 -19348 32308
rect -19292 32252 -19188 32308
rect -19132 32252 -19028 32308
rect -18972 32252 -18868 32308
rect -18812 32252 -18708 32308
rect -18652 32252 -18548 32308
rect -18492 32252 -18388 32308
rect -18332 32252 -18228 32308
rect -18172 32252 -18068 32308
rect -18012 32252 -17908 32308
rect -17852 32252 -17748 32308
rect -17692 32252 -17588 32308
rect -17532 32252 -17428 32308
rect -17372 32252 -17268 32308
rect -17212 32252 -17108 32308
rect -17052 32252 -16948 32308
rect -16892 32252 -16788 32308
rect -16732 32252 -16628 32308
rect -16572 32252 -16468 32308
rect -16412 32252 -16308 32308
rect -16252 32252 -16148 32308
rect -16092 32252 -15988 32308
rect -15932 32252 -15828 32308
rect -15772 32252 -15668 32308
rect -15612 32252 -15508 32308
rect -15452 32252 -15348 32308
rect -15292 32252 -15188 32308
rect -15132 32252 -15028 32308
rect -14972 32252 -14868 32308
rect -14812 32252 -14708 32308
rect -14652 32252 -14548 32308
rect -14492 32252 -14388 32308
rect -14332 32252 -14228 32308
rect -14172 32252 -14068 32308
rect -14012 32252 -13908 32308
rect -13852 32252 -13748 32308
rect -13692 32252 -13588 32308
rect -13532 32252 -13428 32308
rect -13372 32252 -13268 32308
rect -13212 32252 -13108 32308
rect -13052 32252 -12948 32308
rect -12892 32252 -12788 32308
rect -12732 32252 -12628 32308
rect -12572 32252 -12468 32308
rect -12412 32252 -12308 32308
rect -12252 32252 -12148 32308
rect -12092 32252 -11988 32308
rect -11932 32252 -11828 32308
rect -11772 32252 -11668 32308
rect -11612 32252 -11508 32308
rect -11452 32252 -11348 32308
rect -11292 32252 -11188 32308
rect -11132 32252 -10868 32308
rect -10812 32252 -10708 32308
rect -10652 32252 -10548 32308
rect -10492 32252 -10388 32308
rect -10332 32252 -10228 32308
rect -10172 32252 -10068 32308
rect -10012 32252 -9908 32308
rect -9852 32252 -9748 32308
rect -9692 32252 -9588 32308
rect -9532 32252 -9428 32308
rect -9372 32252 -9268 32308
rect -9212 32252 -9108 32308
rect -9052 32252 -8948 32308
rect -8892 32252 -8788 32308
rect -8732 32252 -8628 32308
rect -8572 32252 -8468 32308
rect -8412 32252 -8308 32308
rect -8252 32252 -8148 32308
rect -8092 32252 -7988 32308
rect -7932 32252 -7828 32308
rect -7772 32252 -7668 32308
rect -7612 32252 -7508 32308
rect -7452 32252 -7348 32308
rect -7292 32252 -7188 32308
rect -7132 32252 -7028 32308
rect -6972 32252 -6868 32308
rect -6812 32252 -6708 32308
rect -6652 32252 -6548 32308
rect -6492 32252 -6388 32308
rect -6332 32252 -6228 32308
rect -6172 32252 -6068 32308
rect -6012 32252 -5908 32308
rect -5852 32252 -5748 32308
rect -5692 32252 -5588 32308
rect -5532 32252 -5428 32308
rect -5372 32252 -5268 32308
rect -5212 32252 -5108 32308
rect -5052 32252 -4948 32308
rect -4892 32252 -4788 32308
rect -4732 32252 -4628 32308
rect -4572 32252 -4468 32308
rect -4412 32252 -4308 32308
rect -4252 32252 -4148 32308
rect -4092 32252 -3988 32308
rect -3932 32252 -3668 32308
rect -3612 32252 -3508 32308
rect -3452 32252 -3348 32308
rect -3292 32252 -3188 32308
rect -3132 32252 -3028 32308
rect -2972 32252 -2868 32308
rect -2812 32252 -2708 32308
rect -2652 32252 -2388 32308
rect -2332 32252 -2068 32308
rect -2012 32252 -1748 32308
rect -1692 32252 -1428 32308
rect -1372 32252 -1108 32308
rect -1052 32252 -1040 32308
rect -31040 32240 -1040 32252
rect -31040 32148 -30640 32160
rect -31040 32092 -31028 32148
rect -30972 32092 -30708 32148
rect -30652 32092 -30640 32148
rect -31040 32080 -30640 32092
rect -30560 32148 -2160 32160
rect -30560 32092 -30548 32148
rect -30492 32092 -11028 32148
rect -10972 32092 -2228 32148
rect -2172 32092 -2160 32148
rect -30560 32080 -2160 32092
rect -2080 32080 -2000 32160
rect -1760 32080 -1680 32160
rect -1440 32080 -1360 32160
rect -1120 32080 -1040 32160
rect -31040 31988 -1040 32000
rect -31040 31932 -31028 31988
rect -30972 31932 -30708 31988
rect -30652 31932 -30388 31988
rect -30332 31932 -30068 31988
rect -30012 31932 -29908 31988
rect -29852 31932 -29748 31988
rect -29692 31932 -29588 31988
rect -29532 31932 -29428 31988
rect -29372 31932 -29268 31988
rect -29212 31932 -29108 31988
rect -29052 31932 -28948 31988
rect -28892 31932 -28788 31988
rect -28732 31932 -28628 31988
rect -28572 31932 -28468 31988
rect -28412 31932 -28308 31988
rect -28252 31932 -28148 31988
rect -28092 31932 -27988 31988
rect -27932 31932 -27828 31988
rect -27772 31932 -27668 31988
rect -27612 31932 -27508 31988
rect -27452 31932 -27348 31988
rect -27292 31932 -27188 31988
rect -27132 31932 -27028 31988
rect -26972 31932 -26868 31988
rect -26812 31932 -26708 31988
rect -26652 31932 -26548 31988
rect -26492 31932 -26388 31988
rect -26332 31932 -26228 31988
rect -26172 31932 -26068 31988
rect -26012 31932 -25908 31988
rect -25852 31932 -25748 31988
rect -25692 31932 -25588 31988
rect -25532 31932 -25428 31988
rect -25372 31932 -25268 31988
rect -25212 31932 -25108 31988
rect -25052 31932 -24948 31988
rect -24892 31932 -24788 31988
rect -24732 31932 -24628 31988
rect -24572 31932 -24468 31988
rect -24412 31932 -24308 31988
rect -24252 31932 -24148 31988
rect -24092 31932 -23988 31988
rect -23932 31932 -23828 31988
rect -23772 31932 -23668 31988
rect -23612 31932 -23508 31988
rect -23452 31932 -23348 31988
rect -23292 31932 -23188 31988
rect -23132 31932 -23028 31988
rect -22972 31932 -22868 31988
rect -22812 31932 -22708 31988
rect -22652 31932 -22548 31988
rect -22492 31932 -22388 31988
rect -22332 31932 -22228 31988
rect -22172 31932 -22068 31988
rect -22012 31932 -21908 31988
rect -21852 31932 -21748 31988
rect -21692 31932 -21588 31988
rect -21532 31932 -21428 31988
rect -21372 31932 -21268 31988
rect -21212 31932 -21108 31988
rect -21052 31932 -20948 31988
rect -20892 31932 -20788 31988
rect -20732 31932 -20628 31988
rect -20572 31932 -20468 31988
rect -20412 31932 -20308 31988
rect -20252 31932 -20148 31988
rect -20092 31932 -19988 31988
rect -19932 31932 -19828 31988
rect -19772 31932 -19668 31988
rect -19612 31932 -19508 31988
rect -19452 31932 -19348 31988
rect -19292 31932 -19188 31988
rect -19132 31932 -19028 31988
rect -18972 31932 -18868 31988
rect -18812 31932 -18708 31988
rect -18652 31932 -18548 31988
rect -18492 31932 -18388 31988
rect -18332 31932 -18228 31988
rect -18172 31932 -18068 31988
rect -18012 31932 -17908 31988
rect -17852 31932 -17748 31988
rect -17692 31932 -17588 31988
rect -17532 31932 -17428 31988
rect -17372 31932 -17268 31988
rect -17212 31932 -17108 31988
rect -17052 31932 -16948 31988
rect -16892 31932 -16788 31988
rect -16732 31932 -16628 31988
rect -16572 31932 -16468 31988
rect -16412 31932 -16308 31988
rect -16252 31932 -16148 31988
rect -16092 31932 -15988 31988
rect -15932 31932 -15828 31988
rect -15772 31932 -15668 31988
rect -15612 31932 -15508 31988
rect -15452 31932 -15348 31988
rect -15292 31932 -15188 31988
rect -15132 31932 -15028 31988
rect -14972 31932 -14868 31988
rect -14812 31932 -14708 31988
rect -14652 31932 -14548 31988
rect -14492 31932 -14388 31988
rect -14332 31932 -14228 31988
rect -14172 31932 -14068 31988
rect -14012 31932 -13908 31988
rect -13852 31932 -13748 31988
rect -13692 31932 -13588 31988
rect -13532 31932 -13428 31988
rect -13372 31932 -13268 31988
rect -13212 31932 -13108 31988
rect -13052 31932 -12948 31988
rect -12892 31932 -12788 31988
rect -12732 31932 -12628 31988
rect -12572 31932 -12468 31988
rect -12412 31932 -12308 31988
rect -12252 31932 -12148 31988
rect -12092 31932 -11988 31988
rect -11932 31932 -11828 31988
rect -11772 31932 -11668 31988
rect -11612 31932 -11508 31988
rect -11452 31932 -11348 31988
rect -11292 31932 -11188 31988
rect -11132 31932 -10868 31988
rect -10812 31932 -10708 31988
rect -10652 31932 -10548 31988
rect -10492 31932 -10388 31988
rect -10332 31932 -10228 31988
rect -10172 31932 -10068 31988
rect -10012 31932 -9908 31988
rect -9852 31932 -9748 31988
rect -9692 31932 -9588 31988
rect -9532 31932 -9428 31988
rect -9372 31932 -9268 31988
rect -9212 31932 -9108 31988
rect -9052 31932 -8948 31988
rect -8892 31932 -8788 31988
rect -8732 31932 -8628 31988
rect -8572 31932 -8468 31988
rect -8412 31932 -8308 31988
rect -8252 31932 -8148 31988
rect -8092 31932 -7988 31988
rect -7932 31932 -7828 31988
rect -7772 31932 -7668 31988
rect -7612 31932 -7508 31988
rect -7452 31932 -7348 31988
rect -7292 31932 -7188 31988
rect -7132 31932 -7028 31988
rect -6972 31932 -6868 31988
rect -6812 31932 -6708 31988
rect -6652 31932 -6548 31988
rect -6492 31932 -6388 31988
rect -6332 31932 -6228 31988
rect -6172 31932 -6068 31988
rect -6012 31932 -5908 31988
rect -5852 31932 -5748 31988
rect -5692 31932 -5588 31988
rect -5532 31932 -5428 31988
rect -5372 31932 -5268 31988
rect -5212 31932 -5108 31988
rect -5052 31932 -4948 31988
rect -4892 31932 -4788 31988
rect -4732 31932 -4628 31988
rect -4572 31932 -4468 31988
rect -4412 31932 -4308 31988
rect -4252 31932 -4148 31988
rect -4092 31932 -3988 31988
rect -3932 31932 -3668 31988
rect -3612 31932 -3508 31988
rect -3452 31932 -3348 31988
rect -3292 31932 -3188 31988
rect -3132 31932 -3028 31988
rect -2972 31932 -2868 31988
rect -2812 31932 -2708 31988
rect -2652 31932 -2388 31988
rect -2332 31932 -2068 31988
rect -2012 31932 -1748 31988
rect -1692 31932 -1428 31988
rect -1372 31932 -1108 31988
rect -1052 31932 -1040 31988
rect -31040 31920 -1040 31932
<< via2 >>
rect -31028 42812 -30972 42868
rect -30708 42812 -30652 42868
rect -30388 42812 -30332 42868
rect -30068 42812 -30012 42868
rect -29908 42866 -29852 42868
rect -29908 42814 -29906 42866
rect -29906 42814 -29854 42866
rect -29854 42814 -29852 42866
rect -29908 42812 -29852 42814
rect -29748 42866 -29692 42868
rect -29748 42814 -29746 42866
rect -29746 42814 -29694 42866
rect -29694 42814 -29692 42866
rect -29748 42812 -29692 42814
rect -29588 42866 -29532 42868
rect -29588 42814 -29586 42866
rect -29586 42814 -29534 42866
rect -29534 42814 -29532 42866
rect -29588 42812 -29532 42814
rect -29428 42866 -29372 42868
rect -29428 42814 -29426 42866
rect -29426 42814 -29374 42866
rect -29374 42814 -29372 42866
rect -29428 42812 -29372 42814
rect -29268 42866 -29212 42868
rect -29268 42814 -29266 42866
rect -29266 42814 -29214 42866
rect -29214 42814 -29212 42866
rect -29268 42812 -29212 42814
rect -29108 42866 -29052 42868
rect -29108 42814 -29106 42866
rect -29106 42814 -29054 42866
rect -29054 42814 -29052 42866
rect -29108 42812 -29052 42814
rect -28948 42866 -28892 42868
rect -28948 42814 -28946 42866
rect -28946 42814 -28894 42866
rect -28894 42814 -28892 42866
rect -28948 42812 -28892 42814
rect -28788 42866 -28732 42868
rect -28788 42814 -28786 42866
rect -28786 42814 -28734 42866
rect -28734 42814 -28732 42866
rect -28788 42812 -28732 42814
rect -28628 42866 -28572 42868
rect -28628 42814 -28626 42866
rect -28626 42814 -28574 42866
rect -28574 42814 -28572 42866
rect -28628 42812 -28572 42814
rect -28468 42866 -28412 42868
rect -28468 42814 -28466 42866
rect -28466 42814 -28414 42866
rect -28414 42814 -28412 42866
rect -28468 42812 -28412 42814
rect -28308 42866 -28252 42868
rect -28308 42814 -28306 42866
rect -28306 42814 -28254 42866
rect -28254 42814 -28252 42866
rect -28308 42812 -28252 42814
rect -28148 42866 -28092 42868
rect -28148 42814 -28146 42866
rect -28146 42814 -28094 42866
rect -28094 42814 -28092 42866
rect -28148 42812 -28092 42814
rect -27988 42866 -27932 42868
rect -27988 42814 -27986 42866
rect -27986 42814 -27934 42866
rect -27934 42814 -27932 42866
rect -27988 42812 -27932 42814
rect -27828 42866 -27772 42868
rect -27828 42814 -27826 42866
rect -27826 42814 -27774 42866
rect -27774 42814 -27772 42866
rect -27828 42812 -27772 42814
rect -27668 42866 -27612 42868
rect -27668 42814 -27666 42866
rect -27666 42814 -27614 42866
rect -27614 42814 -27612 42866
rect -27668 42812 -27612 42814
rect -27508 42866 -27452 42868
rect -27508 42814 -27506 42866
rect -27506 42814 -27454 42866
rect -27454 42814 -27452 42866
rect -27508 42812 -27452 42814
rect -27348 42866 -27292 42868
rect -27348 42814 -27346 42866
rect -27346 42814 -27294 42866
rect -27294 42814 -27292 42866
rect -27348 42812 -27292 42814
rect -27188 42866 -27132 42868
rect -27188 42814 -27186 42866
rect -27186 42814 -27134 42866
rect -27134 42814 -27132 42866
rect -27188 42812 -27132 42814
rect -27028 42866 -26972 42868
rect -27028 42814 -27026 42866
rect -27026 42814 -26974 42866
rect -26974 42814 -26972 42866
rect -27028 42812 -26972 42814
rect -26868 42866 -26812 42868
rect -26868 42814 -26866 42866
rect -26866 42814 -26814 42866
rect -26814 42814 -26812 42866
rect -26868 42812 -26812 42814
rect -26708 42866 -26652 42868
rect -26708 42814 -26706 42866
rect -26706 42814 -26654 42866
rect -26654 42814 -26652 42866
rect -26708 42812 -26652 42814
rect -26548 42866 -26492 42868
rect -26548 42814 -26546 42866
rect -26546 42814 -26494 42866
rect -26494 42814 -26492 42866
rect -26548 42812 -26492 42814
rect -26388 42866 -26332 42868
rect -26388 42814 -26386 42866
rect -26386 42814 -26334 42866
rect -26334 42814 -26332 42866
rect -26388 42812 -26332 42814
rect -26228 42866 -26172 42868
rect -26228 42814 -26226 42866
rect -26226 42814 -26174 42866
rect -26174 42814 -26172 42866
rect -26228 42812 -26172 42814
rect -26068 42866 -26012 42868
rect -26068 42814 -26066 42866
rect -26066 42814 -26014 42866
rect -26014 42814 -26012 42866
rect -26068 42812 -26012 42814
rect -25908 42866 -25852 42868
rect -25908 42814 -25906 42866
rect -25906 42814 -25854 42866
rect -25854 42814 -25852 42866
rect -25908 42812 -25852 42814
rect -25748 42866 -25692 42868
rect -25748 42814 -25746 42866
rect -25746 42814 -25694 42866
rect -25694 42814 -25692 42866
rect -25748 42812 -25692 42814
rect -25588 42866 -25532 42868
rect -25588 42814 -25586 42866
rect -25586 42814 -25534 42866
rect -25534 42814 -25532 42866
rect -25588 42812 -25532 42814
rect -25428 42866 -25372 42868
rect -25428 42814 -25426 42866
rect -25426 42814 -25374 42866
rect -25374 42814 -25372 42866
rect -25428 42812 -25372 42814
rect -25268 42866 -25212 42868
rect -25268 42814 -25266 42866
rect -25266 42814 -25214 42866
rect -25214 42814 -25212 42866
rect -25268 42812 -25212 42814
rect -25108 42866 -25052 42868
rect -25108 42814 -25106 42866
rect -25106 42814 -25054 42866
rect -25054 42814 -25052 42866
rect -25108 42812 -25052 42814
rect -24948 42866 -24892 42868
rect -24948 42814 -24946 42866
rect -24946 42814 -24894 42866
rect -24894 42814 -24892 42866
rect -24948 42812 -24892 42814
rect -24788 42866 -24732 42868
rect -24788 42814 -24786 42866
rect -24786 42814 -24734 42866
rect -24734 42814 -24732 42866
rect -24788 42812 -24732 42814
rect -24628 42866 -24572 42868
rect -24628 42814 -24626 42866
rect -24626 42814 -24574 42866
rect -24574 42814 -24572 42866
rect -24628 42812 -24572 42814
rect -24468 42866 -24412 42868
rect -24468 42814 -24466 42866
rect -24466 42814 -24414 42866
rect -24414 42814 -24412 42866
rect -24468 42812 -24412 42814
rect -24308 42866 -24252 42868
rect -24308 42814 -24306 42866
rect -24306 42814 -24254 42866
rect -24254 42814 -24252 42866
rect -24308 42812 -24252 42814
rect -24148 42866 -24092 42868
rect -24148 42814 -24146 42866
rect -24146 42814 -24094 42866
rect -24094 42814 -24092 42866
rect -24148 42812 -24092 42814
rect -23988 42866 -23932 42868
rect -23988 42814 -23986 42866
rect -23986 42814 -23934 42866
rect -23934 42814 -23932 42866
rect -23988 42812 -23932 42814
rect -23828 42866 -23772 42868
rect -23828 42814 -23826 42866
rect -23826 42814 -23774 42866
rect -23774 42814 -23772 42866
rect -23828 42812 -23772 42814
rect -23668 42866 -23612 42868
rect -23668 42814 -23666 42866
rect -23666 42814 -23614 42866
rect -23614 42814 -23612 42866
rect -23668 42812 -23612 42814
rect -23508 42866 -23452 42868
rect -23508 42814 -23506 42866
rect -23506 42814 -23454 42866
rect -23454 42814 -23452 42866
rect -23508 42812 -23452 42814
rect -23348 42866 -23292 42868
rect -23348 42814 -23346 42866
rect -23346 42814 -23294 42866
rect -23294 42814 -23292 42866
rect -23348 42812 -23292 42814
rect -23188 42866 -23132 42868
rect -23188 42814 -23186 42866
rect -23186 42814 -23134 42866
rect -23134 42814 -23132 42866
rect -23188 42812 -23132 42814
rect -23028 42866 -22972 42868
rect -23028 42814 -23026 42866
rect -23026 42814 -22974 42866
rect -22974 42814 -22972 42866
rect -23028 42812 -22972 42814
rect -22868 42866 -22812 42868
rect -22868 42814 -22866 42866
rect -22866 42814 -22814 42866
rect -22814 42814 -22812 42866
rect -22868 42812 -22812 42814
rect -22708 42866 -22652 42868
rect -22708 42814 -22706 42866
rect -22706 42814 -22654 42866
rect -22654 42814 -22652 42866
rect -22708 42812 -22652 42814
rect -22548 42866 -22492 42868
rect -22548 42814 -22546 42866
rect -22546 42814 -22494 42866
rect -22494 42814 -22492 42866
rect -22548 42812 -22492 42814
rect -22388 42866 -22332 42868
rect -22388 42814 -22386 42866
rect -22386 42814 -22334 42866
rect -22334 42814 -22332 42866
rect -22388 42812 -22332 42814
rect -22228 42866 -22172 42868
rect -22228 42814 -22226 42866
rect -22226 42814 -22174 42866
rect -22174 42814 -22172 42866
rect -22228 42812 -22172 42814
rect -22068 42866 -22012 42868
rect -22068 42814 -22066 42866
rect -22066 42814 -22014 42866
rect -22014 42814 -22012 42866
rect -22068 42812 -22012 42814
rect -21908 42866 -21852 42868
rect -21908 42814 -21906 42866
rect -21906 42814 -21854 42866
rect -21854 42814 -21852 42866
rect -21908 42812 -21852 42814
rect -21748 42866 -21692 42868
rect -21748 42814 -21746 42866
rect -21746 42814 -21694 42866
rect -21694 42814 -21692 42866
rect -21748 42812 -21692 42814
rect -21588 42866 -21532 42868
rect -21588 42814 -21586 42866
rect -21586 42814 -21534 42866
rect -21534 42814 -21532 42866
rect -21588 42812 -21532 42814
rect -21428 42866 -21372 42868
rect -21428 42814 -21426 42866
rect -21426 42814 -21374 42866
rect -21374 42814 -21372 42866
rect -21428 42812 -21372 42814
rect -21268 42866 -21212 42868
rect -21268 42814 -21266 42866
rect -21266 42814 -21214 42866
rect -21214 42814 -21212 42866
rect -21268 42812 -21212 42814
rect -21108 42866 -21052 42868
rect -21108 42814 -21106 42866
rect -21106 42814 -21054 42866
rect -21054 42814 -21052 42866
rect -21108 42812 -21052 42814
rect -20948 42866 -20892 42868
rect -20948 42814 -20946 42866
rect -20946 42814 -20894 42866
rect -20894 42814 -20892 42866
rect -20948 42812 -20892 42814
rect -20788 42866 -20732 42868
rect -20788 42814 -20786 42866
rect -20786 42814 -20734 42866
rect -20734 42814 -20732 42866
rect -20788 42812 -20732 42814
rect -20628 42866 -20572 42868
rect -20628 42814 -20626 42866
rect -20626 42814 -20574 42866
rect -20574 42814 -20572 42866
rect -20628 42812 -20572 42814
rect -20468 42866 -20412 42868
rect -20468 42814 -20466 42866
rect -20466 42814 -20414 42866
rect -20414 42814 -20412 42866
rect -20468 42812 -20412 42814
rect -20308 42866 -20252 42868
rect -20308 42814 -20306 42866
rect -20306 42814 -20254 42866
rect -20254 42814 -20252 42866
rect -20308 42812 -20252 42814
rect -20148 42866 -20092 42868
rect -20148 42814 -20146 42866
rect -20146 42814 -20094 42866
rect -20094 42814 -20092 42866
rect -20148 42812 -20092 42814
rect -19988 42866 -19932 42868
rect -19988 42814 -19986 42866
rect -19986 42814 -19934 42866
rect -19934 42814 -19932 42866
rect -19988 42812 -19932 42814
rect -19828 42866 -19772 42868
rect -19828 42814 -19826 42866
rect -19826 42814 -19774 42866
rect -19774 42814 -19772 42866
rect -19828 42812 -19772 42814
rect -19668 42866 -19612 42868
rect -19668 42814 -19666 42866
rect -19666 42814 -19614 42866
rect -19614 42814 -19612 42866
rect -19668 42812 -19612 42814
rect -19508 42866 -19452 42868
rect -19508 42814 -19506 42866
rect -19506 42814 -19454 42866
rect -19454 42814 -19452 42866
rect -19508 42812 -19452 42814
rect -19348 42866 -19292 42868
rect -19348 42814 -19346 42866
rect -19346 42814 -19294 42866
rect -19294 42814 -19292 42866
rect -19348 42812 -19292 42814
rect -19188 42866 -19132 42868
rect -19188 42814 -19186 42866
rect -19186 42814 -19134 42866
rect -19134 42814 -19132 42866
rect -19188 42812 -19132 42814
rect -19028 42866 -18972 42868
rect -19028 42814 -19026 42866
rect -19026 42814 -18974 42866
rect -18974 42814 -18972 42866
rect -19028 42812 -18972 42814
rect -18868 42866 -18812 42868
rect -18868 42814 -18866 42866
rect -18866 42814 -18814 42866
rect -18814 42814 -18812 42866
rect -18868 42812 -18812 42814
rect -18708 42866 -18652 42868
rect -18708 42814 -18706 42866
rect -18706 42814 -18654 42866
rect -18654 42814 -18652 42866
rect -18708 42812 -18652 42814
rect -18548 42866 -18492 42868
rect -18548 42814 -18546 42866
rect -18546 42814 -18494 42866
rect -18494 42814 -18492 42866
rect -18548 42812 -18492 42814
rect -18388 42866 -18332 42868
rect -18388 42814 -18386 42866
rect -18386 42814 -18334 42866
rect -18334 42814 -18332 42866
rect -18388 42812 -18332 42814
rect -18228 42866 -18172 42868
rect -18228 42814 -18226 42866
rect -18226 42814 -18174 42866
rect -18174 42814 -18172 42866
rect -18228 42812 -18172 42814
rect -18068 42866 -18012 42868
rect -18068 42814 -18066 42866
rect -18066 42814 -18014 42866
rect -18014 42814 -18012 42866
rect -18068 42812 -18012 42814
rect -17908 42866 -17852 42868
rect -17908 42814 -17906 42866
rect -17906 42814 -17854 42866
rect -17854 42814 -17852 42866
rect -17908 42812 -17852 42814
rect -17748 42866 -17692 42868
rect -17748 42814 -17746 42866
rect -17746 42814 -17694 42866
rect -17694 42814 -17692 42866
rect -17748 42812 -17692 42814
rect -17588 42866 -17532 42868
rect -17588 42814 -17586 42866
rect -17586 42814 -17534 42866
rect -17534 42814 -17532 42866
rect -17588 42812 -17532 42814
rect -17428 42866 -17372 42868
rect -17428 42814 -17426 42866
rect -17426 42814 -17374 42866
rect -17374 42814 -17372 42866
rect -17428 42812 -17372 42814
rect -17268 42866 -17212 42868
rect -17268 42814 -17266 42866
rect -17266 42814 -17214 42866
rect -17214 42814 -17212 42866
rect -17268 42812 -17212 42814
rect -17108 42866 -17052 42868
rect -17108 42814 -17106 42866
rect -17106 42814 -17054 42866
rect -17054 42814 -17052 42866
rect -17108 42812 -17052 42814
rect -16948 42866 -16892 42868
rect -16948 42814 -16946 42866
rect -16946 42814 -16894 42866
rect -16894 42814 -16892 42866
rect -16948 42812 -16892 42814
rect -16788 42866 -16732 42868
rect -16788 42814 -16786 42866
rect -16786 42814 -16734 42866
rect -16734 42814 -16732 42866
rect -16788 42812 -16732 42814
rect -16628 42866 -16572 42868
rect -16628 42814 -16626 42866
rect -16626 42814 -16574 42866
rect -16574 42814 -16572 42866
rect -16628 42812 -16572 42814
rect -16468 42866 -16412 42868
rect -16468 42814 -16466 42866
rect -16466 42814 -16414 42866
rect -16414 42814 -16412 42866
rect -16468 42812 -16412 42814
rect -16308 42866 -16252 42868
rect -16308 42814 -16306 42866
rect -16306 42814 -16254 42866
rect -16254 42814 -16252 42866
rect -16308 42812 -16252 42814
rect -16148 42866 -16092 42868
rect -16148 42814 -16146 42866
rect -16146 42814 -16094 42866
rect -16094 42814 -16092 42866
rect -16148 42812 -16092 42814
rect -15988 42866 -15932 42868
rect -15988 42814 -15986 42866
rect -15986 42814 -15934 42866
rect -15934 42814 -15932 42866
rect -15988 42812 -15932 42814
rect -15828 42866 -15772 42868
rect -15828 42814 -15826 42866
rect -15826 42814 -15774 42866
rect -15774 42814 -15772 42866
rect -15828 42812 -15772 42814
rect -15668 42866 -15612 42868
rect -15668 42814 -15666 42866
rect -15666 42814 -15614 42866
rect -15614 42814 -15612 42866
rect -15668 42812 -15612 42814
rect -15508 42866 -15452 42868
rect -15508 42814 -15506 42866
rect -15506 42814 -15454 42866
rect -15454 42814 -15452 42866
rect -15508 42812 -15452 42814
rect -15348 42866 -15292 42868
rect -15348 42814 -15346 42866
rect -15346 42814 -15294 42866
rect -15294 42814 -15292 42866
rect -15348 42812 -15292 42814
rect -15188 42866 -15132 42868
rect -15188 42814 -15186 42866
rect -15186 42814 -15134 42866
rect -15134 42814 -15132 42866
rect -15188 42812 -15132 42814
rect -15028 42866 -14972 42868
rect -15028 42814 -15026 42866
rect -15026 42814 -14974 42866
rect -14974 42814 -14972 42866
rect -15028 42812 -14972 42814
rect -14868 42866 -14812 42868
rect -14868 42814 -14866 42866
rect -14866 42814 -14814 42866
rect -14814 42814 -14812 42866
rect -14868 42812 -14812 42814
rect -14708 42866 -14652 42868
rect -14708 42814 -14706 42866
rect -14706 42814 -14654 42866
rect -14654 42814 -14652 42866
rect -14708 42812 -14652 42814
rect -14548 42866 -14492 42868
rect -14548 42814 -14546 42866
rect -14546 42814 -14494 42866
rect -14494 42814 -14492 42866
rect -14548 42812 -14492 42814
rect -14388 42866 -14332 42868
rect -14388 42814 -14386 42866
rect -14386 42814 -14334 42866
rect -14334 42814 -14332 42866
rect -14388 42812 -14332 42814
rect -14228 42866 -14172 42868
rect -14228 42814 -14226 42866
rect -14226 42814 -14174 42866
rect -14174 42814 -14172 42866
rect -14228 42812 -14172 42814
rect -14068 42866 -14012 42868
rect -14068 42814 -14066 42866
rect -14066 42814 -14014 42866
rect -14014 42814 -14012 42866
rect -14068 42812 -14012 42814
rect -13908 42866 -13852 42868
rect -13908 42814 -13906 42866
rect -13906 42814 -13854 42866
rect -13854 42814 -13852 42866
rect -13908 42812 -13852 42814
rect -13748 42866 -13692 42868
rect -13748 42814 -13746 42866
rect -13746 42814 -13694 42866
rect -13694 42814 -13692 42866
rect -13748 42812 -13692 42814
rect -13588 42866 -13532 42868
rect -13588 42814 -13586 42866
rect -13586 42814 -13534 42866
rect -13534 42814 -13532 42866
rect -13588 42812 -13532 42814
rect -13428 42866 -13372 42868
rect -13428 42814 -13426 42866
rect -13426 42814 -13374 42866
rect -13374 42814 -13372 42866
rect -13428 42812 -13372 42814
rect -13268 42866 -13212 42868
rect -13268 42814 -13266 42866
rect -13266 42814 -13214 42866
rect -13214 42814 -13212 42866
rect -13268 42812 -13212 42814
rect -13108 42866 -13052 42868
rect -13108 42814 -13106 42866
rect -13106 42814 -13054 42866
rect -13054 42814 -13052 42866
rect -13108 42812 -13052 42814
rect -12948 42866 -12892 42868
rect -12948 42814 -12946 42866
rect -12946 42814 -12894 42866
rect -12894 42814 -12892 42866
rect -12948 42812 -12892 42814
rect -12788 42866 -12732 42868
rect -12788 42814 -12786 42866
rect -12786 42814 -12734 42866
rect -12734 42814 -12732 42866
rect -12788 42812 -12732 42814
rect -12628 42866 -12572 42868
rect -12628 42814 -12626 42866
rect -12626 42814 -12574 42866
rect -12574 42814 -12572 42866
rect -12628 42812 -12572 42814
rect -12468 42866 -12412 42868
rect -12468 42814 -12466 42866
rect -12466 42814 -12414 42866
rect -12414 42814 -12412 42866
rect -12468 42812 -12412 42814
rect -12308 42866 -12252 42868
rect -12308 42814 -12306 42866
rect -12306 42814 -12254 42866
rect -12254 42814 -12252 42866
rect -12308 42812 -12252 42814
rect -12148 42812 -12092 42868
rect -11828 42812 -11772 42868
rect -11508 42812 -11452 42868
rect -11348 42866 -11292 42868
rect -11348 42814 -11346 42866
rect -11346 42814 -11294 42866
rect -11294 42814 -11292 42866
rect -11348 42812 -11292 42814
rect -11188 42866 -11132 42868
rect -11188 42814 -11186 42866
rect -11186 42814 -11134 42866
rect -11134 42814 -11132 42866
rect -11188 42812 -11132 42814
rect -11028 42866 -10972 42868
rect -11028 42814 -11026 42866
rect -11026 42814 -10974 42866
rect -10974 42814 -10972 42866
rect -11028 42812 -10972 42814
rect -10868 42866 -10812 42868
rect -10868 42814 -10866 42866
rect -10866 42814 -10814 42866
rect -10814 42814 -10812 42866
rect -10868 42812 -10812 42814
rect -10708 42866 -10652 42868
rect -10708 42814 -10706 42866
rect -10706 42814 -10654 42866
rect -10654 42814 -10652 42866
rect -10708 42812 -10652 42814
rect -10548 42866 -10492 42868
rect -10548 42814 -10546 42866
rect -10546 42814 -10494 42866
rect -10494 42814 -10492 42866
rect -10548 42812 -10492 42814
rect -10388 42866 -10332 42868
rect -10388 42814 -10386 42866
rect -10386 42814 -10334 42866
rect -10334 42814 -10332 42866
rect -10388 42812 -10332 42814
rect -10228 42866 -10172 42868
rect -10228 42814 -10226 42866
rect -10226 42814 -10174 42866
rect -10174 42814 -10172 42866
rect -10228 42812 -10172 42814
rect -10068 42866 -10012 42868
rect -10068 42814 -10066 42866
rect -10066 42814 -10014 42866
rect -10014 42814 -10012 42866
rect -10068 42812 -10012 42814
rect -9908 42866 -9852 42868
rect -9908 42814 -9906 42866
rect -9906 42814 -9854 42866
rect -9854 42814 -9852 42866
rect -9908 42812 -9852 42814
rect -9748 42866 -9692 42868
rect -9748 42814 -9746 42866
rect -9746 42814 -9694 42866
rect -9694 42814 -9692 42866
rect -9748 42812 -9692 42814
rect -9588 42866 -9532 42868
rect -9588 42814 -9586 42866
rect -9586 42814 -9534 42866
rect -9534 42814 -9532 42866
rect -9588 42812 -9532 42814
rect -9428 42866 -9372 42868
rect -9428 42814 -9426 42866
rect -9426 42814 -9374 42866
rect -9374 42814 -9372 42866
rect -9428 42812 -9372 42814
rect -9268 42866 -9212 42868
rect -9268 42814 -9266 42866
rect -9266 42814 -9214 42866
rect -9214 42814 -9212 42866
rect -9268 42812 -9212 42814
rect -9108 42866 -9052 42868
rect -9108 42814 -9106 42866
rect -9106 42814 -9054 42866
rect -9054 42814 -9052 42866
rect -9108 42812 -9052 42814
rect -8948 42866 -8892 42868
rect -8948 42814 -8946 42866
rect -8946 42814 -8894 42866
rect -8894 42814 -8892 42866
rect -8948 42812 -8892 42814
rect -8788 42866 -8732 42868
rect -8788 42814 -8786 42866
rect -8786 42814 -8734 42866
rect -8734 42814 -8732 42866
rect -8788 42812 -8732 42814
rect -8628 42866 -8572 42868
rect -8628 42814 -8626 42866
rect -8626 42814 -8574 42866
rect -8574 42814 -8572 42866
rect -8628 42812 -8572 42814
rect -8468 42866 -8412 42868
rect -8468 42814 -8466 42866
rect -8466 42814 -8414 42866
rect -8414 42814 -8412 42866
rect -8468 42812 -8412 42814
rect -8308 42866 -8252 42868
rect -8308 42814 -8306 42866
rect -8306 42814 -8254 42866
rect -8254 42814 -8252 42866
rect -8308 42812 -8252 42814
rect -8148 42866 -8092 42868
rect -8148 42814 -8146 42866
rect -8146 42814 -8094 42866
rect -8094 42814 -8092 42866
rect -8148 42812 -8092 42814
rect -7988 42866 -7932 42868
rect -7988 42814 -7986 42866
rect -7986 42814 -7934 42866
rect -7934 42814 -7932 42866
rect -7988 42812 -7932 42814
rect -7828 42866 -7772 42868
rect -7828 42814 -7826 42866
rect -7826 42814 -7774 42866
rect -7774 42814 -7772 42866
rect -7828 42812 -7772 42814
rect -7668 42866 -7612 42868
rect -7668 42814 -7666 42866
rect -7666 42814 -7614 42866
rect -7614 42814 -7612 42866
rect -7668 42812 -7612 42814
rect -7508 42866 -7452 42868
rect -7508 42814 -7506 42866
rect -7506 42814 -7454 42866
rect -7454 42814 -7452 42866
rect -7508 42812 -7452 42814
rect -7348 42866 -7292 42868
rect -7348 42814 -7346 42866
rect -7346 42814 -7294 42866
rect -7294 42814 -7292 42866
rect -7348 42812 -7292 42814
rect -7188 42866 -7132 42868
rect -7188 42814 -7186 42866
rect -7186 42814 -7134 42866
rect -7134 42814 -7132 42866
rect -7188 42812 -7132 42814
rect -7028 42866 -6972 42868
rect -7028 42814 -7026 42866
rect -7026 42814 -6974 42866
rect -6974 42814 -6972 42866
rect -7028 42812 -6972 42814
rect -6868 42866 -6812 42868
rect -6868 42814 -6866 42866
rect -6866 42814 -6814 42866
rect -6814 42814 -6812 42866
rect -6868 42812 -6812 42814
rect -6708 42866 -6652 42868
rect -6708 42814 -6706 42866
rect -6706 42814 -6654 42866
rect -6654 42814 -6652 42866
rect -6708 42812 -6652 42814
rect -6548 42866 -6492 42868
rect -6548 42814 -6546 42866
rect -6546 42814 -6494 42866
rect -6494 42814 -6492 42866
rect -6548 42812 -6492 42814
rect -6388 42866 -6332 42868
rect -6388 42814 -6386 42866
rect -6386 42814 -6334 42866
rect -6334 42814 -6332 42866
rect -6388 42812 -6332 42814
rect -6228 42866 -6172 42868
rect -6228 42814 -6226 42866
rect -6226 42814 -6174 42866
rect -6174 42814 -6172 42866
rect -6228 42812 -6172 42814
rect -6068 42866 -6012 42868
rect -6068 42814 -6066 42866
rect -6066 42814 -6014 42866
rect -6014 42814 -6012 42866
rect -6068 42812 -6012 42814
rect -5908 42866 -5852 42868
rect -5908 42814 -5906 42866
rect -5906 42814 -5854 42866
rect -5854 42814 -5852 42866
rect -5908 42812 -5852 42814
rect -5748 42866 -5692 42868
rect -5748 42814 -5746 42866
rect -5746 42814 -5694 42866
rect -5694 42814 -5692 42866
rect -5748 42812 -5692 42814
rect -5588 42866 -5532 42868
rect -5588 42814 -5586 42866
rect -5586 42814 -5534 42866
rect -5534 42814 -5532 42866
rect -5588 42812 -5532 42814
rect -5428 42866 -5372 42868
rect -5428 42814 -5426 42866
rect -5426 42814 -5374 42866
rect -5374 42814 -5372 42866
rect -5428 42812 -5372 42814
rect -5268 42866 -5212 42868
rect -5268 42814 -5266 42866
rect -5266 42814 -5214 42866
rect -5214 42814 -5212 42866
rect -5268 42812 -5212 42814
rect -5108 42866 -5052 42868
rect -5108 42814 -5106 42866
rect -5106 42814 -5054 42866
rect -5054 42814 -5052 42866
rect -5108 42812 -5052 42814
rect -4948 42866 -4892 42868
rect -4948 42814 -4946 42866
rect -4946 42814 -4894 42866
rect -4894 42814 -4892 42866
rect -4948 42812 -4892 42814
rect -4788 42866 -4732 42868
rect -4788 42814 -4786 42866
rect -4786 42814 -4734 42866
rect -4734 42814 -4732 42866
rect -4788 42812 -4732 42814
rect -4628 42866 -4572 42868
rect -4628 42814 -4626 42866
rect -4626 42814 -4574 42866
rect -4574 42814 -4572 42866
rect -4628 42812 -4572 42814
rect -4468 42866 -4412 42868
rect -4468 42814 -4466 42866
rect -4466 42814 -4414 42866
rect -4414 42814 -4412 42866
rect -4468 42812 -4412 42814
rect -4308 42866 -4252 42868
rect -4308 42814 -4306 42866
rect -4306 42814 -4254 42866
rect -4254 42814 -4252 42866
rect -4308 42812 -4252 42814
rect -4148 42866 -4092 42868
rect -4148 42814 -4146 42866
rect -4146 42814 -4094 42866
rect -4094 42814 -4092 42866
rect -4148 42812 -4092 42814
rect -3988 42866 -3932 42868
rect -3988 42814 -3986 42866
rect -3986 42814 -3934 42866
rect -3934 42814 -3932 42866
rect -3988 42812 -3932 42814
rect -3668 42866 -3612 42868
rect -3668 42814 -3666 42866
rect -3666 42814 -3614 42866
rect -3614 42814 -3612 42866
rect -3668 42812 -3612 42814
rect -3508 42866 -3452 42868
rect -3508 42814 -3506 42866
rect -3506 42814 -3454 42866
rect -3454 42814 -3452 42866
rect -3508 42812 -3452 42814
rect -3348 42866 -3292 42868
rect -3348 42814 -3346 42866
rect -3346 42814 -3294 42866
rect -3294 42814 -3292 42866
rect -3348 42812 -3292 42814
rect -3188 42812 -3132 42868
rect -3028 42866 -2972 42868
rect -3028 42814 -3026 42866
rect -3026 42814 -2974 42866
rect -2974 42814 -2972 42866
rect -3028 42812 -2972 42814
rect -2708 42866 -2652 42868
rect -2708 42814 -2706 42866
rect -2706 42814 -2654 42866
rect -2654 42814 -2652 42866
rect -2708 42812 -2652 42814
rect -2548 42866 -2492 42868
rect -2548 42814 -2546 42866
rect -2546 42814 -2494 42866
rect -2494 42814 -2492 42866
rect -2548 42812 -2492 42814
rect -2388 42866 -2332 42868
rect -2388 42814 -2386 42866
rect -2386 42814 -2334 42866
rect -2334 42814 -2332 42866
rect -2388 42812 -2332 42814
rect -2228 42866 -2172 42868
rect -2228 42814 -2226 42866
rect -2226 42814 -2174 42866
rect -2174 42814 -2172 42866
rect -2228 42812 -2172 42814
rect -2068 42866 -2012 42868
rect -2068 42814 -2066 42866
rect -2066 42814 -2014 42866
rect -2014 42814 -2012 42866
rect -2068 42812 -2012 42814
rect -1748 42866 -1692 42868
rect -1748 42814 -1746 42866
rect -1746 42814 -1694 42866
rect -1694 42814 -1692 42866
rect -1748 42812 -1692 42814
rect -1428 42866 -1372 42868
rect -1428 42814 -1426 42866
rect -1426 42814 -1374 42866
rect -1374 42814 -1372 42866
rect -1428 42812 -1372 42814
rect -1108 42866 -1052 42868
rect -1108 42814 -1106 42866
rect -1106 42814 -1054 42866
rect -1054 42814 -1052 42866
rect -1108 42812 -1052 42814
rect -31028 42652 -30972 42708
rect -30708 42652 -30652 42708
rect -30388 42652 -30332 42708
rect -30228 42652 -30172 42708
rect -11988 42652 -11932 42708
rect -2868 42652 -2812 42708
rect -31028 42492 -30972 42548
rect -30708 42492 -30652 42548
rect -30388 42492 -30332 42548
rect -30068 42492 -30012 42548
rect -29908 42546 -29852 42548
rect -29908 42494 -29906 42546
rect -29906 42494 -29854 42546
rect -29854 42494 -29852 42546
rect -29908 42492 -29852 42494
rect -29748 42546 -29692 42548
rect -29748 42494 -29746 42546
rect -29746 42494 -29694 42546
rect -29694 42494 -29692 42546
rect -29748 42492 -29692 42494
rect -29588 42546 -29532 42548
rect -29588 42494 -29586 42546
rect -29586 42494 -29534 42546
rect -29534 42494 -29532 42546
rect -29588 42492 -29532 42494
rect -29428 42546 -29372 42548
rect -29428 42494 -29426 42546
rect -29426 42494 -29374 42546
rect -29374 42494 -29372 42546
rect -29428 42492 -29372 42494
rect -29268 42546 -29212 42548
rect -29268 42494 -29266 42546
rect -29266 42494 -29214 42546
rect -29214 42494 -29212 42546
rect -29268 42492 -29212 42494
rect -29108 42546 -29052 42548
rect -29108 42494 -29106 42546
rect -29106 42494 -29054 42546
rect -29054 42494 -29052 42546
rect -29108 42492 -29052 42494
rect -28948 42546 -28892 42548
rect -28948 42494 -28946 42546
rect -28946 42494 -28894 42546
rect -28894 42494 -28892 42546
rect -28948 42492 -28892 42494
rect -28788 42546 -28732 42548
rect -28788 42494 -28786 42546
rect -28786 42494 -28734 42546
rect -28734 42494 -28732 42546
rect -28788 42492 -28732 42494
rect -28628 42546 -28572 42548
rect -28628 42494 -28626 42546
rect -28626 42494 -28574 42546
rect -28574 42494 -28572 42546
rect -28628 42492 -28572 42494
rect -28468 42546 -28412 42548
rect -28468 42494 -28466 42546
rect -28466 42494 -28414 42546
rect -28414 42494 -28412 42546
rect -28468 42492 -28412 42494
rect -28308 42546 -28252 42548
rect -28308 42494 -28306 42546
rect -28306 42494 -28254 42546
rect -28254 42494 -28252 42546
rect -28308 42492 -28252 42494
rect -28148 42546 -28092 42548
rect -28148 42494 -28146 42546
rect -28146 42494 -28094 42546
rect -28094 42494 -28092 42546
rect -28148 42492 -28092 42494
rect -27988 42546 -27932 42548
rect -27988 42494 -27986 42546
rect -27986 42494 -27934 42546
rect -27934 42494 -27932 42546
rect -27988 42492 -27932 42494
rect -27828 42546 -27772 42548
rect -27828 42494 -27826 42546
rect -27826 42494 -27774 42546
rect -27774 42494 -27772 42546
rect -27828 42492 -27772 42494
rect -27668 42546 -27612 42548
rect -27668 42494 -27666 42546
rect -27666 42494 -27614 42546
rect -27614 42494 -27612 42546
rect -27668 42492 -27612 42494
rect -27508 42546 -27452 42548
rect -27508 42494 -27506 42546
rect -27506 42494 -27454 42546
rect -27454 42494 -27452 42546
rect -27508 42492 -27452 42494
rect -27348 42546 -27292 42548
rect -27348 42494 -27346 42546
rect -27346 42494 -27294 42546
rect -27294 42494 -27292 42546
rect -27348 42492 -27292 42494
rect -27188 42546 -27132 42548
rect -27188 42494 -27186 42546
rect -27186 42494 -27134 42546
rect -27134 42494 -27132 42546
rect -27188 42492 -27132 42494
rect -27028 42546 -26972 42548
rect -27028 42494 -27026 42546
rect -27026 42494 -26974 42546
rect -26974 42494 -26972 42546
rect -27028 42492 -26972 42494
rect -26868 42546 -26812 42548
rect -26868 42494 -26866 42546
rect -26866 42494 -26814 42546
rect -26814 42494 -26812 42546
rect -26868 42492 -26812 42494
rect -26708 42546 -26652 42548
rect -26708 42494 -26706 42546
rect -26706 42494 -26654 42546
rect -26654 42494 -26652 42546
rect -26708 42492 -26652 42494
rect -26548 42546 -26492 42548
rect -26548 42494 -26546 42546
rect -26546 42494 -26494 42546
rect -26494 42494 -26492 42546
rect -26548 42492 -26492 42494
rect -26388 42546 -26332 42548
rect -26388 42494 -26386 42546
rect -26386 42494 -26334 42546
rect -26334 42494 -26332 42546
rect -26388 42492 -26332 42494
rect -26228 42546 -26172 42548
rect -26228 42494 -26226 42546
rect -26226 42494 -26174 42546
rect -26174 42494 -26172 42546
rect -26228 42492 -26172 42494
rect -26068 42546 -26012 42548
rect -26068 42494 -26066 42546
rect -26066 42494 -26014 42546
rect -26014 42494 -26012 42546
rect -26068 42492 -26012 42494
rect -25908 42546 -25852 42548
rect -25908 42494 -25906 42546
rect -25906 42494 -25854 42546
rect -25854 42494 -25852 42546
rect -25908 42492 -25852 42494
rect -25748 42546 -25692 42548
rect -25748 42494 -25746 42546
rect -25746 42494 -25694 42546
rect -25694 42494 -25692 42546
rect -25748 42492 -25692 42494
rect -25588 42546 -25532 42548
rect -25588 42494 -25586 42546
rect -25586 42494 -25534 42546
rect -25534 42494 -25532 42546
rect -25588 42492 -25532 42494
rect -25428 42546 -25372 42548
rect -25428 42494 -25426 42546
rect -25426 42494 -25374 42546
rect -25374 42494 -25372 42546
rect -25428 42492 -25372 42494
rect -25268 42546 -25212 42548
rect -25268 42494 -25266 42546
rect -25266 42494 -25214 42546
rect -25214 42494 -25212 42546
rect -25268 42492 -25212 42494
rect -25108 42546 -25052 42548
rect -25108 42494 -25106 42546
rect -25106 42494 -25054 42546
rect -25054 42494 -25052 42546
rect -25108 42492 -25052 42494
rect -24948 42546 -24892 42548
rect -24948 42494 -24946 42546
rect -24946 42494 -24894 42546
rect -24894 42494 -24892 42546
rect -24948 42492 -24892 42494
rect -24788 42546 -24732 42548
rect -24788 42494 -24786 42546
rect -24786 42494 -24734 42546
rect -24734 42494 -24732 42546
rect -24788 42492 -24732 42494
rect -24628 42546 -24572 42548
rect -24628 42494 -24626 42546
rect -24626 42494 -24574 42546
rect -24574 42494 -24572 42546
rect -24628 42492 -24572 42494
rect -24468 42546 -24412 42548
rect -24468 42494 -24466 42546
rect -24466 42494 -24414 42546
rect -24414 42494 -24412 42546
rect -24468 42492 -24412 42494
rect -24308 42546 -24252 42548
rect -24308 42494 -24306 42546
rect -24306 42494 -24254 42546
rect -24254 42494 -24252 42546
rect -24308 42492 -24252 42494
rect -24148 42546 -24092 42548
rect -24148 42494 -24146 42546
rect -24146 42494 -24094 42546
rect -24094 42494 -24092 42546
rect -24148 42492 -24092 42494
rect -23988 42546 -23932 42548
rect -23988 42494 -23986 42546
rect -23986 42494 -23934 42546
rect -23934 42494 -23932 42546
rect -23988 42492 -23932 42494
rect -23828 42546 -23772 42548
rect -23828 42494 -23826 42546
rect -23826 42494 -23774 42546
rect -23774 42494 -23772 42546
rect -23828 42492 -23772 42494
rect -23668 42546 -23612 42548
rect -23668 42494 -23666 42546
rect -23666 42494 -23614 42546
rect -23614 42494 -23612 42546
rect -23668 42492 -23612 42494
rect -23508 42546 -23452 42548
rect -23508 42494 -23506 42546
rect -23506 42494 -23454 42546
rect -23454 42494 -23452 42546
rect -23508 42492 -23452 42494
rect -23348 42546 -23292 42548
rect -23348 42494 -23346 42546
rect -23346 42494 -23294 42546
rect -23294 42494 -23292 42546
rect -23348 42492 -23292 42494
rect -23188 42546 -23132 42548
rect -23188 42494 -23186 42546
rect -23186 42494 -23134 42546
rect -23134 42494 -23132 42546
rect -23188 42492 -23132 42494
rect -23028 42546 -22972 42548
rect -23028 42494 -23026 42546
rect -23026 42494 -22974 42546
rect -22974 42494 -22972 42546
rect -23028 42492 -22972 42494
rect -22868 42546 -22812 42548
rect -22868 42494 -22866 42546
rect -22866 42494 -22814 42546
rect -22814 42494 -22812 42546
rect -22868 42492 -22812 42494
rect -22708 42546 -22652 42548
rect -22708 42494 -22706 42546
rect -22706 42494 -22654 42546
rect -22654 42494 -22652 42546
rect -22708 42492 -22652 42494
rect -22548 42546 -22492 42548
rect -22548 42494 -22546 42546
rect -22546 42494 -22494 42546
rect -22494 42494 -22492 42546
rect -22548 42492 -22492 42494
rect -22388 42546 -22332 42548
rect -22388 42494 -22386 42546
rect -22386 42494 -22334 42546
rect -22334 42494 -22332 42546
rect -22388 42492 -22332 42494
rect -22228 42546 -22172 42548
rect -22228 42494 -22226 42546
rect -22226 42494 -22174 42546
rect -22174 42494 -22172 42546
rect -22228 42492 -22172 42494
rect -22068 42546 -22012 42548
rect -22068 42494 -22066 42546
rect -22066 42494 -22014 42546
rect -22014 42494 -22012 42546
rect -22068 42492 -22012 42494
rect -21908 42546 -21852 42548
rect -21908 42494 -21906 42546
rect -21906 42494 -21854 42546
rect -21854 42494 -21852 42546
rect -21908 42492 -21852 42494
rect -21748 42546 -21692 42548
rect -21748 42494 -21746 42546
rect -21746 42494 -21694 42546
rect -21694 42494 -21692 42546
rect -21748 42492 -21692 42494
rect -21588 42546 -21532 42548
rect -21588 42494 -21586 42546
rect -21586 42494 -21534 42546
rect -21534 42494 -21532 42546
rect -21588 42492 -21532 42494
rect -21428 42546 -21372 42548
rect -21428 42494 -21426 42546
rect -21426 42494 -21374 42546
rect -21374 42494 -21372 42546
rect -21428 42492 -21372 42494
rect -21268 42546 -21212 42548
rect -21268 42494 -21266 42546
rect -21266 42494 -21214 42546
rect -21214 42494 -21212 42546
rect -21268 42492 -21212 42494
rect -21108 42546 -21052 42548
rect -21108 42494 -21106 42546
rect -21106 42494 -21054 42546
rect -21054 42494 -21052 42546
rect -21108 42492 -21052 42494
rect -20948 42546 -20892 42548
rect -20948 42494 -20946 42546
rect -20946 42494 -20894 42546
rect -20894 42494 -20892 42546
rect -20948 42492 -20892 42494
rect -20788 42546 -20732 42548
rect -20788 42494 -20786 42546
rect -20786 42494 -20734 42546
rect -20734 42494 -20732 42546
rect -20788 42492 -20732 42494
rect -20628 42546 -20572 42548
rect -20628 42494 -20626 42546
rect -20626 42494 -20574 42546
rect -20574 42494 -20572 42546
rect -20628 42492 -20572 42494
rect -20468 42546 -20412 42548
rect -20468 42494 -20466 42546
rect -20466 42494 -20414 42546
rect -20414 42494 -20412 42546
rect -20468 42492 -20412 42494
rect -20308 42546 -20252 42548
rect -20308 42494 -20306 42546
rect -20306 42494 -20254 42546
rect -20254 42494 -20252 42546
rect -20308 42492 -20252 42494
rect -20148 42546 -20092 42548
rect -20148 42494 -20146 42546
rect -20146 42494 -20094 42546
rect -20094 42494 -20092 42546
rect -20148 42492 -20092 42494
rect -19988 42546 -19932 42548
rect -19988 42494 -19986 42546
rect -19986 42494 -19934 42546
rect -19934 42494 -19932 42546
rect -19988 42492 -19932 42494
rect -19828 42546 -19772 42548
rect -19828 42494 -19826 42546
rect -19826 42494 -19774 42546
rect -19774 42494 -19772 42546
rect -19828 42492 -19772 42494
rect -19668 42546 -19612 42548
rect -19668 42494 -19666 42546
rect -19666 42494 -19614 42546
rect -19614 42494 -19612 42546
rect -19668 42492 -19612 42494
rect -19508 42546 -19452 42548
rect -19508 42494 -19506 42546
rect -19506 42494 -19454 42546
rect -19454 42494 -19452 42546
rect -19508 42492 -19452 42494
rect -19348 42546 -19292 42548
rect -19348 42494 -19346 42546
rect -19346 42494 -19294 42546
rect -19294 42494 -19292 42546
rect -19348 42492 -19292 42494
rect -19188 42546 -19132 42548
rect -19188 42494 -19186 42546
rect -19186 42494 -19134 42546
rect -19134 42494 -19132 42546
rect -19188 42492 -19132 42494
rect -19028 42546 -18972 42548
rect -19028 42494 -19026 42546
rect -19026 42494 -18974 42546
rect -18974 42494 -18972 42546
rect -19028 42492 -18972 42494
rect -18868 42546 -18812 42548
rect -18868 42494 -18866 42546
rect -18866 42494 -18814 42546
rect -18814 42494 -18812 42546
rect -18868 42492 -18812 42494
rect -18708 42546 -18652 42548
rect -18708 42494 -18706 42546
rect -18706 42494 -18654 42546
rect -18654 42494 -18652 42546
rect -18708 42492 -18652 42494
rect -18548 42546 -18492 42548
rect -18548 42494 -18546 42546
rect -18546 42494 -18494 42546
rect -18494 42494 -18492 42546
rect -18548 42492 -18492 42494
rect -18388 42546 -18332 42548
rect -18388 42494 -18386 42546
rect -18386 42494 -18334 42546
rect -18334 42494 -18332 42546
rect -18388 42492 -18332 42494
rect -18228 42546 -18172 42548
rect -18228 42494 -18226 42546
rect -18226 42494 -18174 42546
rect -18174 42494 -18172 42546
rect -18228 42492 -18172 42494
rect -18068 42546 -18012 42548
rect -18068 42494 -18066 42546
rect -18066 42494 -18014 42546
rect -18014 42494 -18012 42546
rect -18068 42492 -18012 42494
rect -17908 42546 -17852 42548
rect -17908 42494 -17906 42546
rect -17906 42494 -17854 42546
rect -17854 42494 -17852 42546
rect -17908 42492 -17852 42494
rect -17748 42546 -17692 42548
rect -17748 42494 -17746 42546
rect -17746 42494 -17694 42546
rect -17694 42494 -17692 42546
rect -17748 42492 -17692 42494
rect -17588 42546 -17532 42548
rect -17588 42494 -17586 42546
rect -17586 42494 -17534 42546
rect -17534 42494 -17532 42546
rect -17588 42492 -17532 42494
rect -17428 42546 -17372 42548
rect -17428 42494 -17426 42546
rect -17426 42494 -17374 42546
rect -17374 42494 -17372 42546
rect -17428 42492 -17372 42494
rect -17268 42546 -17212 42548
rect -17268 42494 -17266 42546
rect -17266 42494 -17214 42546
rect -17214 42494 -17212 42546
rect -17268 42492 -17212 42494
rect -17108 42546 -17052 42548
rect -17108 42494 -17106 42546
rect -17106 42494 -17054 42546
rect -17054 42494 -17052 42546
rect -17108 42492 -17052 42494
rect -16948 42546 -16892 42548
rect -16948 42494 -16946 42546
rect -16946 42494 -16894 42546
rect -16894 42494 -16892 42546
rect -16948 42492 -16892 42494
rect -16788 42546 -16732 42548
rect -16788 42494 -16786 42546
rect -16786 42494 -16734 42546
rect -16734 42494 -16732 42546
rect -16788 42492 -16732 42494
rect -16628 42546 -16572 42548
rect -16628 42494 -16626 42546
rect -16626 42494 -16574 42546
rect -16574 42494 -16572 42546
rect -16628 42492 -16572 42494
rect -16468 42546 -16412 42548
rect -16468 42494 -16466 42546
rect -16466 42494 -16414 42546
rect -16414 42494 -16412 42546
rect -16468 42492 -16412 42494
rect -16308 42546 -16252 42548
rect -16308 42494 -16306 42546
rect -16306 42494 -16254 42546
rect -16254 42494 -16252 42546
rect -16308 42492 -16252 42494
rect -16148 42546 -16092 42548
rect -16148 42494 -16146 42546
rect -16146 42494 -16094 42546
rect -16094 42494 -16092 42546
rect -16148 42492 -16092 42494
rect -15988 42546 -15932 42548
rect -15988 42494 -15986 42546
rect -15986 42494 -15934 42546
rect -15934 42494 -15932 42546
rect -15988 42492 -15932 42494
rect -15828 42546 -15772 42548
rect -15828 42494 -15826 42546
rect -15826 42494 -15774 42546
rect -15774 42494 -15772 42546
rect -15828 42492 -15772 42494
rect -15668 42546 -15612 42548
rect -15668 42494 -15666 42546
rect -15666 42494 -15614 42546
rect -15614 42494 -15612 42546
rect -15668 42492 -15612 42494
rect -15508 42546 -15452 42548
rect -15508 42494 -15506 42546
rect -15506 42494 -15454 42546
rect -15454 42494 -15452 42546
rect -15508 42492 -15452 42494
rect -15348 42546 -15292 42548
rect -15348 42494 -15346 42546
rect -15346 42494 -15294 42546
rect -15294 42494 -15292 42546
rect -15348 42492 -15292 42494
rect -15188 42546 -15132 42548
rect -15188 42494 -15186 42546
rect -15186 42494 -15134 42546
rect -15134 42494 -15132 42546
rect -15188 42492 -15132 42494
rect -15028 42546 -14972 42548
rect -15028 42494 -15026 42546
rect -15026 42494 -14974 42546
rect -14974 42494 -14972 42546
rect -15028 42492 -14972 42494
rect -14868 42546 -14812 42548
rect -14868 42494 -14866 42546
rect -14866 42494 -14814 42546
rect -14814 42494 -14812 42546
rect -14868 42492 -14812 42494
rect -14708 42546 -14652 42548
rect -14708 42494 -14706 42546
rect -14706 42494 -14654 42546
rect -14654 42494 -14652 42546
rect -14708 42492 -14652 42494
rect -14548 42546 -14492 42548
rect -14548 42494 -14546 42546
rect -14546 42494 -14494 42546
rect -14494 42494 -14492 42546
rect -14548 42492 -14492 42494
rect -14388 42546 -14332 42548
rect -14388 42494 -14386 42546
rect -14386 42494 -14334 42546
rect -14334 42494 -14332 42546
rect -14388 42492 -14332 42494
rect -14228 42546 -14172 42548
rect -14228 42494 -14226 42546
rect -14226 42494 -14174 42546
rect -14174 42494 -14172 42546
rect -14228 42492 -14172 42494
rect -14068 42546 -14012 42548
rect -14068 42494 -14066 42546
rect -14066 42494 -14014 42546
rect -14014 42494 -14012 42546
rect -14068 42492 -14012 42494
rect -13908 42546 -13852 42548
rect -13908 42494 -13906 42546
rect -13906 42494 -13854 42546
rect -13854 42494 -13852 42546
rect -13908 42492 -13852 42494
rect -13748 42546 -13692 42548
rect -13748 42494 -13746 42546
rect -13746 42494 -13694 42546
rect -13694 42494 -13692 42546
rect -13748 42492 -13692 42494
rect -13588 42546 -13532 42548
rect -13588 42494 -13586 42546
rect -13586 42494 -13534 42546
rect -13534 42494 -13532 42546
rect -13588 42492 -13532 42494
rect -13428 42546 -13372 42548
rect -13428 42494 -13426 42546
rect -13426 42494 -13374 42546
rect -13374 42494 -13372 42546
rect -13428 42492 -13372 42494
rect -13268 42546 -13212 42548
rect -13268 42494 -13266 42546
rect -13266 42494 -13214 42546
rect -13214 42494 -13212 42546
rect -13268 42492 -13212 42494
rect -13108 42546 -13052 42548
rect -13108 42494 -13106 42546
rect -13106 42494 -13054 42546
rect -13054 42494 -13052 42546
rect -13108 42492 -13052 42494
rect -12948 42546 -12892 42548
rect -12948 42494 -12946 42546
rect -12946 42494 -12894 42546
rect -12894 42494 -12892 42546
rect -12948 42492 -12892 42494
rect -12788 42546 -12732 42548
rect -12788 42494 -12786 42546
rect -12786 42494 -12734 42546
rect -12734 42494 -12732 42546
rect -12788 42492 -12732 42494
rect -12628 42546 -12572 42548
rect -12628 42494 -12626 42546
rect -12626 42494 -12574 42546
rect -12574 42494 -12572 42546
rect -12628 42492 -12572 42494
rect -12468 42546 -12412 42548
rect -12468 42494 -12466 42546
rect -12466 42494 -12414 42546
rect -12414 42494 -12412 42546
rect -12468 42492 -12412 42494
rect -12308 42546 -12252 42548
rect -12308 42494 -12306 42546
rect -12306 42494 -12254 42546
rect -12254 42494 -12252 42546
rect -12308 42492 -12252 42494
rect -12148 42492 -12092 42548
rect -11828 42492 -11772 42548
rect -11508 42492 -11452 42548
rect -11348 42546 -11292 42548
rect -11348 42494 -11346 42546
rect -11346 42494 -11294 42546
rect -11294 42494 -11292 42546
rect -11348 42492 -11292 42494
rect -11188 42546 -11132 42548
rect -11188 42494 -11186 42546
rect -11186 42494 -11134 42546
rect -11134 42494 -11132 42546
rect -11188 42492 -11132 42494
rect -11028 42546 -10972 42548
rect -11028 42494 -11026 42546
rect -11026 42494 -10974 42546
rect -10974 42494 -10972 42546
rect -11028 42492 -10972 42494
rect -10868 42546 -10812 42548
rect -10868 42494 -10866 42546
rect -10866 42494 -10814 42546
rect -10814 42494 -10812 42546
rect -10868 42492 -10812 42494
rect -10708 42546 -10652 42548
rect -10708 42494 -10706 42546
rect -10706 42494 -10654 42546
rect -10654 42494 -10652 42546
rect -10708 42492 -10652 42494
rect -10548 42546 -10492 42548
rect -10548 42494 -10546 42546
rect -10546 42494 -10494 42546
rect -10494 42494 -10492 42546
rect -10548 42492 -10492 42494
rect -10388 42546 -10332 42548
rect -10388 42494 -10386 42546
rect -10386 42494 -10334 42546
rect -10334 42494 -10332 42546
rect -10388 42492 -10332 42494
rect -10228 42546 -10172 42548
rect -10228 42494 -10226 42546
rect -10226 42494 -10174 42546
rect -10174 42494 -10172 42546
rect -10228 42492 -10172 42494
rect -10068 42546 -10012 42548
rect -10068 42494 -10066 42546
rect -10066 42494 -10014 42546
rect -10014 42494 -10012 42546
rect -10068 42492 -10012 42494
rect -9908 42546 -9852 42548
rect -9908 42494 -9906 42546
rect -9906 42494 -9854 42546
rect -9854 42494 -9852 42546
rect -9908 42492 -9852 42494
rect -9748 42546 -9692 42548
rect -9748 42494 -9746 42546
rect -9746 42494 -9694 42546
rect -9694 42494 -9692 42546
rect -9748 42492 -9692 42494
rect -9588 42546 -9532 42548
rect -9588 42494 -9586 42546
rect -9586 42494 -9534 42546
rect -9534 42494 -9532 42546
rect -9588 42492 -9532 42494
rect -9428 42546 -9372 42548
rect -9428 42494 -9426 42546
rect -9426 42494 -9374 42546
rect -9374 42494 -9372 42546
rect -9428 42492 -9372 42494
rect -9268 42546 -9212 42548
rect -9268 42494 -9266 42546
rect -9266 42494 -9214 42546
rect -9214 42494 -9212 42546
rect -9268 42492 -9212 42494
rect -9108 42546 -9052 42548
rect -9108 42494 -9106 42546
rect -9106 42494 -9054 42546
rect -9054 42494 -9052 42546
rect -9108 42492 -9052 42494
rect -8948 42546 -8892 42548
rect -8948 42494 -8946 42546
rect -8946 42494 -8894 42546
rect -8894 42494 -8892 42546
rect -8948 42492 -8892 42494
rect -8788 42546 -8732 42548
rect -8788 42494 -8786 42546
rect -8786 42494 -8734 42546
rect -8734 42494 -8732 42546
rect -8788 42492 -8732 42494
rect -8628 42546 -8572 42548
rect -8628 42494 -8626 42546
rect -8626 42494 -8574 42546
rect -8574 42494 -8572 42546
rect -8628 42492 -8572 42494
rect -8468 42546 -8412 42548
rect -8468 42494 -8466 42546
rect -8466 42494 -8414 42546
rect -8414 42494 -8412 42546
rect -8468 42492 -8412 42494
rect -8308 42546 -8252 42548
rect -8308 42494 -8306 42546
rect -8306 42494 -8254 42546
rect -8254 42494 -8252 42546
rect -8308 42492 -8252 42494
rect -8148 42546 -8092 42548
rect -8148 42494 -8146 42546
rect -8146 42494 -8094 42546
rect -8094 42494 -8092 42546
rect -8148 42492 -8092 42494
rect -7988 42546 -7932 42548
rect -7988 42494 -7986 42546
rect -7986 42494 -7934 42546
rect -7934 42494 -7932 42546
rect -7988 42492 -7932 42494
rect -7828 42546 -7772 42548
rect -7828 42494 -7826 42546
rect -7826 42494 -7774 42546
rect -7774 42494 -7772 42546
rect -7828 42492 -7772 42494
rect -7668 42546 -7612 42548
rect -7668 42494 -7666 42546
rect -7666 42494 -7614 42546
rect -7614 42494 -7612 42546
rect -7668 42492 -7612 42494
rect -7508 42546 -7452 42548
rect -7508 42494 -7506 42546
rect -7506 42494 -7454 42546
rect -7454 42494 -7452 42546
rect -7508 42492 -7452 42494
rect -7348 42546 -7292 42548
rect -7348 42494 -7346 42546
rect -7346 42494 -7294 42546
rect -7294 42494 -7292 42546
rect -7348 42492 -7292 42494
rect -7188 42546 -7132 42548
rect -7188 42494 -7186 42546
rect -7186 42494 -7134 42546
rect -7134 42494 -7132 42546
rect -7188 42492 -7132 42494
rect -7028 42546 -6972 42548
rect -7028 42494 -7026 42546
rect -7026 42494 -6974 42546
rect -6974 42494 -6972 42546
rect -7028 42492 -6972 42494
rect -6868 42546 -6812 42548
rect -6868 42494 -6866 42546
rect -6866 42494 -6814 42546
rect -6814 42494 -6812 42546
rect -6868 42492 -6812 42494
rect -6708 42546 -6652 42548
rect -6708 42494 -6706 42546
rect -6706 42494 -6654 42546
rect -6654 42494 -6652 42546
rect -6708 42492 -6652 42494
rect -6548 42546 -6492 42548
rect -6548 42494 -6546 42546
rect -6546 42494 -6494 42546
rect -6494 42494 -6492 42546
rect -6548 42492 -6492 42494
rect -6388 42546 -6332 42548
rect -6388 42494 -6386 42546
rect -6386 42494 -6334 42546
rect -6334 42494 -6332 42546
rect -6388 42492 -6332 42494
rect -6228 42546 -6172 42548
rect -6228 42494 -6226 42546
rect -6226 42494 -6174 42546
rect -6174 42494 -6172 42546
rect -6228 42492 -6172 42494
rect -6068 42546 -6012 42548
rect -6068 42494 -6066 42546
rect -6066 42494 -6014 42546
rect -6014 42494 -6012 42546
rect -6068 42492 -6012 42494
rect -5908 42546 -5852 42548
rect -5908 42494 -5906 42546
rect -5906 42494 -5854 42546
rect -5854 42494 -5852 42546
rect -5908 42492 -5852 42494
rect -5748 42546 -5692 42548
rect -5748 42494 -5746 42546
rect -5746 42494 -5694 42546
rect -5694 42494 -5692 42546
rect -5748 42492 -5692 42494
rect -5588 42546 -5532 42548
rect -5588 42494 -5586 42546
rect -5586 42494 -5534 42546
rect -5534 42494 -5532 42546
rect -5588 42492 -5532 42494
rect -5428 42546 -5372 42548
rect -5428 42494 -5426 42546
rect -5426 42494 -5374 42546
rect -5374 42494 -5372 42546
rect -5428 42492 -5372 42494
rect -5268 42546 -5212 42548
rect -5268 42494 -5266 42546
rect -5266 42494 -5214 42546
rect -5214 42494 -5212 42546
rect -5268 42492 -5212 42494
rect -5108 42546 -5052 42548
rect -5108 42494 -5106 42546
rect -5106 42494 -5054 42546
rect -5054 42494 -5052 42546
rect -5108 42492 -5052 42494
rect -4948 42546 -4892 42548
rect -4948 42494 -4946 42546
rect -4946 42494 -4894 42546
rect -4894 42494 -4892 42546
rect -4948 42492 -4892 42494
rect -4788 42546 -4732 42548
rect -4788 42494 -4786 42546
rect -4786 42494 -4734 42546
rect -4734 42494 -4732 42546
rect -4788 42492 -4732 42494
rect -4628 42546 -4572 42548
rect -4628 42494 -4626 42546
rect -4626 42494 -4574 42546
rect -4574 42494 -4572 42546
rect -4628 42492 -4572 42494
rect -4468 42546 -4412 42548
rect -4468 42494 -4466 42546
rect -4466 42494 -4414 42546
rect -4414 42494 -4412 42546
rect -4468 42492 -4412 42494
rect -4308 42546 -4252 42548
rect -4308 42494 -4306 42546
rect -4306 42494 -4254 42546
rect -4254 42494 -4252 42546
rect -4308 42492 -4252 42494
rect -4148 42546 -4092 42548
rect -4148 42494 -4146 42546
rect -4146 42494 -4094 42546
rect -4094 42494 -4092 42546
rect -4148 42492 -4092 42494
rect -3988 42546 -3932 42548
rect -3988 42494 -3986 42546
rect -3986 42494 -3934 42546
rect -3934 42494 -3932 42546
rect -3988 42492 -3932 42494
rect -3668 42546 -3612 42548
rect -3668 42494 -3666 42546
rect -3666 42494 -3614 42546
rect -3614 42494 -3612 42546
rect -3668 42492 -3612 42494
rect -3508 42546 -3452 42548
rect -3508 42494 -3506 42546
rect -3506 42494 -3454 42546
rect -3454 42494 -3452 42546
rect -3508 42492 -3452 42494
rect -3348 42546 -3292 42548
rect -3348 42494 -3346 42546
rect -3346 42494 -3294 42546
rect -3294 42494 -3292 42546
rect -3348 42492 -3292 42494
rect -3188 42492 -3132 42548
rect -3028 42546 -2972 42548
rect -3028 42494 -3026 42546
rect -3026 42494 -2974 42546
rect -2974 42494 -2972 42546
rect -3028 42492 -2972 42494
rect -2708 42546 -2652 42548
rect -2708 42494 -2706 42546
rect -2706 42494 -2654 42546
rect -2654 42494 -2652 42546
rect -2708 42492 -2652 42494
rect -2548 42546 -2492 42548
rect -2548 42494 -2546 42546
rect -2546 42494 -2494 42546
rect -2494 42494 -2492 42546
rect -2548 42492 -2492 42494
rect -2388 42546 -2332 42548
rect -2388 42494 -2386 42546
rect -2386 42494 -2334 42546
rect -2334 42494 -2332 42546
rect -2388 42492 -2332 42494
rect -2228 42546 -2172 42548
rect -2228 42494 -2226 42546
rect -2226 42494 -2174 42546
rect -2174 42494 -2172 42546
rect -2228 42492 -2172 42494
rect -2068 42546 -2012 42548
rect -2068 42494 -2066 42546
rect -2066 42494 -2014 42546
rect -2014 42494 -2012 42546
rect -2068 42492 -2012 42494
rect -1748 42546 -1692 42548
rect -1748 42494 -1746 42546
rect -1746 42494 -1694 42546
rect -1694 42494 -1692 42546
rect -1748 42492 -1692 42494
rect -1428 42546 -1372 42548
rect -1428 42494 -1426 42546
rect -1426 42494 -1374 42546
rect -1374 42494 -1372 42546
rect -1428 42492 -1372 42494
rect -1108 42546 -1052 42548
rect -1108 42494 -1106 42546
rect -1106 42494 -1054 42546
rect -1054 42494 -1052 42546
rect -1108 42492 -1052 42494
rect -31028 42332 -30972 42388
rect -30708 42332 -30652 42388
rect -30548 42332 -30492 42388
rect -11668 42332 -11612 42388
rect -3188 42332 -3132 42388
rect -31028 42172 -30972 42228
rect -30708 42172 -30652 42228
rect -30388 42172 -30332 42228
rect -30068 42172 -30012 42228
rect -29908 42226 -29852 42228
rect -29908 42174 -29906 42226
rect -29906 42174 -29854 42226
rect -29854 42174 -29852 42226
rect -29908 42172 -29852 42174
rect -29748 42226 -29692 42228
rect -29748 42174 -29746 42226
rect -29746 42174 -29694 42226
rect -29694 42174 -29692 42226
rect -29748 42172 -29692 42174
rect -29588 42226 -29532 42228
rect -29588 42174 -29586 42226
rect -29586 42174 -29534 42226
rect -29534 42174 -29532 42226
rect -29588 42172 -29532 42174
rect -29428 42226 -29372 42228
rect -29428 42174 -29426 42226
rect -29426 42174 -29374 42226
rect -29374 42174 -29372 42226
rect -29428 42172 -29372 42174
rect -29268 42226 -29212 42228
rect -29268 42174 -29266 42226
rect -29266 42174 -29214 42226
rect -29214 42174 -29212 42226
rect -29268 42172 -29212 42174
rect -29108 42226 -29052 42228
rect -29108 42174 -29106 42226
rect -29106 42174 -29054 42226
rect -29054 42174 -29052 42226
rect -29108 42172 -29052 42174
rect -28948 42226 -28892 42228
rect -28948 42174 -28946 42226
rect -28946 42174 -28894 42226
rect -28894 42174 -28892 42226
rect -28948 42172 -28892 42174
rect -28788 42226 -28732 42228
rect -28788 42174 -28786 42226
rect -28786 42174 -28734 42226
rect -28734 42174 -28732 42226
rect -28788 42172 -28732 42174
rect -28628 42226 -28572 42228
rect -28628 42174 -28626 42226
rect -28626 42174 -28574 42226
rect -28574 42174 -28572 42226
rect -28628 42172 -28572 42174
rect -28468 42226 -28412 42228
rect -28468 42174 -28466 42226
rect -28466 42174 -28414 42226
rect -28414 42174 -28412 42226
rect -28468 42172 -28412 42174
rect -28308 42226 -28252 42228
rect -28308 42174 -28306 42226
rect -28306 42174 -28254 42226
rect -28254 42174 -28252 42226
rect -28308 42172 -28252 42174
rect -28148 42226 -28092 42228
rect -28148 42174 -28146 42226
rect -28146 42174 -28094 42226
rect -28094 42174 -28092 42226
rect -28148 42172 -28092 42174
rect -27988 42226 -27932 42228
rect -27988 42174 -27986 42226
rect -27986 42174 -27934 42226
rect -27934 42174 -27932 42226
rect -27988 42172 -27932 42174
rect -27828 42226 -27772 42228
rect -27828 42174 -27826 42226
rect -27826 42174 -27774 42226
rect -27774 42174 -27772 42226
rect -27828 42172 -27772 42174
rect -27668 42226 -27612 42228
rect -27668 42174 -27666 42226
rect -27666 42174 -27614 42226
rect -27614 42174 -27612 42226
rect -27668 42172 -27612 42174
rect -27508 42226 -27452 42228
rect -27508 42174 -27506 42226
rect -27506 42174 -27454 42226
rect -27454 42174 -27452 42226
rect -27508 42172 -27452 42174
rect -27348 42226 -27292 42228
rect -27348 42174 -27346 42226
rect -27346 42174 -27294 42226
rect -27294 42174 -27292 42226
rect -27348 42172 -27292 42174
rect -27188 42226 -27132 42228
rect -27188 42174 -27186 42226
rect -27186 42174 -27134 42226
rect -27134 42174 -27132 42226
rect -27188 42172 -27132 42174
rect -27028 42226 -26972 42228
rect -27028 42174 -27026 42226
rect -27026 42174 -26974 42226
rect -26974 42174 -26972 42226
rect -27028 42172 -26972 42174
rect -26868 42226 -26812 42228
rect -26868 42174 -26866 42226
rect -26866 42174 -26814 42226
rect -26814 42174 -26812 42226
rect -26868 42172 -26812 42174
rect -26708 42226 -26652 42228
rect -26708 42174 -26706 42226
rect -26706 42174 -26654 42226
rect -26654 42174 -26652 42226
rect -26708 42172 -26652 42174
rect -26548 42226 -26492 42228
rect -26548 42174 -26546 42226
rect -26546 42174 -26494 42226
rect -26494 42174 -26492 42226
rect -26548 42172 -26492 42174
rect -26388 42226 -26332 42228
rect -26388 42174 -26386 42226
rect -26386 42174 -26334 42226
rect -26334 42174 -26332 42226
rect -26388 42172 -26332 42174
rect -26228 42226 -26172 42228
rect -26228 42174 -26226 42226
rect -26226 42174 -26174 42226
rect -26174 42174 -26172 42226
rect -26228 42172 -26172 42174
rect -26068 42226 -26012 42228
rect -26068 42174 -26066 42226
rect -26066 42174 -26014 42226
rect -26014 42174 -26012 42226
rect -26068 42172 -26012 42174
rect -25908 42226 -25852 42228
rect -25908 42174 -25906 42226
rect -25906 42174 -25854 42226
rect -25854 42174 -25852 42226
rect -25908 42172 -25852 42174
rect -25748 42226 -25692 42228
rect -25748 42174 -25746 42226
rect -25746 42174 -25694 42226
rect -25694 42174 -25692 42226
rect -25748 42172 -25692 42174
rect -25588 42226 -25532 42228
rect -25588 42174 -25586 42226
rect -25586 42174 -25534 42226
rect -25534 42174 -25532 42226
rect -25588 42172 -25532 42174
rect -25428 42226 -25372 42228
rect -25428 42174 -25426 42226
rect -25426 42174 -25374 42226
rect -25374 42174 -25372 42226
rect -25428 42172 -25372 42174
rect -25268 42226 -25212 42228
rect -25268 42174 -25266 42226
rect -25266 42174 -25214 42226
rect -25214 42174 -25212 42226
rect -25268 42172 -25212 42174
rect -25108 42226 -25052 42228
rect -25108 42174 -25106 42226
rect -25106 42174 -25054 42226
rect -25054 42174 -25052 42226
rect -25108 42172 -25052 42174
rect -24948 42226 -24892 42228
rect -24948 42174 -24946 42226
rect -24946 42174 -24894 42226
rect -24894 42174 -24892 42226
rect -24948 42172 -24892 42174
rect -24788 42226 -24732 42228
rect -24788 42174 -24786 42226
rect -24786 42174 -24734 42226
rect -24734 42174 -24732 42226
rect -24788 42172 -24732 42174
rect -24628 42226 -24572 42228
rect -24628 42174 -24626 42226
rect -24626 42174 -24574 42226
rect -24574 42174 -24572 42226
rect -24628 42172 -24572 42174
rect -24468 42226 -24412 42228
rect -24468 42174 -24466 42226
rect -24466 42174 -24414 42226
rect -24414 42174 -24412 42226
rect -24468 42172 -24412 42174
rect -24308 42226 -24252 42228
rect -24308 42174 -24306 42226
rect -24306 42174 -24254 42226
rect -24254 42174 -24252 42226
rect -24308 42172 -24252 42174
rect -24148 42226 -24092 42228
rect -24148 42174 -24146 42226
rect -24146 42174 -24094 42226
rect -24094 42174 -24092 42226
rect -24148 42172 -24092 42174
rect -23988 42226 -23932 42228
rect -23988 42174 -23986 42226
rect -23986 42174 -23934 42226
rect -23934 42174 -23932 42226
rect -23988 42172 -23932 42174
rect -23828 42226 -23772 42228
rect -23828 42174 -23826 42226
rect -23826 42174 -23774 42226
rect -23774 42174 -23772 42226
rect -23828 42172 -23772 42174
rect -23668 42226 -23612 42228
rect -23668 42174 -23666 42226
rect -23666 42174 -23614 42226
rect -23614 42174 -23612 42226
rect -23668 42172 -23612 42174
rect -23508 42226 -23452 42228
rect -23508 42174 -23506 42226
rect -23506 42174 -23454 42226
rect -23454 42174 -23452 42226
rect -23508 42172 -23452 42174
rect -23348 42226 -23292 42228
rect -23348 42174 -23346 42226
rect -23346 42174 -23294 42226
rect -23294 42174 -23292 42226
rect -23348 42172 -23292 42174
rect -23188 42226 -23132 42228
rect -23188 42174 -23186 42226
rect -23186 42174 -23134 42226
rect -23134 42174 -23132 42226
rect -23188 42172 -23132 42174
rect -23028 42226 -22972 42228
rect -23028 42174 -23026 42226
rect -23026 42174 -22974 42226
rect -22974 42174 -22972 42226
rect -23028 42172 -22972 42174
rect -22868 42226 -22812 42228
rect -22868 42174 -22866 42226
rect -22866 42174 -22814 42226
rect -22814 42174 -22812 42226
rect -22868 42172 -22812 42174
rect -22708 42226 -22652 42228
rect -22708 42174 -22706 42226
rect -22706 42174 -22654 42226
rect -22654 42174 -22652 42226
rect -22708 42172 -22652 42174
rect -22548 42226 -22492 42228
rect -22548 42174 -22546 42226
rect -22546 42174 -22494 42226
rect -22494 42174 -22492 42226
rect -22548 42172 -22492 42174
rect -22388 42226 -22332 42228
rect -22388 42174 -22386 42226
rect -22386 42174 -22334 42226
rect -22334 42174 -22332 42226
rect -22388 42172 -22332 42174
rect -22228 42226 -22172 42228
rect -22228 42174 -22226 42226
rect -22226 42174 -22174 42226
rect -22174 42174 -22172 42226
rect -22228 42172 -22172 42174
rect -22068 42226 -22012 42228
rect -22068 42174 -22066 42226
rect -22066 42174 -22014 42226
rect -22014 42174 -22012 42226
rect -22068 42172 -22012 42174
rect -21908 42226 -21852 42228
rect -21908 42174 -21906 42226
rect -21906 42174 -21854 42226
rect -21854 42174 -21852 42226
rect -21908 42172 -21852 42174
rect -21748 42226 -21692 42228
rect -21748 42174 -21746 42226
rect -21746 42174 -21694 42226
rect -21694 42174 -21692 42226
rect -21748 42172 -21692 42174
rect -21588 42226 -21532 42228
rect -21588 42174 -21586 42226
rect -21586 42174 -21534 42226
rect -21534 42174 -21532 42226
rect -21588 42172 -21532 42174
rect -21428 42226 -21372 42228
rect -21428 42174 -21426 42226
rect -21426 42174 -21374 42226
rect -21374 42174 -21372 42226
rect -21428 42172 -21372 42174
rect -21268 42226 -21212 42228
rect -21268 42174 -21266 42226
rect -21266 42174 -21214 42226
rect -21214 42174 -21212 42226
rect -21268 42172 -21212 42174
rect -21108 42226 -21052 42228
rect -21108 42174 -21106 42226
rect -21106 42174 -21054 42226
rect -21054 42174 -21052 42226
rect -21108 42172 -21052 42174
rect -20948 42226 -20892 42228
rect -20948 42174 -20946 42226
rect -20946 42174 -20894 42226
rect -20894 42174 -20892 42226
rect -20948 42172 -20892 42174
rect -20788 42226 -20732 42228
rect -20788 42174 -20786 42226
rect -20786 42174 -20734 42226
rect -20734 42174 -20732 42226
rect -20788 42172 -20732 42174
rect -20628 42226 -20572 42228
rect -20628 42174 -20626 42226
rect -20626 42174 -20574 42226
rect -20574 42174 -20572 42226
rect -20628 42172 -20572 42174
rect -20468 42226 -20412 42228
rect -20468 42174 -20466 42226
rect -20466 42174 -20414 42226
rect -20414 42174 -20412 42226
rect -20468 42172 -20412 42174
rect -20308 42226 -20252 42228
rect -20308 42174 -20306 42226
rect -20306 42174 -20254 42226
rect -20254 42174 -20252 42226
rect -20308 42172 -20252 42174
rect -20148 42226 -20092 42228
rect -20148 42174 -20146 42226
rect -20146 42174 -20094 42226
rect -20094 42174 -20092 42226
rect -20148 42172 -20092 42174
rect -19988 42226 -19932 42228
rect -19988 42174 -19986 42226
rect -19986 42174 -19934 42226
rect -19934 42174 -19932 42226
rect -19988 42172 -19932 42174
rect -19828 42226 -19772 42228
rect -19828 42174 -19826 42226
rect -19826 42174 -19774 42226
rect -19774 42174 -19772 42226
rect -19828 42172 -19772 42174
rect -19668 42226 -19612 42228
rect -19668 42174 -19666 42226
rect -19666 42174 -19614 42226
rect -19614 42174 -19612 42226
rect -19668 42172 -19612 42174
rect -19508 42226 -19452 42228
rect -19508 42174 -19506 42226
rect -19506 42174 -19454 42226
rect -19454 42174 -19452 42226
rect -19508 42172 -19452 42174
rect -19348 42226 -19292 42228
rect -19348 42174 -19346 42226
rect -19346 42174 -19294 42226
rect -19294 42174 -19292 42226
rect -19348 42172 -19292 42174
rect -19188 42226 -19132 42228
rect -19188 42174 -19186 42226
rect -19186 42174 -19134 42226
rect -19134 42174 -19132 42226
rect -19188 42172 -19132 42174
rect -19028 42226 -18972 42228
rect -19028 42174 -19026 42226
rect -19026 42174 -18974 42226
rect -18974 42174 -18972 42226
rect -19028 42172 -18972 42174
rect -18868 42226 -18812 42228
rect -18868 42174 -18866 42226
rect -18866 42174 -18814 42226
rect -18814 42174 -18812 42226
rect -18868 42172 -18812 42174
rect -18708 42226 -18652 42228
rect -18708 42174 -18706 42226
rect -18706 42174 -18654 42226
rect -18654 42174 -18652 42226
rect -18708 42172 -18652 42174
rect -18548 42226 -18492 42228
rect -18548 42174 -18546 42226
rect -18546 42174 -18494 42226
rect -18494 42174 -18492 42226
rect -18548 42172 -18492 42174
rect -18388 42226 -18332 42228
rect -18388 42174 -18386 42226
rect -18386 42174 -18334 42226
rect -18334 42174 -18332 42226
rect -18388 42172 -18332 42174
rect -18228 42226 -18172 42228
rect -18228 42174 -18226 42226
rect -18226 42174 -18174 42226
rect -18174 42174 -18172 42226
rect -18228 42172 -18172 42174
rect -18068 42226 -18012 42228
rect -18068 42174 -18066 42226
rect -18066 42174 -18014 42226
rect -18014 42174 -18012 42226
rect -18068 42172 -18012 42174
rect -17908 42226 -17852 42228
rect -17908 42174 -17906 42226
rect -17906 42174 -17854 42226
rect -17854 42174 -17852 42226
rect -17908 42172 -17852 42174
rect -17748 42226 -17692 42228
rect -17748 42174 -17746 42226
rect -17746 42174 -17694 42226
rect -17694 42174 -17692 42226
rect -17748 42172 -17692 42174
rect -17588 42226 -17532 42228
rect -17588 42174 -17586 42226
rect -17586 42174 -17534 42226
rect -17534 42174 -17532 42226
rect -17588 42172 -17532 42174
rect -17428 42226 -17372 42228
rect -17428 42174 -17426 42226
rect -17426 42174 -17374 42226
rect -17374 42174 -17372 42226
rect -17428 42172 -17372 42174
rect -17268 42226 -17212 42228
rect -17268 42174 -17266 42226
rect -17266 42174 -17214 42226
rect -17214 42174 -17212 42226
rect -17268 42172 -17212 42174
rect -17108 42226 -17052 42228
rect -17108 42174 -17106 42226
rect -17106 42174 -17054 42226
rect -17054 42174 -17052 42226
rect -17108 42172 -17052 42174
rect -16948 42226 -16892 42228
rect -16948 42174 -16946 42226
rect -16946 42174 -16894 42226
rect -16894 42174 -16892 42226
rect -16948 42172 -16892 42174
rect -16788 42226 -16732 42228
rect -16788 42174 -16786 42226
rect -16786 42174 -16734 42226
rect -16734 42174 -16732 42226
rect -16788 42172 -16732 42174
rect -16628 42226 -16572 42228
rect -16628 42174 -16626 42226
rect -16626 42174 -16574 42226
rect -16574 42174 -16572 42226
rect -16628 42172 -16572 42174
rect -16468 42226 -16412 42228
rect -16468 42174 -16466 42226
rect -16466 42174 -16414 42226
rect -16414 42174 -16412 42226
rect -16468 42172 -16412 42174
rect -16308 42226 -16252 42228
rect -16308 42174 -16306 42226
rect -16306 42174 -16254 42226
rect -16254 42174 -16252 42226
rect -16308 42172 -16252 42174
rect -16148 42226 -16092 42228
rect -16148 42174 -16146 42226
rect -16146 42174 -16094 42226
rect -16094 42174 -16092 42226
rect -16148 42172 -16092 42174
rect -15988 42226 -15932 42228
rect -15988 42174 -15986 42226
rect -15986 42174 -15934 42226
rect -15934 42174 -15932 42226
rect -15988 42172 -15932 42174
rect -15828 42226 -15772 42228
rect -15828 42174 -15826 42226
rect -15826 42174 -15774 42226
rect -15774 42174 -15772 42226
rect -15828 42172 -15772 42174
rect -15668 42226 -15612 42228
rect -15668 42174 -15666 42226
rect -15666 42174 -15614 42226
rect -15614 42174 -15612 42226
rect -15668 42172 -15612 42174
rect -15508 42226 -15452 42228
rect -15508 42174 -15506 42226
rect -15506 42174 -15454 42226
rect -15454 42174 -15452 42226
rect -15508 42172 -15452 42174
rect -15348 42226 -15292 42228
rect -15348 42174 -15346 42226
rect -15346 42174 -15294 42226
rect -15294 42174 -15292 42226
rect -15348 42172 -15292 42174
rect -15188 42226 -15132 42228
rect -15188 42174 -15186 42226
rect -15186 42174 -15134 42226
rect -15134 42174 -15132 42226
rect -15188 42172 -15132 42174
rect -15028 42226 -14972 42228
rect -15028 42174 -15026 42226
rect -15026 42174 -14974 42226
rect -14974 42174 -14972 42226
rect -15028 42172 -14972 42174
rect -14868 42226 -14812 42228
rect -14868 42174 -14866 42226
rect -14866 42174 -14814 42226
rect -14814 42174 -14812 42226
rect -14868 42172 -14812 42174
rect -14708 42226 -14652 42228
rect -14708 42174 -14706 42226
rect -14706 42174 -14654 42226
rect -14654 42174 -14652 42226
rect -14708 42172 -14652 42174
rect -14548 42226 -14492 42228
rect -14548 42174 -14546 42226
rect -14546 42174 -14494 42226
rect -14494 42174 -14492 42226
rect -14548 42172 -14492 42174
rect -14388 42226 -14332 42228
rect -14388 42174 -14386 42226
rect -14386 42174 -14334 42226
rect -14334 42174 -14332 42226
rect -14388 42172 -14332 42174
rect -14228 42226 -14172 42228
rect -14228 42174 -14226 42226
rect -14226 42174 -14174 42226
rect -14174 42174 -14172 42226
rect -14228 42172 -14172 42174
rect -14068 42226 -14012 42228
rect -14068 42174 -14066 42226
rect -14066 42174 -14014 42226
rect -14014 42174 -14012 42226
rect -14068 42172 -14012 42174
rect -13908 42226 -13852 42228
rect -13908 42174 -13906 42226
rect -13906 42174 -13854 42226
rect -13854 42174 -13852 42226
rect -13908 42172 -13852 42174
rect -13748 42226 -13692 42228
rect -13748 42174 -13746 42226
rect -13746 42174 -13694 42226
rect -13694 42174 -13692 42226
rect -13748 42172 -13692 42174
rect -13588 42226 -13532 42228
rect -13588 42174 -13586 42226
rect -13586 42174 -13534 42226
rect -13534 42174 -13532 42226
rect -13588 42172 -13532 42174
rect -13428 42226 -13372 42228
rect -13428 42174 -13426 42226
rect -13426 42174 -13374 42226
rect -13374 42174 -13372 42226
rect -13428 42172 -13372 42174
rect -13268 42226 -13212 42228
rect -13268 42174 -13266 42226
rect -13266 42174 -13214 42226
rect -13214 42174 -13212 42226
rect -13268 42172 -13212 42174
rect -13108 42226 -13052 42228
rect -13108 42174 -13106 42226
rect -13106 42174 -13054 42226
rect -13054 42174 -13052 42226
rect -13108 42172 -13052 42174
rect -12948 42226 -12892 42228
rect -12948 42174 -12946 42226
rect -12946 42174 -12894 42226
rect -12894 42174 -12892 42226
rect -12948 42172 -12892 42174
rect -12788 42226 -12732 42228
rect -12788 42174 -12786 42226
rect -12786 42174 -12734 42226
rect -12734 42174 -12732 42226
rect -12788 42172 -12732 42174
rect -12628 42226 -12572 42228
rect -12628 42174 -12626 42226
rect -12626 42174 -12574 42226
rect -12574 42174 -12572 42226
rect -12628 42172 -12572 42174
rect -12468 42226 -12412 42228
rect -12468 42174 -12466 42226
rect -12466 42174 -12414 42226
rect -12414 42174 -12412 42226
rect -12468 42172 -12412 42174
rect -12308 42226 -12252 42228
rect -12308 42174 -12306 42226
rect -12306 42174 -12254 42226
rect -12254 42174 -12252 42226
rect -12308 42172 -12252 42174
rect -12148 42172 -12092 42228
rect -11828 42172 -11772 42228
rect -11508 42172 -11452 42228
rect -11348 42226 -11292 42228
rect -11348 42174 -11346 42226
rect -11346 42174 -11294 42226
rect -11294 42174 -11292 42226
rect -11348 42172 -11292 42174
rect -11188 42226 -11132 42228
rect -11188 42174 -11186 42226
rect -11186 42174 -11134 42226
rect -11134 42174 -11132 42226
rect -11188 42172 -11132 42174
rect -11028 42226 -10972 42228
rect -11028 42174 -11026 42226
rect -11026 42174 -10974 42226
rect -10974 42174 -10972 42226
rect -11028 42172 -10972 42174
rect -10868 42226 -10812 42228
rect -10868 42174 -10866 42226
rect -10866 42174 -10814 42226
rect -10814 42174 -10812 42226
rect -10868 42172 -10812 42174
rect -10708 42226 -10652 42228
rect -10708 42174 -10706 42226
rect -10706 42174 -10654 42226
rect -10654 42174 -10652 42226
rect -10708 42172 -10652 42174
rect -10548 42226 -10492 42228
rect -10548 42174 -10546 42226
rect -10546 42174 -10494 42226
rect -10494 42174 -10492 42226
rect -10548 42172 -10492 42174
rect -10388 42226 -10332 42228
rect -10388 42174 -10386 42226
rect -10386 42174 -10334 42226
rect -10334 42174 -10332 42226
rect -10388 42172 -10332 42174
rect -10228 42226 -10172 42228
rect -10228 42174 -10226 42226
rect -10226 42174 -10174 42226
rect -10174 42174 -10172 42226
rect -10228 42172 -10172 42174
rect -10068 42226 -10012 42228
rect -10068 42174 -10066 42226
rect -10066 42174 -10014 42226
rect -10014 42174 -10012 42226
rect -10068 42172 -10012 42174
rect -9908 42226 -9852 42228
rect -9908 42174 -9906 42226
rect -9906 42174 -9854 42226
rect -9854 42174 -9852 42226
rect -9908 42172 -9852 42174
rect -9748 42226 -9692 42228
rect -9748 42174 -9746 42226
rect -9746 42174 -9694 42226
rect -9694 42174 -9692 42226
rect -9748 42172 -9692 42174
rect -9588 42226 -9532 42228
rect -9588 42174 -9586 42226
rect -9586 42174 -9534 42226
rect -9534 42174 -9532 42226
rect -9588 42172 -9532 42174
rect -9428 42226 -9372 42228
rect -9428 42174 -9426 42226
rect -9426 42174 -9374 42226
rect -9374 42174 -9372 42226
rect -9428 42172 -9372 42174
rect -9268 42226 -9212 42228
rect -9268 42174 -9266 42226
rect -9266 42174 -9214 42226
rect -9214 42174 -9212 42226
rect -9268 42172 -9212 42174
rect -9108 42226 -9052 42228
rect -9108 42174 -9106 42226
rect -9106 42174 -9054 42226
rect -9054 42174 -9052 42226
rect -9108 42172 -9052 42174
rect -8948 42226 -8892 42228
rect -8948 42174 -8946 42226
rect -8946 42174 -8894 42226
rect -8894 42174 -8892 42226
rect -8948 42172 -8892 42174
rect -8788 42226 -8732 42228
rect -8788 42174 -8786 42226
rect -8786 42174 -8734 42226
rect -8734 42174 -8732 42226
rect -8788 42172 -8732 42174
rect -8628 42226 -8572 42228
rect -8628 42174 -8626 42226
rect -8626 42174 -8574 42226
rect -8574 42174 -8572 42226
rect -8628 42172 -8572 42174
rect -8468 42226 -8412 42228
rect -8468 42174 -8466 42226
rect -8466 42174 -8414 42226
rect -8414 42174 -8412 42226
rect -8468 42172 -8412 42174
rect -8308 42226 -8252 42228
rect -8308 42174 -8306 42226
rect -8306 42174 -8254 42226
rect -8254 42174 -8252 42226
rect -8308 42172 -8252 42174
rect -8148 42226 -8092 42228
rect -8148 42174 -8146 42226
rect -8146 42174 -8094 42226
rect -8094 42174 -8092 42226
rect -8148 42172 -8092 42174
rect -7988 42226 -7932 42228
rect -7988 42174 -7986 42226
rect -7986 42174 -7934 42226
rect -7934 42174 -7932 42226
rect -7988 42172 -7932 42174
rect -7828 42226 -7772 42228
rect -7828 42174 -7826 42226
rect -7826 42174 -7774 42226
rect -7774 42174 -7772 42226
rect -7828 42172 -7772 42174
rect -7668 42226 -7612 42228
rect -7668 42174 -7666 42226
rect -7666 42174 -7614 42226
rect -7614 42174 -7612 42226
rect -7668 42172 -7612 42174
rect -7508 42226 -7452 42228
rect -7508 42174 -7506 42226
rect -7506 42174 -7454 42226
rect -7454 42174 -7452 42226
rect -7508 42172 -7452 42174
rect -7348 42226 -7292 42228
rect -7348 42174 -7346 42226
rect -7346 42174 -7294 42226
rect -7294 42174 -7292 42226
rect -7348 42172 -7292 42174
rect -7188 42226 -7132 42228
rect -7188 42174 -7186 42226
rect -7186 42174 -7134 42226
rect -7134 42174 -7132 42226
rect -7188 42172 -7132 42174
rect -7028 42226 -6972 42228
rect -7028 42174 -7026 42226
rect -7026 42174 -6974 42226
rect -6974 42174 -6972 42226
rect -7028 42172 -6972 42174
rect -6868 42226 -6812 42228
rect -6868 42174 -6866 42226
rect -6866 42174 -6814 42226
rect -6814 42174 -6812 42226
rect -6868 42172 -6812 42174
rect -6708 42226 -6652 42228
rect -6708 42174 -6706 42226
rect -6706 42174 -6654 42226
rect -6654 42174 -6652 42226
rect -6708 42172 -6652 42174
rect -6548 42226 -6492 42228
rect -6548 42174 -6546 42226
rect -6546 42174 -6494 42226
rect -6494 42174 -6492 42226
rect -6548 42172 -6492 42174
rect -6388 42226 -6332 42228
rect -6388 42174 -6386 42226
rect -6386 42174 -6334 42226
rect -6334 42174 -6332 42226
rect -6388 42172 -6332 42174
rect -6228 42226 -6172 42228
rect -6228 42174 -6226 42226
rect -6226 42174 -6174 42226
rect -6174 42174 -6172 42226
rect -6228 42172 -6172 42174
rect -6068 42226 -6012 42228
rect -6068 42174 -6066 42226
rect -6066 42174 -6014 42226
rect -6014 42174 -6012 42226
rect -6068 42172 -6012 42174
rect -5908 42226 -5852 42228
rect -5908 42174 -5906 42226
rect -5906 42174 -5854 42226
rect -5854 42174 -5852 42226
rect -5908 42172 -5852 42174
rect -5748 42226 -5692 42228
rect -5748 42174 -5746 42226
rect -5746 42174 -5694 42226
rect -5694 42174 -5692 42226
rect -5748 42172 -5692 42174
rect -5588 42226 -5532 42228
rect -5588 42174 -5586 42226
rect -5586 42174 -5534 42226
rect -5534 42174 -5532 42226
rect -5588 42172 -5532 42174
rect -5428 42226 -5372 42228
rect -5428 42174 -5426 42226
rect -5426 42174 -5374 42226
rect -5374 42174 -5372 42226
rect -5428 42172 -5372 42174
rect -5268 42226 -5212 42228
rect -5268 42174 -5266 42226
rect -5266 42174 -5214 42226
rect -5214 42174 -5212 42226
rect -5268 42172 -5212 42174
rect -5108 42226 -5052 42228
rect -5108 42174 -5106 42226
rect -5106 42174 -5054 42226
rect -5054 42174 -5052 42226
rect -5108 42172 -5052 42174
rect -4948 42226 -4892 42228
rect -4948 42174 -4946 42226
rect -4946 42174 -4894 42226
rect -4894 42174 -4892 42226
rect -4948 42172 -4892 42174
rect -4788 42226 -4732 42228
rect -4788 42174 -4786 42226
rect -4786 42174 -4734 42226
rect -4734 42174 -4732 42226
rect -4788 42172 -4732 42174
rect -4628 42226 -4572 42228
rect -4628 42174 -4626 42226
rect -4626 42174 -4574 42226
rect -4574 42174 -4572 42226
rect -4628 42172 -4572 42174
rect -4468 42226 -4412 42228
rect -4468 42174 -4466 42226
rect -4466 42174 -4414 42226
rect -4414 42174 -4412 42226
rect -4468 42172 -4412 42174
rect -4308 42226 -4252 42228
rect -4308 42174 -4306 42226
rect -4306 42174 -4254 42226
rect -4254 42174 -4252 42226
rect -4308 42172 -4252 42174
rect -4148 42226 -4092 42228
rect -4148 42174 -4146 42226
rect -4146 42174 -4094 42226
rect -4094 42174 -4092 42226
rect -4148 42172 -4092 42174
rect -3988 42226 -3932 42228
rect -3988 42174 -3986 42226
rect -3986 42174 -3934 42226
rect -3934 42174 -3932 42226
rect -3988 42172 -3932 42174
rect -3668 42226 -3612 42228
rect -3668 42174 -3666 42226
rect -3666 42174 -3614 42226
rect -3614 42174 -3612 42226
rect -3668 42172 -3612 42174
rect -3508 42226 -3452 42228
rect -3508 42174 -3506 42226
rect -3506 42174 -3454 42226
rect -3454 42174 -3452 42226
rect -3508 42172 -3452 42174
rect -3348 42226 -3292 42228
rect -3348 42174 -3346 42226
rect -3346 42174 -3294 42226
rect -3294 42174 -3292 42226
rect -3348 42172 -3292 42174
rect -3028 42226 -2972 42228
rect -3028 42174 -3026 42226
rect -3026 42174 -2974 42226
rect -2974 42174 -2972 42226
rect -3028 42172 -2972 42174
rect -2708 42226 -2652 42228
rect -2708 42174 -2706 42226
rect -2706 42174 -2654 42226
rect -2654 42174 -2652 42226
rect -2708 42172 -2652 42174
rect -2548 42226 -2492 42228
rect -2548 42174 -2546 42226
rect -2546 42174 -2494 42226
rect -2494 42174 -2492 42226
rect -2548 42172 -2492 42174
rect -2388 42226 -2332 42228
rect -2388 42174 -2386 42226
rect -2386 42174 -2334 42226
rect -2334 42174 -2332 42226
rect -2388 42172 -2332 42174
rect -2228 42226 -2172 42228
rect -2228 42174 -2226 42226
rect -2226 42174 -2174 42226
rect -2174 42174 -2172 42226
rect -2228 42172 -2172 42174
rect -2068 42226 -2012 42228
rect -2068 42174 -2066 42226
rect -2066 42174 -2014 42226
rect -2014 42174 -2012 42226
rect -2068 42172 -2012 42174
rect -1748 42226 -1692 42228
rect -1748 42174 -1746 42226
rect -1746 42174 -1694 42226
rect -1694 42174 -1692 42226
rect -1748 42172 -1692 42174
rect -1428 42226 -1372 42228
rect -1428 42174 -1426 42226
rect -1426 42174 -1374 42226
rect -1374 42174 -1372 42226
rect -1428 42172 -1372 42174
rect -1108 42226 -1052 42228
rect -1108 42174 -1106 42226
rect -1106 42174 -1054 42226
rect -1054 42174 -1052 42226
rect -1108 42172 -1052 42174
rect -31028 42012 -30972 42068
rect -30708 42012 -30652 42068
rect -30388 42012 -30332 42068
rect -30228 42012 -30172 42068
rect -1268 42012 -1212 42068
rect -31028 41852 -30972 41908
rect -30708 41852 -30652 41908
rect -30388 41852 -30332 41908
rect -30068 41852 -30012 41908
rect -29908 41906 -29852 41908
rect -29908 41854 -29906 41906
rect -29906 41854 -29854 41906
rect -29854 41854 -29852 41906
rect -29908 41852 -29852 41854
rect -29748 41906 -29692 41908
rect -29748 41854 -29746 41906
rect -29746 41854 -29694 41906
rect -29694 41854 -29692 41906
rect -29748 41852 -29692 41854
rect -29588 41906 -29532 41908
rect -29588 41854 -29586 41906
rect -29586 41854 -29534 41906
rect -29534 41854 -29532 41906
rect -29588 41852 -29532 41854
rect -29428 41906 -29372 41908
rect -29428 41854 -29426 41906
rect -29426 41854 -29374 41906
rect -29374 41854 -29372 41906
rect -29428 41852 -29372 41854
rect -29268 41906 -29212 41908
rect -29268 41854 -29266 41906
rect -29266 41854 -29214 41906
rect -29214 41854 -29212 41906
rect -29268 41852 -29212 41854
rect -29108 41906 -29052 41908
rect -29108 41854 -29106 41906
rect -29106 41854 -29054 41906
rect -29054 41854 -29052 41906
rect -29108 41852 -29052 41854
rect -28948 41906 -28892 41908
rect -28948 41854 -28946 41906
rect -28946 41854 -28894 41906
rect -28894 41854 -28892 41906
rect -28948 41852 -28892 41854
rect -28788 41906 -28732 41908
rect -28788 41854 -28786 41906
rect -28786 41854 -28734 41906
rect -28734 41854 -28732 41906
rect -28788 41852 -28732 41854
rect -28628 41906 -28572 41908
rect -28628 41854 -28626 41906
rect -28626 41854 -28574 41906
rect -28574 41854 -28572 41906
rect -28628 41852 -28572 41854
rect -28468 41906 -28412 41908
rect -28468 41854 -28466 41906
rect -28466 41854 -28414 41906
rect -28414 41854 -28412 41906
rect -28468 41852 -28412 41854
rect -28308 41906 -28252 41908
rect -28308 41854 -28306 41906
rect -28306 41854 -28254 41906
rect -28254 41854 -28252 41906
rect -28308 41852 -28252 41854
rect -28148 41906 -28092 41908
rect -28148 41854 -28146 41906
rect -28146 41854 -28094 41906
rect -28094 41854 -28092 41906
rect -28148 41852 -28092 41854
rect -27988 41906 -27932 41908
rect -27988 41854 -27986 41906
rect -27986 41854 -27934 41906
rect -27934 41854 -27932 41906
rect -27988 41852 -27932 41854
rect -27828 41906 -27772 41908
rect -27828 41854 -27826 41906
rect -27826 41854 -27774 41906
rect -27774 41854 -27772 41906
rect -27828 41852 -27772 41854
rect -27668 41906 -27612 41908
rect -27668 41854 -27666 41906
rect -27666 41854 -27614 41906
rect -27614 41854 -27612 41906
rect -27668 41852 -27612 41854
rect -27508 41906 -27452 41908
rect -27508 41854 -27506 41906
rect -27506 41854 -27454 41906
rect -27454 41854 -27452 41906
rect -27508 41852 -27452 41854
rect -27348 41906 -27292 41908
rect -27348 41854 -27346 41906
rect -27346 41854 -27294 41906
rect -27294 41854 -27292 41906
rect -27348 41852 -27292 41854
rect -27188 41906 -27132 41908
rect -27188 41854 -27186 41906
rect -27186 41854 -27134 41906
rect -27134 41854 -27132 41906
rect -27188 41852 -27132 41854
rect -27028 41906 -26972 41908
rect -27028 41854 -27026 41906
rect -27026 41854 -26974 41906
rect -26974 41854 -26972 41906
rect -27028 41852 -26972 41854
rect -26868 41906 -26812 41908
rect -26868 41854 -26866 41906
rect -26866 41854 -26814 41906
rect -26814 41854 -26812 41906
rect -26868 41852 -26812 41854
rect -26708 41906 -26652 41908
rect -26708 41854 -26706 41906
rect -26706 41854 -26654 41906
rect -26654 41854 -26652 41906
rect -26708 41852 -26652 41854
rect -26548 41906 -26492 41908
rect -26548 41854 -26546 41906
rect -26546 41854 -26494 41906
rect -26494 41854 -26492 41906
rect -26548 41852 -26492 41854
rect -26388 41906 -26332 41908
rect -26388 41854 -26386 41906
rect -26386 41854 -26334 41906
rect -26334 41854 -26332 41906
rect -26388 41852 -26332 41854
rect -26228 41906 -26172 41908
rect -26228 41854 -26226 41906
rect -26226 41854 -26174 41906
rect -26174 41854 -26172 41906
rect -26228 41852 -26172 41854
rect -26068 41906 -26012 41908
rect -26068 41854 -26066 41906
rect -26066 41854 -26014 41906
rect -26014 41854 -26012 41906
rect -26068 41852 -26012 41854
rect -25908 41906 -25852 41908
rect -25908 41854 -25906 41906
rect -25906 41854 -25854 41906
rect -25854 41854 -25852 41906
rect -25908 41852 -25852 41854
rect -25748 41906 -25692 41908
rect -25748 41854 -25746 41906
rect -25746 41854 -25694 41906
rect -25694 41854 -25692 41906
rect -25748 41852 -25692 41854
rect -25588 41906 -25532 41908
rect -25588 41854 -25586 41906
rect -25586 41854 -25534 41906
rect -25534 41854 -25532 41906
rect -25588 41852 -25532 41854
rect -25428 41906 -25372 41908
rect -25428 41854 -25426 41906
rect -25426 41854 -25374 41906
rect -25374 41854 -25372 41906
rect -25428 41852 -25372 41854
rect -25268 41906 -25212 41908
rect -25268 41854 -25266 41906
rect -25266 41854 -25214 41906
rect -25214 41854 -25212 41906
rect -25268 41852 -25212 41854
rect -25108 41906 -25052 41908
rect -25108 41854 -25106 41906
rect -25106 41854 -25054 41906
rect -25054 41854 -25052 41906
rect -25108 41852 -25052 41854
rect -24948 41906 -24892 41908
rect -24948 41854 -24946 41906
rect -24946 41854 -24894 41906
rect -24894 41854 -24892 41906
rect -24948 41852 -24892 41854
rect -24788 41906 -24732 41908
rect -24788 41854 -24786 41906
rect -24786 41854 -24734 41906
rect -24734 41854 -24732 41906
rect -24788 41852 -24732 41854
rect -24628 41906 -24572 41908
rect -24628 41854 -24626 41906
rect -24626 41854 -24574 41906
rect -24574 41854 -24572 41906
rect -24628 41852 -24572 41854
rect -24468 41906 -24412 41908
rect -24468 41854 -24466 41906
rect -24466 41854 -24414 41906
rect -24414 41854 -24412 41906
rect -24468 41852 -24412 41854
rect -24308 41906 -24252 41908
rect -24308 41854 -24306 41906
rect -24306 41854 -24254 41906
rect -24254 41854 -24252 41906
rect -24308 41852 -24252 41854
rect -24148 41906 -24092 41908
rect -24148 41854 -24146 41906
rect -24146 41854 -24094 41906
rect -24094 41854 -24092 41906
rect -24148 41852 -24092 41854
rect -23988 41906 -23932 41908
rect -23988 41854 -23986 41906
rect -23986 41854 -23934 41906
rect -23934 41854 -23932 41906
rect -23988 41852 -23932 41854
rect -23828 41906 -23772 41908
rect -23828 41854 -23826 41906
rect -23826 41854 -23774 41906
rect -23774 41854 -23772 41906
rect -23828 41852 -23772 41854
rect -23668 41906 -23612 41908
rect -23668 41854 -23666 41906
rect -23666 41854 -23614 41906
rect -23614 41854 -23612 41906
rect -23668 41852 -23612 41854
rect -23508 41906 -23452 41908
rect -23508 41854 -23506 41906
rect -23506 41854 -23454 41906
rect -23454 41854 -23452 41906
rect -23508 41852 -23452 41854
rect -23348 41906 -23292 41908
rect -23348 41854 -23346 41906
rect -23346 41854 -23294 41906
rect -23294 41854 -23292 41906
rect -23348 41852 -23292 41854
rect -23188 41906 -23132 41908
rect -23188 41854 -23186 41906
rect -23186 41854 -23134 41906
rect -23134 41854 -23132 41906
rect -23188 41852 -23132 41854
rect -23028 41906 -22972 41908
rect -23028 41854 -23026 41906
rect -23026 41854 -22974 41906
rect -22974 41854 -22972 41906
rect -23028 41852 -22972 41854
rect -22868 41906 -22812 41908
rect -22868 41854 -22866 41906
rect -22866 41854 -22814 41906
rect -22814 41854 -22812 41906
rect -22868 41852 -22812 41854
rect -22708 41906 -22652 41908
rect -22708 41854 -22706 41906
rect -22706 41854 -22654 41906
rect -22654 41854 -22652 41906
rect -22708 41852 -22652 41854
rect -22548 41906 -22492 41908
rect -22548 41854 -22546 41906
rect -22546 41854 -22494 41906
rect -22494 41854 -22492 41906
rect -22548 41852 -22492 41854
rect -22388 41906 -22332 41908
rect -22388 41854 -22386 41906
rect -22386 41854 -22334 41906
rect -22334 41854 -22332 41906
rect -22388 41852 -22332 41854
rect -22228 41906 -22172 41908
rect -22228 41854 -22226 41906
rect -22226 41854 -22174 41906
rect -22174 41854 -22172 41906
rect -22228 41852 -22172 41854
rect -22068 41906 -22012 41908
rect -22068 41854 -22066 41906
rect -22066 41854 -22014 41906
rect -22014 41854 -22012 41906
rect -22068 41852 -22012 41854
rect -21908 41906 -21852 41908
rect -21908 41854 -21906 41906
rect -21906 41854 -21854 41906
rect -21854 41854 -21852 41906
rect -21908 41852 -21852 41854
rect -21748 41906 -21692 41908
rect -21748 41854 -21746 41906
rect -21746 41854 -21694 41906
rect -21694 41854 -21692 41906
rect -21748 41852 -21692 41854
rect -21588 41906 -21532 41908
rect -21588 41854 -21586 41906
rect -21586 41854 -21534 41906
rect -21534 41854 -21532 41906
rect -21588 41852 -21532 41854
rect -21428 41906 -21372 41908
rect -21428 41854 -21426 41906
rect -21426 41854 -21374 41906
rect -21374 41854 -21372 41906
rect -21428 41852 -21372 41854
rect -21268 41906 -21212 41908
rect -21268 41854 -21266 41906
rect -21266 41854 -21214 41906
rect -21214 41854 -21212 41906
rect -21268 41852 -21212 41854
rect -21108 41906 -21052 41908
rect -21108 41854 -21106 41906
rect -21106 41854 -21054 41906
rect -21054 41854 -21052 41906
rect -21108 41852 -21052 41854
rect -20948 41906 -20892 41908
rect -20948 41854 -20946 41906
rect -20946 41854 -20894 41906
rect -20894 41854 -20892 41906
rect -20948 41852 -20892 41854
rect -20788 41906 -20732 41908
rect -20788 41854 -20786 41906
rect -20786 41854 -20734 41906
rect -20734 41854 -20732 41906
rect -20788 41852 -20732 41854
rect -20628 41906 -20572 41908
rect -20628 41854 -20626 41906
rect -20626 41854 -20574 41906
rect -20574 41854 -20572 41906
rect -20628 41852 -20572 41854
rect -20468 41906 -20412 41908
rect -20468 41854 -20466 41906
rect -20466 41854 -20414 41906
rect -20414 41854 -20412 41906
rect -20468 41852 -20412 41854
rect -20308 41906 -20252 41908
rect -20308 41854 -20306 41906
rect -20306 41854 -20254 41906
rect -20254 41854 -20252 41906
rect -20308 41852 -20252 41854
rect -20148 41906 -20092 41908
rect -20148 41854 -20146 41906
rect -20146 41854 -20094 41906
rect -20094 41854 -20092 41906
rect -20148 41852 -20092 41854
rect -19988 41906 -19932 41908
rect -19988 41854 -19986 41906
rect -19986 41854 -19934 41906
rect -19934 41854 -19932 41906
rect -19988 41852 -19932 41854
rect -19828 41906 -19772 41908
rect -19828 41854 -19826 41906
rect -19826 41854 -19774 41906
rect -19774 41854 -19772 41906
rect -19828 41852 -19772 41854
rect -19668 41906 -19612 41908
rect -19668 41854 -19666 41906
rect -19666 41854 -19614 41906
rect -19614 41854 -19612 41906
rect -19668 41852 -19612 41854
rect -19508 41906 -19452 41908
rect -19508 41854 -19506 41906
rect -19506 41854 -19454 41906
rect -19454 41854 -19452 41906
rect -19508 41852 -19452 41854
rect -19348 41906 -19292 41908
rect -19348 41854 -19346 41906
rect -19346 41854 -19294 41906
rect -19294 41854 -19292 41906
rect -19348 41852 -19292 41854
rect -19188 41906 -19132 41908
rect -19188 41854 -19186 41906
rect -19186 41854 -19134 41906
rect -19134 41854 -19132 41906
rect -19188 41852 -19132 41854
rect -19028 41906 -18972 41908
rect -19028 41854 -19026 41906
rect -19026 41854 -18974 41906
rect -18974 41854 -18972 41906
rect -19028 41852 -18972 41854
rect -18868 41906 -18812 41908
rect -18868 41854 -18866 41906
rect -18866 41854 -18814 41906
rect -18814 41854 -18812 41906
rect -18868 41852 -18812 41854
rect -18708 41906 -18652 41908
rect -18708 41854 -18706 41906
rect -18706 41854 -18654 41906
rect -18654 41854 -18652 41906
rect -18708 41852 -18652 41854
rect -18548 41906 -18492 41908
rect -18548 41854 -18546 41906
rect -18546 41854 -18494 41906
rect -18494 41854 -18492 41906
rect -18548 41852 -18492 41854
rect -18388 41906 -18332 41908
rect -18388 41854 -18386 41906
rect -18386 41854 -18334 41906
rect -18334 41854 -18332 41906
rect -18388 41852 -18332 41854
rect -18228 41906 -18172 41908
rect -18228 41854 -18226 41906
rect -18226 41854 -18174 41906
rect -18174 41854 -18172 41906
rect -18228 41852 -18172 41854
rect -18068 41906 -18012 41908
rect -18068 41854 -18066 41906
rect -18066 41854 -18014 41906
rect -18014 41854 -18012 41906
rect -18068 41852 -18012 41854
rect -17908 41906 -17852 41908
rect -17908 41854 -17906 41906
rect -17906 41854 -17854 41906
rect -17854 41854 -17852 41906
rect -17908 41852 -17852 41854
rect -17748 41906 -17692 41908
rect -17748 41854 -17746 41906
rect -17746 41854 -17694 41906
rect -17694 41854 -17692 41906
rect -17748 41852 -17692 41854
rect -17588 41906 -17532 41908
rect -17588 41854 -17586 41906
rect -17586 41854 -17534 41906
rect -17534 41854 -17532 41906
rect -17588 41852 -17532 41854
rect -17428 41906 -17372 41908
rect -17428 41854 -17426 41906
rect -17426 41854 -17374 41906
rect -17374 41854 -17372 41906
rect -17428 41852 -17372 41854
rect -17268 41906 -17212 41908
rect -17268 41854 -17266 41906
rect -17266 41854 -17214 41906
rect -17214 41854 -17212 41906
rect -17268 41852 -17212 41854
rect -17108 41906 -17052 41908
rect -17108 41854 -17106 41906
rect -17106 41854 -17054 41906
rect -17054 41854 -17052 41906
rect -17108 41852 -17052 41854
rect -16948 41906 -16892 41908
rect -16948 41854 -16946 41906
rect -16946 41854 -16894 41906
rect -16894 41854 -16892 41906
rect -16948 41852 -16892 41854
rect -16788 41906 -16732 41908
rect -16788 41854 -16786 41906
rect -16786 41854 -16734 41906
rect -16734 41854 -16732 41906
rect -16788 41852 -16732 41854
rect -16628 41906 -16572 41908
rect -16628 41854 -16626 41906
rect -16626 41854 -16574 41906
rect -16574 41854 -16572 41906
rect -16628 41852 -16572 41854
rect -16468 41906 -16412 41908
rect -16468 41854 -16466 41906
rect -16466 41854 -16414 41906
rect -16414 41854 -16412 41906
rect -16468 41852 -16412 41854
rect -16308 41906 -16252 41908
rect -16308 41854 -16306 41906
rect -16306 41854 -16254 41906
rect -16254 41854 -16252 41906
rect -16308 41852 -16252 41854
rect -16148 41906 -16092 41908
rect -16148 41854 -16146 41906
rect -16146 41854 -16094 41906
rect -16094 41854 -16092 41906
rect -16148 41852 -16092 41854
rect -15988 41906 -15932 41908
rect -15988 41854 -15986 41906
rect -15986 41854 -15934 41906
rect -15934 41854 -15932 41906
rect -15988 41852 -15932 41854
rect -15828 41906 -15772 41908
rect -15828 41854 -15826 41906
rect -15826 41854 -15774 41906
rect -15774 41854 -15772 41906
rect -15828 41852 -15772 41854
rect -15668 41906 -15612 41908
rect -15668 41854 -15666 41906
rect -15666 41854 -15614 41906
rect -15614 41854 -15612 41906
rect -15668 41852 -15612 41854
rect -15508 41906 -15452 41908
rect -15508 41854 -15506 41906
rect -15506 41854 -15454 41906
rect -15454 41854 -15452 41906
rect -15508 41852 -15452 41854
rect -15348 41906 -15292 41908
rect -15348 41854 -15346 41906
rect -15346 41854 -15294 41906
rect -15294 41854 -15292 41906
rect -15348 41852 -15292 41854
rect -15188 41906 -15132 41908
rect -15188 41854 -15186 41906
rect -15186 41854 -15134 41906
rect -15134 41854 -15132 41906
rect -15188 41852 -15132 41854
rect -15028 41906 -14972 41908
rect -15028 41854 -15026 41906
rect -15026 41854 -14974 41906
rect -14974 41854 -14972 41906
rect -15028 41852 -14972 41854
rect -14868 41906 -14812 41908
rect -14868 41854 -14866 41906
rect -14866 41854 -14814 41906
rect -14814 41854 -14812 41906
rect -14868 41852 -14812 41854
rect -14708 41906 -14652 41908
rect -14708 41854 -14706 41906
rect -14706 41854 -14654 41906
rect -14654 41854 -14652 41906
rect -14708 41852 -14652 41854
rect -14548 41906 -14492 41908
rect -14548 41854 -14546 41906
rect -14546 41854 -14494 41906
rect -14494 41854 -14492 41906
rect -14548 41852 -14492 41854
rect -14388 41906 -14332 41908
rect -14388 41854 -14386 41906
rect -14386 41854 -14334 41906
rect -14334 41854 -14332 41906
rect -14388 41852 -14332 41854
rect -14228 41906 -14172 41908
rect -14228 41854 -14226 41906
rect -14226 41854 -14174 41906
rect -14174 41854 -14172 41906
rect -14228 41852 -14172 41854
rect -14068 41906 -14012 41908
rect -14068 41854 -14066 41906
rect -14066 41854 -14014 41906
rect -14014 41854 -14012 41906
rect -14068 41852 -14012 41854
rect -13908 41906 -13852 41908
rect -13908 41854 -13906 41906
rect -13906 41854 -13854 41906
rect -13854 41854 -13852 41906
rect -13908 41852 -13852 41854
rect -13748 41906 -13692 41908
rect -13748 41854 -13746 41906
rect -13746 41854 -13694 41906
rect -13694 41854 -13692 41906
rect -13748 41852 -13692 41854
rect -13588 41906 -13532 41908
rect -13588 41854 -13586 41906
rect -13586 41854 -13534 41906
rect -13534 41854 -13532 41906
rect -13588 41852 -13532 41854
rect -13428 41906 -13372 41908
rect -13428 41854 -13426 41906
rect -13426 41854 -13374 41906
rect -13374 41854 -13372 41906
rect -13428 41852 -13372 41854
rect -13268 41906 -13212 41908
rect -13268 41854 -13266 41906
rect -13266 41854 -13214 41906
rect -13214 41854 -13212 41906
rect -13268 41852 -13212 41854
rect -13108 41906 -13052 41908
rect -13108 41854 -13106 41906
rect -13106 41854 -13054 41906
rect -13054 41854 -13052 41906
rect -13108 41852 -13052 41854
rect -12948 41906 -12892 41908
rect -12948 41854 -12946 41906
rect -12946 41854 -12894 41906
rect -12894 41854 -12892 41906
rect -12948 41852 -12892 41854
rect -12788 41906 -12732 41908
rect -12788 41854 -12786 41906
rect -12786 41854 -12734 41906
rect -12734 41854 -12732 41906
rect -12788 41852 -12732 41854
rect -12628 41906 -12572 41908
rect -12628 41854 -12626 41906
rect -12626 41854 -12574 41906
rect -12574 41854 -12572 41906
rect -12628 41852 -12572 41854
rect -12468 41906 -12412 41908
rect -12468 41854 -12466 41906
rect -12466 41854 -12414 41906
rect -12414 41854 -12412 41906
rect -12468 41852 -12412 41854
rect -12308 41906 -12252 41908
rect -12308 41854 -12306 41906
rect -12306 41854 -12254 41906
rect -12254 41854 -12252 41906
rect -12308 41852 -12252 41854
rect -12148 41852 -12092 41908
rect -11828 41852 -11772 41908
rect -11508 41852 -11452 41908
rect -11348 41906 -11292 41908
rect -11348 41854 -11346 41906
rect -11346 41854 -11294 41906
rect -11294 41854 -11292 41906
rect -11348 41852 -11292 41854
rect -11188 41906 -11132 41908
rect -11188 41854 -11186 41906
rect -11186 41854 -11134 41906
rect -11134 41854 -11132 41906
rect -11188 41852 -11132 41854
rect -11028 41906 -10972 41908
rect -11028 41854 -11026 41906
rect -11026 41854 -10974 41906
rect -10974 41854 -10972 41906
rect -11028 41852 -10972 41854
rect -10868 41906 -10812 41908
rect -10868 41854 -10866 41906
rect -10866 41854 -10814 41906
rect -10814 41854 -10812 41906
rect -10868 41852 -10812 41854
rect -10708 41906 -10652 41908
rect -10708 41854 -10706 41906
rect -10706 41854 -10654 41906
rect -10654 41854 -10652 41906
rect -10708 41852 -10652 41854
rect -10548 41906 -10492 41908
rect -10548 41854 -10546 41906
rect -10546 41854 -10494 41906
rect -10494 41854 -10492 41906
rect -10548 41852 -10492 41854
rect -10388 41906 -10332 41908
rect -10388 41854 -10386 41906
rect -10386 41854 -10334 41906
rect -10334 41854 -10332 41906
rect -10388 41852 -10332 41854
rect -10228 41906 -10172 41908
rect -10228 41854 -10226 41906
rect -10226 41854 -10174 41906
rect -10174 41854 -10172 41906
rect -10228 41852 -10172 41854
rect -10068 41906 -10012 41908
rect -10068 41854 -10066 41906
rect -10066 41854 -10014 41906
rect -10014 41854 -10012 41906
rect -10068 41852 -10012 41854
rect -9908 41906 -9852 41908
rect -9908 41854 -9906 41906
rect -9906 41854 -9854 41906
rect -9854 41854 -9852 41906
rect -9908 41852 -9852 41854
rect -9748 41906 -9692 41908
rect -9748 41854 -9746 41906
rect -9746 41854 -9694 41906
rect -9694 41854 -9692 41906
rect -9748 41852 -9692 41854
rect -9588 41906 -9532 41908
rect -9588 41854 -9586 41906
rect -9586 41854 -9534 41906
rect -9534 41854 -9532 41906
rect -9588 41852 -9532 41854
rect -9428 41906 -9372 41908
rect -9428 41854 -9426 41906
rect -9426 41854 -9374 41906
rect -9374 41854 -9372 41906
rect -9428 41852 -9372 41854
rect -9268 41906 -9212 41908
rect -9268 41854 -9266 41906
rect -9266 41854 -9214 41906
rect -9214 41854 -9212 41906
rect -9268 41852 -9212 41854
rect -9108 41906 -9052 41908
rect -9108 41854 -9106 41906
rect -9106 41854 -9054 41906
rect -9054 41854 -9052 41906
rect -9108 41852 -9052 41854
rect -8948 41906 -8892 41908
rect -8948 41854 -8946 41906
rect -8946 41854 -8894 41906
rect -8894 41854 -8892 41906
rect -8948 41852 -8892 41854
rect -8788 41906 -8732 41908
rect -8788 41854 -8786 41906
rect -8786 41854 -8734 41906
rect -8734 41854 -8732 41906
rect -8788 41852 -8732 41854
rect -8628 41906 -8572 41908
rect -8628 41854 -8626 41906
rect -8626 41854 -8574 41906
rect -8574 41854 -8572 41906
rect -8628 41852 -8572 41854
rect -8468 41906 -8412 41908
rect -8468 41854 -8466 41906
rect -8466 41854 -8414 41906
rect -8414 41854 -8412 41906
rect -8468 41852 -8412 41854
rect -8308 41906 -8252 41908
rect -8308 41854 -8306 41906
rect -8306 41854 -8254 41906
rect -8254 41854 -8252 41906
rect -8308 41852 -8252 41854
rect -8148 41906 -8092 41908
rect -8148 41854 -8146 41906
rect -8146 41854 -8094 41906
rect -8094 41854 -8092 41906
rect -8148 41852 -8092 41854
rect -7988 41906 -7932 41908
rect -7988 41854 -7986 41906
rect -7986 41854 -7934 41906
rect -7934 41854 -7932 41906
rect -7988 41852 -7932 41854
rect -7828 41906 -7772 41908
rect -7828 41854 -7826 41906
rect -7826 41854 -7774 41906
rect -7774 41854 -7772 41906
rect -7828 41852 -7772 41854
rect -7668 41906 -7612 41908
rect -7668 41854 -7666 41906
rect -7666 41854 -7614 41906
rect -7614 41854 -7612 41906
rect -7668 41852 -7612 41854
rect -7508 41906 -7452 41908
rect -7508 41854 -7506 41906
rect -7506 41854 -7454 41906
rect -7454 41854 -7452 41906
rect -7508 41852 -7452 41854
rect -7348 41906 -7292 41908
rect -7348 41854 -7346 41906
rect -7346 41854 -7294 41906
rect -7294 41854 -7292 41906
rect -7348 41852 -7292 41854
rect -7188 41906 -7132 41908
rect -7188 41854 -7186 41906
rect -7186 41854 -7134 41906
rect -7134 41854 -7132 41906
rect -7188 41852 -7132 41854
rect -7028 41906 -6972 41908
rect -7028 41854 -7026 41906
rect -7026 41854 -6974 41906
rect -6974 41854 -6972 41906
rect -7028 41852 -6972 41854
rect -6868 41906 -6812 41908
rect -6868 41854 -6866 41906
rect -6866 41854 -6814 41906
rect -6814 41854 -6812 41906
rect -6868 41852 -6812 41854
rect -6708 41906 -6652 41908
rect -6708 41854 -6706 41906
rect -6706 41854 -6654 41906
rect -6654 41854 -6652 41906
rect -6708 41852 -6652 41854
rect -6548 41906 -6492 41908
rect -6548 41854 -6546 41906
rect -6546 41854 -6494 41906
rect -6494 41854 -6492 41906
rect -6548 41852 -6492 41854
rect -6388 41906 -6332 41908
rect -6388 41854 -6386 41906
rect -6386 41854 -6334 41906
rect -6334 41854 -6332 41906
rect -6388 41852 -6332 41854
rect -6228 41906 -6172 41908
rect -6228 41854 -6226 41906
rect -6226 41854 -6174 41906
rect -6174 41854 -6172 41906
rect -6228 41852 -6172 41854
rect -6068 41906 -6012 41908
rect -6068 41854 -6066 41906
rect -6066 41854 -6014 41906
rect -6014 41854 -6012 41906
rect -6068 41852 -6012 41854
rect -5908 41906 -5852 41908
rect -5908 41854 -5906 41906
rect -5906 41854 -5854 41906
rect -5854 41854 -5852 41906
rect -5908 41852 -5852 41854
rect -5748 41906 -5692 41908
rect -5748 41854 -5746 41906
rect -5746 41854 -5694 41906
rect -5694 41854 -5692 41906
rect -5748 41852 -5692 41854
rect -5588 41906 -5532 41908
rect -5588 41854 -5586 41906
rect -5586 41854 -5534 41906
rect -5534 41854 -5532 41906
rect -5588 41852 -5532 41854
rect -5428 41906 -5372 41908
rect -5428 41854 -5426 41906
rect -5426 41854 -5374 41906
rect -5374 41854 -5372 41906
rect -5428 41852 -5372 41854
rect -5268 41906 -5212 41908
rect -5268 41854 -5266 41906
rect -5266 41854 -5214 41906
rect -5214 41854 -5212 41906
rect -5268 41852 -5212 41854
rect -5108 41906 -5052 41908
rect -5108 41854 -5106 41906
rect -5106 41854 -5054 41906
rect -5054 41854 -5052 41906
rect -5108 41852 -5052 41854
rect -4948 41906 -4892 41908
rect -4948 41854 -4946 41906
rect -4946 41854 -4894 41906
rect -4894 41854 -4892 41906
rect -4948 41852 -4892 41854
rect -4788 41906 -4732 41908
rect -4788 41854 -4786 41906
rect -4786 41854 -4734 41906
rect -4734 41854 -4732 41906
rect -4788 41852 -4732 41854
rect -4628 41906 -4572 41908
rect -4628 41854 -4626 41906
rect -4626 41854 -4574 41906
rect -4574 41854 -4572 41906
rect -4628 41852 -4572 41854
rect -4468 41906 -4412 41908
rect -4468 41854 -4466 41906
rect -4466 41854 -4414 41906
rect -4414 41854 -4412 41906
rect -4468 41852 -4412 41854
rect -4308 41906 -4252 41908
rect -4308 41854 -4306 41906
rect -4306 41854 -4254 41906
rect -4254 41854 -4252 41906
rect -4308 41852 -4252 41854
rect -4148 41906 -4092 41908
rect -4148 41854 -4146 41906
rect -4146 41854 -4094 41906
rect -4094 41854 -4092 41906
rect -4148 41852 -4092 41854
rect -3988 41906 -3932 41908
rect -3988 41854 -3986 41906
rect -3986 41854 -3934 41906
rect -3934 41854 -3932 41906
rect -3988 41852 -3932 41854
rect -3668 41906 -3612 41908
rect -3668 41854 -3666 41906
rect -3666 41854 -3614 41906
rect -3614 41854 -3612 41906
rect -3668 41852 -3612 41854
rect -3508 41906 -3452 41908
rect -3508 41854 -3506 41906
rect -3506 41854 -3454 41906
rect -3454 41854 -3452 41906
rect -3508 41852 -3452 41854
rect -3348 41906 -3292 41908
rect -3348 41854 -3346 41906
rect -3346 41854 -3294 41906
rect -3294 41854 -3292 41906
rect -3348 41852 -3292 41854
rect -3028 41906 -2972 41908
rect -3028 41854 -3026 41906
rect -3026 41854 -2974 41906
rect -2974 41854 -2972 41906
rect -3028 41852 -2972 41854
rect -2708 41906 -2652 41908
rect -2708 41854 -2706 41906
rect -2706 41854 -2654 41906
rect -2654 41854 -2652 41906
rect -2708 41852 -2652 41854
rect -2548 41906 -2492 41908
rect -2548 41854 -2546 41906
rect -2546 41854 -2494 41906
rect -2494 41854 -2492 41906
rect -2548 41852 -2492 41854
rect -2388 41906 -2332 41908
rect -2388 41854 -2386 41906
rect -2386 41854 -2334 41906
rect -2334 41854 -2332 41906
rect -2388 41852 -2332 41854
rect -2228 41906 -2172 41908
rect -2228 41854 -2226 41906
rect -2226 41854 -2174 41906
rect -2174 41854 -2172 41906
rect -2228 41852 -2172 41854
rect -2068 41906 -2012 41908
rect -2068 41854 -2066 41906
rect -2066 41854 -2014 41906
rect -2014 41854 -2012 41906
rect -2068 41852 -2012 41854
rect -1748 41906 -1692 41908
rect -1748 41854 -1746 41906
rect -1746 41854 -1694 41906
rect -1694 41854 -1692 41906
rect -1748 41852 -1692 41854
rect -1428 41906 -1372 41908
rect -1428 41854 -1426 41906
rect -1426 41854 -1374 41906
rect -1374 41854 -1372 41906
rect -1428 41852 -1372 41854
rect -1108 41906 -1052 41908
rect -1108 41854 -1106 41906
rect -1106 41854 -1054 41906
rect -1054 41854 -1052 41906
rect -1108 41852 -1052 41854
rect -31028 41692 -30972 41748
rect -30708 41692 -30652 41748
rect -30388 41692 -30332 41748
rect -30068 41692 -30012 41748
rect -12148 41692 -12092 41748
rect -11828 41692 -11772 41748
rect -11508 41692 -11452 41748
rect -3348 41692 -3292 41748
rect -3028 41692 -2972 41748
rect -2708 41692 -2652 41748
rect -2388 41692 -2332 41748
rect -2068 41692 -2012 41748
rect -1748 41692 -1692 41748
rect -1428 41692 -1372 41748
rect -1108 41692 -1052 41748
rect -31028 41532 -30972 41588
rect -30708 41532 -30652 41588
rect -30388 41532 -30332 41588
rect -30068 41532 -30012 41588
rect -12148 41532 -12092 41588
rect -11828 41532 -11772 41588
rect -11508 41532 -11452 41588
rect -3348 41532 -3292 41588
rect -3028 41532 -2972 41588
rect -2708 41532 -2652 41588
rect -2388 41532 -2332 41588
rect -2068 41532 -2012 41588
rect -1748 41532 -1692 41588
rect -1428 41532 -1372 41588
rect -1108 41532 -1052 41588
rect -33108 41346 -33052 41348
rect -33108 41294 -33106 41346
rect -33106 41294 -33054 41346
rect -33054 41294 -33052 41346
rect -33108 41292 -33052 41294
rect -32948 41346 -32892 41348
rect -32948 41294 -32946 41346
rect -32946 41294 -32894 41346
rect -32894 41294 -32892 41346
rect -32948 41292 -32892 41294
rect -32788 41346 -32732 41348
rect -32788 41294 -32786 41346
rect -32786 41294 -32734 41346
rect -32734 41294 -32732 41346
rect -32788 41292 -32732 41294
rect -32628 41346 -32572 41348
rect -32628 41294 -32626 41346
rect -32626 41294 -32574 41346
rect -32574 41294 -32572 41346
rect -32628 41292 -32572 41294
rect -32468 41346 -32412 41348
rect -32468 41294 -32466 41346
rect -32466 41294 -32414 41346
rect -32414 41294 -32412 41346
rect -32468 41292 -32412 41294
rect -32308 41346 -32252 41348
rect -32308 41294 -32306 41346
rect -32306 41294 -32254 41346
rect -32254 41294 -32252 41346
rect -32308 41292 -32252 41294
rect -32148 41346 -32092 41348
rect -32148 41294 -32146 41346
rect -32146 41294 -32094 41346
rect -32094 41294 -32092 41346
rect -32148 41292 -32092 41294
rect -31988 41346 -31932 41348
rect -31988 41294 -31986 41346
rect -31986 41294 -31934 41346
rect -31934 41294 -31932 41346
rect -31988 41292 -31932 41294
rect -31828 41346 -31772 41348
rect -31828 41294 -31826 41346
rect -31826 41294 -31774 41346
rect -31774 41294 -31772 41346
rect -31828 41292 -31772 41294
rect -31668 41346 -31612 41348
rect -31668 41294 -31666 41346
rect -31666 41294 -31614 41346
rect -31614 41294 -31612 41346
rect -31668 41292 -31612 41294
rect -31508 41346 -31452 41348
rect -31508 41294 -31506 41346
rect -31506 41294 -31454 41346
rect -31454 41294 -31452 41346
rect -31508 41292 -31452 41294
rect -31348 41346 -31292 41348
rect -31348 41294 -31346 41346
rect -31346 41294 -31294 41346
rect -31294 41294 -31292 41346
rect -31348 41292 -31292 41294
rect -31188 41346 -31132 41348
rect -31188 41294 -31186 41346
rect -31186 41294 -31134 41346
rect -31134 41294 -31132 41346
rect -31188 41292 -31132 41294
rect -29908 41346 -29852 41348
rect -29908 41294 -29906 41346
rect -29906 41294 -29854 41346
rect -29854 41294 -29852 41346
rect -29908 41292 -29852 41294
rect -29748 41346 -29692 41348
rect -29748 41294 -29746 41346
rect -29746 41294 -29694 41346
rect -29694 41294 -29692 41346
rect -29748 41292 -29692 41294
rect -29588 41346 -29532 41348
rect -29588 41294 -29586 41346
rect -29586 41294 -29534 41346
rect -29534 41294 -29532 41346
rect -29588 41292 -29532 41294
rect -29428 41346 -29372 41348
rect -29428 41294 -29426 41346
rect -29426 41294 -29374 41346
rect -29374 41294 -29372 41346
rect -29428 41292 -29372 41294
rect -29268 41346 -29212 41348
rect -29268 41294 -29266 41346
rect -29266 41294 -29214 41346
rect -29214 41294 -29212 41346
rect -29268 41292 -29212 41294
rect -29108 41346 -29052 41348
rect -29108 41294 -29106 41346
rect -29106 41294 -29054 41346
rect -29054 41294 -29052 41346
rect -29108 41292 -29052 41294
rect -28948 41346 -28892 41348
rect -28948 41294 -28946 41346
rect -28946 41294 -28894 41346
rect -28894 41294 -28892 41346
rect -28948 41292 -28892 41294
rect -28788 41346 -28732 41348
rect -28788 41294 -28786 41346
rect -28786 41294 -28734 41346
rect -28734 41294 -28732 41346
rect -28788 41292 -28732 41294
rect -28628 41346 -28572 41348
rect -28628 41294 -28626 41346
rect -28626 41294 -28574 41346
rect -28574 41294 -28572 41346
rect -28628 41292 -28572 41294
rect -28468 41346 -28412 41348
rect -28468 41294 -28466 41346
rect -28466 41294 -28414 41346
rect -28414 41294 -28412 41346
rect -28468 41292 -28412 41294
rect -28308 41346 -28252 41348
rect -28308 41294 -28306 41346
rect -28306 41294 -28254 41346
rect -28254 41294 -28252 41346
rect -28308 41292 -28252 41294
rect -28148 41346 -28092 41348
rect -28148 41294 -28146 41346
rect -28146 41294 -28094 41346
rect -28094 41294 -28092 41346
rect -28148 41292 -28092 41294
rect -27988 41346 -27932 41348
rect -27988 41294 -27986 41346
rect -27986 41294 -27934 41346
rect -27934 41294 -27932 41346
rect -27988 41292 -27932 41294
rect -27828 41346 -27772 41348
rect -27828 41294 -27826 41346
rect -27826 41294 -27774 41346
rect -27774 41294 -27772 41346
rect -27828 41292 -27772 41294
rect -27668 41346 -27612 41348
rect -27668 41294 -27666 41346
rect -27666 41294 -27614 41346
rect -27614 41294 -27612 41346
rect -27668 41292 -27612 41294
rect -27508 41346 -27452 41348
rect -27508 41294 -27506 41346
rect -27506 41294 -27454 41346
rect -27454 41294 -27452 41346
rect -27508 41292 -27452 41294
rect -27348 41346 -27292 41348
rect -27348 41294 -27346 41346
rect -27346 41294 -27294 41346
rect -27294 41294 -27292 41346
rect -27348 41292 -27292 41294
rect -27188 41346 -27132 41348
rect -27188 41294 -27186 41346
rect -27186 41294 -27134 41346
rect -27134 41294 -27132 41346
rect -27188 41292 -27132 41294
rect -27028 41346 -26972 41348
rect -27028 41294 -27026 41346
rect -27026 41294 -26974 41346
rect -26974 41294 -26972 41346
rect -27028 41292 -26972 41294
rect -26868 41346 -26812 41348
rect -26868 41294 -26866 41346
rect -26866 41294 -26814 41346
rect -26814 41294 -26812 41346
rect -26868 41292 -26812 41294
rect -26708 41346 -26652 41348
rect -26708 41294 -26706 41346
rect -26706 41294 -26654 41346
rect -26654 41294 -26652 41346
rect -26708 41292 -26652 41294
rect -26548 41346 -26492 41348
rect -26548 41294 -26546 41346
rect -26546 41294 -26494 41346
rect -26494 41294 -26492 41346
rect -26548 41292 -26492 41294
rect -26388 41346 -26332 41348
rect -26388 41294 -26386 41346
rect -26386 41294 -26334 41346
rect -26334 41294 -26332 41346
rect -26388 41292 -26332 41294
rect -26228 41346 -26172 41348
rect -26228 41294 -26226 41346
rect -26226 41294 -26174 41346
rect -26174 41294 -26172 41346
rect -26228 41292 -26172 41294
rect -26068 41346 -26012 41348
rect -26068 41294 -26066 41346
rect -26066 41294 -26014 41346
rect -26014 41294 -26012 41346
rect -26068 41292 -26012 41294
rect -25908 41346 -25852 41348
rect -25908 41294 -25906 41346
rect -25906 41294 -25854 41346
rect -25854 41294 -25852 41346
rect -25908 41292 -25852 41294
rect -25748 41346 -25692 41348
rect -25748 41294 -25746 41346
rect -25746 41294 -25694 41346
rect -25694 41294 -25692 41346
rect -25748 41292 -25692 41294
rect -25588 41346 -25532 41348
rect -25588 41294 -25586 41346
rect -25586 41294 -25534 41346
rect -25534 41294 -25532 41346
rect -25588 41292 -25532 41294
rect -25428 41346 -25372 41348
rect -25428 41294 -25426 41346
rect -25426 41294 -25374 41346
rect -25374 41294 -25372 41346
rect -25428 41292 -25372 41294
rect -25268 41346 -25212 41348
rect -25268 41294 -25266 41346
rect -25266 41294 -25214 41346
rect -25214 41294 -25212 41346
rect -25268 41292 -25212 41294
rect -25108 41346 -25052 41348
rect -25108 41294 -25106 41346
rect -25106 41294 -25054 41346
rect -25054 41294 -25052 41346
rect -25108 41292 -25052 41294
rect -24948 41346 -24892 41348
rect -24948 41294 -24946 41346
rect -24946 41294 -24894 41346
rect -24894 41294 -24892 41346
rect -24948 41292 -24892 41294
rect -24788 41346 -24732 41348
rect -24788 41294 -24786 41346
rect -24786 41294 -24734 41346
rect -24734 41294 -24732 41346
rect -24788 41292 -24732 41294
rect -24628 41346 -24572 41348
rect -24628 41294 -24626 41346
rect -24626 41294 -24574 41346
rect -24574 41294 -24572 41346
rect -24628 41292 -24572 41294
rect -24468 41346 -24412 41348
rect -24468 41294 -24466 41346
rect -24466 41294 -24414 41346
rect -24414 41294 -24412 41346
rect -24468 41292 -24412 41294
rect -24308 41346 -24252 41348
rect -24308 41294 -24306 41346
rect -24306 41294 -24254 41346
rect -24254 41294 -24252 41346
rect -24308 41292 -24252 41294
rect -24148 41346 -24092 41348
rect -24148 41294 -24146 41346
rect -24146 41294 -24094 41346
rect -24094 41294 -24092 41346
rect -24148 41292 -24092 41294
rect -23988 41346 -23932 41348
rect -23988 41294 -23986 41346
rect -23986 41294 -23934 41346
rect -23934 41294 -23932 41346
rect -23988 41292 -23932 41294
rect -23828 41346 -23772 41348
rect -23828 41294 -23826 41346
rect -23826 41294 -23774 41346
rect -23774 41294 -23772 41346
rect -23828 41292 -23772 41294
rect -23668 41346 -23612 41348
rect -23668 41294 -23666 41346
rect -23666 41294 -23614 41346
rect -23614 41294 -23612 41346
rect -23668 41292 -23612 41294
rect -23508 41346 -23452 41348
rect -23508 41294 -23506 41346
rect -23506 41294 -23454 41346
rect -23454 41294 -23452 41346
rect -23508 41292 -23452 41294
rect -23348 41346 -23292 41348
rect -23348 41294 -23346 41346
rect -23346 41294 -23294 41346
rect -23294 41294 -23292 41346
rect -23348 41292 -23292 41294
rect -23188 41346 -23132 41348
rect -23188 41294 -23186 41346
rect -23186 41294 -23134 41346
rect -23134 41294 -23132 41346
rect -23188 41292 -23132 41294
rect -23028 41346 -22972 41348
rect -23028 41294 -23026 41346
rect -23026 41294 -22974 41346
rect -22974 41294 -22972 41346
rect -23028 41292 -22972 41294
rect -22868 41346 -22812 41348
rect -22868 41294 -22866 41346
rect -22866 41294 -22814 41346
rect -22814 41294 -22812 41346
rect -22868 41292 -22812 41294
rect -22708 41346 -22652 41348
rect -22708 41294 -22706 41346
rect -22706 41294 -22654 41346
rect -22654 41294 -22652 41346
rect -22708 41292 -22652 41294
rect -22548 41346 -22492 41348
rect -22548 41294 -22546 41346
rect -22546 41294 -22494 41346
rect -22494 41294 -22492 41346
rect -22548 41292 -22492 41294
rect -22388 41346 -22332 41348
rect -22388 41294 -22386 41346
rect -22386 41294 -22334 41346
rect -22334 41294 -22332 41346
rect -22388 41292 -22332 41294
rect -22228 41346 -22172 41348
rect -22228 41294 -22226 41346
rect -22226 41294 -22174 41346
rect -22174 41294 -22172 41346
rect -22228 41292 -22172 41294
rect -22068 41346 -22012 41348
rect -22068 41294 -22066 41346
rect -22066 41294 -22014 41346
rect -22014 41294 -22012 41346
rect -22068 41292 -22012 41294
rect -21908 41346 -21852 41348
rect -21908 41294 -21906 41346
rect -21906 41294 -21854 41346
rect -21854 41294 -21852 41346
rect -21908 41292 -21852 41294
rect -21748 41346 -21692 41348
rect -21748 41294 -21746 41346
rect -21746 41294 -21694 41346
rect -21694 41294 -21692 41346
rect -21748 41292 -21692 41294
rect -21588 41346 -21532 41348
rect -21588 41294 -21586 41346
rect -21586 41294 -21534 41346
rect -21534 41294 -21532 41346
rect -21588 41292 -21532 41294
rect -21428 41346 -21372 41348
rect -21428 41294 -21426 41346
rect -21426 41294 -21374 41346
rect -21374 41294 -21372 41346
rect -21428 41292 -21372 41294
rect -21268 41346 -21212 41348
rect -21268 41294 -21266 41346
rect -21266 41294 -21214 41346
rect -21214 41294 -21212 41346
rect -21268 41292 -21212 41294
rect -21108 41346 -21052 41348
rect -21108 41294 -21106 41346
rect -21106 41294 -21054 41346
rect -21054 41294 -21052 41346
rect -21108 41292 -21052 41294
rect -20948 41346 -20892 41348
rect -20948 41294 -20946 41346
rect -20946 41294 -20894 41346
rect -20894 41294 -20892 41346
rect -20948 41292 -20892 41294
rect -20788 41346 -20732 41348
rect -20788 41294 -20786 41346
rect -20786 41294 -20734 41346
rect -20734 41294 -20732 41346
rect -20788 41292 -20732 41294
rect -20628 41346 -20572 41348
rect -20628 41294 -20626 41346
rect -20626 41294 -20574 41346
rect -20574 41294 -20572 41346
rect -20628 41292 -20572 41294
rect -20468 41346 -20412 41348
rect -20468 41294 -20466 41346
rect -20466 41294 -20414 41346
rect -20414 41294 -20412 41346
rect -20468 41292 -20412 41294
rect -20308 41346 -20252 41348
rect -20308 41294 -20306 41346
rect -20306 41294 -20254 41346
rect -20254 41294 -20252 41346
rect -20308 41292 -20252 41294
rect -20148 41346 -20092 41348
rect -20148 41294 -20146 41346
rect -20146 41294 -20094 41346
rect -20094 41294 -20092 41346
rect -20148 41292 -20092 41294
rect -19988 41346 -19932 41348
rect -19988 41294 -19986 41346
rect -19986 41294 -19934 41346
rect -19934 41294 -19932 41346
rect -19988 41292 -19932 41294
rect -19828 41346 -19772 41348
rect -19828 41294 -19826 41346
rect -19826 41294 -19774 41346
rect -19774 41294 -19772 41346
rect -19828 41292 -19772 41294
rect -19668 41346 -19612 41348
rect -19668 41294 -19666 41346
rect -19666 41294 -19614 41346
rect -19614 41294 -19612 41346
rect -19668 41292 -19612 41294
rect -19508 41346 -19452 41348
rect -19508 41294 -19506 41346
rect -19506 41294 -19454 41346
rect -19454 41294 -19452 41346
rect -19508 41292 -19452 41294
rect -19348 41346 -19292 41348
rect -19348 41294 -19346 41346
rect -19346 41294 -19294 41346
rect -19294 41294 -19292 41346
rect -19348 41292 -19292 41294
rect -19188 41346 -19132 41348
rect -19188 41294 -19186 41346
rect -19186 41294 -19134 41346
rect -19134 41294 -19132 41346
rect -19188 41292 -19132 41294
rect -19028 41346 -18972 41348
rect -19028 41294 -19026 41346
rect -19026 41294 -18974 41346
rect -18974 41294 -18972 41346
rect -19028 41292 -18972 41294
rect -18868 41346 -18812 41348
rect -18868 41294 -18866 41346
rect -18866 41294 -18814 41346
rect -18814 41294 -18812 41346
rect -18868 41292 -18812 41294
rect -18708 41346 -18652 41348
rect -18708 41294 -18706 41346
rect -18706 41294 -18654 41346
rect -18654 41294 -18652 41346
rect -18708 41292 -18652 41294
rect -18548 41346 -18492 41348
rect -18548 41294 -18546 41346
rect -18546 41294 -18494 41346
rect -18494 41294 -18492 41346
rect -18548 41292 -18492 41294
rect -18388 41346 -18332 41348
rect -18388 41294 -18386 41346
rect -18386 41294 -18334 41346
rect -18334 41294 -18332 41346
rect -18388 41292 -18332 41294
rect -18228 41346 -18172 41348
rect -18228 41294 -18226 41346
rect -18226 41294 -18174 41346
rect -18174 41294 -18172 41346
rect -18228 41292 -18172 41294
rect -18068 41346 -18012 41348
rect -18068 41294 -18066 41346
rect -18066 41294 -18014 41346
rect -18014 41294 -18012 41346
rect -18068 41292 -18012 41294
rect -17908 41346 -17852 41348
rect -17908 41294 -17906 41346
rect -17906 41294 -17854 41346
rect -17854 41294 -17852 41346
rect -17908 41292 -17852 41294
rect -17748 41346 -17692 41348
rect -17748 41294 -17746 41346
rect -17746 41294 -17694 41346
rect -17694 41294 -17692 41346
rect -17748 41292 -17692 41294
rect -17588 41346 -17532 41348
rect -17588 41294 -17586 41346
rect -17586 41294 -17534 41346
rect -17534 41294 -17532 41346
rect -17588 41292 -17532 41294
rect -17428 41346 -17372 41348
rect -17428 41294 -17426 41346
rect -17426 41294 -17374 41346
rect -17374 41294 -17372 41346
rect -17428 41292 -17372 41294
rect -17268 41346 -17212 41348
rect -17268 41294 -17266 41346
rect -17266 41294 -17214 41346
rect -17214 41294 -17212 41346
rect -17268 41292 -17212 41294
rect -17108 41346 -17052 41348
rect -17108 41294 -17106 41346
rect -17106 41294 -17054 41346
rect -17054 41294 -17052 41346
rect -17108 41292 -17052 41294
rect -16948 41346 -16892 41348
rect -16948 41294 -16946 41346
rect -16946 41294 -16894 41346
rect -16894 41294 -16892 41346
rect -16948 41292 -16892 41294
rect -16788 41346 -16732 41348
rect -16788 41294 -16786 41346
rect -16786 41294 -16734 41346
rect -16734 41294 -16732 41346
rect -16788 41292 -16732 41294
rect -16628 41346 -16572 41348
rect -16628 41294 -16626 41346
rect -16626 41294 -16574 41346
rect -16574 41294 -16572 41346
rect -16628 41292 -16572 41294
rect -16468 41346 -16412 41348
rect -16468 41294 -16466 41346
rect -16466 41294 -16414 41346
rect -16414 41294 -16412 41346
rect -16468 41292 -16412 41294
rect -16308 41346 -16252 41348
rect -16308 41294 -16306 41346
rect -16306 41294 -16254 41346
rect -16254 41294 -16252 41346
rect -16308 41292 -16252 41294
rect -16148 41346 -16092 41348
rect -16148 41294 -16146 41346
rect -16146 41294 -16094 41346
rect -16094 41294 -16092 41346
rect -16148 41292 -16092 41294
rect -15988 41346 -15932 41348
rect -15988 41294 -15986 41346
rect -15986 41294 -15934 41346
rect -15934 41294 -15932 41346
rect -15988 41292 -15932 41294
rect -15828 41346 -15772 41348
rect -15828 41294 -15826 41346
rect -15826 41294 -15774 41346
rect -15774 41294 -15772 41346
rect -15828 41292 -15772 41294
rect -15668 41346 -15612 41348
rect -15668 41294 -15666 41346
rect -15666 41294 -15614 41346
rect -15614 41294 -15612 41346
rect -15668 41292 -15612 41294
rect -15508 41346 -15452 41348
rect -15508 41294 -15506 41346
rect -15506 41294 -15454 41346
rect -15454 41294 -15452 41346
rect -15508 41292 -15452 41294
rect -15348 41346 -15292 41348
rect -15348 41294 -15346 41346
rect -15346 41294 -15294 41346
rect -15294 41294 -15292 41346
rect -15348 41292 -15292 41294
rect -15188 41346 -15132 41348
rect -15188 41294 -15186 41346
rect -15186 41294 -15134 41346
rect -15134 41294 -15132 41346
rect -15188 41292 -15132 41294
rect -15028 41346 -14972 41348
rect -15028 41294 -15026 41346
rect -15026 41294 -14974 41346
rect -14974 41294 -14972 41346
rect -15028 41292 -14972 41294
rect -14868 41346 -14812 41348
rect -14868 41294 -14866 41346
rect -14866 41294 -14814 41346
rect -14814 41294 -14812 41346
rect -14868 41292 -14812 41294
rect -14708 41346 -14652 41348
rect -14708 41294 -14706 41346
rect -14706 41294 -14654 41346
rect -14654 41294 -14652 41346
rect -14708 41292 -14652 41294
rect -14548 41346 -14492 41348
rect -14548 41294 -14546 41346
rect -14546 41294 -14494 41346
rect -14494 41294 -14492 41346
rect -14548 41292 -14492 41294
rect -14388 41346 -14332 41348
rect -14388 41294 -14386 41346
rect -14386 41294 -14334 41346
rect -14334 41294 -14332 41346
rect -14388 41292 -14332 41294
rect -14228 41346 -14172 41348
rect -14228 41294 -14226 41346
rect -14226 41294 -14174 41346
rect -14174 41294 -14172 41346
rect -14228 41292 -14172 41294
rect -14068 41346 -14012 41348
rect -14068 41294 -14066 41346
rect -14066 41294 -14014 41346
rect -14014 41294 -14012 41346
rect -14068 41292 -14012 41294
rect -13908 41346 -13852 41348
rect -13908 41294 -13906 41346
rect -13906 41294 -13854 41346
rect -13854 41294 -13852 41346
rect -13908 41292 -13852 41294
rect -13748 41346 -13692 41348
rect -13748 41294 -13746 41346
rect -13746 41294 -13694 41346
rect -13694 41294 -13692 41346
rect -13748 41292 -13692 41294
rect -13588 41346 -13532 41348
rect -13588 41294 -13586 41346
rect -13586 41294 -13534 41346
rect -13534 41294 -13532 41346
rect -13588 41292 -13532 41294
rect -13428 41346 -13372 41348
rect -13428 41294 -13426 41346
rect -13426 41294 -13374 41346
rect -13374 41294 -13372 41346
rect -13428 41292 -13372 41294
rect -13268 41346 -13212 41348
rect -13268 41294 -13266 41346
rect -13266 41294 -13214 41346
rect -13214 41294 -13212 41346
rect -13268 41292 -13212 41294
rect -13108 41346 -13052 41348
rect -13108 41294 -13106 41346
rect -13106 41294 -13054 41346
rect -13054 41294 -13052 41346
rect -13108 41292 -13052 41294
rect -12948 41346 -12892 41348
rect -12948 41294 -12946 41346
rect -12946 41294 -12894 41346
rect -12894 41294 -12892 41346
rect -12948 41292 -12892 41294
rect -12788 41346 -12732 41348
rect -12788 41294 -12786 41346
rect -12786 41294 -12734 41346
rect -12734 41294 -12732 41346
rect -12788 41292 -12732 41294
rect -12628 41346 -12572 41348
rect -12628 41294 -12626 41346
rect -12626 41294 -12574 41346
rect -12574 41294 -12572 41346
rect -12628 41292 -12572 41294
rect -12468 41346 -12412 41348
rect -12468 41294 -12466 41346
rect -12466 41294 -12414 41346
rect -12414 41294 -12412 41346
rect -12468 41292 -12412 41294
rect -12308 41346 -12252 41348
rect -12308 41294 -12306 41346
rect -12306 41294 -12254 41346
rect -12254 41294 -12252 41346
rect -12308 41292 -12252 41294
rect -11348 41346 -11292 41348
rect -11348 41294 -11346 41346
rect -11346 41294 -11294 41346
rect -11294 41294 -11292 41346
rect -11348 41292 -11292 41294
rect -11188 41346 -11132 41348
rect -11188 41294 -11186 41346
rect -11186 41294 -11134 41346
rect -11134 41294 -11132 41346
rect -11188 41292 -11132 41294
rect -11028 41346 -10972 41348
rect -11028 41294 -11026 41346
rect -11026 41294 -10974 41346
rect -10974 41294 -10972 41346
rect -11028 41292 -10972 41294
rect -10868 41346 -10812 41348
rect -10868 41294 -10866 41346
rect -10866 41294 -10814 41346
rect -10814 41294 -10812 41346
rect -10868 41292 -10812 41294
rect -10708 41346 -10652 41348
rect -10708 41294 -10706 41346
rect -10706 41294 -10654 41346
rect -10654 41294 -10652 41346
rect -10708 41292 -10652 41294
rect -10548 41346 -10492 41348
rect -10548 41294 -10546 41346
rect -10546 41294 -10494 41346
rect -10494 41294 -10492 41346
rect -10548 41292 -10492 41294
rect -10388 41346 -10332 41348
rect -10388 41294 -10386 41346
rect -10386 41294 -10334 41346
rect -10334 41294 -10332 41346
rect -10388 41292 -10332 41294
rect -10228 41346 -10172 41348
rect -10228 41294 -10226 41346
rect -10226 41294 -10174 41346
rect -10174 41294 -10172 41346
rect -10228 41292 -10172 41294
rect -10068 41346 -10012 41348
rect -10068 41294 -10066 41346
rect -10066 41294 -10014 41346
rect -10014 41294 -10012 41346
rect -10068 41292 -10012 41294
rect -9908 41346 -9852 41348
rect -9908 41294 -9906 41346
rect -9906 41294 -9854 41346
rect -9854 41294 -9852 41346
rect -9908 41292 -9852 41294
rect -9748 41346 -9692 41348
rect -9748 41294 -9746 41346
rect -9746 41294 -9694 41346
rect -9694 41294 -9692 41346
rect -9748 41292 -9692 41294
rect -9588 41346 -9532 41348
rect -9588 41294 -9586 41346
rect -9586 41294 -9534 41346
rect -9534 41294 -9532 41346
rect -9588 41292 -9532 41294
rect -9428 41346 -9372 41348
rect -9428 41294 -9426 41346
rect -9426 41294 -9374 41346
rect -9374 41294 -9372 41346
rect -9428 41292 -9372 41294
rect -9268 41346 -9212 41348
rect -9268 41294 -9266 41346
rect -9266 41294 -9214 41346
rect -9214 41294 -9212 41346
rect -9268 41292 -9212 41294
rect -9108 41346 -9052 41348
rect -9108 41294 -9106 41346
rect -9106 41294 -9054 41346
rect -9054 41294 -9052 41346
rect -9108 41292 -9052 41294
rect -8948 41346 -8892 41348
rect -8948 41294 -8946 41346
rect -8946 41294 -8894 41346
rect -8894 41294 -8892 41346
rect -8948 41292 -8892 41294
rect -8788 41346 -8732 41348
rect -8788 41294 -8786 41346
rect -8786 41294 -8734 41346
rect -8734 41294 -8732 41346
rect -8788 41292 -8732 41294
rect -8628 41346 -8572 41348
rect -8628 41294 -8626 41346
rect -8626 41294 -8574 41346
rect -8574 41294 -8572 41346
rect -8628 41292 -8572 41294
rect -8468 41346 -8412 41348
rect -8468 41294 -8466 41346
rect -8466 41294 -8414 41346
rect -8414 41294 -8412 41346
rect -8468 41292 -8412 41294
rect -8308 41346 -8252 41348
rect -8308 41294 -8306 41346
rect -8306 41294 -8254 41346
rect -8254 41294 -8252 41346
rect -8308 41292 -8252 41294
rect -8148 41346 -8092 41348
rect -8148 41294 -8146 41346
rect -8146 41294 -8094 41346
rect -8094 41294 -8092 41346
rect -8148 41292 -8092 41294
rect -7988 41346 -7932 41348
rect -7988 41294 -7986 41346
rect -7986 41294 -7934 41346
rect -7934 41294 -7932 41346
rect -7988 41292 -7932 41294
rect -7828 41346 -7772 41348
rect -7828 41294 -7826 41346
rect -7826 41294 -7774 41346
rect -7774 41294 -7772 41346
rect -7828 41292 -7772 41294
rect -7668 41346 -7612 41348
rect -7668 41294 -7666 41346
rect -7666 41294 -7614 41346
rect -7614 41294 -7612 41346
rect -7668 41292 -7612 41294
rect -7508 41346 -7452 41348
rect -7508 41294 -7506 41346
rect -7506 41294 -7454 41346
rect -7454 41294 -7452 41346
rect -7508 41292 -7452 41294
rect -7348 41346 -7292 41348
rect -7348 41294 -7346 41346
rect -7346 41294 -7294 41346
rect -7294 41294 -7292 41346
rect -7348 41292 -7292 41294
rect -7188 41346 -7132 41348
rect -7188 41294 -7186 41346
rect -7186 41294 -7134 41346
rect -7134 41294 -7132 41346
rect -7188 41292 -7132 41294
rect -7028 41346 -6972 41348
rect -7028 41294 -7026 41346
rect -7026 41294 -6974 41346
rect -6974 41294 -6972 41346
rect -7028 41292 -6972 41294
rect -6868 41346 -6812 41348
rect -6868 41294 -6866 41346
rect -6866 41294 -6814 41346
rect -6814 41294 -6812 41346
rect -6868 41292 -6812 41294
rect -6708 41346 -6652 41348
rect -6708 41294 -6706 41346
rect -6706 41294 -6654 41346
rect -6654 41294 -6652 41346
rect -6708 41292 -6652 41294
rect -6548 41346 -6492 41348
rect -6548 41294 -6546 41346
rect -6546 41294 -6494 41346
rect -6494 41294 -6492 41346
rect -6548 41292 -6492 41294
rect -6388 41346 -6332 41348
rect -6388 41294 -6386 41346
rect -6386 41294 -6334 41346
rect -6334 41294 -6332 41346
rect -6388 41292 -6332 41294
rect -6228 41346 -6172 41348
rect -6228 41294 -6226 41346
rect -6226 41294 -6174 41346
rect -6174 41294 -6172 41346
rect -6228 41292 -6172 41294
rect -6068 41346 -6012 41348
rect -6068 41294 -6066 41346
rect -6066 41294 -6014 41346
rect -6014 41294 -6012 41346
rect -6068 41292 -6012 41294
rect -5908 41346 -5852 41348
rect -5908 41294 -5906 41346
rect -5906 41294 -5854 41346
rect -5854 41294 -5852 41346
rect -5908 41292 -5852 41294
rect -5748 41346 -5692 41348
rect -5748 41294 -5746 41346
rect -5746 41294 -5694 41346
rect -5694 41294 -5692 41346
rect -5748 41292 -5692 41294
rect -5588 41346 -5532 41348
rect -5588 41294 -5586 41346
rect -5586 41294 -5534 41346
rect -5534 41294 -5532 41346
rect -5588 41292 -5532 41294
rect -5428 41346 -5372 41348
rect -5428 41294 -5426 41346
rect -5426 41294 -5374 41346
rect -5374 41294 -5372 41346
rect -5428 41292 -5372 41294
rect -5268 41346 -5212 41348
rect -5268 41294 -5266 41346
rect -5266 41294 -5214 41346
rect -5214 41294 -5212 41346
rect -5268 41292 -5212 41294
rect -5108 41346 -5052 41348
rect -5108 41294 -5106 41346
rect -5106 41294 -5054 41346
rect -5054 41294 -5052 41346
rect -5108 41292 -5052 41294
rect -4948 41346 -4892 41348
rect -4948 41294 -4946 41346
rect -4946 41294 -4894 41346
rect -4894 41294 -4892 41346
rect -4948 41292 -4892 41294
rect -4788 41346 -4732 41348
rect -4788 41294 -4786 41346
rect -4786 41294 -4734 41346
rect -4734 41294 -4732 41346
rect -4788 41292 -4732 41294
rect -4628 41346 -4572 41348
rect -4628 41294 -4626 41346
rect -4626 41294 -4574 41346
rect -4574 41294 -4572 41346
rect -4628 41292 -4572 41294
rect -4468 41346 -4412 41348
rect -4468 41294 -4466 41346
rect -4466 41294 -4414 41346
rect -4414 41294 -4412 41346
rect -4468 41292 -4412 41294
rect -4308 41346 -4252 41348
rect -4308 41294 -4306 41346
rect -4306 41294 -4254 41346
rect -4254 41294 -4252 41346
rect -4308 41292 -4252 41294
rect -4148 41346 -4092 41348
rect -4148 41294 -4146 41346
rect -4146 41294 -4094 41346
rect -4094 41294 -4092 41346
rect -4148 41292 -4092 41294
rect -3988 41346 -3932 41348
rect -3988 41294 -3986 41346
rect -3986 41294 -3934 41346
rect -3934 41294 -3932 41346
rect -3988 41292 -3932 41294
rect -3828 41292 -3772 41348
rect -3668 41346 -3612 41348
rect -3668 41294 -3666 41346
rect -3666 41294 -3614 41346
rect -3614 41294 -3612 41346
rect -3668 41292 -3612 41294
rect -3508 41346 -3452 41348
rect -3508 41294 -3506 41346
rect -3506 41294 -3454 41346
rect -3454 41294 -3452 41346
rect -3508 41292 -3452 41294
rect 41052 41346 41108 41348
rect 41052 41294 41054 41346
rect 41054 41294 41106 41346
rect 41106 41294 41108 41346
rect 41052 41292 41108 41294
rect 41212 41346 41268 41348
rect 41212 41294 41214 41346
rect 41214 41294 41266 41346
rect 41266 41294 41268 41346
rect 41212 41292 41268 41294
rect 41372 41346 41428 41348
rect 41372 41294 41374 41346
rect 41374 41294 41426 41346
rect 41426 41294 41428 41346
rect 41372 41292 41428 41294
rect 41532 41346 41588 41348
rect 41532 41294 41534 41346
rect 41534 41294 41586 41346
rect 41586 41294 41588 41346
rect 41532 41292 41588 41294
rect 41692 41346 41748 41348
rect 41692 41294 41694 41346
rect 41694 41294 41746 41346
rect 41746 41294 41748 41346
rect 41692 41292 41748 41294
rect 41852 41346 41908 41348
rect 41852 41294 41854 41346
rect 41854 41294 41906 41346
rect 41906 41294 41908 41346
rect 41852 41292 41908 41294
rect 42012 41346 42068 41348
rect 42012 41294 42014 41346
rect 42014 41294 42066 41346
rect 42066 41294 42068 41346
rect 42012 41292 42068 41294
rect 42172 41346 42228 41348
rect 42172 41294 42174 41346
rect 42174 41294 42226 41346
rect 42226 41294 42228 41346
rect 42172 41292 42228 41294
rect 42332 41346 42388 41348
rect 42332 41294 42334 41346
rect 42334 41294 42386 41346
rect 42386 41294 42388 41346
rect 42332 41292 42388 41294
rect 42492 41346 42548 41348
rect 42492 41294 42494 41346
rect 42494 41294 42546 41346
rect 42546 41294 42548 41346
rect 42492 41292 42548 41294
rect 42652 41346 42708 41348
rect 42652 41294 42654 41346
rect 42654 41294 42706 41346
rect 42706 41294 42708 41346
rect 42652 41292 42708 41294
rect 42812 41346 42868 41348
rect 42812 41294 42814 41346
rect 42814 41294 42866 41346
rect 42866 41294 42868 41346
rect 42812 41292 42868 41294
rect 42972 41346 43028 41348
rect 42972 41294 42974 41346
rect 42974 41294 43026 41346
rect 43026 41294 43028 41346
rect 42972 41292 43028 41294
rect 43132 41346 43188 41348
rect 43132 41294 43134 41346
rect 43134 41294 43186 41346
rect 43186 41294 43188 41346
rect 43132 41292 43188 41294
rect -33108 41026 -33052 41028
rect -33108 40974 -33106 41026
rect -33106 40974 -33054 41026
rect -33054 40974 -33052 41026
rect -33108 40972 -33052 40974
rect -32948 41026 -32892 41028
rect -32948 40974 -32946 41026
rect -32946 40974 -32894 41026
rect -32894 40974 -32892 41026
rect -32948 40972 -32892 40974
rect -32788 41026 -32732 41028
rect -32788 40974 -32786 41026
rect -32786 40974 -32734 41026
rect -32734 40974 -32732 41026
rect -32788 40972 -32732 40974
rect -32628 41026 -32572 41028
rect -32628 40974 -32626 41026
rect -32626 40974 -32574 41026
rect -32574 40974 -32572 41026
rect -32628 40972 -32572 40974
rect -32468 41026 -32412 41028
rect -32468 40974 -32466 41026
rect -32466 40974 -32414 41026
rect -32414 40974 -32412 41026
rect -32468 40972 -32412 40974
rect -32308 41026 -32252 41028
rect -32308 40974 -32306 41026
rect -32306 40974 -32254 41026
rect -32254 40974 -32252 41026
rect -32308 40972 -32252 40974
rect -32148 41026 -32092 41028
rect -32148 40974 -32146 41026
rect -32146 40974 -32094 41026
rect -32094 40974 -32092 41026
rect -32148 40972 -32092 40974
rect -31988 41026 -31932 41028
rect -31988 40974 -31986 41026
rect -31986 40974 -31934 41026
rect -31934 40974 -31932 41026
rect -31988 40972 -31932 40974
rect -31828 41026 -31772 41028
rect -31828 40974 -31826 41026
rect -31826 40974 -31774 41026
rect -31774 40974 -31772 41026
rect -31828 40972 -31772 40974
rect -31668 41026 -31612 41028
rect -31668 40974 -31666 41026
rect -31666 40974 -31614 41026
rect -31614 40974 -31612 41026
rect -31668 40972 -31612 40974
rect -31508 41026 -31452 41028
rect -31508 40974 -31506 41026
rect -31506 40974 -31454 41026
rect -31454 40974 -31452 41026
rect -31508 40972 -31452 40974
rect -31348 41026 -31292 41028
rect -31348 40974 -31346 41026
rect -31346 40974 -31294 41026
rect -31294 40974 -31292 41026
rect -31348 40972 -31292 40974
rect -31188 41026 -31132 41028
rect -31188 40974 -31186 41026
rect -31186 40974 -31134 41026
rect -31134 40974 -31132 41026
rect -31188 40972 -31132 40974
rect -29908 41026 -29852 41028
rect -29908 40974 -29906 41026
rect -29906 40974 -29854 41026
rect -29854 40974 -29852 41026
rect -29908 40972 -29852 40974
rect -29748 41026 -29692 41028
rect -29748 40974 -29746 41026
rect -29746 40974 -29694 41026
rect -29694 40974 -29692 41026
rect -29748 40972 -29692 40974
rect -29588 41026 -29532 41028
rect -29588 40974 -29586 41026
rect -29586 40974 -29534 41026
rect -29534 40974 -29532 41026
rect -29588 40972 -29532 40974
rect -29428 41026 -29372 41028
rect -29428 40974 -29426 41026
rect -29426 40974 -29374 41026
rect -29374 40974 -29372 41026
rect -29428 40972 -29372 40974
rect -29268 41026 -29212 41028
rect -29268 40974 -29266 41026
rect -29266 40974 -29214 41026
rect -29214 40974 -29212 41026
rect -29268 40972 -29212 40974
rect -29108 41026 -29052 41028
rect -29108 40974 -29106 41026
rect -29106 40974 -29054 41026
rect -29054 40974 -29052 41026
rect -29108 40972 -29052 40974
rect -28948 41026 -28892 41028
rect -28948 40974 -28946 41026
rect -28946 40974 -28894 41026
rect -28894 40974 -28892 41026
rect -28948 40972 -28892 40974
rect -28788 41026 -28732 41028
rect -28788 40974 -28786 41026
rect -28786 40974 -28734 41026
rect -28734 40974 -28732 41026
rect -28788 40972 -28732 40974
rect -28628 41026 -28572 41028
rect -28628 40974 -28626 41026
rect -28626 40974 -28574 41026
rect -28574 40974 -28572 41026
rect -28628 40972 -28572 40974
rect -28468 41026 -28412 41028
rect -28468 40974 -28466 41026
rect -28466 40974 -28414 41026
rect -28414 40974 -28412 41026
rect -28468 40972 -28412 40974
rect -28308 41026 -28252 41028
rect -28308 40974 -28306 41026
rect -28306 40974 -28254 41026
rect -28254 40974 -28252 41026
rect -28308 40972 -28252 40974
rect -28148 41026 -28092 41028
rect -28148 40974 -28146 41026
rect -28146 40974 -28094 41026
rect -28094 40974 -28092 41026
rect -28148 40972 -28092 40974
rect -27988 41026 -27932 41028
rect -27988 40974 -27986 41026
rect -27986 40974 -27934 41026
rect -27934 40974 -27932 41026
rect -27988 40972 -27932 40974
rect -27828 41026 -27772 41028
rect -27828 40974 -27826 41026
rect -27826 40974 -27774 41026
rect -27774 40974 -27772 41026
rect -27828 40972 -27772 40974
rect -27668 41026 -27612 41028
rect -27668 40974 -27666 41026
rect -27666 40974 -27614 41026
rect -27614 40974 -27612 41026
rect -27668 40972 -27612 40974
rect -27508 41026 -27452 41028
rect -27508 40974 -27506 41026
rect -27506 40974 -27454 41026
rect -27454 40974 -27452 41026
rect -27508 40972 -27452 40974
rect -27348 41026 -27292 41028
rect -27348 40974 -27346 41026
rect -27346 40974 -27294 41026
rect -27294 40974 -27292 41026
rect -27348 40972 -27292 40974
rect -27188 41026 -27132 41028
rect -27188 40974 -27186 41026
rect -27186 40974 -27134 41026
rect -27134 40974 -27132 41026
rect -27188 40972 -27132 40974
rect -27028 41026 -26972 41028
rect -27028 40974 -27026 41026
rect -27026 40974 -26974 41026
rect -26974 40974 -26972 41026
rect -27028 40972 -26972 40974
rect -26868 41026 -26812 41028
rect -26868 40974 -26866 41026
rect -26866 40974 -26814 41026
rect -26814 40974 -26812 41026
rect -26868 40972 -26812 40974
rect -26708 41026 -26652 41028
rect -26708 40974 -26706 41026
rect -26706 40974 -26654 41026
rect -26654 40974 -26652 41026
rect -26708 40972 -26652 40974
rect -26548 41026 -26492 41028
rect -26548 40974 -26546 41026
rect -26546 40974 -26494 41026
rect -26494 40974 -26492 41026
rect -26548 40972 -26492 40974
rect -26388 41026 -26332 41028
rect -26388 40974 -26386 41026
rect -26386 40974 -26334 41026
rect -26334 40974 -26332 41026
rect -26388 40972 -26332 40974
rect -26228 41026 -26172 41028
rect -26228 40974 -26226 41026
rect -26226 40974 -26174 41026
rect -26174 40974 -26172 41026
rect -26228 40972 -26172 40974
rect -26068 41026 -26012 41028
rect -26068 40974 -26066 41026
rect -26066 40974 -26014 41026
rect -26014 40974 -26012 41026
rect -26068 40972 -26012 40974
rect -25908 41026 -25852 41028
rect -25908 40974 -25906 41026
rect -25906 40974 -25854 41026
rect -25854 40974 -25852 41026
rect -25908 40972 -25852 40974
rect -25748 41026 -25692 41028
rect -25748 40974 -25746 41026
rect -25746 40974 -25694 41026
rect -25694 40974 -25692 41026
rect -25748 40972 -25692 40974
rect -25588 41026 -25532 41028
rect -25588 40974 -25586 41026
rect -25586 40974 -25534 41026
rect -25534 40974 -25532 41026
rect -25588 40972 -25532 40974
rect -25428 41026 -25372 41028
rect -25428 40974 -25426 41026
rect -25426 40974 -25374 41026
rect -25374 40974 -25372 41026
rect -25428 40972 -25372 40974
rect -25268 41026 -25212 41028
rect -25268 40974 -25266 41026
rect -25266 40974 -25214 41026
rect -25214 40974 -25212 41026
rect -25268 40972 -25212 40974
rect -25108 41026 -25052 41028
rect -25108 40974 -25106 41026
rect -25106 40974 -25054 41026
rect -25054 40974 -25052 41026
rect -25108 40972 -25052 40974
rect -24948 41026 -24892 41028
rect -24948 40974 -24946 41026
rect -24946 40974 -24894 41026
rect -24894 40974 -24892 41026
rect -24948 40972 -24892 40974
rect -24788 41026 -24732 41028
rect -24788 40974 -24786 41026
rect -24786 40974 -24734 41026
rect -24734 40974 -24732 41026
rect -24788 40972 -24732 40974
rect -24628 41026 -24572 41028
rect -24628 40974 -24626 41026
rect -24626 40974 -24574 41026
rect -24574 40974 -24572 41026
rect -24628 40972 -24572 40974
rect -24468 41026 -24412 41028
rect -24468 40974 -24466 41026
rect -24466 40974 -24414 41026
rect -24414 40974 -24412 41026
rect -24468 40972 -24412 40974
rect -24308 41026 -24252 41028
rect -24308 40974 -24306 41026
rect -24306 40974 -24254 41026
rect -24254 40974 -24252 41026
rect -24308 40972 -24252 40974
rect -24148 41026 -24092 41028
rect -24148 40974 -24146 41026
rect -24146 40974 -24094 41026
rect -24094 40974 -24092 41026
rect -24148 40972 -24092 40974
rect -23988 41026 -23932 41028
rect -23988 40974 -23986 41026
rect -23986 40974 -23934 41026
rect -23934 40974 -23932 41026
rect -23988 40972 -23932 40974
rect -23828 41026 -23772 41028
rect -23828 40974 -23826 41026
rect -23826 40974 -23774 41026
rect -23774 40974 -23772 41026
rect -23828 40972 -23772 40974
rect -23668 41026 -23612 41028
rect -23668 40974 -23666 41026
rect -23666 40974 -23614 41026
rect -23614 40974 -23612 41026
rect -23668 40972 -23612 40974
rect -23508 41026 -23452 41028
rect -23508 40974 -23506 41026
rect -23506 40974 -23454 41026
rect -23454 40974 -23452 41026
rect -23508 40972 -23452 40974
rect -23348 41026 -23292 41028
rect -23348 40974 -23346 41026
rect -23346 40974 -23294 41026
rect -23294 40974 -23292 41026
rect -23348 40972 -23292 40974
rect -23188 41026 -23132 41028
rect -23188 40974 -23186 41026
rect -23186 40974 -23134 41026
rect -23134 40974 -23132 41026
rect -23188 40972 -23132 40974
rect -23028 41026 -22972 41028
rect -23028 40974 -23026 41026
rect -23026 40974 -22974 41026
rect -22974 40974 -22972 41026
rect -23028 40972 -22972 40974
rect -22868 41026 -22812 41028
rect -22868 40974 -22866 41026
rect -22866 40974 -22814 41026
rect -22814 40974 -22812 41026
rect -22868 40972 -22812 40974
rect -22708 41026 -22652 41028
rect -22708 40974 -22706 41026
rect -22706 40974 -22654 41026
rect -22654 40974 -22652 41026
rect -22708 40972 -22652 40974
rect -22548 41026 -22492 41028
rect -22548 40974 -22546 41026
rect -22546 40974 -22494 41026
rect -22494 40974 -22492 41026
rect -22548 40972 -22492 40974
rect -22388 41026 -22332 41028
rect -22388 40974 -22386 41026
rect -22386 40974 -22334 41026
rect -22334 40974 -22332 41026
rect -22388 40972 -22332 40974
rect -22228 41026 -22172 41028
rect -22228 40974 -22226 41026
rect -22226 40974 -22174 41026
rect -22174 40974 -22172 41026
rect -22228 40972 -22172 40974
rect -22068 41026 -22012 41028
rect -22068 40974 -22066 41026
rect -22066 40974 -22014 41026
rect -22014 40974 -22012 41026
rect -22068 40972 -22012 40974
rect -21908 41026 -21852 41028
rect -21908 40974 -21906 41026
rect -21906 40974 -21854 41026
rect -21854 40974 -21852 41026
rect -21908 40972 -21852 40974
rect -21748 41026 -21692 41028
rect -21748 40974 -21746 41026
rect -21746 40974 -21694 41026
rect -21694 40974 -21692 41026
rect -21748 40972 -21692 40974
rect -21588 41026 -21532 41028
rect -21588 40974 -21586 41026
rect -21586 40974 -21534 41026
rect -21534 40974 -21532 41026
rect -21588 40972 -21532 40974
rect -21428 41026 -21372 41028
rect -21428 40974 -21426 41026
rect -21426 40974 -21374 41026
rect -21374 40974 -21372 41026
rect -21428 40972 -21372 40974
rect -21268 41026 -21212 41028
rect -21268 40974 -21266 41026
rect -21266 40974 -21214 41026
rect -21214 40974 -21212 41026
rect -21268 40972 -21212 40974
rect -21108 41026 -21052 41028
rect -21108 40974 -21106 41026
rect -21106 40974 -21054 41026
rect -21054 40974 -21052 41026
rect -21108 40972 -21052 40974
rect -20948 41026 -20892 41028
rect -20948 40974 -20946 41026
rect -20946 40974 -20894 41026
rect -20894 40974 -20892 41026
rect -20948 40972 -20892 40974
rect -20788 41026 -20732 41028
rect -20788 40974 -20786 41026
rect -20786 40974 -20734 41026
rect -20734 40974 -20732 41026
rect -20788 40972 -20732 40974
rect -20628 41026 -20572 41028
rect -20628 40974 -20626 41026
rect -20626 40974 -20574 41026
rect -20574 40974 -20572 41026
rect -20628 40972 -20572 40974
rect -20468 41026 -20412 41028
rect -20468 40974 -20466 41026
rect -20466 40974 -20414 41026
rect -20414 40974 -20412 41026
rect -20468 40972 -20412 40974
rect -20308 41026 -20252 41028
rect -20308 40974 -20306 41026
rect -20306 40974 -20254 41026
rect -20254 40974 -20252 41026
rect -20308 40972 -20252 40974
rect -20148 41026 -20092 41028
rect -20148 40974 -20146 41026
rect -20146 40974 -20094 41026
rect -20094 40974 -20092 41026
rect -20148 40972 -20092 40974
rect -19988 41026 -19932 41028
rect -19988 40974 -19986 41026
rect -19986 40974 -19934 41026
rect -19934 40974 -19932 41026
rect -19988 40972 -19932 40974
rect -19828 41026 -19772 41028
rect -19828 40974 -19826 41026
rect -19826 40974 -19774 41026
rect -19774 40974 -19772 41026
rect -19828 40972 -19772 40974
rect -19668 41026 -19612 41028
rect -19668 40974 -19666 41026
rect -19666 40974 -19614 41026
rect -19614 40974 -19612 41026
rect -19668 40972 -19612 40974
rect -19508 41026 -19452 41028
rect -19508 40974 -19506 41026
rect -19506 40974 -19454 41026
rect -19454 40974 -19452 41026
rect -19508 40972 -19452 40974
rect -19348 41026 -19292 41028
rect -19348 40974 -19346 41026
rect -19346 40974 -19294 41026
rect -19294 40974 -19292 41026
rect -19348 40972 -19292 40974
rect -19188 41026 -19132 41028
rect -19188 40974 -19186 41026
rect -19186 40974 -19134 41026
rect -19134 40974 -19132 41026
rect -19188 40972 -19132 40974
rect -19028 41026 -18972 41028
rect -19028 40974 -19026 41026
rect -19026 40974 -18974 41026
rect -18974 40974 -18972 41026
rect -19028 40972 -18972 40974
rect -18868 41026 -18812 41028
rect -18868 40974 -18866 41026
rect -18866 40974 -18814 41026
rect -18814 40974 -18812 41026
rect -18868 40972 -18812 40974
rect -18708 41026 -18652 41028
rect -18708 40974 -18706 41026
rect -18706 40974 -18654 41026
rect -18654 40974 -18652 41026
rect -18708 40972 -18652 40974
rect -18548 41026 -18492 41028
rect -18548 40974 -18546 41026
rect -18546 40974 -18494 41026
rect -18494 40974 -18492 41026
rect -18548 40972 -18492 40974
rect -18388 41026 -18332 41028
rect -18388 40974 -18386 41026
rect -18386 40974 -18334 41026
rect -18334 40974 -18332 41026
rect -18388 40972 -18332 40974
rect -18228 41026 -18172 41028
rect -18228 40974 -18226 41026
rect -18226 40974 -18174 41026
rect -18174 40974 -18172 41026
rect -18228 40972 -18172 40974
rect -18068 41026 -18012 41028
rect -18068 40974 -18066 41026
rect -18066 40974 -18014 41026
rect -18014 40974 -18012 41026
rect -18068 40972 -18012 40974
rect -17908 41026 -17852 41028
rect -17908 40974 -17906 41026
rect -17906 40974 -17854 41026
rect -17854 40974 -17852 41026
rect -17908 40972 -17852 40974
rect -17748 41026 -17692 41028
rect -17748 40974 -17746 41026
rect -17746 40974 -17694 41026
rect -17694 40974 -17692 41026
rect -17748 40972 -17692 40974
rect -17588 41026 -17532 41028
rect -17588 40974 -17586 41026
rect -17586 40974 -17534 41026
rect -17534 40974 -17532 41026
rect -17588 40972 -17532 40974
rect -17428 41026 -17372 41028
rect -17428 40974 -17426 41026
rect -17426 40974 -17374 41026
rect -17374 40974 -17372 41026
rect -17428 40972 -17372 40974
rect -17268 41026 -17212 41028
rect -17268 40974 -17266 41026
rect -17266 40974 -17214 41026
rect -17214 40974 -17212 41026
rect -17268 40972 -17212 40974
rect -17108 41026 -17052 41028
rect -17108 40974 -17106 41026
rect -17106 40974 -17054 41026
rect -17054 40974 -17052 41026
rect -17108 40972 -17052 40974
rect -16948 41026 -16892 41028
rect -16948 40974 -16946 41026
rect -16946 40974 -16894 41026
rect -16894 40974 -16892 41026
rect -16948 40972 -16892 40974
rect -16788 41026 -16732 41028
rect -16788 40974 -16786 41026
rect -16786 40974 -16734 41026
rect -16734 40974 -16732 41026
rect -16788 40972 -16732 40974
rect -16628 41026 -16572 41028
rect -16628 40974 -16626 41026
rect -16626 40974 -16574 41026
rect -16574 40974 -16572 41026
rect -16628 40972 -16572 40974
rect -16468 41026 -16412 41028
rect -16468 40974 -16466 41026
rect -16466 40974 -16414 41026
rect -16414 40974 -16412 41026
rect -16468 40972 -16412 40974
rect -16308 41026 -16252 41028
rect -16308 40974 -16306 41026
rect -16306 40974 -16254 41026
rect -16254 40974 -16252 41026
rect -16308 40972 -16252 40974
rect -16148 41026 -16092 41028
rect -16148 40974 -16146 41026
rect -16146 40974 -16094 41026
rect -16094 40974 -16092 41026
rect -16148 40972 -16092 40974
rect -15988 41026 -15932 41028
rect -15988 40974 -15986 41026
rect -15986 40974 -15934 41026
rect -15934 40974 -15932 41026
rect -15988 40972 -15932 40974
rect -15828 41026 -15772 41028
rect -15828 40974 -15826 41026
rect -15826 40974 -15774 41026
rect -15774 40974 -15772 41026
rect -15828 40972 -15772 40974
rect -15668 41026 -15612 41028
rect -15668 40974 -15666 41026
rect -15666 40974 -15614 41026
rect -15614 40974 -15612 41026
rect -15668 40972 -15612 40974
rect -15508 41026 -15452 41028
rect -15508 40974 -15506 41026
rect -15506 40974 -15454 41026
rect -15454 40974 -15452 41026
rect -15508 40972 -15452 40974
rect -15348 41026 -15292 41028
rect -15348 40974 -15346 41026
rect -15346 40974 -15294 41026
rect -15294 40974 -15292 41026
rect -15348 40972 -15292 40974
rect -15188 41026 -15132 41028
rect -15188 40974 -15186 41026
rect -15186 40974 -15134 41026
rect -15134 40974 -15132 41026
rect -15188 40972 -15132 40974
rect -15028 41026 -14972 41028
rect -15028 40974 -15026 41026
rect -15026 40974 -14974 41026
rect -14974 40974 -14972 41026
rect -15028 40972 -14972 40974
rect -14868 41026 -14812 41028
rect -14868 40974 -14866 41026
rect -14866 40974 -14814 41026
rect -14814 40974 -14812 41026
rect -14868 40972 -14812 40974
rect -14708 41026 -14652 41028
rect -14708 40974 -14706 41026
rect -14706 40974 -14654 41026
rect -14654 40974 -14652 41026
rect -14708 40972 -14652 40974
rect -14548 41026 -14492 41028
rect -14548 40974 -14546 41026
rect -14546 40974 -14494 41026
rect -14494 40974 -14492 41026
rect -14548 40972 -14492 40974
rect -14388 41026 -14332 41028
rect -14388 40974 -14386 41026
rect -14386 40974 -14334 41026
rect -14334 40974 -14332 41026
rect -14388 40972 -14332 40974
rect -14228 41026 -14172 41028
rect -14228 40974 -14226 41026
rect -14226 40974 -14174 41026
rect -14174 40974 -14172 41026
rect -14228 40972 -14172 40974
rect -14068 41026 -14012 41028
rect -14068 40974 -14066 41026
rect -14066 40974 -14014 41026
rect -14014 40974 -14012 41026
rect -14068 40972 -14012 40974
rect -13908 41026 -13852 41028
rect -13908 40974 -13906 41026
rect -13906 40974 -13854 41026
rect -13854 40974 -13852 41026
rect -13908 40972 -13852 40974
rect -13748 41026 -13692 41028
rect -13748 40974 -13746 41026
rect -13746 40974 -13694 41026
rect -13694 40974 -13692 41026
rect -13748 40972 -13692 40974
rect -13588 41026 -13532 41028
rect -13588 40974 -13586 41026
rect -13586 40974 -13534 41026
rect -13534 40974 -13532 41026
rect -13588 40972 -13532 40974
rect -13428 41026 -13372 41028
rect -13428 40974 -13426 41026
rect -13426 40974 -13374 41026
rect -13374 40974 -13372 41026
rect -13428 40972 -13372 40974
rect -13268 41026 -13212 41028
rect -13268 40974 -13266 41026
rect -13266 40974 -13214 41026
rect -13214 40974 -13212 41026
rect -13268 40972 -13212 40974
rect -13108 41026 -13052 41028
rect -13108 40974 -13106 41026
rect -13106 40974 -13054 41026
rect -13054 40974 -13052 41026
rect -13108 40972 -13052 40974
rect -12948 41026 -12892 41028
rect -12948 40974 -12946 41026
rect -12946 40974 -12894 41026
rect -12894 40974 -12892 41026
rect -12948 40972 -12892 40974
rect -12788 41026 -12732 41028
rect -12788 40974 -12786 41026
rect -12786 40974 -12734 41026
rect -12734 40974 -12732 41026
rect -12788 40972 -12732 40974
rect -12628 41026 -12572 41028
rect -12628 40974 -12626 41026
rect -12626 40974 -12574 41026
rect -12574 40974 -12572 41026
rect -12628 40972 -12572 40974
rect -12468 41026 -12412 41028
rect -12468 40974 -12466 41026
rect -12466 40974 -12414 41026
rect -12414 40974 -12412 41026
rect -12468 40972 -12412 40974
rect -12308 41026 -12252 41028
rect -12308 40974 -12306 41026
rect -12306 40974 -12254 41026
rect -12254 40974 -12252 41026
rect -12308 40972 -12252 40974
rect -11348 41026 -11292 41028
rect -11348 40974 -11346 41026
rect -11346 40974 -11294 41026
rect -11294 40974 -11292 41026
rect -11348 40972 -11292 40974
rect -11188 41026 -11132 41028
rect -11188 40974 -11186 41026
rect -11186 40974 -11134 41026
rect -11134 40974 -11132 41026
rect -11188 40972 -11132 40974
rect -11028 41026 -10972 41028
rect -11028 40974 -11026 41026
rect -11026 40974 -10974 41026
rect -10974 40974 -10972 41026
rect -11028 40972 -10972 40974
rect -10868 41026 -10812 41028
rect -10868 40974 -10866 41026
rect -10866 40974 -10814 41026
rect -10814 40974 -10812 41026
rect -10868 40972 -10812 40974
rect -10708 41026 -10652 41028
rect -10708 40974 -10706 41026
rect -10706 40974 -10654 41026
rect -10654 40974 -10652 41026
rect -10708 40972 -10652 40974
rect -10548 41026 -10492 41028
rect -10548 40974 -10546 41026
rect -10546 40974 -10494 41026
rect -10494 40974 -10492 41026
rect -10548 40972 -10492 40974
rect -10388 41026 -10332 41028
rect -10388 40974 -10386 41026
rect -10386 40974 -10334 41026
rect -10334 40974 -10332 41026
rect -10388 40972 -10332 40974
rect -10228 41026 -10172 41028
rect -10228 40974 -10226 41026
rect -10226 40974 -10174 41026
rect -10174 40974 -10172 41026
rect -10228 40972 -10172 40974
rect -10068 41026 -10012 41028
rect -10068 40974 -10066 41026
rect -10066 40974 -10014 41026
rect -10014 40974 -10012 41026
rect -10068 40972 -10012 40974
rect -9908 41026 -9852 41028
rect -9908 40974 -9906 41026
rect -9906 40974 -9854 41026
rect -9854 40974 -9852 41026
rect -9908 40972 -9852 40974
rect -9748 41026 -9692 41028
rect -9748 40974 -9746 41026
rect -9746 40974 -9694 41026
rect -9694 40974 -9692 41026
rect -9748 40972 -9692 40974
rect -9588 41026 -9532 41028
rect -9588 40974 -9586 41026
rect -9586 40974 -9534 41026
rect -9534 40974 -9532 41026
rect -9588 40972 -9532 40974
rect -9428 41026 -9372 41028
rect -9428 40974 -9426 41026
rect -9426 40974 -9374 41026
rect -9374 40974 -9372 41026
rect -9428 40972 -9372 40974
rect -9268 41026 -9212 41028
rect -9268 40974 -9266 41026
rect -9266 40974 -9214 41026
rect -9214 40974 -9212 41026
rect -9268 40972 -9212 40974
rect -9108 41026 -9052 41028
rect -9108 40974 -9106 41026
rect -9106 40974 -9054 41026
rect -9054 40974 -9052 41026
rect -9108 40972 -9052 40974
rect -8948 41026 -8892 41028
rect -8948 40974 -8946 41026
rect -8946 40974 -8894 41026
rect -8894 40974 -8892 41026
rect -8948 40972 -8892 40974
rect -8788 41026 -8732 41028
rect -8788 40974 -8786 41026
rect -8786 40974 -8734 41026
rect -8734 40974 -8732 41026
rect -8788 40972 -8732 40974
rect -8628 41026 -8572 41028
rect -8628 40974 -8626 41026
rect -8626 40974 -8574 41026
rect -8574 40974 -8572 41026
rect -8628 40972 -8572 40974
rect -8468 41026 -8412 41028
rect -8468 40974 -8466 41026
rect -8466 40974 -8414 41026
rect -8414 40974 -8412 41026
rect -8468 40972 -8412 40974
rect -8308 41026 -8252 41028
rect -8308 40974 -8306 41026
rect -8306 40974 -8254 41026
rect -8254 40974 -8252 41026
rect -8308 40972 -8252 40974
rect -8148 41026 -8092 41028
rect -8148 40974 -8146 41026
rect -8146 40974 -8094 41026
rect -8094 40974 -8092 41026
rect -8148 40972 -8092 40974
rect -7988 41026 -7932 41028
rect -7988 40974 -7986 41026
rect -7986 40974 -7934 41026
rect -7934 40974 -7932 41026
rect -7988 40972 -7932 40974
rect -7828 41026 -7772 41028
rect -7828 40974 -7826 41026
rect -7826 40974 -7774 41026
rect -7774 40974 -7772 41026
rect -7828 40972 -7772 40974
rect -7668 41026 -7612 41028
rect -7668 40974 -7666 41026
rect -7666 40974 -7614 41026
rect -7614 40974 -7612 41026
rect -7668 40972 -7612 40974
rect -7508 41026 -7452 41028
rect -7508 40974 -7506 41026
rect -7506 40974 -7454 41026
rect -7454 40974 -7452 41026
rect -7508 40972 -7452 40974
rect -7348 41026 -7292 41028
rect -7348 40974 -7346 41026
rect -7346 40974 -7294 41026
rect -7294 40974 -7292 41026
rect -7348 40972 -7292 40974
rect -7188 41026 -7132 41028
rect -7188 40974 -7186 41026
rect -7186 40974 -7134 41026
rect -7134 40974 -7132 41026
rect -7188 40972 -7132 40974
rect -7028 41026 -6972 41028
rect -7028 40974 -7026 41026
rect -7026 40974 -6974 41026
rect -6974 40974 -6972 41026
rect -7028 40972 -6972 40974
rect -6868 41026 -6812 41028
rect -6868 40974 -6866 41026
rect -6866 40974 -6814 41026
rect -6814 40974 -6812 41026
rect -6868 40972 -6812 40974
rect -6708 41026 -6652 41028
rect -6708 40974 -6706 41026
rect -6706 40974 -6654 41026
rect -6654 40974 -6652 41026
rect -6708 40972 -6652 40974
rect -6548 41026 -6492 41028
rect -6548 40974 -6546 41026
rect -6546 40974 -6494 41026
rect -6494 40974 -6492 41026
rect -6548 40972 -6492 40974
rect -6388 41026 -6332 41028
rect -6388 40974 -6386 41026
rect -6386 40974 -6334 41026
rect -6334 40974 -6332 41026
rect -6388 40972 -6332 40974
rect -6228 41026 -6172 41028
rect -6228 40974 -6226 41026
rect -6226 40974 -6174 41026
rect -6174 40974 -6172 41026
rect -6228 40972 -6172 40974
rect -6068 41026 -6012 41028
rect -6068 40974 -6066 41026
rect -6066 40974 -6014 41026
rect -6014 40974 -6012 41026
rect -6068 40972 -6012 40974
rect -5908 41026 -5852 41028
rect -5908 40974 -5906 41026
rect -5906 40974 -5854 41026
rect -5854 40974 -5852 41026
rect -5908 40972 -5852 40974
rect -5748 41026 -5692 41028
rect -5748 40974 -5746 41026
rect -5746 40974 -5694 41026
rect -5694 40974 -5692 41026
rect -5748 40972 -5692 40974
rect -5588 41026 -5532 41028
rect -5588 40974 -5586 41026
rect -5586 40974 -5534 41026
rect -5534 40974 -5532 41026
rect -5588 40972 -5532 40974
rect -5428 41026 -5372 41028
rect -5428 40974 -5426 41026
rect -5426 40974 -5374 41026
rect -5374 40974 -5372 41026
rect -5428 40972 -5372 40974
rect -5268 41026 -5212 41028
rect -5268 40974 -5266 41026
rect -5266 40974 -5214 41026
rect -5214 40974 -5212 41026
rect -5268 40972 -5212 40974
rect -5108 41026 -5052 41028
rect -5108 40974 -5106 41026
rect -5106 40974 -5054 41026
rect -5054 40974 -5052 41026
rect -5108 40972 -5052 40974
rect -4948 41026 -4892 41028
rect -4948 40974 -4946 41026
rect -4946 40974 -4894 41026
rect -4894 40974 -4892 41026
rect -4948 40972 -4892 40974
rect -4788 41026 -4732 41028
rect -4788 40974 -4786 41026
rect -4786 40974 -4734 41026
rect -4734 40974 -4732 41026
rect -4788 40972 -4732 40974
rect -4628 41026 -4572 41028
rect -4628 40974 -4626 41026
rect -4626 40974 -4574 41026
rect -4574 40974 -4572 41026
rect -4628 40972 -4572 40974
rect -4468 41026 -4412 41028
rect -4468 40974 -4466 41026
rect -4466 40974 -4414 41026
rect -4414 40974 -4412 41026
rect -4468 40972 -4412 40974
rect -4308 41026 -4252 41028
rect -4308 40974 -4306 41026
rect -4306 40974 -4254 41026
rect -4254 40974 -4252 41026
rect -4308 40972 -4252 40974
rect -4148 41026 -4092 41028
rect -4148 40974 -4146 41026
rect -4146 40974 -4094 41026
rect -4094 40974 -4092 41026
rect -4148 40972 -4092 40974
rect -3988 41026 -3932 41028
rect -3988 40974 -3986 41026
rect -3986 40974 -3934 41026
rect -3934 40974 -3932 41026
rect -3988 40972 -3932 40974
rect -3828 40972 -3772 41028
rect -3668 41026 -3612 41028
rect -3668 40974 -3666 41026
rect -3666 40974 -3614 41026
rect -3614 40974 -3612 41026
rect -3668 40972 -3612 40974
rect -3508 41026 -3452 41028
rect -3508 40974 -3506 41026
rect -3506 40974 -3454 41026
rect -3454 40974 -3452 41026
rect -3508 40972 -3452 40974
rect 41052 41026 41108 41028
rect 41052 40974 41054 41026
rect 41054 40974 41106 41026
rect 41106 40974 41108 41026
rect 41052 40972 41108 40974
rect 41212 41026 41268 41028
rect 41212 40974 41214 41026
rect 41214 40974 41266 41026
rect 41266 40974 41268 41026
rect 41212 40972 41268 40974
rect 41372 41026 41428 41028
rect 41372 40974 41374 41026
rect 41374 40974 41426 41026
rect 41426 40974 41428 41026
rect 41372 40972 41428 40974
rect 41532 41026 41588 41028
rect 41532 40974 41534 41026
rect 41534 40974 41586 41026
rect 41586 40974 41588 41026
rect 41532 40972 41588 40974
rect 41692 41026 41748 41028
rect 41692 40974 41694 41026
rect 41694 40974 41746 41026
rect 41746 40974 41748 41026
rect 41692 40972 41748 40974
rect 41852 41026 41908 41028
rect 41852 40974 41854 41026
rect 41854 40974 41906 41026
rect 41906 40974 41908 41026
rect 41852 40972 41908 40974
rect 42012 41026 42068 41028
rect 42012 40974 42014 41026
rect 42014 40974 42066 41026
rect 42066 40974 42068 41026
rect 42012 40972 42068 40974
rect 42172 41026 42228 41028
rect 42172 40974 42174 41026
rect 42174 40974 42226 41026
rect 42226 40974 42228 41026
rect 42172 40972 42228 40974
rect 42332 41026 42388 41028
rect 42332 40974 42334 41026
rect 42334 40974 42386 41026
rect 42386 40974 42388 41026
rect 42332 40972 42388 40974
rect 42492 41026 42548 41028
rect 42492 40974 42494 41026
rect 42494 40974 42546 41026
rect 42546 40974 42548 41026
rect 42492 40972 42548 40974
rect 42652 41026 42708 41028
rect 42652 40974 42654 41026
rect 42654 40974 42706 41026
rect 42706 40974 42708 41026
rect 42652 40972 42708 40974
rect 42812 41026 42868 41028
rect 42812 40974 42814 41026
rect 42814 40974 42866 41026
rect 42866 40974 42868 41026
rect 42812 40972 42868 40974
rect 42972 41026 43028 41028
rect 42972 40974 42974 41026
rect 42974 40974 43026 41026
rect 43026 40974 43028 41026
rect 42972 40972 43028 40974
rect 43132 41026 43188 41028
rect 43132 40974 43134 41026
rect 43134 40974 43186 41026
rect 43186 40974 43188 41026
rect 43132 40972 43188 40974
rect -12148 40812 -12092 40868
rect -11828 40812 -11772 40868
rect -11508 40812 -11452 40868
rect -3348 40812 -3292 40868
rect -3028 40812 -2972 40868
rect -2708 40812 -2652 40868
rect -2388 40812 -2332 40868
rect -2068 40812 -2012 40868
rect -1748 40812 -1692 40868
rect -1428 40812 -1372 40868
rect -1108 40812 -1052 40868
rect -31028 40732 -30972 40788
rect -30708 40732 -30652 40788
rect -30388 40732 -30332 40788
rect -30068 40732 -30012 40788
rect -12148 40652 -12092 40708
rect -11828 40652 -11772 40708
rect -11508 40652 -11452 40708
rect -10548 40706 -10492 40708
rect -10548 40654 -10546 40706
rect -10546 40654 -10494 40706
rect -10494 40654 -10492 40706
rect -10548 40652 -10492 40654
rect -10228 40706 -10172 40708
rect -10228 40654 -10226 40706
rect -10226 40654 -10174 40706
rect -10174 40654 -10172 40706
rect -10228 40652 -10172 40654
rect -10068 40706 -10012 40708
rect -10068 40654 -10066 40706
rect -10066 40654 -10014 40706
rect -10014 40654 -10012 40706
rect -10068 40652 -10012 40654
rect -9908 40706 -9852 40708
rect -9908 40654 -9906 40706
rect -9906 40654 -9854 40706
rect -9854 40654 -9852 40706
rect -9908 40652 -9852 40654
rect -9748 40706 -9692 40708
rect -9748 40654 -9746 40706
rect -9746 40654 -9694 40706
rect -9694 40654 -9692 40706
rect -9748 40652 -9692 40654
rect -9588 40706 -9532 40708
rect -9588 40654 -9586 40706
rect -9586 40654 -9534 40706
rect -9534 40654 -9532 40706
rect -9588 40652 -9532 40654
rect -9428 40706 -9372 40708
rect -9428 40654 -9426 40706
rect -9426 40654 -9374 40706
rect -9374 40654 -9372 40706
rect -9428 40652 -9372 40654
rect -9268 40706 -9212 40708
rect -9268 40654 -9266 40706
rect -9266 40654 -9214 40706
rect -9214 40654 -9212 40706
rect -9268 40652 -9212 40654
rect -9108 40706 -9052 40708
rect -9108 40654 -9106 40706
rect -9106 40654 -9054 40706
rect -9054 40654 -9052 40706
rect -9108 40652 -9052 40654
rect -8948 40706 -8892 40708
rect -8948 40654 -8946 40706
rect -8946 40654 -8894 40706
rect -8894 40654 -8892 40706
rect -8948 40652 -8892 40654
rect -8788 40706 -8732 40708
rect -8788 40654 -8786 40706
rect -8786 40654 -8734 40706
rect -8734 40654 -8732 40706
rect -8788 40652 -8732 40654
rect -8628 40706 -8572 40708
rect -8628 40654 -8626 40706
rect -8626 40654 -8574 40706
rect -8574 40654 -8572 40706
rect -8628 40652 -8572 40654
rect -8468 40706 -8412 40708
rect -8468 40654 -8466 40706
rect -8466 40654 -8414 40706
rect -8414 40654 -8412 40706
rect -8468 40652 -8412 40654
rect -8308 40706 -8252 40708
rect -8308 40654 -8306 40706
rect -8306 40654 -8254 40706
rect -8254 40654 -8252 40706
rect -8308 40652 -8252 40654
rect -8148 40706 -8092 40708
rect -8148 40654 -8146 40706
rect -8146 40654 -8094 40706
rect -8094 40654 -8092 40706
rect -8148 40652 -8092 40654
rect -7988 40706 -7932 40708
rect -7988 40654 -7986 40706
rect -7986 40654 -7934 40706
rect -7934 40654 -7932 40706
rect -7988 40652 -7932 40654
rect -7828 40706 -7772 40708
rect -7828 40654 -7826 40706
rect -7826 40654 -7774 40706
rect -7774 40654 -7772 40706
rect -7828 40652 -7772 40654
rect -7668 40706 -7612 40708
rect -7668 40654 -7666 40706
rect -7666 40654 -7614 40706
rect -7614 40654 -7612 40706
rect -7668 40652 -7612 40654
rect -7508 40706 -7452 40708
rect -7508 40654 -7506 40706
rect -7506 40654 -7454 40706
rect -7454 40654 -7452 40706
rect -7508 40652 -7452 40654
rect -7348 40706 -7292 40708
rect -7348 40654 -7346 40706
rect -7346 40654 -7294 40706
rect -7294 40654 -7292 40706
rect -7348 40652 -7292 40654
rect -7188 40706 -7132 40708
rect -7188 40654 -7186 40706
rect -7186 40654 -7134 40706
rect -7134 40654 -7132 40706
rect -7188 40652 -7132 40654
rect -7028 40706 -6972 40708
rect -7028 40654 -7026 40706
rect -7026 40654 -6974 40706
rect -6974 40654 -6972 40706
rect -7028 40652 -6972 40654
rect -6868 40706 -6812 40708
rect -6868 40654 -6866 40706
rect -6866 40654 -6814 40706
rect -6814 40654 -6812 40706
rect -6868 40652 -6812 40654
rect -6708 40706 -6652 40708
rect -6708 40654 -6706 40706
rect -6706 40654 -6654 40706
rect -6654 40654 -6652 40706
rect -6708 40652 -6652 40654
rect -6548 40706 -6492 40708
rect -6548 40654 -6546 40706
rect -6546 40654 -6494 40706
rect -6494 40654 -6492 40706
rect -6548 40652 -6492 40654
rect -6388 40706 -6332 40708
rect -6388 40654 -6386 40706
rect -6386 40654 -6334 40706
rect -6334 40654 -6332 40706
rect -6388 40652 -6332 40654
rect -6228 40706 -6172 40708
rect -6228 40654 -6226 40706
rect -6226 40654 -6174 40706
rect -6174 40654 -6172 40706
rect -6228 40652 -6172 40654
rect -6068 40706 -6012 40708
rect -6068 40654 -6066 40706
rect -6066 40654 -6014 40706
rect -6014 40654 -6012 40706
rect -6068 40652 -6012 40654
rect -5908 40706 -5852 40708
rect -5908 40654 -5906 40706
rect -5906 40654 -5854 40706
rect -5854 40654 -5852 40706
rect -5908 40652 -5852 40654
rect -5748 40706 -5692 40708
rect -5748 40654 -5746 40706
rect -5746 40654 -5694 40706
rect -5694 40654 -5692 40706
rect -5748 40652 -5692 40654
rect -5588 40706 -5532 40708
rect -5588 40654 -5586 40706
rect -5586 40654 -5534 40706
rect -5534 40654 -5532 40706
rect -5588 40652 -5532 40654
rect -5428 40706 -5372 40708
rect -5428 40654 -5426 40706
rect -5426 40654 -5374 40706
rect -5374 40654 -5372 40706
rect -5428 40652 -5372 40654
rect -5268 40706 -5212 40708
rect -5268 40654 -5266 40706
rect -5266 40654 -5214 40706
rect -5214 40654 -5212 40706
rect -5268 40652 -5212 40654
rect -5108 40706 -5052 40708
rect -5108 40654 -5106 40706
rect -5106 40654 -5054 40706
rect -5054 40654 -5052 40706
rect -5108 40652 -5052 40654
rect -4948 40706 -4892 40708
rect -4948 40654 -4946 40706
rect -4946 40654 -4894 40706
rect -4894 40654 -4892 40706
rect -4948 40652 -4892 40654
rect -4788 40706 -4732 40708
rect -4788 40654 -4786 40706
rect -4786 40654 -4734 40706
rect -4734 40654 -4732 40706
rect -4788 40652 -4732 40654
rect -4628 40706 -4572 40708
rect -4628 40654 -4626 40706
rect -4626 40654 -4574 40706
rect -4574 40654 -4572 40706
rect -4628 40652 -4572 40654
rect -4468 40706 -4412 40708
rect -4468 40654 -4466 40706
rect -4466 40654 -4414 40706
rect -4414 40654 -4412 40706
rect -4468 40652 -4412 40654
rect -4308 40706 -4252 40708
rect -4308 40654 -4306 40706
rect -4306 40654 -4254 40706
rect -4254 40654 -4252 40706
rect -4308 40652 -4252 40654
rect -4148 40706 -4092 40708
rect -4148 40654 -4146 40706
rect -4146 40654 -4094 40706
rect -4094 40654 -4092 40706
rect -4148 40652 -4092 40654
rect -3988 40706 -3932 40708
rect -3988 40654 -3986 40706
rect -3986 40654 -3934 40706
rect -3934 40654 -3932 40706
rect -3988 40652 -3932 40654
rect -3668 40706 -3612 40708
rect -3668 40654 -3666 40706
rect -3666 40654 -3614 40706
rect -3614 40654 -3612 40706
rect -3668 40652 -3612 40654
rect -3508 40706 -3452 40708
rect -3508 40654 -3506 40706
rect -3506 40654 -3454 40706
rect -3454 40654 -3452 40706
rect -3508 40652 -3452 40654
rect -3348 40652 -3292 40708
rect -3028 40652 -2972 40708
rect -2708 40652 -2652 40708
rect -2388 40652 -2332 40708
rect -2068 40652 -2012 40708
rect -1748 40652 -1692 40708
rect -1428 40652 -1372 40708
rect -1108 40652 -1052 40708
rect -31028 40572 -30972 40628
rect -30708 40572 -30652 40628
rect -30388 40572 -30332 40628
rect -30068 40572 -30012 40628
rect -10388 40492 -10332 40548
rect -1268 40492 -1212 40548
rect -31028 40412 -30972 40468
rect -30708 40412 -30652 40468
rect -30388 40412 -30332 40468
rect -30068 40412 -30012 40468
rect -12148 40332 -12092 40388
rect -11828 40332 -11772 40388
rect -11508 40332 -11452 40388
rect -10548 40386 -10492 40388
rect -10548 40334 -10546 40386
rect -10546 40334 -10494 40386
rect -10494 40334 -10492 40386
rect -10548 40332 -10492 40334
rect -10228 40386 -10172 40388
rect -10228 40334 -10226 40386
rect -10226 40334 -10174 40386
rect -10174 40334 -10172 40386
rect -10228 40332 -10172 40334
rect -10068 40386 -10012 40388
rect -10068 40334 -10066 40386
rect -10066 40334 -10014 40386
rect -10014 40334 -10012 40386
rect -10068 40332 -10012 40334
rect -9908 40386 -9852 40388
rect -9908 40334 -9906 40386
rect -9906 40334 -9854 40386
rect -9854 40334 -9852 40386
rect -9908 40332 -9852 40334
rect -9748 40386 -9692 40388
rect -9748 40334 -9746 40386
rect -9746 40334 -9694 40386
rect -9694 40334 -9692 40386
rect -9748 40332 -9692 40334
rect -9588 40386 -9532 40388
rect -9588 40334 -9586 40386
rect -9586 40334 -9534 40386
rect -9534 40334 -9532 40386
rect -9588 40332 -9532 40334
rect -9428 40386 -9372 40388
rect -9428 40334 -9426 40386
rect -9426 40334 -9374 40386
rect -9374 40334 -9372 40386
rect -9428 40332 -9372 40334
rect -9268 40386 -9212 40388
rect -9268 40334 -9266 40386
rect -9266 40334 -9214 40386
rect -9214 40334 -9212 40386
rect -9268 40332 -9212 40334
rect -9108 40386 -9052 40388
rect -9108 40334 -9106 40386
rect -9106 40334 -9054 40386
rect -9054 40334 -9052 40386
rect -9108 40332 -9052 40334
rect -8948 40386 -8892 40388
rect -8948 40334 -8946 40386
rect -8946 40334 -8894 40386
rect -8894 40334 -8892 40386
rect -8948 40332 -8892 40334
rect -8788 40386 -8732 40388
rect -8788 40334 -8786 40386
rect -8786 40334 -8734 40386
rect -8734 40334 -8732 40386
rect -8788 40332 -8732 40334
rect -8628 40386 -8572 40388
rect -8628 40334 -8626 40386
rect -8626 40334 -8574 40386
rect -8574 40334 -8572 40386
rect -8628 40332 -8572 40334
rect -8468 40386 -8412 40388
rect -8468 40334 -8466 40386
rect -8466 40334 -8414 40386
rect -8414 40334 -8412 40386
rect -8468 40332 -8412 40334
rect -8308 40386 -8252 40388
rect -8308 40334 -8306 40386
rect -8306 40334 -8254 40386
rect -8254 40334 -8252 40386
rect -8308 40332 -8252 40334
rect -8148 40386 -8092 40388
rect -8148 40334 -8146 40386
rect -8146 40334 -8094 40386
rect -8094 40334 -8092 40386
rect -8148 40332 -8092 40334
rect -7988 40386 -7932 40388
rect -7988 40334 -7986 40386
rect -7986 40334 -7934 40386
rect -7934 40334 -7932 40386
rect -7988 40332 -7932 40334
rect -7828 40386 -7772 40388
rect -7828 40334 -7826 40386
rect -7826 40334 -7774 40386
rect -7774 40334 -7772 40386
rect -7828 40332 -7772 40334
rect -7668 40386 -7612 40388
rect -7668 40334 -7666 40386
rect -7666 40334 -7614 40386
rect -7614 40334 -7612 40386
rect -7668 40332 -7612 40334
rect -7508 40386 -7452 40388
rect -7508 40334 -7506 40386
rect -7506 40334 -7454 40386
rect -7454 40334 -7452 40386
rect -7508 40332 -7452 40334
rect -7348 40386 -7292 40388
rect -7348 40334 -7346 40386
rect -7346 40334 -7294 40386
rect -7294 40334 -7292 40386
rect -7348 40332 -7292 40334
rect -7188 40386 -7132 40388
rect -7188 40334 -7186 40386
rect -7186 40334 -7134 40386
rect -7134 40334 -7132 40386
rect -7188 40332 -7132 40334
rect -7028 40386 -6972 40388
rect -7028 40334 -7026 40386
rect -7026 40334 -6974 40386
rect -6974 40334 -6972 40386
rect -7028 40332 -6972 40334
rect -6868 40386 -6812 40388
rect -6868 40334 -6866 40386
rect -6866 40334 -6814 40386
rect -6814 40334 -6812 40386
rect -6868 40332 -6812 40334
rect -6708 40386 -6652 40388
rect -6708 40334 -6706 40386
rect -6706 40334 -6654 40386
rect -6654 40334 -6652 40386
rect -6708 40332 -6652 40334
rect -6548 40386 -6492 40388
rect -6548 40334 -6546 40386
rect -6546 40334 -6494 40386
rect -6494 40334 -6492 40386
rect -6548 40332 -6492 40334
rect -6388 40386 -6332 40388
rect -6388 40334 -6386 40386
rect -6386 40334 -6334 40386
rect -6334 40334 -6332 40386
rect -6388 40332 -6332 40334
rect -6228 40386 -6172 40388
rect -6228 40334 -6226 40386
rect -6226 40334 -6174 40386
rect -6174 40334 -6172 40386
rect -6228 40332 -6172 40334
rect -6068 40386 -6012 40388
rect -6068 40334 -6066 40386
rect -6066 40334 -6014 40386
rect -6014 40334 -6012 40386
rect -6068 40332 -6012 40334
rect -5908 40386 -5852 40388
rect -5908 40334 -5906 40386
rect -5906 40334 -5854 40386
rect -5854 40334 -5852 40386
rect -5908 40332 -5852 40334
rect -5748 40386 -5692 40388
rect -5748 40334 -5746 40386
rect -5746 40334 -5694 40386
rect -5694 40334 -5692 40386
rect -5748 40332 -5692 40334
rect -5588 40386 -5532 40388
rect -5588 40334 -5586 40386
rect -5586 40334 -5534 40386
rect -5534 40334 -5532 40386
rect -5588 40332 -5532 40334
rect -5428 40386 -5372 40388
rect -5428 40334 -5426 40386
rect -5426 40334 -5374 40386
rect -5374 40334 -5372 40386
rect -5428 40332 -5372 40334
rect -5268 40386 -5212 40388
rect -5268 40334 -5266 40386
rect -5266 40334 -5214 40386
rect -5214 40334 -5212 40386
rect -5268 40332 -5212 40334
rect -5108 40386 -5052 40388
rect -5108 40334 -5106 40386
rect -5106 40334 -5054 40386
rect -5054 40334 -5052 40386
rect -5108 40332 -5052 40334
rect -4948 40386 -4892 40388
rect -4948 40334 -4946 40386
rect -4946 40334 -4894 40386
rect -4894 40334 -4892 40386
rect -4948 40332 -4892 40334
rect -4788 40386 -4732 40388
rect -4788 40334 -4786 40386
rect -4786 40334 -4734 40386
rect -4734 40334 -4732 40386
rect -4788 40332 -4732 40334
rect -4628 40386 -4572 40388
rect -4628 40334 -4626 40386
rect -4626 40334 -4574 40386
rect -4574 40334 -4572 40386
rect -4628 40332 -4572 40334
rect -4468 40386 -4412 40388
rect -4468 40334 -4466 40386
rect -4466 40334 -4414 40386
rect -4414 40334 -4412 40386
rect -4468 40332 -4412 40334
rect -4308 40386 -4252 40388
rect -4308 40334 -4306 40386
rect -4306 40334 -4254 40386
rect -4254 40334 -4252 40386
rect -4308 40332 -4252 40334
rect -4148 40386 -4092 40388
rect -4148 40334 -4146 40386
rect -4146 40334 -4094 40386
rect -4094 40334 -4092 40386
rect -4148 40332 -4092 40334
rect -3988 40386 -3932 40388
rect -3988 40334 -3986 40386
rect -3986 40334 -3934 40386
rect -3934 40334 -3932 40386
rect -3988 40332 -3932 40334
rect -3668 40386 -3612 40388
rect -3668 40334 -3666 40386
rect -3666 40334 -3614 40386
rect -3614 40334 -3612 40386
rect -3668 40332 -3612 40334
rect -3508 40386 -3452 40388
rect -3508 40334 -3506 40386
rect -3506 40334 -3454 40386
rect -3454 40334 -3452 40386
rect -3508 40332 -3452 40334
rect -3348 40332 -3292 40388
rect -3028 40332 -2972 40388
rect -2708 40332 -2652 40388
rect -2388 40332 -2332 40388
rect -2068 40332 -2012 40388
rect -1748 40332 -1692 40388
rect -1428 40332 -1372 40388
rect -1108 40332 -1052 40388
rect -31028 40252 -30972 40308
rect -30708 40252 -30652 40308
rect -30388 40252 -30332 40308
rect -30068 40252 -30012 40308
rect -3348 40172 -3292 40228
rect -3028 40172 -2972 40228
rect -2708 40172 -2652 40228
rect -2548 40172 -2492 40228
rect -1908 40172 -1852 40228
rect -31028 40092 -30972 40148
rect -30708 40092 -30652 40148
rect -30388 40092 -30332 40148
rect -30068 40092 -30012 40148
rect -3348 40012 -3292 40068
rect -3028 40012 -2972 40068
rect -2708 40012 -2652 40068
rect -2388 40012 -2332 40068
rect -2068 40012 -2012 40068
rect -1748 40012 -1692 40068
rect -1428 40012 -1372 40068
rect -1108 40012 -1052 40068
rect 41052 40066 41108 40068
rect 41052 40014 41054 40066
rect 41054 40014 41106 40066
rect 41106 40014 41108 40066
rect 41052 40012 41108 40014
rect 41212 40066 41268 40068
rect 41212 40014 41214 40066
rect 41214 40014 41266 40066
rect 41266 40014 41268 40066
rect 41212 40012 41268 40014
rect 41372 40066 41428 40068
rect 41372 40014 41374 40066
rect 41374 40014 41426 40066
rect 41426 40014 41428 40066
rect 41372 40012 41428 40014
rect 41532 40066 41588 40068
rect 41532 40014 41534 40066
rect 41534 40014 41586 40066
rect 41586 40014 41588 40066
rect 41532 40012 41588 40014
rect 41692 40066 41748 40068
rect 41692 40014 41694 40066
rect 41694 40014 41746 40066
rect 41746 40014 41748 40066
rect 41692 40012 41748 40014
rect 41852 40066 41908 40068
rect 41852 40014 41854 40066
rect 41854 40014 41906 40066
rect 41906 40014 41908 40066
rect 41852 40012 41908 40014
rect 42012 40066 42068 40068
rect 42012 40014 42014 40066
rect 42014 40014 42066 40066
rect 42066 40014 42068 40066
rect 42012 40012 42068 40014
rect 42172 40066 42228 40068
rect 42172 40014 42174 40066
rect 42174 40014 42226 40066
rect 42226 40014 42228 40066
rect 42172 40012 42228 40014
rect 42332 40066 42388 40068
rect 42332 40014 42334 40066
rect 42334 40014 42386 40066
rect 42386 40014 42388 40066
rect 42332 40012 42388 40014
rect 42492 40066 42548 40068
rect 42492 40014 42494 40066
rect 42494 40014 42546 40066
rect 42546 40014 42548 40066
rect 42492 40012 42548 40014
rect 42652 40066 42708 40068
rect 42652 40014 42654 40066
rect 42654 40014 42706 40066
rect 42706 40014 42708 40066
rect 42652 40012 42708 40014
rect 42812 40066 42868 40068
rect 42812 40014 42814 40066
rect 42814 40014 42866 40066
rect 42866 40014 42868 40066
rect 42812 40012 42868 40014
rect 42972 40066 43028 40068
rect 42972 40014 42974 40066
rect 42974 40014 43026 40066
rect 43026 40014 43028 40066
rect 42972 40012 43028 40014
rect 43132 40066 43188 40068
rect 43132 40014 43134 40066
rect 43134 40014 43186 40066
rect 43186 40014 43188 40066
rect 43132 40012 43188 40014
rect -31028 39932 -30972 39988
rect -30708 39932 -30652 39988
rect -30388 39932 -30332 39988
rect -30068 39932 -30012 39988
rect -3348 39852 -3292 39908
rect -3028 39852 -2972 39908
rect -2708 39852 -2652 39908
rect -2388 39852 -2332 39908
rect -2228 39852 -2172 39908
rect -1588 39852 -1532 39908
rect -31028 39772 -30972 39828
rect -30708 39772 -30652 39828
rect -30388 39772 -30332 39828
rect -30068 39772 -30012 39828
rect -3348 39692 -3292 39748
rect -3028 39692 -2972 39748
rect -2708 39692 -2652 39748
rect -2388 39692 -2332 39748
rect -2068 39692 -2012 39748
rect -1748 39692 -1692 39748
rect -1428 39692 -1372 39748
rect -1108 39692 -1052 39748
rect 41052 39746 41108 39748
rect 41052 39694 41054 39746
rect 41054 39694 41106 39746
rect 41106 39694 41108 39746
rect 41052 39692 41108 39694
rect 41212 39746 41268 39748
rect 41212 39694 41214 39746
rect 41214 39694 41266 39746
rect 41266 39694 41268 39746
rect 41212 39692 41268 39694
rect 41372 39746 41428 39748
rect 41372 39694 41374 39746
rect 41374 39694 41426 39746
rect 41426 39694 41428 39746
rect 41372 39692 41428 39694
rect 41532 39746 41588 39748
rect 41532 39694 41534 39746
rect 41534 39694 41586 39746
rect 41586 39694 41588 39746
rect 41532 39692 41588 39694
rect 41692 39746 41748 39748
rect 41692 39694 41694 39746
rect 41694 39694 41746 39746
rect 41746 39694 41748 39746
rect 41692 39692 41748 39694
rect 41852 39746 41908 39748
rect 41852 39694 41854 39746
rect 41854 39694 41906 39746
rect 41906 39694 41908 39746
rect 41852 39692 41908 39694
rect 42012 39746 42068 39748
rect 42012 39694 42014 39746
rect 42014 39694 42066 39746
rect 42066 39694 42068 39746
rect 42012 39692 42068 39694
rect 42172 39746 42228 39748
rect 42172 39694 42174 39746
rect 42174 39694 42226 39746
rect 42226 39694 42228 39746
rect 42172 39692 42228 39694
rect 42332 39746 42388 39748
rect 42332 39694 42334 39746
rect 42334 39694 42386 39746
rect 42386 39694 42388 39746
rect 42332 39692 42388 39694
rect 42492 39746 42548 39748
rect 42492 39694 42494 39746
rect 42494 39694 42546 39746
rect 42546 39694 42548 39746
rect 42492 39692 42548 39694
rect 42652 39746 42708 39748
rect 42652 39694 42654 39746
rect 42654 39694 42706 39746
rect 42706 39694 42708 39746
rect 42652 39692 42708 39694
rect 42812 39746 42868 39748
rect 42812 39694 42814 39746
rect 42814 39694 42866 39746
rect 42866 39694 42868 39746
rect 42812 39692 42868 39694
rect 42972 39746 43028 39748
rect 42972 39694 42974 39746
rect 42974 39694 43026 39746
rect 43026 39694 43028 39746
rect 42972 39692 43028 39694
rect 43132 39746 43188 39748
rect 43132 39694 43134 39746
rect 43134 39694 43186 39746
rect 43186 39694 43188 39746
rect 43132 39692 43188 39694
rect -31028 39612 -30972 39668
rect -30708 39612 -30652 39668
rect -30388 39612 -30332 39668
rect -30068 39612 -30012 39668
rect -3348 39532 -3292 39588
rect -3028 39532 -2972 39588
rect -2708 39532 -2652 39588
rect -2388 39532 -2332 39588
rect -2068 39532 -2012 39588
rect -1748 39532 -1692 39588
rect -1428 39532 -1372 39588
rect -1108 39532 -1052 39588
rect -31028 39452 -30972 39508
rect -30708 39452 -30652 39508
rect -30388 39452 -30332 39508
rect -30068 39452 -30012 39508
rect -3348 39372 -3292 39428
rect -3028 39372 -2972 39428
rect -2708 39372 -2652 39428
rect -2388 39372 -2332 39428
rect -2068 39372 -2012 39428
rect -1748 39372 -1692 39428
rect -1428 39372 -1372 39428
rect -1108 39372 -1052 39428
rect -31028 39292 -30972 39348
rect -30708 39292 -30652 39348
rect -30388 39292 -30332 39348
rect -30068 39292 -30012 39348
rect -3348 39212 -3292 39268
rect -3028 39212 -2972 39268
rect -2708 39212 -2652 39268
rect -2388 39212 -2332 39268
rect -2068 39212 -2012 39268
rect -1748 39212 -1692 39268
rect -1428 39212 -1372 39268
rect -1108 39212 -1052 39268
rect -31028 39132 -30972 39188
rect -30708 39132 -30652 39188
rect -30388 39132 -30332 39188
rect -30068 39132 -30012 39188
rect -3348 39052 -3292 39108
rect -3028 39052 -2972 39108
rect -2708 39052 -2652 39108
rect -2388 39052 -2332 39108
rect -2068 39052 -2012 39108
rect -1748 39052 -1692 39108
rect -1428 39052 -1372 39108
rect -1108 39052 -1052 39108
rect -31028 38972 -30972 39028
rect -30708 38972 -30652 39028
rect -30388 38972 -30332 39028
rect -30068 38972 -30012 39028
rect -3348 38892 -3292 38948
rect -3028 38892 -2972 38948
rect -2708 38892 -2652 38948
rect -2388 38892 -2332 38948
rect -2068 38892 -2012 38948
rect -1748 38892 -1692 38948
rect -1428 38892 -1372 38948
rect -1108 38892 -1052 38948
rect -31028 38812 -30972 38868
rect -30708 38812 -30652 38868
rect -30388 38812 -30332 38868
rect -30068 38812 -30012 38868
rect -3348 38732 -3292 38788
rect -3028 38732 -2972 38788
rect -2708 38732 -2652 38788
rect -2388 38732 -2332 38788
rect -2068 38732 -2012 38788
rect -1748 38732 -1692 38788
rect -1428 38732 -1372 38788
rect -1108 38732 -1052 38788
rect -31028 38652 -30972 38708
rect -30708 38652 -30652 38708
rect -30388 38652 -30332 38708
rect -30068 38652 -30012 38708
rect -3348 38572 -3292 38628
rect -3028 38572 -2972 38628
rect -2708 38572 -2652 38628
rect -2388 38572 -2332 38628
rect -2068 38572 -2012 38628
rect -1748 38572 -1692 38628
rect -1428 38572 -1372 38628
rect -1108 38572 -1052 38628
rect -31028 38492 -30972 38548
rect -30708 38492 -30652 38548
rect -30388 38492 -30332 38548
rect -30068 38492 -30012 38548
rect -3348 38412 -3292 38468
rect -3028 38412 -2972 38468
rect -2708 38412 -2652 38468
rect -2388 38412 -2332 38468
rect -2068 38412 -2012 38468
rect -1748 38412 -1692 38468
rect -1428 38412 -1372 38468
rect -1108 38412 -1052 38468
rect -31028 38332 -30972 38388
rect -30708 38332 -30652 38388
rect -30388 38332 -30332 38388
rect -30068 38332 -30012 38388
rect -3348 38252 -3292 38308
rect -3028 38252 -2972 38308
rect -2708 38252 -2652 38308
rect -2388 38252 -2332 38308
rect -2068 38252 -2012 38308
rect -1748 38252 -1692 38308
rect -1428 38252 -1372 38308
rect -1108 38252 -1052 38308
rect -31028 38172 -30972 38228
rect -30708 38172 -30652 38228
rect -30388 38172 -30332 38228
rect -30068 38172 -30012 38228
rect -3348 38092 -3292 38148
rect -3028 38092 -2972 38148
rect -2708 38092 -2652 38148
rect -2388 38092 -2332 38148
rect -2068 38092 -2012 38148
rect -1748 38092 -1692 38148
rect -1428 38092 -1372 38148
rect -1108 38092 -1052 38148
rect -31028 38012 -30972 38068
rect -30708 38012 -30652 38068
rect -30388 38012 -30332 38068
rect -30068 38012 -30012 38068
rect -3348 37932 -3292 37988
rect -3028 37932 -2972 37988
rect -2708 37932 -2652 37988
rect -2388 37932 -2332 37988
rect -2068 37932 -2012 37988
rect -1748 37932 -1692 37988
rect -1428 37932 -1372 37988
rect -1108 37932 -1052 37988
rect -31028 37852 -30972 37908
rect -30708 37852 -30652 37908
rect -30388 37852 -30332 37908
rect -30068 37852 -30012 37908
rect -3348 37772 -3292 37828
rect -3028 37772 -2972 37828
rect -2708 37772 -2652 37828
rect -2388 37772 -2332 37828
rect -2068 37772 -2012 37828
rect -1748 37772 -1692 37828
rect -1428 37772 -1372 37828
rect -1108 37772 -1052 37828
rect -33108 37746 -33052 37748
rect -33108 37694 -33106 37746
rect -33106 37694 -33054 37746
rect -33054 37694 -33052 37746
rect -33108 37692 -33052 37694
rect -32948 37746 -32892 37748
rect -32948 37694 -32946 37746
rect -32946 37694 -32894 37746
rect -32894 37694 -32892 37746
rect -32948 37692 -32892 37694
rect -32788 37746 -32732 37748
rect -32788 37694 -32786 37746
rect -32786 37694 -32734 37746
rect -32734 37694 -32732 37746
rect -32788 37692 -32732 37694
rect -32628 37746 -32572 37748
rect -32628 37694 -32626 37746
rect -32626 37694 -32574 37746
rect -32574 37694 -32572 37746
rect -32628 37692 -32572 37694
rect -32468 37746 -32412 37748
rect -32468 37694 -32466 37746
rect -32466 37694 -32414 37746
rect -32414 37694 -32412 37746
rect -32468 37692 -32412 37694
rect -32308 37746 -32252 37748
rect -32308 37694 -32306 37746
rect -32306 37694 -32254 37746
rect -32254 37694 -32252 37746
rect -32308 37692 -32252 37694
rect -32148 37746 -32092 37748
rect -32148 37694 -32146 37746
rect -32146 37694 -32094 37746
rect -32094 37694 -32092 37746
rect -32148 37692 -32092 37694
rect -31988 37746 -31932 37748
rect -31988 37694 -31986 37746
rect -31986 37694 -31934 37746
rect -31934 37694 -31932 37746
rect -31988 37692 -31932 37694
rect -31828 37746 -31772 37748
rect -31828 37694 -31826 37746
rect -31826 37694 -31774 37746
rect -31774 37694 -31772 37746
rect -31828 37692 -31772 37694
rect -31668 37746 -31612 37748
rect -31668 37694 -31666 37746
rect -31666 37694 -31614 37746
rect -31614 37694 -31612 37746
rect -31668 37692 -31612 37694
rect -31508 37746 -31452 37748
rect -31508 37694 -31506 37746
rect -31506 37694 -31454 37746
rect -31454 37694 -31452 37746
rect -31508 37692 -31452 37694
rect -31348 37746 -31292 37748
rect -31348 37694 -31346 37746
rect -31346 37694 -31294 37746
rect -31294 37694 -31292 37746
rect -31348 37692 -31292 37694
rect -31188 37746 -31132 37748
rect -31188 37694 -31186 37746
rect -31186 37694 -31134 37746
rect -31134 37694 -31132 37746
rect -31188 37692 -31132 37694
rect -31028 37692 -30972 37748
rect -30708 37692 -30652 37748
rect -30388 37692 -30332 37748
rect -30068 37692 -30012 37748
rect -3348 37612 -3292 37668
rect -3028 37612 -2972 37668
rect -2708 37612 -2652 37668
rect -2388 37612 -2332 37668
rect -2068 37612 -2012 37668
rect -1748 37612 -1692 37668
rect -1428 37612 -1372 37668
rect -1268 37612 -1212 37668
rect -30868 37532 -30812 37588
rect -30548 37532 -30492 37588
rect -3348 37452 -3292 37508
rect -3028 37452 -2972 37508
rect -2708 37452 -2652 37508
rect -2388 37452 -2332 37508
rect -2068 37452 -2012 37508
rect -1748 37452 -1692 37508
rect -1428 37452 -1372 37508
rect -1108 37452 -1052 37508
rect -33108 37426 -33052 37428
rect -33108 37374 -33106 37426
rect -33106 37374 -33054 37426
rect -33054 37374 -33052 37426
rect -33108 37372 -33052 37374
rect -32948 37426 -32892 37428
rect -32948 37374 -32946 37426
rect -32946 37374 -32894 37426
rect -32894 37374 -32892 37426
rect -32948 37372 -32892 37374
rect -32788 37426 -32732 37428
rect -32788 37374 -32786 37426
rect -32786 37374 -32734 37426
rect -32734 37374 -32732 37426
rect -32788 37372 -32732 37374
rect -32628 37426 -32572 37428
rect -32628 37374 -32626 37426
rect -32626 37374 -32574 37426
rect -32574 37374 -32572 37426
rect -32628 37372 -32572 37374
rect -32468 37426 -32412 37428
rect -32468 37374 -32466 37426
rect -32466 37374 -32414 37426
rect -32414 37374 -32412 37426
rect -32468 37372 -32412 37374
rect -32308 37426 -32252 37428
rect -32308 37374 -32306 37426
rect -32306 37374 -32254 37426
rect -32254 37374 -32252 37426
rect -32308 37372 -32252 37374
rect -32148 37426 -32092 37428
rect -32148 37374 -32146 37426
rect -32146 37374 -32094 37426
rect -32094 37374 -32092 37426
rect -32148 37372 -32092 37374
rect -31988 37426 -31932 37428
rect -31988 37374 -31986 37426
rect -31986 37374 -31934 37426
rect -31934 37374 -31932 37426
rect -31988 37372 -31932 37374
rect -31828 37426 -31772 37428
rect -31828 37374 -31826 37426
rect -31826 37374 -31774 37426
rect -31774 37374 -31772 37426
rect -31828 37372 -31772 37374
rect -31668 37426 -31612 37428
rect -31668 37374 -31666 37426
rect -31666 37374 -31614 37426
rect -31614 37374 -31612 37426
rect -31668 37372 -31612 37374
rect -31508 37426 -31452 37428
rect -31508 37374 -31506 37426
rect -31506 37374 -31454 37426
rect -31454 37374 -31452 37426
rect -31508 37372 -31452 37374
rect -31348 37426 -31292 37428
rect -31348 37374 -31346 37426
rect -31346 37374 -31294 37426
rect -31294 37374 -31292 37426
rect -31348 37372 -31292 37374
rect -31188 37426 -31132 37428
rect -31188 37374 -31186 37426
rect -31186 37374 -31134 37426
rect -31134 37374 -31132 37426
rect -31188 37372 -31132 37374
rect -31028 37372 -30972 37428
rect -30708 37372 -30652 37428
rect -30388 37372 -30332 37428
rect -30068 37372 -30012 37428
rect -3348 37292 -3292 37348
rect -3028 37292 -2972 37348
rect -2708 37292 -2652 37348
rect -2388 37292 -2332 37348
rect -2068 37292 -2012 37348
rect -1748 37292 -1692 37348
rect -1428 37292 -1372 37348
rect -1108 37292 -1052 37348
rect -30868 37212 -30812 37268
rect -30228 37212 -30172 37268
rect -3348 37132 -3292 37188
rect -3028 37132 -2972 37188
rect -2708 37132 -2652 37188
rect -2388 37132 -2332 37188
rect -2068 37132 -2012 37188
rect -1748 37132 -1692 37188
rect -1428 37132 -1372 37188
rect -1108 37132 -1052 37188
rect -33108 37106 -33052 37108
rect -33108 37054 -33106 37106
rect -33106 37054 -33054 37106
rect -33054 37054 -33052 37106
rect -33108 37052 -33052 37054
rect -32948 37106 -32892 37108
rect -32948 37054 -32946 37106
rect -32946 37054 -32894 37106
rect -32894 37054 -32892 37106
rect -32948 37052 -32892 37054
rect -32788 37106 -32732 37108
rect -32788 37054 -32786 37106
rect -32786 37054 -32734 37106
rect -32734 37054 -32732 37106
rect -32788 37052 -32732 37054
rect -32628 37106 -32572 37108
rect -32628 37054 -32626 37106
rect -32626 37054 -32574 37106
rect -32574 37054 -32572 37106
rect -32628 37052 -32572 37054
rect -32468 37106 -32412 37108
rect -32468 37054 -32466 37106
rect -32466 37054 -32414 37106
rect -32414 37054 -32412 37106
rect -32468 37052 -32412 37054
rect -32308 37106 -32252 37108
rect -32308 37054 -32306 37106
rect -32306 37054 -32254 37106
rect -32254 37054 -32252 37106
rect -32308 37052 -32252 37054
rect -32148 37106 -32092 37108
rect -32148 37054 -32146 37106
rect -32146 37054 -32094 37106
rect -32094 37054 -32092 37106
rect -32148 37052 -32092 37054
rect -31988 37106 -31932 37108
rect -31988 37054 -31986 37106
rect -31986 37054 -31934 37106
rect -31934 37054 -31932 37106
rect -31988 37052 -31932 37054
rect -31828 37106 -31772 37108
rect -31828 37054 -31826 37106
rect -31826 37054 -31774 37106
rect -31774 37054 -31772 37106
rect -31828 37052 -31772 37054
rect -31668 37106 -31612 37108
rect -31668 37054 -31666 37106
rect -31666 37054 -31614 37106
rect -31614 37054 -31612 37106
rect -31668 37052 -31612 37054
rect -31508 37106 -31452 37108
rect -31508 37054 -31506 37106
rect -31506 37054 -31454 37106
rect -31454 37054 -31452 37106
rect -31508 37052 -31452 37054
rect -31348 37106 -31292 37108
rect -31348 37054 -31346 37106
rect -31346 37054 -31294 37106
rect -31294 37054 -31292 37106
rect -31348 37052 -31292 37054
rect -31188 37106 -31132 37108
rect -31188 37054 -31186 37106
rect -31186 37054 -31134 37106
rect -31134 37054 -31132 37106
rect -31188 37052 -31132 37054
rect -31028 37052 -30972 37108
rect -30708 37052 -30652 37108
rect -30388 37052 -30332 37108
rect -30068 37052 -30012 37108
rect -3348 36972 -3292 37028
rect -3028 36972 -2972 37028
rect -2708 36972 -2652 37028
rect -2388 36972 -2332 37028
rect -2068 36972 -2012 37028
rect -1748 36972 -1692 37028
rect -1428 36972 -1372 37028
rect -1108 36972 -1052 37028
rect -31028 36892 -30972 36948
rect -30708 36892 -30652 36948
rect -30388 36892 -30332 36948
rect -30068 36892 -30012 36948
rect -3348 36812 -3292 36868
rect -3028 36812 -2972 36868
rect -2708 36812 -2652 36868
rect -2388 36812 -2332 36868
rect -2068 36812 -2012 36868
rect -1748 36812 -1692 36868
rect -1428 36812 -1372 36868
rect -1108 36812 -1052 36868
rect -31028 36732 -30972 36788
rect -30708 36732 -30652 36788
rect -30388 36732 -30332 36788
rect -30068 36732 -30012 36788
rect -3348 36652 -3292 36708
rect -3028 36652 -2972 36708
rect -2708 36652 -2652 36708
rect -2388 36652 -2332 36708
rect -2068 36652 -2012 36708
rect -1748 36652 -1692 36708
rect -1428 36652 -1372 36708
rect -1108 36652 -1052 36708
rect -31028 36572 -30972 36628
rect -30708 36572 -30652 36628
rect -30388 36572 -30332 36628
rect -30068 36572 -30012 36628
rect -3348 36492 -3292 36548
rect -3028 36492 -2972 36548
rect -2708 36492 -2652 36548
rect -2388 36492 -2332 36548
rect -2068 36492 -2012 36548
rect -1748 36492 -1692 36548
rect -1428 36492 -1372 36548
rect -1108 36492 -1052 36548
rect -31028 36412 -30972 36468
rect -30708 36412 -30652 36468
rect -30388 36412 -30332 36468
rect -30068 36412 -30012 36468
rect -3348 36332 -3292 36388
rect -3028 36332 -2972 36388
rect -2708 36332 -2652 36388
rect -2388 36332 -2332 36388
rect -2068 36332 -2012 36388
rect -1748 36332 -1692 36388
rect -1428 36332 -1372 36388
rect -1108 36332 -1052 36388
rect -31028 36252 -30972 36308
rect -30708 36252 -30652 36308
rect -30388 36252 -30332 36308
rect -30068 36252 -30012 36308
rect -3348 36172 -3292 36228
rect -3028 36172 -2972 36228
rect -2868 36172 -2812 36228
rect -1908 36172 -1852 36228
rect -31028 36092 -30972 36148
rect -30708 36092 -30652 36148
rect -30388 36092 -30332 36148
rect -30068 36092 -30012 36148
rect -3348 36012 -3292 36068
rect -3028 36012 -2972 36068
rect -2708 36012 -2652 36068
rect -2388 36012 -2332 36068
rect -2068 36012 -2012 36068
rect -1748 36012 -1692 36068
rect -1428 36012 -1372 36068
rect -1108 36012 -1052 36068
rect 41052 36066 41108 36068
rect 41052 36014 41054 36066
rect 41054 36014 41106 36066
rect 41106 36014 41108 36066
rect 41052 36012 41108 36014
rect 41212 36066 41268 36068
rect 41212 36014 41214 36066
rect 41214 36014 41266 36066
rect 41266 36014 41268 36066
rect 41212 36012 41268 36014
rect 41372 36066 41428 36068
rect 41372 36014 41374 36066
rect 41374 36014 41426 36066
rect 41426 36014 41428 36066
rect 41372 36012 41428 36014
rect 41532 36066 41588 36068
rect 41532 36014 41534 36066
rect 41534 36014 41586 36066
rect 41586 36014 41588 36066
rect 41532 36012 41588 36014
rect 41692 36066 41748 36068
rect 41692 36014 41694 36066
rect 41694 36014 41746 36066
rect 41746 36014 41748 36066
rect 41692 36012 41748 36014
rect 41852 36066 41908 36068
rect 41852 36014 41854 36066
rect 41854 36014 41906 36066
rect 41906 36014 41908 36066
rect 41852 36012 41908 36014
rect 42012 36066 42068 36068
rect 42012 36014 42014 36066
rect 42014 36014 42066 36066
rect 42066 36014 42068 36066
rect 42012 36012 42068 36014
rect 42172 36066 42228 36068
rect 42172 36014 42174 36066
rect 42174 36014 42226 36066
rect 42226 36014 42228 36066
rect 42172 36012 42228 36014
rect 42332 36066 42388 36068
rect 42332 36014 42334 36066
rect 42334 36014 42386 36066
rect 42386 36014 42388 36066
rect 42332 36012 42388 36014
rect 42492 36066 42548 36068
rect 42492 36014 42494 36066
rect 42494 36014 42546 36066
rect 42546 36014 42548 36066
rect 42492 36012 42548 36014
rect 42652 36066 42708 36068
rect 42652 36014 42654 36066
rect 42654 36014 42706 36066
rect 42706 36014 42708 36066
rect 42652 36012 42708 36014
rect 42812 36066 42868 36068
rect 42812 36014 42814 36066
rect 42814 36014 42866 36066
rect 42866 36014 42868 36066
rect 42812 36012 42868 36014
rect 42972 36066 43028 36068
rect 42972 36014 42974 36066
rect 42974 36014 43026 36066
rect 43026 36014 43028 36066
rect 42972 36012 43028 36014
rect 43132 36066 43188 36068
rect 43132 36014 43134 36066
rect 43134 36014 43186 36066
rect 43186 36014 43188 36066
rect 43132 36012 43188 36014
rect -31028 35932 -30972 35988
rect -30708 35932 -30652 35988
rect -30388 35932 -30332 35988
rect -30068 35932 -30012 35988
rect -3188 35852 -3132 35908
rect -1588 35852 -1532 35908
rect -31028 35772 -30972 35828
rect -30708 35772 -30652 35828
rect -30388 35772 -30332 35828
rect -30068 35772 -30012 35828
rect -3348 35692 -3292 35748
rect -3028 35692 -2972 35748
rect -2708 35692 -2652 35748
rect -2388 35692 -2332 35748
rect -2068 35692 -2012 35748
rect -1748 35692 -1692 35748
rect -1428 35692 -1372 35748
rect -1108 35692 -1052 35748
rect 41052 35746 41108 35748
rect 41052 35694 41054 35746
rect 41054 35694 41106 35746
rect 41106 35694 41108 35746
rect 41052 35692 41108 35694
rect 41212 35746 41268 35748
rect 41212 35694 41214 35746
rect 41214 35694 41266 35746
rect 41266 35694 41268 35746
rect 41212 35692 41268 35694
rect 41372 35746 41428 35748
rect 41372 35694 41374 35746
rect 41374 35694 41426 35746
rect 41426 35694 41428 35746
rect 41372 35692 41428 35694
rect 41532 35746 41588 35748
rect 41532 35694 41534 35746
rect 41534 35694 41586 35746
rect 41586 35694 41588 35746
rect 41532 35692 41588 35694
rect 41692 35746 41748 35748
rect 41692 35694 41694 35746
rect 41694 35694 41746 35746
rect 41746 35694 41748 35746
rect 41692 35692 41748 35694
rect 41852 35746 41908 35748
rect 41852 35694 41854 35746
rect 41854 35694 41906 35746
rect 41906 35694 41908 35746
rect 41852 35692 41908 35694
rect 42012 35746 42068 35748
rect 42012 35694 42014 35746
rect 42014 35694 42066 35746
rect 42066 35694 42068 35746
rect 42012 35692 42068 35694
rect 42172 35746 42228 35748
rect 42172 35694 42174 35746
rect 42174 35694 42226 35746
rect 42226 35694 42228 35746
rect 42172 35692 42228 35694
rect 42332 35746 42388 35748
rect 42332 35694 42334 35746
rect 42334 35694 42386 35746
rect 42386 35694 42388 35746
rect 42332 35692 42388 35694
rect 42492 35746 42548 35748
rect 42492 35694 42494 35746
rect 42494 35694 42546 35746
rect 42546 35694 42548 35746
rect 42492 35692 42548 35694
rect 42652 35746 42708 35748
rect 42652 35694 42654 35746
rect 42654 35694 42706 35746
rect 42706 35694 42708 35746
rect 42652 35692 42708 35694
rect 42812 35746 42868 35748
rect 42812 35694 42814 35746
rect 42814 35694 42866 35746
rect 42866 35694 42868 35746
rect 42812 35692 42868 35694
rect 42972 35746 43028 35748
rect 42972 35694 42974 35746
rect 42974 35694 43026 35746
rect 43026 35694 43028 35746
rect 42972 35692 43028 35694
rect 43132 35746 43188 35748
rect 43132 35694 43134 35746
rect 43134 35694 43186 35746
rect 43186 35694 43188 35746
rect 43132 35692 43188 35694
rect -31028 35612 -30972 35668
rect -30708 35612 -30652 35668
rect -30388 35612 -30332 35668
rect -30068 35612 -30012 35668
rect -3348 35532 -3292 35588
rect -3028 35532 -2972 35588
rect -2708 35532 -2652 35588
rect -2388 35532 -2332 35588
rect -2068 35532 -2012 35588
rect -1748 35532 -1692 35588
rect -1428 35532 -1372 35588
rect -1108 35532 -1052 35588
rect -31028 35452 -30972 35508
rect -30708 35452 -30652 35508
rect -30388 35452 -30332 35508
rect -30068 35452 -30012 35508
rect -3348 35372 -3292 35428
rect -3028 35372 -2972 35428
rect -2708 35372 -2652 35428
rect -2388 35372 -2332 35428
rect -2068 35372 -2012 35428
rect -1748 35372 -1692 35428
rect -1428 35372 -1372 35428
rect -1108 35372 -1052 35428
rect -31028 35292 -30972 35348
rect -30708 35292 -30652 35348
rect -30388 35292 -30332 35348
rect -30068 35292 -30012 35348
rect -3348 35212 -3292 35268
rect -3028 35212 -2972 35268
rect -2708 35212 -2652 35268
rect -2388 35212 -2332 35268
rect -2068 35212 -2012 35268
rect -1748 35212 -1692 35268
rect -1428 35212 -1372 35268
rect -1108 35212 -1052 35268
rect -31028 35132 -30972 35188
rect -30708 35132 -30652 35188
rect -30388 35132 -30332 35188
rect -30068 35132 -30012 35188
rect -3348 35052 -3292 35108
rect -3028 35052 -2972 35108
rect -2708 35052 -2652 35108
rect -2388 35052 -2332 35108
rect -2068 35052 -2012 35108
rect -1748 35052 -1692 35108
rect -1428 35052 -1372 35108
rect -1108 35052 -1052 35108
rect -31028 34972 -30972 35028
rect -30708 34972 -30652 35028
rect -30388 34972 -30332 35028
rect -30068 34972 -30012 35028
rect -3348 34892 -3292 34948
rect -3028 34892 -2972 34948
rect -2708 34892 -2652 34948
rect -2388 34892 -2332 34948
rect -2068 34892 -2012 34948
rect -1748 34892 -1692 34948
rect -1428 34892 -1372 34948
rect -1108 34892 -1052 34948
rect -31028 34812 -30972 34868
rect -30708 34812 -30652 34868
rect -30388 34812 -30332 34868
rect -30068 34812 -30012 34868
rect -3348 34732 -3292 34788
rect -3028 34732 -2972 34788
rect -2708 34732 -2652 34788
rect -2388 34732 -2332 34788
rect -2068 34732 -2012 34788
rect -1748 34732 -1692 34788
rect -1428 34732 -1372 34788
rect -1108 34732 -1052 34788
rect -33108 34706 -33052 34708
rect -33108 34654 -33106 34706
rect -33106 34654 -33054 34706
rect -33054 34654 -33052 34706
rect -33108 34652 -33052 34654
rect -32948 34706 -32892 34708
rect -32948 34654 -32946 34706
rect -32946 34654 -32894 34706
rect -32894 34654 -32892 34706
rect -32948 34652 -32892 34654
rect -32788 34706 -32732 34708
rect -32788 34654 -32786 34706
rect -32786 34654 -32734 34706
rect -32734 34654 -32732 34706
rect -32788 34652 -32732 34654
rect -32628 34706 -32572 34708
rect -32628 34654 -32626 34706
rect -32626 34654 -32574 34706
rect -32574 34654 -32572 34706
rect -32628 34652 -32572 34654
rect -32468 34706 -32412 34708
rect -32468 34654 -32466 34706
rect -32466 34654 -32414 34706
rect -32414 34654 -32412 34706
rect -32468 34652 -32412 34654
rect -32308 34706 -32252 34708
rect -32308 34654 -32306 34706
rect -32306 34654 -32254 34706
rect -32254 34654 -32252 34706
rect -32308 34652 -32252 34654
rect -32148 34706 -32092 34708
rect -32148 34654 -32146 34706
rect -32146 34654 -32094 34706
rect -32094 34654 -32092 34706
rect -32148 34652 -32092 34654
rect -31988 34706 -31932 34708
rect -31988 34654 -31986 34706
rect -31986 34654 -31934 34706
rect -31934 34654 -31932 34706
rect -31988 34652 -31932 34654
rect -31828 34706 -31772 34708
rect -31828 34654 -31826 34706
rect -31826 34654 -31774 34706
rect -31774 34654 -31772 34706
rect -31828 34652 -31772 34654
rect -31668 34706 -31612 34708
rect -31668 34654 -31666 34706
rect -31666 34654 -31614 34706
rect -31614 34654 -31612 34706
rect -31668 34652 -31612 34654
rect -31508 34706 -31452 34708
rect -31508 34654 -31506 34706
rect -31506 34654 -31454 34706
rect -31454 34654 -31452 34706
rect -31508 34652 -31452 34654
rect -31348 34706 -31292 34708
rect -31348 34654 -31346 34706
rect -31346 34654 -31294 34706
rect -31294 34654 -31292 34706
rect -31348 34652 -31292 34654
rect -31188 34706 -31132 34708
rect -31188 34654 -31186 34706
rect -31186 34654 -31134 34706
rect -31134 34654 -31132 34706
rect -31188 34652 -31132 34654
rect -31028 34652 -30972 34708
rect -30708 34652 -30652 34708
rect -30388 34652 -30332 34708
rect -30068 34652 -30012 34708
rect -29908 34706 -29852 34708
rect -29908 34654 -29906 34706
rect -29906 34654 -29854 34706
rect -29854 34654 -29852 34706
rect -29908 34652 -29852 34654
rect -29748 34706 -29692 34708
rect -29748 34654 -29746 34706
rect -29746 34654 -29694 34706
rect -29694 34654 -29692 34706
rect -29748 34652 -29692 34654
rect -29588 34706 -29532 34708
rect -29588 34654 -29586 34706
rect -29586 34654 -29534 34706
rect -29534 34654 -29532 34706
rect -29588 34652 -29532 34654
rect -29428 34706 -29372 34708
rect -29428 34654 -29426 34706
rect -29426 34654 -29374 34706
rect -29374 34654 -29372 34706
rect -29428 34652 -29372 34654
rect -29268 34706 -29212 34708
rect -29268 34654 -29266 34706
rect -29266 34654 -29214 34706
rect -29214 34654 -29212 34706
rect -29268 34652 -29212 34654
rect -29108 34706 -29052 34708
rect -29108 34654 -29106 34706
rect -29106 34654 -29054 34706
rect -29054 34654 -29052 34706
rect -29108 34652 -29052 34654
rect -28948 34706 -28892 34708
rect -28948 34654 -28946 34706
rect -28946 34654 -28894 34706
rect -28894 34654 -28892 34706
rect -28948 34652 -28892 34654
rect -28788 34706 -28732 34708
rect -28788 34654 -28786 34706
rect -28786 34654 -28734 34706
rect -28734 34654 -28732 34706
rect -28788 34652 -28732 34654
rect -28628 34706 -28572 34708
rect -28628 34654 -28626 34706
rect -28626 34654 -28574 34706
rect -28574 34654 -28572 34706
rect -28628 34652 -28572 34654
rect -28468 34706 -28412 34708
rect -28468 34654 -28466 34706
rect -28466 34654 -28414 34706
rect -28414 34654 -28412 34706
rect -28468 34652 -28412 34654
rect -28308 34706 -28252 34708
rect -28308 34654 -28306 34706
rect -28306 34654 -28254 34706
rect -28254 34654 -28252 34706
rect -28308 34652 -28252 34654
rect -28148 34706 -28092 34708
rect -28148 34654 -28146 34706
rect -28146 34654 -28094 34706
rect -28094 34654 -28092 34706
rect -28148 34652 -28092 34654
rect -27988 34706 -27932 34708
rect -27988 34654 -27986 34706
rect -27986 34654 -27934 34706
rect -27934 34654 -27932 34706
rect -27988 34652 -27932 34654
rect -27828 34706 -27772 34708
rect -27828 34654 -27826 34706
rect -27826 34654 -27774 34706
rect -27774 34654 -27772 34706
rect -27828 34652 -27772 34654
rect -27668 34706 -27612 34708
rect -27668 34654 -27666 34706
rect -27666 34654 -27614 34706
rect -27614 34654 -27612 34706
rect -27668 34652 -27612 34654
rect -27508 34706 -27452 34708
rect -27508 34654 -27506 34706
rect -27506 34654 -27454 34706
rect -27454 34654 -27452 34706
rect -27508 34652 -27452 34654
rect -27348 34706 -27292 34708
rect -27348 34654 -27346 34706
rect -27346 34654 -27294 34706
rect -27294 34654 -27292 34706
rect -27348 34652 -27292 34654
rect -27188 34706 -27132 34708
rect -27188 34654 -27186 34706
rect -27186 34654 -27134 34706
rect -27134 34654 -27132 34706
rect -27188 34652 -27132 34654
rect -27028 34706 -26972 34708
rect -27028 34654 -27026 34706
rect -27026 34654 -26974 34706
rect -26974 34654 -26972 34706
rect -27028 34652 -26972 34654
rect -26868 34706 -26812 34708
rect -26868 34654 -26866 34706
rect -26866 34654 -26814 34706
rect -26814 34654 -26812 34706
rect -26868 34652 -26812 34654
rect -26708 34706 -26652 34708
rect -26708 34654 -26706 34706
rect -26706 34654 -26654 34706
rect -26654 34654 -26652 34706
rect -26708 34652 -26652 34654
rect -26548 34706 -26492 34708
rect -26548 34654 -26546 34706
rect -26546 34654 -26494 34706
rect -26494 34654 -26492 34706
rect -26548 34652 -26492 34654
rect -26388 34706 -26332 34708
rect -26388 34654 -26386 34706
rect -26386 34654 -26334 34706
rect -26334 34654 -26332 34706
rect -26388 34652 -26332 34654
rect -26228 34706 -26172 34708
rect -26228 34654 -26226 34706
rect -26226 34654 -26174 34706
rect -26174 34654 -26172 34706
rect -26228 34652 -26172 34654
rect -26068 34706 -26012 34708
rect -26068 34654 -26066 34706
rect -26066 34654 -26014 34706
rect -26014 34654 -26012 34706
rect -26068 34652 -26012 34654
rect -25908 34706 -25852 34708
rect -25908 34654 -25906 34706
rect -25906 34654 -25854 34706
rect -25854 34654 -25852 34706
rect -25908 34652 -25852 34654
rect -25748 34706 -25692 34708
rect -25748 34654 -25746 34706
rect -25746 34654 -25694 34706
rect -25694 34654 -25692 34706
rect -25748 34652 -25692 34654
rect -25588 34706 -25532 34708
rect -25588 34654 -25586 34706
rect -25586 34654 -25534 34706
rect -25534 34654 -25532 34706
rect -25588 34652 -25532 34654
rect -25428 34706 -25372 34708
rect -25428 34654 -25426 34706
rect -25426 34654 -25374 34706
rect -25374 34654 -25372 34706
rect -25428 34652 -25372 34654
rect -25268 34706 -25212 34708
rect -25268 34654 -25266 34706
rect -25266 34654 -25214 34706
rect -25214 34654 -25212 34706
rect -25268 34652 -25212 34654
rect -25108 34706 -25052 34708
rect -25108 34654 -25106 34706
rect -25106 34654 -25054 34706
rect -25054 34654 -25052 34706
rect -25108 34652 -25052 34654
rect -24948 34706 -24892 34708
rect -24948 34654 -24946 34706
rect -24946 34654 -24894 34706
rect -24894 34654 -24892 34706
rect -24948 34652 -24892 34654
rect -24788 34706 -24732 34708
rect -24788 34654 -24786 34706
rect -24786 34654 -24734 34706
rect -24734 34654 -24732 34706
rect -24788 34652 -24732 34654
rect -24628 34706 -24572 34708
rect -24628 34654 -24626 34706
rect -24626 34654 -24574 34706
rect -24574 34654 -24572 34706
rect -24628 34652 -24572 34654
rect -24468 34706 -24412 34708
rect -24468 34654 -24466 34706
rect -24466 34654 -24414 34706
rect -24414 34654 -24412 34706
rect -24468 34652 -24412 34654
rect -24308 34706 -24252 34708
rect -24308 34654 -24306 34706
rect -24306 34654 -24254 34706
rect -24254 34654 -24252 34706
rect -24308 34652 -24252 34654
rect -24148 34706 -24092 34708
rect -24148 34654 -24146 34706
rect -24146 34654 -24094 34706
rect -24094 34654 -24092 34706
rect -24148 34652 -24092 34654
rect -23988 34706 -23932 34708
rect -23988 34654 -23986 34706
rect -23986 34654 -23934 34706
rect -23934 34654 -23932 34706
rect -23988 34652 -23932 34654
rect -23828 34706 -23772 34708
rect -23828 34654 -23826 34706
rect -23826 34654 -23774 34706
rect -23774 34654 -23772 34706
rect -23828 34652 -23772 34654
rect -23668 34706 -23612 34708
rect -23668 34654 -23666 34706
rect -23666 34654 -23614 34706
rect -23614 34654 -23612 34706
rect -23668 34652 -23612 34654
rect -23508 34706 -23452 34708
rect -23508 34654 -23506 34706
rect -23506 34654 -23454 34706
rect -23454 34654 -23452 34706
rect -23508 34652 -23452 34654
rect -23348 34706 -23292 34708
rect -23348 34654 -23346 34706
rect -23346 34654 -23294 34706
rect -23294 34654 -23292 34706
rect -23348 34652 -23292 34654
rect -23188 34706 -23132 34708
rect -23188 34654 -23186 34706
rect -23186 34654 -23134 34706
rect -23134 34654 -23132 34706
rect -23188 34652 -23132 34654
rect -23028 34706 -22972 34708
rect -23028 34654 -23026 34706
rect -23026 34654 -22974 34706
rect -22974 34654 -22972 34706
rect -23028 34652 -22972 34654
rect -22868 34706 -22812 34708
rect -22868 34654 -22866 34706
rect -22866 34654 -22814 34706
rect -22814 34654 -22812 34706
rect -22868 34652 -22812 34654
rect -22708 34706 -22652 34708
rect -22708 34654 -22706 34706
rect -22706 34654 -22654 34706
rect -22654 34654 -22652 34706
rect -22708 34652 -22652 34654
rect -22548 34706 -22492 34708
rect -22548 34654 -22546 34706
rect -22546 34654 -22494 34706
rect -22494 34654 -22492 34706
rect -22548 34652 -22492 34654
rect -22388 34706 -22332 34708
rect -22388 34654 -22386 34706
rect -22386 34654 -22334 34706
rect -22334 34654 -22332 34706
rect -22388 34652 -22332 34654
rect -22228 34706 -22172 34708
rect -22228 34654 -22226 34706
rect -22226 34654 -22174 34706
rect -22174 34654 -22172 34706
rect -22228 34652 -22172 34654
rect -22068 34706 -22012 34708
rect -22068 34654 -22066 34706
rect -22066 34654 -22014 34706
rect -22014 34654 -22012 34706
rect -22068 34652 -22012 34654
rect -21908 34706 -21852 34708
rect -21908 34654 -21906 34706
rect -21906 34654 -21854 34706
rect -21854 34654 -21852 34706
rect -21908 34652 -21852 34654
rect -21748 34706 -21692 34708
rect -21748 34654 -21746 34706
rect -21746 34654 -21694 34706
rect -21694 34654 -21692 34706
rect -21748 34652 -21692 34654
rect -21588 34706 -21532 34708
rect -21588 34654 -21586 34706
rect -21586 34654 -21534 34706
rect -21534 34654 -21532 34706
rect -21588 34652 -21532 34654
rect -21428 34706 -21372 34708
rect -21428 34654 -21426 34706
rect -21426 34654 -21374 34706
rect -21374 34654 -21372 34706
rect -21428 34652 -21372 34654
rect -21268 34706 -21212 34708
rect -21268 34654 -21266 34706
rect -21266 34654 -21214 34706
rect -21214 34654 -21212 34706
rect -21268 34652 -21212 34654
rect -21108 34706 -21052 34708
rect -21108 34654 -21106 34706
rect -21106 34654 -21054 34706
rect -21054 34654 -21052 34706
rect -21108 34652 -21052 34654
rect -20948 34706 -20892 34708
rect -20948 34654 -20946 34706
rect -20946 34654 -20894 34706
rect -20894 34654 -20892 34706
rect -20948 34652 -20892 34654
rect -20788 34706 -20732 34708
rect -20788 34654 -20786 34706
rect -20786 34654 -20734 34706
rect -20734 34654 -20732 34706
rect -20788 34652 -20732 34654
rect -20628 34706 -20572 34708
rect -20628 34654 -20626 34706
rect -20626 34654 -20574 34706
rect -20574 34654 -20572 34706
rect -20628 34652 -20572 34654
rect -20468 34706 -20412 34708
rect -20468 34654 -20466 34706
rect -20466 34654 -20414 34706
rect -20414 34654 -20412 34706
rect -20468 34652 -20412 34654
rect -20308 34706 -20252 34708
rect -20308 34654 -20306 34706
rect -20306 34654 -20254 34706
rect -20254 34654 -20252 34706
rect -20308 34652 -20252 34654
rect -20148 34706 -20092 34708
rect -20148 34654 -20146 34706
rect -20146 34654 -20094 34706
rect -20094 34654 -20092 34706
rect -20148 34652 -20092 34654
rect -19988 34706 -19932 34708
rect -19988 34654 -19986 34706
rect -19986 34654 -19934 34706
rect -19934 34654 -19932 34706
rect -19988 34652 -19932 34654
rect -19828 34706 -19772 34708
rect -19828 34654 -19826 34706
rect -19826 34654 -19774 34706
rect -19774 34654 -19772 34706
rect -19828 34652 -19772 34654
rect -19668 34706 -19612 34708
rect -19668 34654 -19666 34706
rect -19666 34654 -19614 34706
rect -19614 34654 -19612 34706
rect -19668 34652 -19612 34654
rect -19508 34706 -19452 34708
rect -19508 34654 -19506 34706
rect -19506 34654 -19454 34706
rect -19454 34654 -19452 34706
rect -19508 34652 -19452 34654
rect -19348 34706 -19292 34708
rect -19348 34654 -19346 34706
rect -19346 34654 -19294 34706
rect -19294 34654 -19292 34706
rect -19348 34652 -19292 34654
rect -19188 34706 -19132 34708
rect -19188 34654 -19186 34706
rect -19186 34654 -19134 34706
rect -19134 34654 -19132 34706
rect -19188 34652 -19132 34654
rect -19028 34706 -18972 34708
rect -19028 34654 -19026 34706
rect -19026 34654 -18974 34706
rect -18974 34654 -18972 34706
rect -19028 34652 -18972 34654
rect -18868 34706 -18812 34708
rect -18868 34654 -18866 34706
rect -18866 34654 -18814 34706
rect -18814 34654 -18812 34706
rect -18868 34652 -18812 34654
rect -18708 34706 -18652 34708
rect -18708 34654 -18706 34706
rect -18706 34654 -18654 34706
rect -18654 34654 -18652 34706
rect -18708 34652 -18652 34654
rect -18548 34706 -18492 34708
rect -18548 34654 -18546 34706
rect -18546 34654 -18494 34706
rect -18494 34654 -18492 34706
rect -18548 34652 -18492 34654
rect -18388 34706 -18332 34708
rect -18388 34654 -18386 34706
rect -18386 34654 -18334 34706
rect -18334 34654 -18332 34706
rect -18388 34652 -18332 34654
rect -18228 34706 -18172 34708
rect -18228 34654 -18226 34706
rect -18226 34654 -18174 34706
rect -18174 34654 -18172 34706
rect -18228 34652 -18172 34654
rect -18068 34706 -18012 34708
rect -18068 34654 -18066 34706
rect -18066 34654 -18014 34706
rect -18014 34654 -18012 34706
rect -18068 34652 -18012 34654
rect -17908 34706 -17852 34708
rect -17908 34654 -17906 34706
rect -17906 34654 -17854 34706
rect -17854 34654 -17852 34706
rect -17908 34652 -17852 34654
rect -17748 34706 -17692 34708
rect -17748 34654 -17746 34706
rect -17746 34654 -17694 34706
rect -17694 34654 -17692 34706
rect -17748 34652 -17692 34654
rect -17588 34706 -17532 34708
rect -17588 34654 -17586 34706
rect -17586 34654 -17534 34706
rect -17534 34654 -17532 34706
rect -17588 34652 -17532 34654
rect -17428 34706 -17372 34708
rect -17428 34654 -17426 34706
rect -17426 34654 -17374 34706
rect -17374 34654 -17372 34706
rect -17428 34652 -17372 34654
rect -17268 34706 -17212 34708
rect -17268 34654 -17266 34706
rect -17266 34654 -17214 34706
rect -17214 34654 -17212 34706
rect -17268 34652 -17212 34654
rect -17108 34706 -17052 34708
rect -17108 34654 -17106 34706
rect -17106 34654 -17054 34706
rect -17054 34654 -17052 34706
rect -17108 34652 -17052 34654
rect -16948 34706 -16892 34708
rect -16948 34654 -16946 34706
rect -16946 34654 -16894 34706
rect -16894 34654 -16892 34706
rect -16948 34652 -16892 34654
rect -16788 34706 -16732 34708
rect -16788 34654 -16786 34706
rect -16786 34654 -16734 34706
rect -16734 34654 -16732 34706
rect -16788 34652 -16732 34654
rect -16628 34706 -16572 34708
rect -16628 34654 -16626 34706
rect -16626 34654 -16574 34706
rect -16574 34654 -16572 34706
rect -16628 34652 -16572 34654
rect -16468 34706 -16412 34708
rect -16468 34654 -16466 34706
rect -16466 34654 -16414 34706
rect -16414 34654 -16412 34706
rect -16468 34652 -16412 34654
rect -16308 34706 -16252 34708
rect -16308 34654 -16306 34706
rect -16306 34654 -16254 34706
rect -16254 34654 -16252 34706
rect -16308 34652 -16252 34654
rect -16148 34706 -16092 34708
rect -16148 34654 -16146 34706
rect -16146 34654 -16094 34706
rect -16094 34654 -16092 34706
rect -16148 34652 -16092 34654
rect -15988 34706 -15932 34708
rect -15988 34654 -15986 34706
rect -15986 34654 -15934 34706
rect -15934 34654 -15932 34706
rect -15988 34652 -15932 34654
rect -15828 34706 -15772 34708
rect -15828 34654 -15826 34706
rect -15826 34654 -15774 34706
rect -15774 34654 -15772 34706
rect -15828 34652 -15772 34654
rect -15668 34706 -15612 34708
rect -15668 34654 -15666 34706
rect -15666 34654 -15614 34706
rect -15614 34654 -15612 34706
rect -15668 34652 -15612 34654
rect -15508 34706 -15452 34708
rect -15508 34654 -15506 34706
rect -15506 34654 -15454 34706
rect -15454 34654 -15452 34706
rect -15508 34652 -15452 34654
rect -15348 34706 -15292 34708
rect -15348 34654 -15346 34706
rect -15346 34654 -15294 34706
rect -15294 34654 -15292 34706
rect -15348 34652 -15292 34654
rect -15188 34706 -15132 34708
rect -15188 34654 -15186 34706
rect -15186 34654 -15134 34706
rect -15134 34654 -15132 34706
rect -15188 34652 -15132 34654
rect -15028 34706 -14972 34708
rect -15028 34654 -15026 34706
rect -15026 34654 -14974 34706
rect -14974 34654 -14972 34706
rect -15028 34652 -14972 34654
rect -14868 34706 -14812 34708
rect -14868 34654 -14866 34706
rect -14866 34654 -14814 34706
rect -14814 34654 -14812 34706
rect -14868 34652 -14812 34654
rect -14708 34706 -14652 34708
rect -14708 34654 -14706 34706
rect -14706 34654 -14654 34706
rect -14654 34654 -14652 34706
rect -14708 34652 -14652 34654
rect -14548 34706 -14492 34708
rect -14548 34654 -14546 34706
rect -14546 34654 -14494 34706
rect -14494 34654 -14492 34706
rect -14548 34652 -14492 34654
rect -14388 34706 -14332 34708
rect -14388 34654 -14386 34706
rect -14386 34654 -14334 34706
rect -14334 34654 -14332 34706
rect -14388 34652 -14332 34654
rect -14228 34706 -14172 34708
rect -14228 34654 -14226 34706
rect -14226 34654 -14174 34706
rect -14174 34654 -14172 34706
rect -14228 34652 -14172 34654
rect -14068 34706 -14012 34708
rect -14068 34654 -14066 34706
rect -14066 34654 -14014 34706
rect -14014 34654 -14012 34706
rect -14068 34652 -14012 34654
rect -13908 34706 -13852 34708
rect -13908 34654 -13906 34706
rect -13906 34654 -13854 34706
rect -13854 34654 -13852 34706
rect -13908 34652 -13852 34654
rect -13748 34706 -13692 34708
rect -13748 34654 -13746 34706
rect -13746 34654 -13694 34706
rect -13694 34654 -13692 34706
rect -13748 34652 -13692 34654
rect -13588 34706 -13532 34708
rect -13588 34654 -13586 34706
rect -13586 34654 -13534 34706
rect -13534 34654 -13532 34706
rect -13588 34652 -13532 34654
rect -13428 34706 -13372 34708
rect -13428 34654 -13426 34706
rect -13426 34654 -13374 34706
rect -13374 34654 -13372 34706
rect -13428 34652 -13372 34654
rect -13268 34706 -13212 34708
rect -13268 34654 -13266 34706
rect -13266 34654 -13214 34706
rect -13214 34654 -13212 34706
rect -13268 34652 -13212 34654
rect -13108 34706 -13052 34708
rect -13108 34654 -13106 34706
rect -13106 34654 -13054 34706
rect -13054 34654 -13052 34706
rect -13108 34652 -13052 34654
rect -12948 34706 -12892 34708
rect -12948 34654 -12946 34706
rect -12946 34654 -12894 34706
rect -12894 34654 -12892 34706
rect -12948 34652 -12892 34654
rect -12788 34706 -12732 34708
rect -12788 34654 -12786 34706
rect -12786 34654 -12734 34706
rect -12734 34654 -12732 34706
rect -12788 34652 -12732 34654
rect -12628 34706 -12572 34708
rect -12628 34654 -12626 34706
rect -12626 34654 -12574 34706
rect -12574 34654 -12572 34706
rect -12628 34652 -12572 34654
rect -12468 34706 -12412 34708
rect -12468 34654 -12466 34706
rect -12466 34654 -12414 34706
rect -12414 34654 -12412 34706
rect -12468 34652 -12412 34654
rect -12308 34706 -12252 34708
rect -12308 34654 -12306 34706
rect -12306 34654 -12254 34706
rect -12254 34654 -12252 34706
rect -12308 34652 -12252 34654
rect -12148 34706 -12092 34708
rect -12148 34654 -12146 34706
rect -12146 34654 -12094 34706
rect -12094 34654 -12092 34706
rect -12148 34652 -12092 34654
rect -11988 34706 -11932 34708
rect -11988 34654 -11986 34706
rect -11986 34654 -11934 34706
rect -11934 34654 -11932 34706
rect -11988 34652 -11932 34654
rect -11828 34706 -11772 34708
rect -11828 34654 -11826 34706
rect -11826 34654 -11774 34706
rect -11774 34654 -11772 34706
rect -11828 34652 -11772 34654
rect -11668 34706 -11612 34708
rect -11668 34654 -11666 34706
rect -11666 34654 -11614 34706
rect -11614 34654 -11612 34706
rect -11668 34652 -11612 34654
rect -11508 34706 -11452 34708
rect -11508 34654 -11506 34706
rect -11506 34654 -11454 34706
rect -11454 34654 -11452 34706
rect -11508 34652 -11452 34654
rect -11188 34652 -11132 34708
rect -10868 34706 -10812 34708
rect -10868 34654 -10866 34706
rect -10866 34654 -10814 34706
rect -10814 34654 -10812 34706
rect -10868 34652 -10812 34654
rect -10548 34706 -10492 34708
rect -10548 34654 -10546 34706
rect -10546 34654 -10494 34706
rect -10494 34654 -10492 34706
rect -10548 34652 -10492 34654
rect -3348 34572 -3292 34628
rect -3028 34572 -2972 34628
rect -2708 34572 -2652 34628
rect -2388 34572 -2332 34628
rect -2068 34572 -2012 34628
rect -1748 34572 -1692 34628
rect -1428 34572 -1372 34628
rect -1108 34572 -1052 34628
rect -10708 34492 -10652 34548
rect -3348 34412 -3292 34468
rect -3028 34412 -2972 34468
rect -2708 34412 -2652 34468
rect -2388 34412 -2332 34468
rect -2068 34412 -2012 34468
rect -1748 34412 -1692 34468
rect -1428 34412 -1372 34468
rect -1108 34412 -1052 34468
rect -33108 34386 -33052 34388
rect -33108 34334 -33106 34386
rect -33106 34334 -33054 34386
rect -33054 34334 -33052 34386
rect -33108 34332 -33052 34334
rect -32948 34386 -32892 34388
rect -32948 34334 -32946 34386
rect -32946 34334 -32894 34386
rect -32894 34334 -32892 34386
rect -32948 34332 -32892 34334
rect -32788 34386 -32732 34388
rect -32788 34334 -32786 34386
rect -32786 34334 -32734 34386
rect -32734 34334 -32732 34386
rect -32788 34332 -32732 34334
rect -32628 34386 -32572 34388
rect -32628 34334 -32626 34386
rect -32626 34334 -32574 34386
rect -32574 34334 -32572 34386
rect -32628 34332 -32572 34334
rect -32468 34386 -32412 34388
rect -32468 34334 -32466 34386
rect -32466 34334 -32414 34386
rect -32414 34334 -32412 34386
rect -32468 34332 -32412 34334
rect -32308 34386 -32252 34388
rect -32308 34334 -32306 34386
rect -32306 34334 -32254 34386
rect -32254 34334 -32252 34386
rect -32308 34332 -32252 34334
rect -32148 34386 -32092 34388
rect -32148 34334 -32146 34386
rect -32146 34334 -32094 34386
rect -32094 34334 -32092 34386
rect -32148 34332 -32092 34334
rect -31988 34386 -31932 34388
rect -31988 34334 -31986 34386
rect -31986 34334 -31934 34386
rect -31934 34334 -31932 34386
rect -31988 34332 -31932 34334
rect -31828 34386 -31772 34388
rect -31828 34334 -31826 34386
rect -31826 34334 -31774 34386
rect -31774 34334 -31772 34386
rect -31828 34332 -31772 34334
rect -31668 34386 -31612 34388
rect -31668 34334 -31666 34386
rect -31666 34334 -31614 34386
rect -31614 34334 -31612 34386
rect -31668 34332 -31612 34334
rect -31508 34386 -31452 34388
rect -31508 34334 -31506 34386
rect -31506 34334 -31454 34386
rect -31454 34334 -31452 34386
rect -31508 34332 -31452 34334
rect -31348 34386 -31292 34388
rect -31348 34334 -31346 34386
rect -31346 34334 -31294 34386
rect -31294 34334 -31292 34386
rect -31348 34332 -31292 34334
rect -31188 34386 -31132 34388
rect -31188 34334 -31186 34386
rect -31186 34334 -31134 34386
rect -31134 34334 -31132 34386
rect -31188 34332 -31132 34334
rect -31028 34332 -30972 34388
rect -30708 34332 -30652 34388
rect -30388 34332 -30332 34388
rect -30068 34332 -30012 34388
rect -29908 34386 -29852 34388
rect -29908 34334 -29906 34386
rect -29906 34334 -29854 34386
rect -29854 34334 -29852 34386
rect -29908 34332 -29852 34334
rect -29748 34386 -29692 34388
rect -29748 34334 -29746 34386
rect -29746 34334 -29694 34386
rect -29694 34334 -29692 34386
rect -29748 34332 -29692 34334
rect -29588 34386 -29532 34388
rect -29588 34334 -29586 34386
rect -29586 34334 -29534 34386
rect -29534 34334 -29532 34386
rect -29588 34332 -29532 34334
rect -29428 34386 -29372 34388
rect -29428 34334 -29426 34386
rect -29426 34334 -29374 34386
rect -29374 34334 -29372 34386
rect -29428 34332 -29372 34334
rect -29268 34386 -29212 34388
rect -29268 34334 -29266 34386
rect -29266 34334 -29214 34386
rect -29214 34334 -29212 34386
rect -29268 34332 -29212 34334
rect -29108 34386 -29052 34388
rect -29108 34334 -29106 34386
rect -29106 34334 -29054 34386
rect -29054 34334 -29052 34386
rect -29108 34332 -29052 34334
rect -28948 34386 -28892 34388
rect -28948 34334 -28946 34386
rect -28946 34334 -28894 34386
rect -28894 34334 -28892 34386
rect -28948 34332 -28892 34334
rect -28788 34386 -28732 34388
rect -28788 34334 -28786 34386
rect -28786 34334 -28734 34386
rect -28734 34334 -28732 34386
rect -28788 34332 -28732 34334
rect -28628 34386 -28572 34388
rect -28628 34334 -28626 34386
rect -28626 34334 -28574 34386
rect -28574 34334 -28572 34386
rect -28628 34332 -28572 34334
rect -28468 34386 -28412 34388
rect -28468 34334 -28466 34386
rect -28466 34334 -28414 34386
rect -28414 34334 -28412 34386
rect -28468 34332 -28412 34334
rect -28308 34386 -28252 34388
rect -28308 34334 -28306 34386
rect -28306 34334 -28254 34386
rect -28254 34334 -28252 34386
rect -28308 34332 -28252 34334
rect -28148 34386 -28092 34388
rect -28148 34334 -28146 34386
rect -28146 34334 -28094 34386
rect -28094 34334 -28092 34386
rect -28148 34332 -28092 34334
rect -27988 34386 -27932 34388
rect -27988 34334 -27986 34386
rect -27986 34334 -27934 34386
rect -27934 34334 -27932 34386
rect -27988 34332 -27932 34334
rect -27828 34386 -27772 34388
rect -27828 34334 -27826 34386
rect -27826 34334 -27774 34386
rect -27774 34334 -27772 34386
rect -27828 34332 -27772 34334
rect -27668 34386 -27612 34388
rect -27668 34334 -27666 34386
rect -27666 34334 -27614 34386
rect -27614 34334 -27612 34386
rect -27668 34332 -27612 34334
rect -27508 34386 -27452 34388
rect -27508 34334 -27506 34386
rect -27506 34334 -27454 34386
rect -27454 34334 -27452 34386
rect -27508 34332 -27452 34334
rect -27348 34386 -27292 34388
rect -27348 34334 -27346 34386
rect -27346 34334 -27294 34386
rect -27294 34334 -27292 34386
rect -27348 34332 -27292 34334
rect -27188 34386 -27132 34388
rect -27188 34334 -27186 34386
rect -27186 34334 -27134 34386
rect -27134 34334 -27132 34386
rect -27188 34332 -27132 34334
rect -27028 34386 -26972 34388
rect -27028 34334 -27026 34386
rect -27026 34334 -26974 34386
rect -26974 34334 -26972 34386
rect -27028 34332 -26972 34334
rect -26868 34386 -26812 34388
rect -26868 34334 -26866 34386
rect -26866 34334 -26814 34386
rect -26814 34334 -26812 34386
rect -26868 34332 -26812 34334
rect -26708 34386 -26652 34388
rect -26708 34334 -26706 34386
rect -26706 34334 -26654 34386
rect -26654 34334 -26652 34386
rect -26708 34332 -26652 34334
rect -26548 34386 -26492 34388
rect -26548 34334 -26546 34386
rect -26546 34334 -26494 34386
rect -26494 34334 -26492 34386
rect -26548 34332 -26492 34334
rect -26388 34386 -26332 34388
rect -26388 34334 -26386 34386
rect -26386 34334 -26334 34386
rect -26334 34334 -26332 34386
rect -26388 34332 -26332 34334
rect -26228 34386 -26172 34388
rect -26228 34334 -26226 34386
rect -26226 34334 -26174 34386
rect -26174 34334 -26172 34386
rect -26228 34332 -26172 34334
rect -26068 34386 -26012 34388
rect -26068 34334 -26066 34386
rect -26066 34334 -26014 34386
rect -26014 34334 -26012 34386
rect -26068 34332 -26012 34334
rect -25908 34386 -25852 34388
rect -25908 34334 -25906 34386
rect -25906 34334 -25854 34386
rect -25854 34334 -25852 34386
rect -25908 34332 -25852 34334
rect -25748 34386 -25692 34388
rect -25748 34334 -25746 34386
rect -25746 34334 -25694 34386
rect -25694 34334 -25692 34386
rect -25748 34332 -25692 34334
rect -25588 34386 -25532 34388
rect -25588 34334 -25586 34386
rect -25586 34334 -25534 34386
rect -25534 34334 -25532 34386
rect -25588 34332 -25532 34334
rect -25428 34386 -25372 34388
rect -25428 34334 -25426 34386
rect -25426 34334 -25374 34386
rect -25374 34334 -25372 34386
rect -25428 34332 -25372 34334
rect -25268 34386 -25212 34388
rect -25268 34334 -25266 34386
rect -25266 34334 -25214 34386
rect -25214 34334 -25212 34386
rect -25268 34332 -25212 34334
rect -25108 34386 -25052 34388
rect -25108 34334 -25106 34386
rect -25106 34334 -25054 34386
rect -25054 34334 -25052 34386
rect -25108 34332 -25052 34334
rect -24948 34386 -24892 34388
rect -24948 34334 -24946 34386
rect -24946 34334 -24894 34386
rect -24894 34334 -24892 34386
rect -24948 34332 -24892 34334
rect -24788 34386 -24732 34388
rect -24788 34334 -24786 34386
rect -24786 34334 -24734 34386
rect -24734 34334 -24732 34386
rect -24788 34332 -24732 34334
rect -24628 34386 -24572 34388
rect -24628 34334 -24626 34386
rect -24626 34334 -24574 34386
rect -24574 34334 -24572 34386
rect -24628 34332 -24572 34334
rect -24468 34386 -24412 34388
rect -24468 34334 -24466 34386
rect -24466 34334 -24414 34386
rect -24414 34334 -24412 34386
rect -24468 34332 -24412 34334
rect -24308 34386 -24252 34388
rect -24308 34334 -24306 34386
rect -24306 34334 -24254 34386
rect -24254 34334 -24252 34386
rect -24308 34332 -24252 34334
rect -24148 34386 -24092 34388
rect -24148 34334 -24146 34386
rect -24146 34334 -24094 34386
rect -24094 34334 -24092 34386
rect -24148 34332 -24092 34334
rect -23988 34386 -23932 34388
rect -23988 34334 -23986 34386
rect -23986 34334 -23934 34386
rect -23934 34334 -23932 34386
rect -23988 34332 -23932 34334
rect -23828 34386 -23772 34388
rect -23828 34334 -23826 34386
rect -23826 34334 -23774 34386
rect -23774 34334 -23772 34386
rect -23828 34332 -23772 34334
rect -23668 34386 -23612 34388
rect -23668 34334 -23666 34386
rect -23666 34334 -23614 34386
rect -23614 34334 -23612 34386
rect -23668 34332 -23612 34334
rect -23508 34386 -23452 34388
rect -23508 34334 -23506 34386
rect -23506 34334 -23454 34386
rect -23454 34334 -23452 34386
rect -23508 34332 -23452 34334
rect -23348 34386 -23292 34388
rect -23348 34334 -23346 34386
rect -23346 34334 -23294 34386
rect -23294 34334 -23292 34386
rect -23348 34332 -23292 34334
rect -23188 34386 -23132 34388
rect -23188 34334 -23186 34386
rect -23186 34334 -23134 34386
rect -23134 34334 -23132 34386
rect -23188 34332 -23132 34334
rect -23028 34386 -22972 34388
rect -23028 34334 -23026 34386
rect -23026 34334 -22974 34386
rect -22974 34334 -22972 34386
rect -23028 34332 -22972 34334
rect -22868 34386 -22812 34388
rect -22868 34334 -22866 34386
rect -22866 34334 -22814 34386
rect -22814 34334 -22812 34386
rect -22868 34332 -22812 34334
rect -22708 34386 -22652 34388
rect -22708 34334 -22706 34386
rect -22706 34334 -22654 34386
rect -22654 34334 -22652 34386
rect -22708 34332 -22652 34334
rect -22548 34386 -22492 34388
rect -22548 34334 -22546 34386
rect -22546 34334 -22494 34386
rect -22494 34334 -22492 34386
rect -22548 34332 -22492 34334
rect -22388 34386 -22332 34388
rect -22388 34334 -22386 34386
rect -22386 34334 -22334 34386
rect -22334 34334 -22332 34386
rect -22388 34332 -22332 34334
rect -22228 34386 -22172 34388
rect -22228 34334 -22226 34386
rect -22226 34334 -22174 34386
rect -22174 34334 -22172 34386
rect -22228 34332 -22172 34334
rect -22068 34386 -22012 34388
rect -22068 34334 -22066 34386
rect -22066 34334 -22014 34386
rect -22014 34334 -22012 34386
rect -22068 34332 -22012 34334
rect -21908 34386 -21852 34388
rect -21908 34334 -21906 34386
rect -21906 34334 -21854 34386
rect -21854 34334 -21852 34386
rect -21908 34332 -21852 34334
rect -21748 34386 -21692 34388
rect -21748 34334 -21746 34386
rect -21746 34334 -21694 34386
rect -21694 34334 -21692 34386
rect -21748 34332 -21692 34334
rect -21588 34386 -21532 34388
rect -21588 34334 -21586 34386
rect -21586 34334 -21534 34386
rect -21534 34334 -21532 34386
rect -21588 34332 -21532 34334
rect -21428 34386 -21372 34388
rect -21428 34334 -21426 34386
rect -21426 34334 -21374 34386
rect -21374 34334 -21372 34386
rect -21428 34332 -21372 34334
rect -21268 34386 -21212 34388
rect -21268 34334 -21266 34386
rect -21266 34334 -21214 34386
rect -21214 34334 -21212 34386
rect -21268 34332 -21212 34334
rect -21108 34386 -21052 34388
rect -21108 34334 -21106 34386
rect -21106 34334 -21054 34386
rect -21054 34334 -21052 34386
rect -21108 34332 -21052 34334
rect -20948 34386 -20892 34388
rect -20948 34334 -20946 34386
rect -20946 34334 -20894 34386
rect -20894 34334 -20892 34386
rect -20948 34332 -20892 34334
rect -20788 34386 -20732 34388
rect -20788 34334 -20786 34386
rect -20786 34334 -20734 34386
rect -20734 34334 -20732 34386
rect -20788 34332 -20732 34334
rect -20628 34386 -20572 34388
rect -20628 34334 -20626 34386
rect -20626 34334 -20574 34386
rect -20574 34334 -20572 34386
rect -20628 34332 -20572 34334
rect -20468 34386 -20412 34388
rect -20468 34334 -20466 34386
rect -20466 34334 -20414 34386
rect -20414 34334 -20412 34386
rect -20468 34332 -20412 34334
rect -20308 34386 -20252 34388
rect -20308 34334 -20306 34386
rect -20306 34334 -20254 34386
rect -20254 34334 -20252 34386
rect -20308 34332 -20252 34334
rect -20148 34386 -20092 34388
rect -20148 34334 -20146 34386
rect -20146 34334 -20094 34386
rect -20094 34334 -20092 34386
rect -20148 34332 -20092 34334
rect -19988 34386 -19932 34388
rect -19988 34334 -19986 34386
rect -19986 34334 -19934 34386
rect -19934 34334 -19932 34386
rect -19988 34332 -19932 34334
rect -19828 34386 -19772 34388
rect -19828 34334 -19826 34386
rect -19826 34334 -19774 34386
rect -19774 34334 -19772 34386
rect -19828 34332 -19772 34334
rect -19668 34386 -19612 34388
rect -19668 34334 -19666 34386
rect -19666 34334 -19614 34386
rect -19614 34334 -19612 34386
rect -19668 34332 -19612 34334
rect -19508 34386 -19452 34388
rect -19508 34334 -19506 34386
rect -19506 34334 -19454 34386
rect -19454 34334 -19452 34386
rect -19508 34332 -19452 34334
rect -19348 34386 -19292 34388
rect -19348 34334 -19346 34386
rect -19346 34334 -19294 34386
rect -19294 34334 -19292 34386
rect -19348 34332 -19292 34334
rect -19188 34386 -19132 34388
rect -19188 34334 -19186 34386
rect -19186 34334 -19134 34386
rect -19134 34334 -19132 34386
rect -19188 34332 -19132 34334
rect -19028 34386 -18972 34388
rect -19028 34334 -19026 34386
rect -19026 34334 -18974 34386
rect -18974 34334 -18972 34386
rect -19028 34332 -18972 34334
rect -18868 34386 -18812 34388
rect -18868 34334 -18866 34386
rect -18866 34334 -18814 34386
rect -18814 34334 -18812 34386
rect -18868 34332 -18812 34334
rect -18708 34386 -18652 34388
rect -18708 34334 -18706 34386
rect -18706 34334 -18654 34386
rect -18654 34334 -18652 34386
rect -18708 34332 -18652 34334
rect -18548 34386 -18492 34388
rect -18548 34334 -18546 34386
rect -18546 34334 -18494 34386
rect -18494 34334 -18492 34386
rect -18548 34332 -18492 34334
rect -18388 34386 -18332 34388
rect -18388 34334 -18386 34386
rect -18386 34334 -18334 34386
rect -18334 34334 -18332 34386
rect -18388 34332 -18332 34334
rect -18228 34386 -18172 34388
rect -18228 34334 -18226 34386
rect -18226 34334 -18174 34386
rect -18174 34334 -18172 34386
rect -18228 34332 -18172 34334
rect -18068 34386 -18012 34388
rect -18068 34334 -18066 34386
rect -18066 34334 -18014 34386
rect -18014 34334 -18012 34386
rect -18068 34332 -18012 34334
rect -17908 34386 -17852 34388
rect -17908 34334 -17906 34386
rect -17906 34334 -17854 34386
rect -17854 34334 -17852 34386
rect -17908 34332 -17852 34334
rect -17748 34386 -17692 34388
rect -17748 34334 -17746 34386
rect -17746 34334 -17694 34386
rect -17694 34334 -17692 34386
rect -17748 34332 -17692 34334
rect -17588 34386 -17532 34388
rect -17588 34334 -17586 34386
rect -17586 34334 -17534 34386
rect -17534 34334 -17532 34386
rect -17588 34332 -17532 34334
rect -17428 34386 -17372 34388
rect -17428 34334 -17426 34386
rect -17426 34334 -17374 34386
rect -17374 34334 -17372 34386
rect -17428 34332 -17372 34334
rect -17268 34386 -17212 34388
rect -17268 34334 -17266 34386
rect -17266 34334 -17214 34386
rect -17214 34334 -17212 34386
rect -17268 34332 -17212 34334
rect -17108 34386 -17052 34388
rect -17108 34334 -17106 34386
rect -17106 34334 -17054 34386
rect -17054 34334 -17052 34386
rect -17108 34332 -17052 34334
rect -16948 34386 -16892 34388
rect -16948 34334 -16946 34386
rect -16946 34334 -16894 34386
rect -16894 34334 -16892 34386
rect -16948 34332 -16892 34334
rect -16788 34386 -16732 34388
rect -16788 34334 -16786 34386
rect -16786 34334 -16734 34386
rect -16734 34334 -16732 34386
rect -16788 34332 -16732 34334
rect -16628 34386 -16572 34388
rect -16628 34334 -16626 34386
rect -16626 34334 -16574 34386
rect -16574 34334 -16572 34386
rect -16628 34332 -16572 34334
rect -16468 34386 -16412 34388
rect -16468 34334 -16466 34386
rect -16466 34334 -16414 34386
rect -16414 34334 -16412 34386
rect -16468 34332 -16412 34334
rect -16308 34386 -16252 34388
rect -16308 34334 -16306 34386
rect -16306 34334 -16254 34386
rect -16254 34334 -16252 34386
rect -16308 34332 -16252 34334
rect -16148 34386 -16092 34388
rect -16148 34334 -16146 34386
rect -16146 34334 -16094 34386
rect -16094 34334 -16092 34386
rect -16148 34332 -16092 34334
rect -15988 34386 -15932 34388
rect -15988 34334 -15986 34386
rect -15986 34334 -15934 34386
rect -15934 34334 -15932 34386
rect -15988 34332 -15932 34334
rect -15828 34386 -15772 34388
rect -15828 34334 -15826 34386
rect -15826 34334 -15774 34386
rect -15774 34334 -15772 34386
rect -15828 34332 -15772 34334
rect -15668 34386 -15612 34388
rect -15668 34334 -15666 34386
rect -15666 34334 -15614 34386
rect -15614 34334 -15612 34386
rect -15668 34332 -15612 34334
rect -15508 34386 -15452 34388
rect -15508 34334 -15506 34386
rect -15506 34334 -15454 34386
rect -15454 34334 -15452 34386
rect -15508 34332 -15452 34334
rect -15348 34386 -15292 34388
rect -15348 34334 -15346 34386
rect -15346 34334 -15294 34386
rect -15294 34334 -15292 34386
rect -15348 34332 -15292 34334
rect -15188 34386 -15132 34388
rect -15188 34334 -15186 34386
rect -15186 34334 -15134 34386
rect -15134 34334 -15132 34386
rect -15188 34332 -15132 34334
rect -15028 34386 -14972 34388
rect -15028 34334 -15026 34386
rect -15026 34334 -14974 34386
rect -14974 34334 -14972 34386
rect -15028 34332 -14972 34334
rect -14868 34386 -14812 34388
rect -14868 34334 -14866 34386
rect -14866 34334 -14814 34386
rect -14814 34334 -14812 34386
rect -14868 34332 -14812 34334
rect -14708 34386 -14652 34388
rect -14708 34334 -14706 34386
rect -14706 34334 -14654 34386
rect -14654 34334 -14652 34386
rect -14708 34332 -14652 34334
rect -14548 34386 -14492 34388
rect -14548 34334 -14546 34386
rect -14546 34334 -14494 34386
rect -14494 34334 -14492 34386
rect -14548 34332 -14492 34334
rect -14388 34386 -14332 34388
rect -14388 34334 -14386 34386
rect -14386 34334 -14334 34386
rect -14334 34334 -14332 34386
rect -14388 34332 -14332 34334
rect -14228 34386 -14172 34388
rect -14228 34334 -14226 34386
rect -14226 34334 -14174 34386
rect -14174 34334 -14172 34386
rect -14228 34332 -14172 34334
rect -14068 34386 -14012 34388
rect -14068 34334 -14066 34386
rect -14066 34334 -14014 34386
rect -14014 34334 -14012 34386
rect -14068 34332 -14012 34334
rect -13908 34386 -13852 34388
rect -13908 34334 -13906 34386
rect -13906 34334 -13854 34386
rect -13854 34334 -13852 34386
rect -13908 34332 -13852 34334
rect -13748 34386 -13692 34388
rect -13748 34334 -13746 34386
rect -13746 34334 -13694 34386
rect -13694 34334 -13692 34386
rect -13748 34332 -13692 34334
rect -13588 34386 -13532 34388
rect -13588 34334 -13586 34386
rect -13586 34334 -13534 34386
rect -13534 34334 -13532 34386
rect -13588 34332 -13532 34334
rect -13428 34386 -13372 34388
rect -13428 34334 -13426 34386
rect -13426 34334 -13374 34386
rect -13374 34334 -13372 34386
rect -13428 34332 -13372 34334
rect -13268 34386 -13212 34388
rect -13268 34334 -13266 34386
rect -13266 34334 -13214 34386
rect -13214 34334 -13212 34386
rect -13268 34332 -13212 34334
rect -13108 34386 -13052 34388
rect -13108 34334 -13106 34386
rect -13106 34334 -13054 34386
rect -13054 34334 -13052 34386
rect -13108 34332 -13052 34334
rect -12948 34386 -12892 34388
rect -12948 34334 -12946 34386
rect -12946 34334 -12894 34386
rect -12894 34334 -12892 34386
rect -12948 34332 -12892 34334
rect -12788 34386 -12732 34388
rect -12788 34334 -12786 34386
rect -12786 34334 -12734 34386
rect -12734 34334 -12732 34386
rect -12788 34332 -12732 34334
rect -12628 34386 -12572 34388
rect -12628 34334 -12626 34386
rect -12626 34334 -12574 34386
rect -12574 34334 -12572 34386
rect -12628 34332 -12572 34334
rect -12468 34386 -12412 34388
rect -12468 34334 -12466 34386
rect -12466 34334 -12414 34386
rect -12414 34334 -12412 34386
rect -12468 34332 -12412 34334
rect -12308 34386 -12252 34388
rect -12308 34334 -12306 34386
rect -12306 34334 -12254 34386
rect -12254 34334 -12252 34386
rect -12308 34332 -12252 34334
rect -12148 34386 -12092 34388
rect -12148 34334 -12146 34386
rect -12146 34334 -12094 34386
rect -12094 34334 -12092 34386
rect -12148 34332 -12092 34334
rect -11988 34386 -11932 34388
rect -11988 34334 -11986 34386
rect -11986 34334 -11934 34386
rect -11934 34334 -11932 34386
rect -11988 34332 -11932 34334
rect -11828 34386 -11772 34388
rect -11828 34334 -11826 34386
rect -11826 34334 -11774 34386
rect -11774 34334 -11772 34386
rect -11828 34332 -11772 34334
rect -11668 34386 -11612 34388
rect -11668 34334 -11666 34386
rect -11666 34334 -11614 34386
rect -11614 34334 -11612 34386
rect -11668 34332 -11612 34334
rect -11508 34386 -11452 34388
rect -11508 34334 -11506 34386
rect -11506 34334 -11454 34386
rect -11454 34334 -11452 34386
rect -11508 34332 -11452 34334
rect -11188 34332 -11132 34388
rect -10868 34386 -10812 34388
rect -10868 34334 -10866 34386
rect -10866 34334 -10814 34386
rect -10814 34334 -10812 34386
rect -10868 34332 -10812 34334
rect -10548 34386 -10492 34388
rect -10548 34334 -10546 34386
rect -10546 34334 -10494 34386
rect -10494 34334 -10492 34386
rect -10548 34332 -10492 34334
rect -3348 34252 -3292 34308
rect -3028 34252 -2972 34308
rect -2708 34252 -2652 34308
rect -2388 34252 -2332 34308
rect -2068 34252 -2012 34308
rect -1748 34252 -1692 34308
rect -1428 34252 -1372 34308
rect -1108 34252 -1052 34308
rect -31028 34172 -30972 34228
rect -30708 34172 -30652 34228
rect -30388 34172 -30332 34228
rect -30068 34172 -30012 34228
rect -3348 34092 -3292 34148
rect -3028 34092 -2972 34148
rect -2708 34092 -2652 34148
rect -2388 34092 -2332 34148
rect -2068 34092 -2012 34148
rect -1748 34092 -1692 34148
rect -1428 34092 -1372 34148
rect -1108 34092 -1052 34148
rect -31028 34012 -30972 34068
rect -30708 34012 -30652 34068
rect -30388 34012 -30332 34068
rect -30068 34012 -30012 34068
rect -3348 33932 -3292 33988
rect -3028 33932 -2972 33988
rect -2708 33932 -2652 33988
rect -2388 33932 -2332 33988
rect -2068 33932 -2012 33988
rect -1748 33932 -1692 33988
rect -1428 33932 -1372 33988
rect -1108 33932 -1052 33988
rect -31028 33852 -30972 33908
rect -30708 33852 -30652 33908
rect -30388 33852 -30332 33908
rect -30068 33852 -30012 33908
rect -3348 33772 -3292 33828
rect -3028 33772 -2972 33828
rect -2708 33772 -2652 33828
rect -2388 33772 -2332 33828
rect -2068 33772 -2012 33828
rect -1748 33772 -1692 33828
rect -1428 33772 -1372 33828
rect -1108 33772 -1052 33828
rect -31028 33692 -30972 33748
rect -30708 33692 -30652 33748
rect -30388 33692 -30332 33748
rect -30068 33692 -30012 33748
rect -3348 33612 -3292 33668
rect -3028 33612 -2972 33668
rect -2708 33612 -2652 33668
rect -2388 33612 -2332 33668
rect -2068 33612 -2012 33668
rect -1748 33612 -1692 33668
rect -1428 33612 -1372 33668
rect -1108 33612 -1052 33668
rect -31028 33532 -30972 33588
rect -30708 33532 -30652 33588
rect -30388 33532 -30332 33588
rect -30068 33532 -30012 33588
rect -3348 33452 -3292 33508
rect -3028 33452 -2972 33508
rect -2708 33452 -2652 33508
rect -2388 33452 -2332 33508
rect -2068 33452 -2012 33508
rect -1748 33452 -1692 33508
rect -1428 33452 -1372 33508
rect -1108 33452 -1052 33508
rect -31028 33372 -30972 33428
rect -30708 33372 -30652 33428
rect -30388 33372 -30332 33428
rect -30068 33372 -30012 33428
rect -31028 33212 -30972 33268
rect -30708 33212 -30652 33268
rect -30388 33212 -30332 33268
rect -30068 33212 -30012 33268
rect -3348 33212 -3292 33268
rect -3028 33212 -2972 33268
rect -2708 33212 -2652 33268
rect -2388 33212 -2332 33268
rect -2068 33212 -2012 33268
rect -1748 33212 -1692 33268
rect -1428 33212 -1372 33268
rect -1108 33212 -1052 33268
rect -31028 33052 -30972 33108
rect -30708 33052 -30652 33108
rect -30388 33052 -30332 33108
rect -30068 33052 -30012 33108
rect -3348 33052 -3292 33108
rect -3028 33052 -2972 33108
rect -2708 33052 -2652 33108
rect -2388 33052 -2332 33108
rect -2068 33052 -2012 33108
rect -1748 33052 -1692 33108
rect -1428 33052 -1372 33108
rect -1108 33052 -1052 33108
rect -31028 32892 -30972 32948
rect -30708 32892 -30652 32948
rect -30388 32892 -30332 32948
rect -30068 32892 -30012 32948
rect -29908 32946 -29852 32948
rect -29908 32894 -29906 32946
rect -29906 32894 -29854 32946
rect -29854 32894 -29852 32946
rect -29908 32892 -29852 32894
rect -29748 32946 -29692 32948
rect -29748 32894 -29746 32946
rect -29746 32894 -29694 32946
rect -29694 32894 -29692 32946
rect -29748 32892 -29692 32894
rect -29588 32946 -29532 32948
rect -29588 32894 -29586 32946
rect -29586 32894 -29534 32946
rect -29534 32894 -29532 32946
rect -29588 32892 -29532 32894
rect -29428 32946 -29372 32948
rect -29428 32894 -29426 32946
rect -29426 32894 -29374 32946
rect -29374 32894 -29372 32946
rect -29428 32892 -29372 32894
rect -29268 32946 -29212 32948
rect -29268 32894 -29266 32946
rect -29266 32894 -29214 32946
rect -29214 32894 -29212 32946
rect -29268 32892 -29212 32894
rect -29108 32946 -29052 32948
rect -29108 32894 -29106 32946
rect -29106 32894 -29054 32946
rect -29054 32894 -29052 32946
rect -29108 32892 -29052 32894
rect -28948 32946 -28892 32948
rect -28948 32894 -28946 32946
rect -28946 32894 -28894 32946
rect -28894 32894 -28892 32946
rect -28948 32892 -28892 32894
rect -28788 32946 -28732 32948
rect -28788 32894 -28786 32946
rect -28786 32894 -28734 32946
rect -28734 32894 -28732 32946
rect -28788 32892 -28732 32894
rect -28628 32946 -28572 32948
rect -28628 32894 -28626 32946
rect -28626 32894 -28574 32946
rect -28574 32894 -28572 32946
rect -28628 32892 -28572 32894
rect -28468 32946 -28412 32948
rect -28468 32894 -28466 32946
rect -28466 32894 -28414 32946
rect -28414 32894 -28412 32946
rect -28468 32892 -28412 32894
rect -28308 32946 -28252 32948
rect -28308 32894 -28306 32946
rect -28306 32894 -28254 32946
rect -28254 32894 -28252 32946
rect -28308 32892 -28252 32894
rect -28148 32946 -28092 32948
rect -28148 32894 -28146 32946
rect -28146 32894 -28094 32946
rect -28094 32894 -28092 32946
rect -28148 32892 -28092 32894
rect -27988 32946 -27932 32948
rect -27988 32894 -27986 32946
rect -27986 32894 -27934 32946
rect -27934 32894 -27932 32946
rect -27988 32892 -27932 32894
rect -27828 32946 -27772 32948
rect -27828 32894 -27826 32946
rect -27826 32894 -27774 32946
rect -27774 32894 -27772 32946
rect -27828 32892 -27772 32894
rect -27668 32946 -27612 32948
rect -27668 32894 -27666 32946
rect -27666 32894 -27614 32946
rect -27614 32894 -27612 32946
rect -27668 32892 -27612 32894
rect -27508 32946 -27452 32948
rect -27508 32894 -27506 32946
rect -27506 32894 -27454 32946
rect -27454 32894 -27452 32946
rect -27508 32892 -27452 32894
rect -27348 32946 -27292 32948
rect -27348 32894 -27346 32946
rect -27346 32894 -27294 32946
rect -27294 32894 -27292 32946
rect -27348 32892 -27292 32894
rect -27188 32946 -27132 32948
rect -27188 32894 -27186 32946
rect -27186 32894 -27134 32946
rect -27134 32894 -27132 32946
rect -27188 32892 -27132 32894
rect -27028 32946 -26972 32948
rect -27028 32894 -27026 32946
rect -27026 32894 -26974 32946
rect -26974 32894 -26972 32946
rect -27028 32892 -26972 32894
rect -26868 32946 -26812 32948
rect -26868 32894 -26866 32946
rect -26866 32894 -26814 32946
rect -26814 32894 -26812 32946
rect -26868 32892 -26812 32894
rect -26708 32946 -26652 32948
rect -26708 32894 -26706 32946
rect -26706 32894 -26654 32946
rect -26654 32894 -26652 32946
rect -26708 32892 -26652 32894
rect -26548 32946 -26492 32948
rect -26548 32894 -26546 32946
rect -26546 32894 -26494 32946
rect -26494 32894 -26492 32946
rect -26548 32892 -26492 32894
rect -26388 32946 -26332 32948
rect -26388 32894 -26386 32946
rect -26386 32894 -26334 32946
rect -26334 32894 -26332 32946
rect -26388 32892 -26332 32894
rect -26228 32946 -26172 32948
rect -26228 32894 -26226 32946
rect -26226 32894 -26174 32946
rect -26174 32894 -26172 32946
rect -26228 32892 -26172 32894
rect -26068 32946 -26012 32948
rect -26068 32894 -26066 32946
rect -26066 32894 -26014 32946
rect -26014 32894 -26012 32946
rect -26068 32892 -26012 32894
rect -25908 32946 -25852 32948
rect -25908 32894 -25906 32946
rect -25906 32894 -25854 32946
rect -25854 32894 -25852 32946
rect -25908 32892 -25852 32894
rect -25748 32946 -25692 32948
rect -25748 32894 -25746 32946
rect -25746 32894 -25694 32946
rect -25694 32894 -25692 32946
rect -25748 32892 -25692 32894
rect -25588 32946 -25532 32948
rect -25588 32894 -25586 32946
rect -25586 32894 -25534 32946
rect -25534 32894 -25532 32946
rect -25588 32892 -25532 32894
rect -25428 32946 -25372 32948
rect -25428 32894 -25426 32946
rect -25426 32894 -25374 32946
rect -25374 32894 -25372 32946
rect -25428 32892 -25372 32894
rect -25268 32946 -25212 32948
rect -25268 32894 -25266 32946
rect -25266 32894 -25214 32946
rect -25214 32894 -25212 32946
rect -25268 32892 -25212 32894
rect -25108 32946 -25052 32948
rect -25108 32894 -25106 32946
rect -25106 32894 -25054 32946
rect -25054 32894 -25052 32946
rect -25108 32892 -25052 32894
rect -24948 32946 -24892 32948
rect -24948 32894 -24946 32946
rect -24946 32894 -24894 32946
rect -24894 32894 -24892 32946
rect -24948 32892 -24892 32894
rect -24788 32946 -24732 32948
rect -24788 32894 -24786 32946
rect -24786 32894 -24734 32946
rect -24734 32894 -24732 32946
rect -24788 32892 -24732 32894
rect -24628 32946 -24572 32948
rect -24628 32894 -24626 32946
rect -24626 32894 -24574 32946
rect -24574 32894 -24572 32946
rect -24628 32892 -24572 32894
rect -24468 32946 -24412 32948
rect -24468 32894 -24466 32946
rect -24466 32894 -24414 32946
rect -24414 32894 -24412 32946
rect -24468 32892 -24412 32894
rect -24308 32946 -24252 32948
rect -24308 32894 -24306 32946
rect -24306 32894 -24254 32946
rect -24254 32894 -24252 32946
rect -24308 32892 -24252 32894
rect -24148 32946 -24092 32948
rect -24148 32894 -24146 32946
rect -24146 32894 -24094 32946
rect -24094 32894 -24092 32946
rect -24148 32892 -24092 32894
rect -23988 32946 -23932 32948
rect -23988 32894 -23986 32946
rect -23986 32894 -23934 32946
rect -23934 32894 -23932 32946
rect -23988 32892 -23932 32894
rect -23828 32946 -23772 32948
rect -23828 32894 -23826 32946
rect -23826 32894 -23774 32946
rect -23774 32894 -23772 32946
rect -23828 32892 -23772 32894
rect -23668 32946 -23612 32948
rect -23668 32894 -23666 32946
rect -23666 32894 -23614 32946
rect -23614 32894 -23612 32946
rect -23668 32892 -23612 32894
rect -23508 32946 -23452 32948
rect -23508 32894 -23506 32946
rect -23506 32894 -23454 32946
rect -23454 32894 -23452 32946
rect -23508 32892 -23452 32894
rect -23348 32946 -23292 32948
rect -23348 32894 -23346 32946
rect -23346 32894 -23294 32946
rect -23294 32894 -23292 32946
rect -23348 32892 -23292 32894
rect -23188 32946 -23132 32948
rect -23188 32894 -23186 32946
rect -23186 32894 -23134 32946
rect -23134 32894 -23132 32946
rect -23188 32892 -23132 32894
rect -23028 32946 -22972 32948
rect -23028 32894 -23026 32946
rect -23026 32894 -22974 32946
rect -22974 32894 -22972 32946
rect -23028 32892 -22972 32894
rect -22868 32946 -22812 32948
rect -22868 32894 -22866 32946
rect -22866 32894 -22814 32946
rect -22814 32894 -22812 32946
rect -22868 32892 -22812 32894
rect -22708 32946 -22652 32948
rect -22708 32894 -22706 32946
rect -22706 32894 -22654 32946
rect -22654 32894 -22652 32946
rect -22708 32892 -22652 32894
rect -22548 32946 -22492 32948
rect -22548 32894 -22546 32946
rect -22546 32894 -22494 32946
rect -22494 32894 -22492 32946
rect -22548 32892 -22492 32894
rect -22388 32946 -22332 32948
rect -22388 32894 -22386 32946
rect -22386 32894 -22334 32946
rect -22334 32894 -22332 32946
rect -22388 32892 -22332 32894
rect -22228 32946 -22172 32948
rect -22228 32894 -22226 32946
rect -22226 32894 -22174 32946
rect -22174 32894 -22172 32946
rect -22228 32892 -22172 32894
rect -22068 32946 -22012 32948
rect -22068 32894 -22066 32946
rect -22066 32894 -22014 32946
rect -22014 32894 -22012 32946
rect -22068 32892 -22012 32894
rect -21908 32946 -21852 32948
rect -21908 32894 -21906 32946
rect -21906 32894 -21854 32946
rect -21854 32894 -21852 32946
rect -21908 32892 -21852 32894
rect -21748 32946 -21692 32948
rect -21748 32894 -21746 32946
rect -21746 32894 -21694 32946
rect -21694 32894 -21692 32946
rect -21748 32892 -21692 32894
rect -21588 32946 -21532 32948
rect -21588 32894 -21586 32946
rect -21586 32894 -21534 32946
rect -21534 32894 -21532 32946
rect -21588 32892 -21532 32894
rect -21428 32946 -21372 32948
rect -21428 32894 -21426 32946
rect -21426 32894 -21374 32946
rect -21374 32894 -21372 32946
rect -21428 32892 -21372 32894
rect -21268 32946 -21212 32948
rect -21268 32894 -21266 32946
rect -21266 32894 -21214 32946
rect -21214 32894 -21212 32946
rect -21268 32892 -21212 32894
rect -21108 32946 -21052 32948
rect -21108 32894 -21106 32946
rect -21106 32894 -21054 32946
rect -21054 32894 -21052 32946
rect -21108 32892 -21052 32894
rect -20948 32946 -20892 32948
rect -20948 32894 -20946 32946
rect -20946 32894 -20894 32946
rect -20894 32894 -20892 32946
rect -20948 32892 -20892 32894
rect -20788 32946 -20732 32948
rect -20788 32894 -20786 32946
rect -20786 32894 -20734 32946
rect -20734 32894 -20732 32946
rect -20788 32892 -20732 32894
rect -20628 32946 -20572 32948
rect -20628 32894 -20626 32946
rect -20626 32894 -20574 32946
rect -20574 32894 -20572 32946
rect -20628 32892 -20572 32894
rect -20468 32946 -20412 32948
rect -20468 32894 -20466 32946
rect -20466 32894 -20414 32946
rect -20414 32894 -20412 32946
rect -20468 32892 -20412 32894
rect -20308 32946 -20252 32948
rect -20308 32894 -20306 32946
rect -20306 32894 -20254 32946
rect -20254 32894 -20252 32946
rect -20308 32892 -20252 32894
rect -20148 32946 -20092 32948
rect -20148 32894 -20146 32946
rect -20146 32894 -20094 32946
rect -20094 32894 -20092 32946
rect -20148 32892 -20092 32894
rect -19988 32946 -19932 32948
rect -19988 32894 -19986 32946
rect -19986 32894 -19934 32946
rect -19934 32894 -19932 32946
rect -19988 32892 -19932 32894
rect -19828 32946 -19772 32948
rect -19828 32894 -19826 32946
rect -19826 32894 -19774 32946
rect -19774 32894 -19772 32946
rect -19828 32892 -19772 32894
rect -19668 32946 -19612 32948
rect -19668 32894 -19666 32946
rect -19666 32894 -19614 32946
rect -19614 32894 -19612 32946
rect -19668 32892 -19612 32894
rect -19508 32946 -19452 32948
rect -19508 32894 -19506 32946
rect -19506 32894 -19454 32946
rect -19454 32894 -19452 32946
rect -19508 32892 -19452 32894
rect -19348 32946 -19292 32948
rect -19348 32894 -19346 32946
rect -19346 32894 -19294 32946
rect -19294 32894 -19292 32946
rect -19348 32892 -19292 32894
rect -19188 32946 -19132 32948
rect -19188 32894 -19186 32946
rect -19186 32894 -19134 32946
rect -19134 32894 -19132 32946
rect -19188 32892 -19132 32894
rect -19028 32946 -18972 32948
rect -19028 32894 -19026 32946
rect -19026 32894 -18974 32946
rect -18974 32894 -18972 32946
rect -19028 32892 -18972 32894
rect -18868 32946 -18812 32948
rect -18868 32894 -18866 32946
rect -18866 32894 -18814 32946
rect -18814 32894 -18812 32946
rect -18868 32892 -18812 32894
rect -18708 32946 -18652 32948
rect -18708 32894 -18706 32946
rect -18706 32894 -18654 32946
rect -18654 32894 -18652 32946
rect -18708 32892 -18652 32894
rect -18548 32946 -18492 32948
rect -18548 32894 -18546 32946
rect -18546 32894 -18494 32946
rect -18494 32894 -18492 32946
rect -18548 32892 -18492 32894
rect -18388 32946 -18332 32948
rect -18388 32894 -18386 32946
rect -18386 32894 -18334 32946
rect -18334 32894 -18332 32946
rect -18388 32892 -18332 32894
rect -18228 32946 -18172 32948
rect -18228 32894 -18226 32946
rect -18226 32894 -18174 32946
rect -18174 32894 -18172 32946
rect -18228 32892 -18172 32894
rect -18068 32946 -18012 32948
rect -18068 32894 -18066 32946
rect -18066 32894 -18014 32946
rect -18014 32894 -18012 32946
rect -18068 32892 -18012 32894
rect -17908 32946 -17852 32948
rect -17908 32894 -17906 32946
rect -17906 32894 -17854 32946
rect -17854 32894 -17852 32946
rect -17908 32892 -17852 32894
rect -17748 32946 -17692 32948
rect -17748 32894 -17746 32946
rect -17746 32894 -17694 32946
rect -17694 32894 -17692 32946
rect -17748 32892 -17692 32894
rect -17588 32946 -17532 32948
rect -17588 32894 -17586 32946
rect -17586 32894 -17534 32946
rect -17534 32894 -17532 32946
rect -17588 32892 -17532 32894
rect -17428 32946 -17372 32948
rect -17428 32894 -17426 32946
rect -17426 32894 -17374 32946
rect -17374 32894 -17372 32946
rect -17428 32892 -17372 32894
rect -17268 32946 -17212 32948
rect -17268 32894 -17266 32946
rect -17266 32894 -17214 32946
rect -17214 32894 -17212 32946
rect -17268 32892 -17212 32894
rect -17108 32946 -17052 32948
rect -17108 32894 -17106 32946
rect -17106 32894 -17054 32946
rect -17054 32894 -17052 32946
rect -17108 32892 -17052 32894
rect -16948 32946 -16892 32948
rect -16948 32894 -16946 32946
rect -16946 32894 -16894 32946
rect -16894 32894 -16892 32946
rect -16948 32892 -16892 32894
rect -16788 32946 -16732 32948
rect -16788 32894 -16786 32946
rect -16786 32894 -16734 32946
rect -16734 32894 -16732 32946
rect -16788 32892 -16732 32894
rect -16628 32946 -16572 32948
rect -16628 32894 -16626 32946
rect -16626 32894 -16574 32946
rect -16574 32894 -16572 32946
rect -16628 32892 -16572 32894
rect -16468 32946 -16412 32948
rect -16468 32894 -16466 32946
rect -16466 32894 -16414 32946
rect -16414 32894 -16412 32946
rect -16468 32892 -16412 32894
rect -16308 32946 -16252 32948
rect -16308 32894 -16306 32946
rect -16306 32894 -16254 32946
rect -16254 32894 -16252 32946
rect -16308 32892 -16252 32894
rect -16148 32946 -16092 32948
rect -16148 32894 -16146 32946
rect -16146 32894 -16094 32946
rect -16094 32894 -16092 32946
rect -16148 32892 -16092 32894
rect -15988 32946 -15932 32948
rect -15988 32894 -15986 32946
rect -15986 32894 -15934 32946
rect -15934 32894 -15932 32946
rect -15988 32892 -15932 32894
rect -15828 32946 -15772 32948
rect -15828 32894 -15826 32946
rect -15826 32894 -15774 32946
rect -15774 32894 -15772 32946
rect -15828 32892 -15772 32894
rect -15668 32946 -15612 32948
rect -15668 32894 -15666 32946
rect -15666 32894 -15614 32946
rect -15614 32894 -15612 32946
rect -15668 32892 -15612 32894
rect -15508 32946 -15452 32948
rect -15508 32894 -15506 32946
rect -15506 32894 -15454 32946
rect -15454 32894 -15452 32946
rect -15508 32892 -15452 32894
rect -15348 32946 -15292 32948
rect -15348 32894 -15346 32946
rect -15346 32894 -15294 32946
rect -15294 32894 -15292 32946
rect -15348 32892 -15292 32894
rect -15188 32946 -15132 32948
rect -15188 32894 -15186 32946
rect -15186 32894 -15134 32946
rect -15134 32894 -15132 32946
rect -15188 32892 -15132 32894
rect -15028 32946 -14972 32948
rect -15028 32894 -15026 32946
rect -15026 32894 -14974 32946
rect -14974 32894 -14972 32946
rect -15028 32892 -14972 32894
rect -14868 32946 -14812 32948
rect -14868 32894 -14866 32946
rect -14866 32894 -14814 32946
rect -14814 32894 -14812 32946
rect -14868 32892 -14812 32894
rect -14708 32946 -14652 32948
rect -14708 32894 -14706 32946
rect -14706 32894 -14654 32946
rect -14654 32894 -14652 32946
rect -14708 32892 -14652 32894
rect -14548 32946 -14492 32948
rect -14548 32894 -14546 32946
rect -14546 32894 -14494 32946
rect -14494 32894 -14492 32946
rect -14548 32892 -14492 32894
rect -14388 32946 -14332 32948
rect -14388 32894 -14386 32946
rect -14386 32894 -14334 32946
rect -14334 32894 -14332 32946
rect -14388 32892 -14332 32894
rect -14228 32946 -14172 32948
rect -14228 32894 -14226 32946
rect -14226 32894 -14174 32946
rect -14174 32894 -14172 32946
rect -14228 32892 -14172 32894
rect -14068 32946 -14012 32948
rect -14068 32894 -14066 32946
rect -14066 32894 -14014 32946
rect -14014 32894 -14012 32946
rect -14068 32892 -14012 32894
rect -13908 32946 -13852 32948
rect -13908 32894 -13906 32946
rect -13906 32894 -13854 32946
rect -13854 32894 -13852 32946
rect -13908 32892 -13852 32894
rect -13748 32946 -13692 32948
rect -13748 32894 -13746 32946
rect -13746 32894 -13694 32946
rect -13694 32894 -13692 32946
rect -13748 32892 -13692 32894
rect -13588 32946 -13532 32948
rect -13588 32894 -13586 32946
rect -13586 32894 -13534 32946
rect -13534 32894 -13532 32946
rect -13588 32892 -13532 32894
rect -13428 32946 -13372 32948
rect -13428 32894 -13426 32946
rect -13426 32894 -13374 32946
rect -13374 32894 -13372 32946
rect -13428 32892 -13372 32894
rect -13268 32946 -13212 32948
rect -13268 32894 -13266 32946
rect -13266 32894 -13214 32946
rect -13214 32894 -13212 32946
rect -13268 32892 -13212 32894
rect -13108 32946 -13052 32948
rect -13108 32894 -13106 32946
rect -13106 32894 -13054 32946
rect -13054 32894 -13052 32946
rect -13108 32892 -13052 32894
rect -12948 32946 -12892 32948
rect -12948 32894 -12946 32946
rect -12946 32894 -12894 32946
rect -12894 32894 -12892 32946
rect -12948 32892 -12892 32894
rect -12788 32946 -12732 32948
rect -12788 32894 -12786 32946
rect -12786 32894 -12734 32946
rect -12734 32894 -12732 32946
rect -12788 32892 -12732 32894
rect -12628 32946 -12572 32948
rect -12628 32894 -12626 32946
rect -12626 32894 -12574 32946
rect -12574 32894 -12572 32946
rect -12628 32892 -12572 32894
rect -12468 32946 -12412 32948
rect -12468 32894 -12466 32946
rect -12466 32894 -12414 32946
rect -12414 32894 -12412 32946
rect -12468 32892 -12412 32894
rect -12308 32946 -12252 32948
rect -12308 32894 -12306 32946
rect -12306 32894 -12254 32946
rect -12254 32894 -12252 32946
rect -12308 32892 -12252 32894
rect -12148 32946 -12092 32948
rect -12148 32894 -12146 32946
rect -12146 32894 -12094 32946
rect -12094 32894 -12092 32946
rect -12148 32892 -12092 32894
rect -11988 32946 -11932 32948
rect -11988 32894 -11986 32946
rect -11986 32894 -11934 32946
rect -11934 32894 -11932 32946
rect -11988 32892 -11932 32894
rect -11828 32946 -11772 32948
rect -11828 32894 -11826 32946
rect -11826 32894 -11774 32946
rect -11774 32894 -11772 32946
rect -11828 32892 -11772 32894
rect -11668 32946 -11612 32948
rect -11668 32894 -11666 32946
rect -11666 32894 -11614 32946
rect -11614 32894 -11612 32946
rect -11668 32892 -11612 32894
rect -11508 32946 -11452 32948
rect -11508 32894 -11506 32946
rect -11506 32894 -11454 32946
rect -11454 32894 -11452 32946
rect -11508 32892 -11452 32894
rect -11188 32946 -11132 32948
rect -11188 32894 -11186 32946
rect -11186 32894 -11134 32946
rect -11134 32894 -11132 32946
rect -11188 32892 -11132 32894
rect -10868 32946 -10812 32948
rect -10868 32894 -10866 32946
rect -10866 32894 -10814 32946
rect -10814 32894 -10812 32946
rect -10868 32892 -10812 32894
rect -10708 32946 -10652 32948
rect -10708 32894 -10706 32946
rect -10706 32894 -10654 32946
rect -10654 32894 -10652 32946
rect -10708 32892 -10652 32894
rect -10548 32946 -10492 32948
rect -10548 32894 -10546 32946
rect -10546 32894 -10494 32946
rect -10494 32894 -10492 32946
rect -10548 32892 -10492 32894
rect -10388 32946 -10332 32948
rect -10388 32894 -10386 32946
rect -10386 32894 -10334 32946
rect -10334 32894 -10332 32946
rect -10388 32892 -10332 32894
rect -10228 32946 -10172 32948
rect -10228 32894 -10226 32946
rect -10226 32894 -10174 32946
rect -10174 32894 -10172 32946
rect -10228 32892 -10172 32894
rect -10068 32946 -10012 32948
rect -10068 32894 -10066 32946
rect -10066 32894 -10014 32946
rect -10014 32894 -10012 32946
rect -10068 32892 -10012 32894
rect -9908 32946 -9852 32948
rect -9908 32894 -9906 32946
rect -9906 32894 -9854 32946
rect -9854 32894 -9852 32946
rect -9908 32892 -9852 32894
rect -9748 32946 -9692 32948
rect -9748 32894 -9746 32946
rect -9746 32894 -9694 32946
rect -9694 32894 -9692 32946
rect -9748 32892 -9692 32894
rect -9588 32946 -9532 32948
rect -9588 32894 -9586 32946
rect -9586 32894 -9534 32946
rect -9534 32894 -9532 32946
rect -9588 32892 -9532 32894
rect -9428 32946 -9372 32948
rect -9428 32894 -9426 32946
rect -9426 32894 -9374 32946
rect -9374 32894 -9372 32946
rect -9428 32892 -9372 32894
rect -9268 32946 -9212 32948
rect -9268 32894 -9266 32946
rect -9266 32894 -9214 32946
rect -9214 32894 -9212 32946
rect -9268 32892 -9212 32894
rect -9108 32946 -9052 32948
rect -9108 32894 -9106 32946
rect -9106 32894 -9054 32946
rect -9054 32894 -9052 32946
rect -9108 32892 -9052 32894
rect -8948 32946 -8892 32948
rect -8948 32894 -8946 32946
rect -8946 32894 -8894 32946
rect -8894 32894 -8892 32946
rect -8948 32892 -8892 32894
rect -8788 32946 -8732 32948
rect -8788 32894 -8786 32946
rect -8786 32894 -8734 32946
rect -8734 32894 -8732 32946
rect -8788 32892 -8732 32894
rect -8628 32946 -8572 32948
rect -8628 32894 -8626 32946
rect -8626 32894 -8574 32946
rect -8574 32894 -8572 32946
rect -8628 32892 -8572 32894
rect -8468 32946 -8412 32948
rect -8468 32894 -8466 32946
rect -8466 32894 -8414 32946
rect -8414 32894 -8412 32946
rect -8468 32892 -8412 32894
rect -8308 32946 -8252 32948
rect -8308 32894 -8306 32946
rect -8306 32894 -8254 32946
rect -8254 32894 -8252 32946
rect -8308 32892 -8252 32894
rect -8148 32946 -8092 32948
rect -8148 32894 -8146 32946
rect -8146 32894 -8094 32946
rect -8094 32894 -8092 32946
rect -8148 32892 -8092 32894
rect -7988 32946 -7932 32948
rect -7988 32894 -7986 32946
rect -7986 32894 -7934 32946
rect -7934 32894 -7932 32946
rect -7988 32892 -7932 32894
rect -7828 32946 -7772 32948
rect -7828 32894 -7826 32946
rect -7826 32894 -7774 32946
rect -7774 32894 -7772 32946
rect -7828 32892 -7772 32894
rect -7668 32946 -7612 32948
rect -7668 32894 -7666 32946
rect -7666 32894 -7614 32946
rect -7614 32894 -7612 32946
rect -7668 32892 -7612 32894
rect -7508 32946 -7452 32948
rect -7508 32894 -7506 32946
rect -7506 32894 -7454 32946
rect -7454 32894 -7452 32946
rect -7508 32892 -7452 32894
rect -7348 32946 -7292 32948
rect -7348 32894 -7346 32946
rect -7346 32894 -7294 32946
rect -7294 32894 -7292 32946
rect -7348 32892 -7292 32894
rect -7188 32946 -7132 32948
rect -7188 32894 -7186 32946
rect -7186 32894 -7134 32946
rect -7134 32894 -7132 32946
rect -7188 32892 -7132 32894
rect -7028 32946 -6972 32948
rect -7028 32894 -7026 32946
rect -7026 32894 -6974 32946
rect -6974 32894 -6972 32946
rect -7028 32892 -6972 32894
rect -6868 32946 -6812 32948
rect -6868 32894 -6866 32946
rect -6866 32894 -6814 32946
rect -6814 32894 -6812 32946
rect -6868 32892 -6812 32894
rect -6708 32946 -6652 32948
rect -6708 32894 -6706 32946
rect -6706 32894 -6654 32946
rect -6654 32894 -6652 32946
rect -6708 32892 -6652 32894
rect -6548 32946 -6492 32948
rect -6548 32894 -6546 32946
rect -6546 32894 -6494 32946
rect -6494 32894 -6492 32946
rect -6548 32892 -6492 32894
rect -6388 32946 -6332 32948
rect -6388 32894 -6386 32946
rect -6386 32894 -6334 32946
rect -6334 32894 -6332 32946
rect -6388 32892 -6332 32894
rect -6228 32946 -6172 32948
rect -6228 32894 -6226 32946
rect -6226 32894 -6174 32946
rect -6174 32894 -6172 32946
rect -6228 32892 -6172 32894
rect -6068 32946 -6012 32948
rect -6068 32894 -6066 32946
rect -6066 32894 -6014 32946
rect -6014 32894 -6012 32946
rect -6068 32892 -6012 32894
rect -5908 32946 -5852 32948
rect -5908 32894 -5906 32946
rect -5906 32894 -5854 32946
rect -5854 32894 -5852 32946
rect -5908 32892 -5852 32894
rect -5748 32946 -5692 32948
rect -5748 32894 -5746 32946
rect -5746 32894 -5694 32946
rect -5694 32894 -5692 32946
rect -5748 32892 -5692 32894
rect -5588 32946 -5532 32948
rect -5588 32894 -5586 32946
rect -5586 32894 -5534 32946
rect -5534 32894 -5532 32946
rect -5588 32892 -5532 32894
rect -5428 32946 -5372 32948
rect -5428 32894 -5426 32946
rect -5426 32894 -5374 32946
rect -5374 32894 -5372 32946
rect -5428 32892 -5372 32894
rect -5268 32946 -5212 32948
rect -5268 32894 -5266 32946
rect -5266 32894 -5214 32946
rect -5214 32894 -5212 32946
rect -5268 32892 -5212 32894
rect -5108 32946 -5052 32948
rect -5108 32894 -5106 32946
rect -5106 32894 -5054 32946
rect -5054 32894 -5052 32946
rect -5108 32892 -5052 32894
rect -4948 32946 -4892 32948
rect -4948 32894 -4946 32946
rect -4946 32894 -4894 32946
rect -4894 32894 -4892 32946
rect -4948 32892 -4892 32894
rect -4788 32946 -4732 32948
rect -4788 32894 -4786 32946
rect -4786 32894 -4734 32946
rect -4734 32894 -4732 32946
rect -4788 32892 -4732 32894
rect -4628 32946 -4572 32948
rect -4628 32894 -4626 32946
rect -4626 32894 -4574 32946
rect -4574 32894 -4572 32946
rect -4628 32892 -4572 32894
rect -4468 32946 -4412 32948
rect -4468 32894 -4466 32946
rect -4466 32894 -4414 32946
rect -4414 32894 -4412 32946
rect -4468 32892 -4412 32894
rect -4308 32946 -4252 32948
rect -4308 32894 -4306 32946
rect -4306 32894 -4254 32946
rect -4254 32894 -4252 32946
rect -4308 32892 -4252 32894
rect -4148 32946 -4092 32948
rect -4148 32894 -4146 32946
rect -4146 32894 -4094 32946
rect -4094 32894 -4092 32946
rect -4148 32892 -4092 32894
rect -3988 32946 -3932 32948
rect -3988 32894 -3986 32946
rect -3986 32894 -3934 32946
rect -3934 32894 -3932 32946
rect -3988 32892 -3932 32894
rect -3668 32946 -3612 32948
rect -3668 32894 -3666 32946
rect -3666 32894 -3614 32946
rect -3614 32894 -3612 32946
rect -3668 32892 -3612 32894
rect -3508 32946 -3452 32948
rect -3508 32894 -3506 32946
rect -3506 32894 -3454 32946
rect -3454 32894 -3452 32946
rect -3508 32892 -3452 32894
rect -3348 32946 -3292 32948
rect -3348 32894 -3346 32946
rect -3346 32894 -3294 32946
rect -3294 32894 -3292 32946
rect -3348 32892 -3292 32894
rect -3188 32946 -3132 32948
rect -3188 32894 -3186 32946
rect -3186 32894 -3134 32946
rect -3134 32894 -3132 32946
rect -3188 32892 -3132 32894
rect -3028 32946 -2972 32948
rect -3028 32894 -3026 32946
rect -3026 32894 -2974 32946
rect -2974 32894 -2972 32946
rect -3028 32892 -2972 32894
rect -2868 32946 -2812 32948
rect -2868 32894 -2866 32946
rect -2866 32894 -2814 32946
rect -2814 32894 -2812 32946
rect -2868 32892 -2812 32894
rect -2708 32946 -2652 32948
rect -2708 32894 -2706 32946
rect -2706 32894 -2654 32946
rect -2654 32894 -2652 32946
rect -2708 32892 -2652 32894
rect -2388 32946 -2332 32948
rect -2388 32894 -2386 32946
rect -2386 32894 -2334 32946
rect -2334 32894 -2332 32946
rect -2388 32892 -2332 32894
rect -2068 32946 -2012 32948
rect -2068 32894 -2066 32946
rect -2066 32894 -2014 32946
rect -2014 32894 -2012 32946
rect -2068 32892 -2012 32894
rect -1748 32946 -1692 32948
rect -1748 32894 -1746 32946
rect -1746 32894 -1694 32946
rect -1694 32894 -1692 32946
rect -1748 32892 -1692 32894
rect -1428 32946 -1372 32948
rect -1428 32894 -1426 32946
rect -1426 32894 -1374 32946
rect -1374 32894 -1372 32946
rect -1428 32892 -1372 32894
rect -1108 32946 -1052 32948
rect -1108 32894 -1106 32946
rect -1106 32894 -1054 32946
rect -1054 32894 -1052 32946
rect -1108 32892 -1052 32894
rect -31028 32732 -30972 32788
rect -30708 32732 -30652 32788
rect -30548 32732 -30492 32788
rect -1268 32732 -1212 32788
rect -31028 32572 -30972 32628
rect -30708 32572 -30652 32628
rect -30388 32572 -30332 32628
rect -30068 32572 -30012 32628
rect -29908 32626 -29852 32628
rect -29908 32574 -29906 32626
rect -29906 32574 -29854 32626
rect -29854 32574 -29852 32626
rect -29908 32572 -29852 32574
rect -29748 32626 -29692 32628
rect -29748 32574 -29746 32626
rect -29746 32574 -29694 32626
rect -29694 32574 -29692 32626
rect -29748 32572 -29692 32574
rect -29588 32626 -29532 32628
rect -29588 32574 -29586 32626
rect -29586 32574 -29534 32626
rect -29534 32574 -29532 32626
rect -29588 32572 -29532 32574
rect -29428 32626 -29372 32628
rect -29428 32574 -29426 32626
rect -29426 32574 -29374 32626
rect -29374 32574 -29372 32626
rect -29428 32572 -29372 32574
rect -29268 32626 -29212 32628
rect -29268 32574 -29266 32626
rect -29266 32574 -29214 32626
rect -29214 32574 -29212 32626
rect -29268 32572 -29212 32574
rect -29108 32626 -29052 32628
rect -29108 32574 -29106 32626
rect -29106 32574 -29054 32626
rect -29054 32574 -29052 32626
rect -29108 32572 -29052 32574
rect -28948 32626 -28892 32628
rect -28948 32574 -28946 32626
rect -28946 32574 -28894 32626
rect -28894 32574 -28892 32626
rect -28948 32572 -28892 32574
rect -28788 32626 -28732 32628
rect -28788 32574 -28786 32626
rect -28786 32574 -28734 32626
rect -28734 32574 -28732 32626
rect -28788 32572 -28732 32574
rect -28628 32626 -28572 32628
rect -28628 32574 -28626 32626
rect -28626 32574 -28574 32626
rect -28574 32574 -28572 32626
rect -28628 32572 -28572 32574
rect -28468 32626 -28412 32628
rect -28468 32574 -28466 32626
rect -28466 32574 -28414 32626
rect -28414 32574 -28412 32626
rect -28468 32572 -28412 32574
rect -28308 32626 -28252 32628
rect -28308 32574 -28306 32626
rect -28306 32574 -28254 32626
rect -28254 32574 -28252 32626
rect -28308 32572 -28252 32574
rect -28148 32626 -28092 32628
rect -28148 32574 -28146 32626
rect -28146 32574 -28094 32626
rect -28094 32574 -28092 32626
rect -28148 32572 -28092 32574
rect -27988 32626 -27932 32628
rect -27988 32574 -27986 32626
rect -27986 32574 -27934 32626
rect -27934 32574 -27932 32626
rect -27988 32572 -27932 32574
rect -27828 32626 -27772 32628
rect -27828 32574 -27826 32626
rect -27826 32574 -27774 32626
rect -27774 32574 -27772 32626
rect -27828 32572 -27772 32574
rect -27668 32626 -27612 32628
rect -27668 32574 -27666 32626
rect -27666 32574 -27614 32626
rect -27614 32574 -27612 32626
rect -27668 32572 -27612 32574
rect -27508 32626 -27452 32628
rect -27508 32574 -27506 32626
rect -27506 32574 -27454 32626
rect -27454 32574 -27452 32626
rect -27508 32572 -27452 32574
rect -27348 32626 -27292 32628
rect -27348 32574 -27346 32626
rect -27346 32574 -27294 32626
rect -27294 32574 -27292 32626
rect -27348 32572 -27292 32574
rect -27188 32626 -27132 32628
rect -27188 32574 -27186 32626
rect -27186 32574 -27134 32626
rect -27134 32574 -27132 32626
rect -27188 32572 -27132 32574
rect -27028 32626 -26972 32628
rect -27028 32574 -27026 32626
rect -27026 32574 -26974 32626
rect -26974 32574 -26972 32626
rect -27028 32572 -26972 32574
rect -26868 32626 -26812 32628
rect -26868 32574 -26866 32626
rect -26866 32574 -26814 32626
rect -26814 32574 -26812 32626
rect -26868 32572 -26812 32574
rect -26708 32626 -26652 32628
rect -26708 32574 -26706 32626
rect -26706 32574 -26654 32626
rect -26654 32574 -26652 32626
rect -26708 32572 -26652 32574
rect -26548 32626 -26492 32628
rect -26548 32574 -26546 32626
rect -26546 32574 -26494 32626
rect -26494 32574 -26492 32626
rect -26548 32572 -26492 32574
rect -26388 32626 -26332 32628
rect -26388 32574 -26386 32626
rect -26386 32574 -26334 32626
rect -26334 32574 -26332 32626
rect -26388 32572 -26332 32574
rect -26228 32626 -26172 32628
rect -26228 32574 -26226 32626
rect -26226 32574 -26174 32626
rect -26174 32574 -26172 32626
rect -26228 32572 -26172 32574
rect -26068 32626 -26012 32628
rect -26068 32574 -26066 32626
rect -26066 32574 -26014 32626
rect -26014 32574 -26012 32626
rect -26068 32572 -26012 32574
rect -25908 32626 -25852 32628
rect -25908 32574 -25906 32626
rect -25906 32574 -25854 32626
rect -25854 32574 -25852 32626
rect -25908 32572 -25852 32574
rect -25748 32626 -25692 32628
rect -25748 32574 -25746 32626
rect -25746 32574 -25694 32626
rect -25694 32574 -25692 32626
rect -25748 32572 -25692 32574
rect -25588 32626 -25532 32628
rect -25588 32574 -25586 32626
rect -25586 32574 -25534 32626
rect -25534 32574 -25532 32626
rect -25588 32572 -25532 32574
rect -25428 32626 -25372 32628
rect -25428 32574 -25426 32626
rect -25426 32574 -25374 32626
rect -25374 32574 -25372 32626
rect -25428 32572 -25372 32574
rect -25268 32626 -25212 32628
rect -25268 32574 -25266 32626
rect -25266 32574 -25214 32626
rect -25214 32574 -25212 32626
rect -25268 32572 -25212 32574
rect -25108 32626 -25052 32628
rect -25108 32574 -25106 32626
rect -25106 32574 -25054 32626
rect -25054 32574 -25052 32626
rect -25108 32572 -25052 32574
rect -24948 32626 -24892 32628
rect -24948 32574 -24946 32626
rect -24946 32574 -24894 32626
rect -24894 32574 -24892 32626
rect -24948 32572 -24892 32574
rect -24788 32626 -24732 32628
rect -24788 32574 -24786 32626
rect -24786 32574 -24734 32626
rect -24734 32574 -24732 32626
rect -24788 32572 -24732 32574
rect -24628 32626 -24572 32628
rect -24628 32574 -24626 32626
rect -24626 32574 -24574 32626
rect -24574 32574 -24572 32626
rect -24628 32572 -24572 32574
rect -24468 32626 -24412 32628
rect -24468 32574 -24466 32626
rect -24466 32574 -24414 32626
rect -24414 32574 -24412 32626
rect -24468 32572 -24412 32574
rect -24308 32626 -24252 32628
rect -24308 32574 -24306 32626
rect -24306 32574 -24254 32626
rect -24254 32574 -24252 32626
rect -24308 32572 -24252 32574
rect -24148 32626 -24092 32628
rect -24148 32574 -24146 32626
rect -24146 32574 -24094 32626
rect -24094 32574 -24092 32626
rect -24148 32572 -24092 32574
rect -23988 32626 -23932 32628
rect -23988 32574 -23986 32626
rect -23986 32574 -23934 32626
rect -23934 32574 -23932 32626
rect -23988 32572 -23932 32574
rect -23828 32626 -23772 32628
rect -23828 32574 -23826 32626
rect -23826 32574 -23774 32626
rect -23774 32574 -23772 32626
rect -23828 32572 -23772 32574
rect -23668 32626 -23612 32628
rect -23668 32574 -23666 32626
rect -23666 32574 -23614 32626
rect -23614 32574 -23612 32626
rect -23668 32572 -23612 32574
rect -23508 32626 -23452 32628
rect -23508 32574 -23506 32626
rect -23506 32574 -23454 32626
rect -23454 32574 -23452 32626
rect -23508 32572 -23452 32574
rect -23348 32626 -23292 32628
rect -23348 32574 -23346 32626
rect -23346 32574 -23294 32626
rect -23294 32574 -23292 32626
rect -23348 32572 -23292 32574
rect -23188 32626 -23132 32628
rect -23188 32574 -23186 32626
rect -23186 32574 -23134 32626
rect -23134 32574 -23132 32626
rect -23188 32572 -23132 32574
rect -23028 32626 -22972 32628
rect -23028 32574 -23026 32626
rect -23026 32574 -22974 32626
rect -22974 32574 -22972 32626
rect -23028 32572 -22972 32574
rect -22868 32626 -22812 32628
rect -22868 32574 -22866 32626
rect -22866 32574 -22814 32626
rect -22814 32574 -22812 32626
rect -22868 32572 -22812 32574
rect -22708 32626 -22652 32628
rect -22708 32574 -22706 32626
rect -22706 32574 -22654 32626
rect -22654 32574 -22652 32626
rect -22708 32572 -22652 32574
rect -22548 32626 -22492 32628
rect -22548 32574 -22546 32626
rect -22546 32574 -22494 32626
rect -22494 32574 -22492 32626
rect -22548 32572 -22492 32574
rect -22388 32626 -22332 32628
rect -22388 32574 -22386 32626
rect -22386 32574 -22334 32626
rect -22334 32574 -22332 32626
rect -22388 32572 -22332 32574
rect -22228 32626 -22172 32628
rect -22228 32574 -22226 32626
rect -22226 32574 -22174 32626
rect -22174 32574 -22172 32626
rect -22228 32572 -22172 32574
rect -22068 32626 -22012 32628
rect -22068 32574 -22066 32626
rect -22066 32574 -22014 32626
rect -22014 32574 -22012 32626
rect -22068 32572 -22012 32574
rect -21908 32626 -21852 32628
rect -21908 32574 -21906 32626
rect -21906 32574 -21854 32626
rect -21854 32574 -21852 32626
rect -21908 32572 -21852 32574
rect -21748 32626 -21692 32628
rect -21748 32574 -21746 32626
rect -21746 32574 -21694 32626
rect -21694 32574 -21692 32626
rect -21748 32572 -21692 32574
rect -21588 32626 -21532 32628
rect -21588 32574 -21586 32626
rect -21586 32574 -21534 32626
rect -21534 32574 -21532 32626
rect -21588 32572 -21532 32574
rect -21428 32626 -21372 32628
rect -21428 32574 -21426 32626
rect -21426 32574 -21374 32626
rect -21374 32574 -21372 32626
rect -21428 32572 -21372 32574
rect -21268 32626 -21212 32628
rect -21268 32574 -21266 32626
rect -21266 32574 -21214 32626
rect -21214 32574 -21212 32626
rect -21268 32572 -21212 32574
rect -21108 32626 -21052 32628
rect -21108 32574 -21106 32626
rect -21106 32574 -21054 32626
rect -21054 32574 -21052 32626
rect -21108 32572 -21052 32574
rect -20948 32626 -20892 32628
rect -20948 32574 -20946 32626
rect -20946 32574 -20894 32626
rect -20894 32574 -20892 32626
rect -20948 32572 -20892 32574
rect -20788 32626 -20732 32628
rect -20788 32574 -20786 32626
rect -20786 32574 -20734 32626
rect -20734 32574 -20732 32626
rect -20788 32572 -20732 32574
rect -20628 32626 -20572 32628
rect -20628 32574 -20626 32626
rect -20626 32574 -20574 32626
rect -20574 32574 -20572 32626
rect -20628 32572 -20572 32574
rect -20468 32626 -20412 32628
rect -20468 32574 -20466 32626
rect -20466 32574 -20414 32626
rect -20414 32574 -20412 32626
rect -20468 32572 -20412 32574
rect -20308 32626 -20252 32628
rect -20308 32574 -20306 32626
rect -20306 32574 -20254 32626
rect -20254 32574 -20252 32626
rect -20308 32572 -20252 32574
rect -20148 32626 -20092 32628
rect -20148 32574 -20146 32626
rect -20146 32574 -20094 32626
rect -20094 32574 -20092 32626
rect -20148 32572 -20092 32574
rect -19988 32626 -19932 32628
rect -19988 32574 -19986 32626
rect -19986 32574 -19934 32626
rect -19934 32574 -19932 32626
rect -19988 32572 -19932 32574
rect -19828 32626 -19772 32628
rect -19828 32574 -19826 32626
rect -19826 32574 -19774 32626
rect -19774 32574 -19772 32626
rect -19828 32572 -19772 32574
rect -19668 32626 -19612 32628
rect -19668 32574 -19666 32626
rect -19666 32574 -19614 32626
rect -19614 32574 -19612 32626
rect -19668 32572 -19612 32574
rect -19508 32626 -19452 32628
rect -19508 32574 -19506 32626
rect -19506 32574 -19454 32626
rect -19454 32574 -19452 32626
rect -19508 32572 -19452 32574
rect -19348 32626 -19292 32628
rect -19348 32574 -19346 32626
rect -19346 32574 -19294 32626
rect -19294 32574 -19292 32626
rect -19348 32572 -19292 32574
rect -19188 32626 -19132 32628
rect -19188 32574 -19186 32626
rect -19186 32574 -19134 32626
rect -19134 32574 -19132 32626
rect -19188 32572 -19132 32574
rect -19028 32626 -18972 32628
rect -19028 32574 -19026 32626
rect -19026 32574 -18974 32626
rect -18974 32574 -18972 32626
rect -19028 32572 -18972 32574
rect -18868 32626 -18812 32628
rect -18868 32574 -18866 32626
rect -18866 32574 -18814 32626
rect -18814 32574 -18812 32626
rect -18868 32572 -18812 32574
rect -18708 32626 -18652 32628
rect -18708 32574 -18706 32626
rect -18706 32574 -18654 32626
rect -18654 32574 -18652 32626
rect -18708 32572 -18652 32574
rect -18548 32626 -18492 32628
rect -18548 32574 -18546 32626
rect -18546 32574 -18494 32626
rect -18494 32574 -18492 32626
rect -18548 32572 -18492 32574
rect -18388 32626 -18332 32628
rect -18388 32574 -18386 32626
rect -18386 32574 -18334 32626
rect -18334 32574 -18332 32626
rect -18388 32572 -18332 32574
rect -18228 32626 -18172 32628
rect -18228 32574 -18226 32626
rect -18226 32574 -18174 32626
rect -18174 32574 -18172 32626
rect -18228 32572 -18172 32574
rect -18068 32626 -18012 32628
rect -18068 32574 -18066 32626
rect -18066 32574 -18014 32626
rect -18014 32574 -18012 32626
rect -18068 32572 -18012 32574
rect -17908 32626 -17852 32628
rect -17908 32574 -17906 32626
rect -17906 32574 -17854 32626
rect -17854 32574 -17852 32626
rect -17908 32572 -17852 32574
rect -17748 32626 -17692 32628
rect -17748 32574 -17746 32626
rect -17746 32574 -17694 32626
rect -17694 32574 -17692 32626
rect -17748 32572 -17692 32574
rect -17588 32626 -17532 32628
rect -17588 32574 -17586 32626
rect -17586 32574 -17534 32626
rect -17534 32574 -17532 32626
rect -17588 32572 -17532 32574
rect -17428 32626 -17372 32628
rect -17428 32574 -17426 32626
rect -17426 32574 -17374 32626
rect -17374 32574 -17372 32626
rect -17428 32572 -17372 32574
rect -17268 32626 -17212 32628
rect -17268 32574 -17266 32626
rect -17266 32574 -17214 32626
rect -17214 32574 -17212 32626
rect -17268 32572 -17212 32574
rect -17108 32626 -17052 32628
rect -17108 32574 -17106 32626
rect -17106 32574 -17054 32626
rect -17054 32574 -17052 32626
rect -17108 32572 -17052 32574
rect -16948 32626 -16892 32628
rect -16948 32574 -16946 32626
rect -16946 32574 -16894 32626
rect -16894 32574 -16892 32626
rect -16948 32572 -16892 32574
rect -16788 32626 -16732 32628
rect -16788 32574 -16786 32626
rect -16786 32574 -16734 32626
rect -16734 32574 -16732 32626
rect -16788 32572 -16732 32574
rect -16628 32626 -16572 32628
rect -16628 32574 -16626 32626
rect -16626 32574 -16574 32626
rect -16574 32574 -16572 32626
rect -16628 32572 -16572 32574
rect -16468 32626 -16412 32628
rect -16468 32574 -16466 32626
rect -16466 32574 -16414 32626
rect -16414 32574 -16412 32626
rect -16468 32572 -16412 32574
rect -16308 32626 -16252 32628
rect -16308 32574 -16306 32626
rect -16306 32574 -16254 32626
rect -16254 32574 -16252 32626
rect -16308 32572 -16252 32574
rect -16148 32626 -16092 32628
rect -16148 32574 -16146 32626
rect -16146 32574 -16094 32626
rect -16094 32574 -16092 32626
rect -16148 32572 -16092 32574
rect -15988 32626 -15932 32628
rect -15988 32574 -15986 32626
rect -15986 32574 -15934 32626
rect -15934 32574 -15932 32626
rect -15988 32572 -15932 32574
rect -15828 32626 -15772 32628
rect -15828 32574 -15826 32626
rect -15826 32574 -15774 32626
rect -15774 32574 -15772 32626
rect -15828 32572 -15772 32574
rect -15668 32626 -15612 32628
rect -15668 32574 -15666 32626
rect -15666 32574 -15614 32626
rect -15614 32574 -15612 32626
rect -15668 32572 -15612 32574
rect -15508 32626 -15452 32628
rect -15508 32574 -15506 32626
rect -15506 32574 -15454 32626
rect -15454 32574 -15452 32626
rect -15508 32572 -15452 32574
rect -15348 32626 -15292 32628
rect -15348 32574 -15346 32626
rect -15346 32574 -15294 32626
rect -15294 32574 -15292 32626
rect -15348 32572 -15292 32574
rect -15188 32626 -15132 32628
rect -15188 32574 -15186 32626
rect -15186 32574 -15134 32626
rect -15134 32574 -15132 32626
rect -15188 32572 -15132 32574
rect -15028 32626 -14972 32628
rect -15028 32574 -15026 32626
rect -15026 32574 -14974 32626
rect -14974 32574 -14972 32626
rect -15028 32572 -14972 32574
rect -14868 32626 -14812 32628
rect -14868 32574 -14866 32626
rect -14866 32574 -14814 32626
rect -14814 32574 -14812 32626
rect -14868 32572 -14812 32574
rect -14708 32626 -14652 32628
rect -14708 32574 -14706 32626
rect -14706 32574 -14654 32626
rect -14654 32574 -14652 32626
rect -14708 32572 -14652 32574
rect -14548 32626 -14492 32628
rect -14548 32574 -14546 32626
rect -14546 32574 -14494 32626
rect -14494 32574 -14492 32626
rect -14548 32572 -14492 32574
rect -14388 32626 -14332 32628
rect -14388 32574 -14386 32626
rect -14386 32574 -14334 32626
rect -14334 32574 -14332 32626
rect -14388 32572 -14332 32574
rect -14228 32626 -14172 32628
rect -14228 32574 -14226 32626
rect -14226 32574 -14174 32626
rect -14174 32574 -14172 32626
rect -14228 32572 -14172 32574
rect -14068 32626 -14012 32628
rect -14068 32574 -14066 32626
rect -14066 32574 -14014 32626
rect -14014 32574 -14012 32626
rect -14068 32572 -14012 32574
rect -13908 32626 -13852 32628
rect -13908 32574 -13906 32626
rect -13906 32574 -13854 32626
rect -13854 32574 -13852 32626
rect -13908 32572 -13852 32574
rect -13748 32626 -13692 32628
rect -13748 32574 -13746 32626
rect -13746 32574 -13694 32626
rect -13694 32574 -13692 32626
rect -13748 32572 -13692 32574
rect -13588 32626 -13532 32628
rect -13588 32574 -13586 32626
rect -13586 32574 -13534 32626
rect -13534 32574 -13532 32626
rect -13588 32572 -13532 32574
rect -13428 32626 -13372 32628
rect -13428 32574 -13426 32626
rect -13426 32574 -13374 32626
rect -13374 32574 -13372 32626
rect -13428 32572 -13372 32574
rect -13268 32626 -13212 32628
rect -13268 32574 -13266 32626
rect -13266 32574 -13214 32626
rect -13214 32574 -13212 32626
rect -13268 32572 -13212 32574
rect -13108 32626 -13052 32628
rect -13108 32574 -13106 32626
rect -13106 32574 -13054 32626
rect -13054 32574 -13052 32626
rect -13108 32572 -13052 32574
rect -12948 32626 -12892 32628
rect -12948 32574 -12946 32626
rect -12946 32574 -12894 32626
rect -12894 32574 -12892 32626
rect -12948 32572 -12892 32574
rect -12788 32626 -12732 32628
rect -12788 32574 -12786 32626
rect -12786 32574 -12734 32626
rect -12734 32574 -12732 32626
rect -12788 32572 -12732 32574
rect -12628 32626 -12572 32628
rect -12628 32574 -12626 32626
rect -12626 32574 -12574 32626
rect -12574 32574 -12572 32626
rect -12628 32572 -12572 32574
rect -12468 32626 -12412 32628
rect -12468 32574 -12466 32626
rect -12466 32574 -12414 32626
rect -12414 32574 -12412 32626
rect -12468 32572 -12412 32574
rect -12308 32626 -12252 32628
rect -12308 32574 -12306 32626
rect -12306 32574 -12254 32626
rect -12254 32574 -12252 32626
rect -12308 32572 -12252 32574
rect -12148 32626 -12092 32628
rect -12148 32574 -12146 32626
rect -12146 32574 -12094 32626
rect -12094 32574 -12092 32626
rect -12148 32572 -12092 32574
rect -11988 32626 -11932 32628
rect -11988 32574 -11986 32626
rect -11986 32574 -11934 32626
rect -11934 32574 -11932 32626
rect -11988 32572 -11932 32574
rect -11828 32626 -11772 32628
rect -11828 32574 -11826 32626
rect -11826 32574 -11774 32626
rect -11774 32574 -11772 32626
rect -11828 32572 -11772 32574
rect -11668 32626 -11612 32628
rect -11668 32574 -11666 32626
rect -11666 32574 -11614 32626
rect -11614 32574 -11612 32626
rect -11668 32572 -11612 32574
rect -11508 32626 -11452 32628
rect -11508 32574 -11506 32626
rect -11506 32574 -11454 32626
rect -11454 32574 -11452 32626
rect -11508 32572 -11452 32574
rect -11188 32626 -11132 32628
rect -11188 32574 -11186 32626
rect -11186 32574 -11134 32626
rect -11134 32574 -11132 32626
rect -11188 32572 -11132 32574
rect -10868 32626 -10812 32628
rect -10868 32574 -10866 32626
rect -10866 32574 -10814 32626
rect -10814 32574 -10812 32626
rect -10868 32572 -10812 32574
rect -10708 32626 -10652 32628
rect -10708 32574 -10706 32626
rect -10706 32574 -10654 32626
rect -10654 32574 -10652 32626
rect -10708 32572 -10652 32574
rect -10548 32626 -10492 32628
rect -10548 32574 -10546 32626
rect -10546 32574 -10494 32626
rect -10494 32574 -10492 32626
rect -10548 32572 -10492 32574
rect -10388 32626 -10332 32628
rect -10388 32574 -10386 32626
rect -10386 32574 -10334 32626
rect -10334 32574 -10332 32626
rect -10388 32572 -10332 32574
rect -10228 32626 -10172 32628
rect -10228 32574 -10226 32626
rect -10226 32574 -10174 32626
rect -10174 32574 -10172 32626
rect -10228 32572 -10172 32574
rect -10068 32626 -10012 32628
rect -10068 32574 -10066 32626
rect -10066 32574 -10014 32626
rect -10014 32574 -10012 32626
rect -10068 32572 -10012 32574
rect -9908 32626 -9852 32628
rect -9908 32574 -9906 32626
rect -9906 32574 -9854 32626
rect -9854 32574 -9852 32626
rect -9908 32572 -9852 32574
rect -9748 32626 -9692 32628
rect -9748 32574 -9746 32626
rect -9746 32574 -9694 32626
rect -9694 32574 -9692 32626
rect -9748 32572 -9692 32574
rect -9588 32626 -9532 32628
rect -9588 32574 -9586 32626
rect -9586 32574 -9534 32626
rect -9534 32574 -9532 32626
rect -9588 32572 -9532 32574
rect -9428 32626 -9372 32628
rect -9428 32574 -9426 32626
rect -9426 32574 -9374 32626
rect -9374 32574 -9372 32626
rect -9428 32572 -9372 32574
rect -9268 32626 -9212 32628
rect -9268 32574 -9266 32626
rect -9266 32574 -9214 32626
rect -9214 32574 -9212 32626
rect -9268 32572 -9212 32574
rect -9108 32626 -9052 32628
rect -9108 32574 -9106 32626
rect -9106 32574 -9054 32626
rect -9054 32574 -9052 32626
rect -9108 32572 -9052 32574
rect -8948 32626 -8892 32628
rect -8948 32574 -8946 32626
rect -8946 32574 -8894 32626
rect -8894 32574 -8892 32626
rect -8948 32572 -8892 32574
rect -8788 32626 -8732 32628
rect -8788 32574 -8786 32626
rect -8786 32574 -8734 32626
rect -8734 32574 -8732 32626
rect -8788 32572 -8732 32574
rect -8628 32626 -8572 32628
rect -8628 32574 -8626 32626
rect -8626 32574 -8574 32626
rect -8574 32574 -8572 32626
rect -8628 32572 -8572 32574
rect -8468 32626 -8412 32628
rect -8468 32574 -8466 32626
rect -8466 32574 -8414 32626
rect -8414 32574 -8412 32626
rect -8468 32572 -8412 32574
rect -8308 32626 -8252 32628
rect -8308 32574 -8306 32626
rect -8306 32574 -8254 32626
rect -8254 32574 -8252 32626
rect -8308 32572 -8252 32574
rect -8148 32626 -8092 32628
rect -8148 32574 -8146 32626
rect -8146 32574 -8094 32626
rect -8094 32574 -8092 32626
rect -8148 32572 -8092 32574
rect -7988 32626 -7932 32628
rect -7988 32574 -7986 32626
rect -7986 32574 -7934 32626
rect -7934 32574 -7932 32626
rect -7988 32572 -7932 32574
rect -7828 32626 -7772 32628
rect -7828 32574 -7826 32626
rect -7826 32574 -7774 32626
rect -7774 32574 -7772 32626
rect -7828 32572 -7772 32574
rect -7668 32626 -7612 32628
rect -7668 32574 -7666 32626
rect -7666 32574 -7614 32626
rect -7614 32574 -7612 32626
rect -7668 32572 -7612 32574
rect -7508 32626 -7452 32628
rect -7508 32574 -7506 32626
rect -7506 32574 -7454 32626
rect -7454 32574 -7452 32626
rect -7508 32572 -7452 32574
rect -7348 32626 -7292 32628
rect -7348 32574 -7346 32626
rect -7346 32574 -7294 32626
rect -7294 32574 -7292 32626
rect -7348 32572 -7292 32574
rect -7188 32626 -7132 32628
rect -7188 32574 -7186 32626
rect -7186 32574 -7134 32626
rect -7134 32574 -7132 32626
rect -7188 32572 -7132 32574
rect -7028 32626 -6972 32628
rect -7028 32574 -7026 32626
rect -7026 32574 -6974 32626
rect -6974 32574 -6972 32626
rect -7028 32572 -6972 32574
rect -6868 32626 -6812 32628
rect -6868 32574 -6866 32626
rect -6866 32574 -6814 32626
rect -6814 32574 -6812 32626
rect -6868 32572 -6812 32574
rect -6708 32626 -6652 32628
rect -6708 32574 -6706 32626
rect -6706 32574 -6654 32626
rect -6654 32574 -6652 32626
rect -6708 32572 -6652 32574
rect -6548 32626 -6492 32628
rect -6548 32574 -6546 32626
rect -6546 32574 -6494 32626
rect -6494 32574 -6492 32626
rect -6548 32572 -6492 32574
rect -6388 32626 -6332 32628
rect -6388 32574 -6386 32626
rect -6386 32574 -6334 32626
rect -6334 32574 -6332 32626
rect -6388 32572 -6332 32574
rect -6228 32626 -6172 32628
rect -6228 32574 -6226 32626
rect -6226 32574 -6174 32626
rect -6174 32574 -6172 32626
rect -6228 32572 -6172 32574
rect -6068 32626 -6012 32628
rect -6068 32574 -6066 32626
rect -6066 32574 -6014 32626
rect -6014 32574 -6012 32626
rect -6068 32572 -6012 32574
rect -5908 32626 -5852 32628
rect -5908 32574 -5906 32626
rect -5906 32574 -5854 32626
rect -5854 32574 -5852 32626
rect -5908 32572 -5852 32574
rect -5748 32626 -5692 32628
rect -5748 32574 -5746 32626
rect -5746 32574 -5694 32626
rect -5694 32574 -5692 32626
rect -5748 32572 -5692 32574
rect -5588 32626 -5532 32628
rect -5588 32574 -5586 32626
rect -5586 32574 -5534 32626
rect -5534 32574 -5532 32626
rect -5588 32572 -5532 32574
rect -5428 32626 -5372 32628
rect -5428 32574 -5426 32626
rect -5426 32574 -5374 32626
rect -5374 32574 -5372 32626
rect -5428 32572 -5372 32574
rect -5268 32626 -5212 32628
rect -5268 32574 -5266 32626
rect -5266 32574 -5214 32626
rect -5214 32574 -5212 32626
rect -5268 32572 -5212 32574
rect -5108 32626 -5052 32628
rect -5108 32574 -5106 32626
rect -5106 32574 -5054 32626
rect -5054 32574 -5052 32626
rect -5108 32572 -5052 32574
rect -4948 32626 -4892 32628
rect -4948 32574 -4946 32626
rect -4946 32574 -4894 32626
rect -4894 32574 -4892 32626
rect -4948 32572 -4892 32574
rect -4788 32626 -4732 32628
rect -4788 32574 -4786 32626
rect -4786 32574 -4734 32626
rect -4734 32574 -4732 32626
rect -4788 32572 -4732 32574
rect -4628 32626 -4572 32628
rect -4628 32574 -4626 32626
rect -4626 32574 -4574 32626
rect -4574 32574 -4572 32626
rect -4628 32572 -4572 32574
rect -4468 32626 -4412 32628
rect -4468 32574 -4466 32626
rect -4466 32574 -4414 32626
rect -4414 32574 -4412 32626
rect -4468 32572 -4412 32574
rect -4308 32626 -4252 32628
rect -4308 32574 -4306 32626
rect -4306 32574 -4254 32626
rect -4254 32574 -4252 32626
rect -4308 32572 -4252 32574
rect -4148 32626 -4092 32628
rect -4148 32574 -4146 32626
rect -4146 32574 -4094 32626
rect -4094 32574 -4092 32626
rect -4148 32572 -4092 32574
rect -3988 32626 -3932 32628
rect -3988 32574 -3986 32626
rect -3986 32574 -3934 32626
rect -3934 32574 -3932 32626
rect -3988 32572 -3932 32574
rect -3668 32626 -3612 32628
rect -3668 32574 -3666 32626
rect -3666 32574 -3614 32626
rect -3614 32574 -3612 32626
rect -3668 32572 -3612 32574
rect -3508 32626 -3452 32628
rect -3508 32574 -3506 32626
rect -3506 32574 -3454 32626
rect -3454 32574 -3452 32626
rect -3508 32572 -3452 32574
rect -3348 32626 -3292 32628
rect -3348 32574 -3346 32626
rect -3346 32574 -3294 32626
rect -3294 32574 -3292 32626
rect -3348 32572 -3292 32574
rect -3188 32626 -3132 32628
rect -3188 32574 -3186 32626
rect -3186 32574 -3134 32626
rect -3134 32574 -3132 32626
rect -3188 32572 -3132 32574
rect -3028 32626 -2972 32628
rect -3028 32574 -3026 32626
rect -3026 32574 -2974 32626
rect -2974 32574 -2972 32626
rect -3028 32572 -2972 32574
rect -2868 32626 -2812 32628
rect -2868 32574 -2866 32626
rect -2866 32574 -2814 32626
rect -2814 32574 -2812 32626
rect -2868 32572 -2812 32574
rect -2708 32626 -2652 32628
rect -2708 32574 -2706 32626
rect -2706 32574 -2654 32626
rect -2654 32574 -2652 32626
rect -2708 32572 -2652 32574
rect -2388 32626 -2332 32628
rect -2388 32574 -2386 32626
rect -2386 32574 -2334 32626
rect -2334 32574 -2332 32626
rect -2388 32572 -2332 32574
rect -2068 32626 -2012 32628
rect -2068 32574 -2066 32626
rect -2066 32574 -2014 32626
rect -2014 32574 -2012 32626
rect -2068 32572 -2012 32574
rect -1748 32626 -1692 32628
rect -1748 32574 -1746 32626
rect -1746 32574 -1694 32626
rect -1694 32574 -1692 32626
rect -1748 32572 -1692 32574
rect -1428 32626 -1372 32628
rect -1428 32574 -1426 32626
rect -1426 32574 -1374 32626
rect -1374 32574 -1372 32626
rect -1428 32572 -1372 32574
rect -1108 32626 -1052 32628
rect -1108 32574 -1106 32626
rect -1106 32574 -1054 32626
rect -1054 32574 -1052 32626
rect -1108 32572 -1052 32574
rect -31028 32412 -30972 32468
rect -30708 32412 -30652 32468
rect -30228 32412 -30172 32468
rect -11348 32412 -11292 32468
rect -2548 32412 -2492 32468
rect -31028 32252 -30972 32308
rect -30708 32252 -30652 32308
rect -30388 32252 -30332 32308
rect -30068 32252 -30012 32308
rect -29908 32306 -29852 32308
rect -29908 32254 -29906 32306
rect -29906 32254 -29854 32306
rect -29854 32254 -29852 32306
rect -29908 32252 -29852 32254
rect -29748 32306 -29692 32308
rect -29748 32254 -29746 32306
rect -29746 32254 -29694 32306
rect -29694 32254 -29692 32306
rect -29748 32252 -29692 32254
rect -29588 32306 -29532 32308
rect -29588 32254 -29586 32306
rect -29586 32254 -29534 32306
rect -29534 32254 -29532 32306
rect -29588 32252 -29532 32254
rect -29428 32306 -29372 32308
rect -29428 32254 -29426 32306
rect -29426 32254 -29374 32306
rect -29374 32254 -29372 32306
rect -29428 32252 -29372 32254
rect -29268 32306 -29212 32308
rect -29268 32254 -29266 32306
rect -29266 32254 -29214 32306
rect -29214 32254 -29212 32306
rect -29268 32252 -29212 32254
rect -29108 32306 -29052 32308
rect -29108 32254 -29106 32306
rect -29106 32254 -29054 32306
rect -29054 32254 -29052 32306
rect -29108 32252 -29052 32254
rect -28948 32306 -28892 32308
rect -28948 32254 -28946 32306
rect -28946 32254 -28894 32306
rect -28894 32254 -28892 32306
rect -28948 32252 -28892 32254
rect -28788 32306 -28732 32308
rect -28788 32254 -28786 32306
rect -28786 32254 -28734 32306
rect -28734 32254 -28732 32306
rect -28788 32252 -28732 32254
rect -28628 32306 -28572 32308
rect -28628 32254 -28626 32306
rect -28626 32254 -28574 32306
rect -28574 32254 -28572 32306
rect -28628 32252 -28572 32254
rect -28468 32306 -28412 32308
rect -28468 32254 -28466 32306
rect -28466 32254 -28414 32306
rect -28414 32254 -28412 32306
rect -28468 32252 -28412 32254
rect -28308 32306 -28252 32308
rect -28308 32254 -28306 32306
rect -28306 32254 -28254 32306
rect -28254 32254 -28252 32306
rect -28308 32252 -28252 32254
rect -28148 32306 -28092 32308
rect -28148 32254 -28146 32306
rect -28146 32254 -28094 32306
rect -28094 32254 -28092 32306
rect -28148 32252 -28092 32254
rect -27988 32306 -27932 32308
rect -27988 32254 -27986 32306
rect -27986 32254 -27934 32306
rect -27934 32254 -27932 32306
rect -27988 32252 -27932 32254
rect -27828 32306 -27772 32308
rect -27828 32254 -27826 32306
rect -27826 32254 -27774 32306
rect -27774 32254 -27772 32306
rect -27828 32252 -27772 32254
rect -27668 32306 -27612 32308
rect -27668 32254 -27666 32306
rect -27666 32254 -27614 32306
rect -27614 32254 -27612 32306
rect -27668 32252 -27612 32254
rect -27508 32306 -27452 32308
rect -27508 32254 -27506 32306
rect -27506 32254 -27454 32306
rect -27454 32254 -27452 32306
rect -27508 32252 -27452 32254
rect -27348 32306 -27292 32308
rect -27348 32254 -27346 32306
rect -27346 32254 -27294 32306
rect -27294 32254 -27292 32306
rect -27348 32252 -27292 32254
rect -27188 32306 -27132 32308
rect -27188 32254 -27186 32306
rect -27186 32254 -27134 32306
rect -27134 32254 -27132 32306
rect -27188 32252 -27132 32254
rect -27028 32306 -26972 32308
rect -27028 32254 -27026 32306
rect -27026 32254 -26974 32306
rect -26974 32254 -26972 32306
rect -27028 32252 -26972 32254
rect -26868 32306 -26812 32308
rect -26868 32254 -26866 32306
rect -26866 32254 -26814 32306
rect -26814 32254 -26812 32306
rect -26868 32252 -26812 32254
rect -26708 32306 -26652 32308
rect -26708 32254 -26706 32306
rect -26706 32254 -26654 32306
rect -26654 32254 -26652 32306
rect -26708 32252 -26652 32254
rect -26548 32306 -26492 32308
rect -26548 32254 -26546 32306
rect -26546 32254 -26494 32306
rect -26494 32254 -26492 32306
rect -26548 32252 -26492 32254
rect -26388 32306 -26332 32308
rect -26388 32254 -26386 32306
rect -26386 32254 -26334 32306
rect -26334 32254 -26332 32306
rect -26388 32252 -26332 32254
rect -26228 32306 -26172 32308
rect -26228 32254 -26226 32306
rect -26226 32254 -26174 32306
rect -26174 32254 -26172 32306
rect -26228 32252 -26172 32254
rect -26068 32306 -26012 32308
rect -26068 32254 -26066 32306
rect -26066 32254 -26014 32306
rect -26014 32254 -26012 32306
rect -26068 32252 -26012 32254
rect -25908 32306 -25852 32308
rect -25908 32254 -25906 32306
rect -25906 32254 -25854 32306
rect -25854 32254 -25852 32306
rect -25908 32252 -25852 32254
rect -25748 32306 -25692 32308
rect -25748 32254 -25746 32306
rect -25746 32254 -25694 32306
rect -25694 32254 -25692 32306
rect -25748 32252 -25692 32254
rect -25588 32306 -25532 32308
rect -25588 32254 -25586 32306
rect -25586 32254 -25534 32306
rect -25534 32254 -25532 32306
rect -25588 32252 -25532 32254
rect -25428 32306 -25372 32308
rect -25428 32254 -25426 32306
rect -25426 32254 -25374 32306
rect -25374 32254 -25372 32306
rect -25428 32252 -25372 32254
rect -25268 32306 -25212 32308
rect -25268 32254 -25266 32306
rect -25266 32254 -25214 32306
rect -25214 32254 -25212 32306
rect -25268 32252 -25212 32254
rect -25108 32306 -25052 32308
rect -25108 32254 -25106 32306
rect -25106 32254 -25054 32306
rect -25054 32254 -25052 32306
rect -25108 32252 -25052 32254
rect -24948 32306 -24892 32308
rect -24948 32254 -24946 32306
rect -24946 32254 -24894 32306
rect -24894 32254 -24892 32306
rect -24948 32252 -24892 32254
rect -24788 32306 -24732 32308
rect -24788 32254 -24786 32306
rect -24786 32254 -24734 32306
rect -24734 32254 -24732 32306
rect -24788 32252 -24732 32254
rect -24628 32306 -24572 32308
rect -24628 32254 -24626 32306
rect -24626 32254 -24574 32306
rect -24574 32254 -24572 32306
rect -24628 32252 -24572 32254
rect -24468 32306 -24412 32308
rect -24468 32254 -24466 32306
rect -24466 32254 -24414 32306
rect -24414 32254 -24412 32306
rect -24468 32252 -24412 32254
rect -24308 32306 -24252 32308
rect -24308 32254 -24306 32306
rect -24306 32254 -24254 32306
rect -24254 32254 -24252 32306
rect -24308 32252 -24252 32254
rect -24148 32306 -24092 32308
rect -24148 32254 -24146 32306
rect -24146 32254 -24094 32306
rect -24094 32254 -24092 32306
rect -24148 32252 -24092 32254
rect -23988 32306 -23932 32308
rect -23988 32254 -23986 32306
rect -23986 32254 -23934 32306
rect -23934 32254 -23932 32306
rect -23988 32252 -23932 32254
rect -23828 32306 -23772 32308
rect -23828 32254 -23826 32306
rect -23826 32254 -23774 32306
rect -23774 32254 -23772 32306
rect -23828 32252 -23772 32254
rect -23668 32306 -23612 32308
rect -23668 32254 -23666 32306
rect -23666 32254 -23614 32306
rect -23614 32254 -23612 32306
rect -23668 32252 -23612 32254
rect -23508 32306 -23452 32308
rect -23508 32254 -23506 32306
rect -23506 32254 -23454 32306
rect -23454 32254 -23452 32306
rect -23508 32252 -23452 32254
rect -23348 32306 -23292 32308
rect -23348 32254 -23346 32306
rect -23346 32254 -23294 32306
rect -23294 32254 -23292 32306
rect -23348 32252 -23292 32254
rect -23188 32306 -23132 32308
rect -23188 32254 -23186 32306
rect -23186 32254 -23134 32306
rect -23134 32254 -23132 32306
rect -23188 32252 -23132 32254
rect -23028 32306 -22972 32308
rect -23028 32254 -23026 32306
rect -23026 32254 -22974 32306
rect -22974 32254 -22972 32306
rect -23028 32252 -22972 32254
rect -22868 32306 -22812 32308
rect -22868 32254 -22866 32306
rect -22866 32254 -22814 32306
rect -22814 32254 -22812 32306
rect -22868 32252 -22812 32254
rect -22708 32306 -22652 32308
rect -22708 32254 -22706 32306
rect -22706 32254 -22654 32306
rect -22654 32254 -22652 32306
rect -22708 32252 -22652 32254
rect -22548 32306 -22492 32308
rect -22548 32254 -22546 32306
rect -22546 32254 -22494 32306
rect -22494 32254 -22492 32306
rect -22548 32252 -22492 32254
rect -22388 32306 -22332 32308
rect -22388 32254 -22386 32306
rect -22386 32254 -22334 32306
rect -22334 32254 -22332 32306
rect -22388 32252 -22332 32254
rect -22228 32306 -22172 32308
rect -22228 32254 -22226 32306
rect -22226 32254 -22174 32306
rect -22174 32254 -22172 32306
rect -22228 32252 -22172 32254
rect -22068 32306 -22012 32308
rect -22068 32254 -22066 32306
rect -22066 32254 -22014 32306
rect -22014 32254 -22012 32306
rect -22068 32252 -22012 32254
rect -21908 32306 -21852 32308
rect -21908 32254 -21906 32306
rect -21906 32254 -21854 32306
rect -21854 32254 -21852 32306
rect -21908 32252 -21852 32254
rect -21748 32306 -21692 32308
rect -21748 32254 -21746 32306
rect -21746 32254 -21694 32306
rect -21694 32254 -21692 32306
rect -21748 32252 -21692 32254
rect -21588 32306 -21532 32308
rect -21588 32254 -21586 32306
rect -21586 32254 -21534 32306
rect -21534 32254 -21532 32306
rect -21588 32252 -21532 32254
rect -21428 32306 -21372 32308
rect -21428 32254 -21426 32306
rect -21426 32254 -21374 32306
rect -21374 32254 -21372 32306
rect -21428 32252 -21372 32254
rect -21268 32306 -21212 32308
rect -21268 32254 -21266 32306
rect -21266 32254 -21214 32306
rect -21214 32254 -21212 32306
rect -21268 32252 -21212 32254
rect -21108 32306 -21052 32308
rect -21108 32254 -21106 32306
rect -21106 32254 -21054 32306
rect -21054 32254 -21052 32306
rect -21108 32252 -21052 32254
rect -20948 32306 -20892 32308
rect -20948 32254 -20946 32306
rect -20946 32254 -20894 32306
rect -20894 32254 -20892 32306
rect -20948 32252 -20892 32254
rect -20788 32306 -20732 32308
rect -20788 32254 -20786 32306
rect -20786 32254 -20734 32306
rect -20734 32254 -20732 32306
rect -20788 32252 -20732 32254
rect -20628 32306 -20572 32308
rect -20628 32254 -20626 32306
rect -20626 32254 -20574 32306
rect -20574 32254 -20572 32306
rect -20628 32252 -20572 32254
rect -20468 32306 -20412 32308
rect -20468 32254 -20466 32306
rect -20466 32254 -20414 32306
rect -20414 32254 -20412 32306
rect -20468 32252 -20412 32254
rect -20308 32306 -20252 32308
rect -20308 32254 -20306 32306
rect -20306 32254 -20254 32306
rect -20254 32254 -20252 32306
rect -20308 32252 -20252 32254
rect -20148 32306 -20092 32308
rect -20148 32254 -20146 32306
rect -20146 32254 -20094 32306
rect -20094 32254 -20092 32306
rect -20148 32252 -20092 32254
rect -19988 32306 -19932 32308
rect -19988 32254 -19986 32306
rect -19986 32254 -19934 32306
rect -19934 32254 -19932 32306
rect -19988 32252 -19932 32254
rect -19828 32306 -19772 32308
rect -19828 32254 -19826 32306
rect -19826 32254 -19774 32306
rect -19774 32254 -19772 32306
rect -19828 32252 -19772 32254
rect -19668 32306 -19612 32308
rect -19668 32254 -19666 32306
rect -19666 32254 -19614 32306
rect -19614 32254 -19612 32306
rect -19668 32252 -19612 32254
rect -19508 32306 -19452 32308
rect -19508 32254 -19506 32306
rect -19506 32254 -19454 32306
rect -19454 32254 -19452 32306
rect -19508 32252 -19452 32254
rect -19348 32306 -19292 32308
rect -19348 32254 -19346 32306
rect -19346 32254 -19294 32306
rect -19294 32254 -19292 32306
rect -19348 32252 -19292 32254
rect -19188 32306 -19132 32308
rect -19188 32254 -19186 32306
rect -19186 32254 -19134 32306
rect -19134 32254 -19132 32306
rect -19188 32252 -19132 32254
rect -19028 32306 -18972 32308
rect -19028 32254 -19026 32306
rect -19026 32254 -18974 32306
rect -18974 32254 -18972 32306
rect -19028 32252 -18972 32254
rect -18868 32306 -18812 32308
rect -18868 32254 -18866 32306
rect -18866 32254 -18814 32306
rect -18814 32254 -18812 32306
rect -18868 32252 -18812 32254
rect -18708 32306 -18652 32308
rect -18708 32254 -18706 32306
rect -18706 32254 -18654 32306
rect -18654 32254 -18652 32306
rect -18708 32252 -18652 32254
rect -18548 32306 -18492 32308
rect -18548 32254 -18546 32306
rect -18546 32254 -18494 32306
rect -18494 32254 -18492 32306
rect -18548 32252 -18492 32254
rect -18388 32306 -18332 32308
rect -18388 32254 -18386 32306
rect -18386 32254 -18334 32306
rect -18334 32254 -18332 32306
rect -18388 32252 -18332 32254
rect -18228 32306 -18172 32308
rect -18228 32254 -18226 32306
rect -18226 32254 -18174 32306
rect -18174 32254 -18172 32306
rect -18228 32252 -18172 32254
rect -18068 32306 -18012 32308
rect -18068 32254 -18066 32306
rect -18066 32254 -18014 32306
rect -18014 32254 -18012 32306
rect -18068 32252 -18012 32254
rect -17908 32306 -17852 32308
rect -17908 32254 -17906 32306
rect -17906 32254 -17854 32306
rect -17854 32254 -17852 32306
rect -17908 32252 -17852 32254
rect -17748 32306 -17692 32308
rect -17748 32254 -17746 32306
rect -17746 32254 -17694 32306
rect -17694 32254 -17692 32306
rect -17748 32252 -17692 32254
rect -17588 32306 -17532 32308
rect -17588 32254 -17586 32306
rect -17586 32254 -17534 32306
rect -17534 32254 -17532 32306
rect -17588 32252 -17532 32254
rect -17428 32306 -17372 32308
rect -17428 32254 -17426 32306
rect -17426 32254 -17374 32306
rect -17374 32254 -17372 32306
rect -17428 32252 -17372 32254
rect -17268 32306 -17212 32308
rect -17268 32254 -17266 32306
rect -17266 32254 -17214 32306
rect -17214 32254 -17212 32306
rect -17268 32252 -17212 32254
rect -17108 32306 -17052 32308
rect -17108 32254 -17106 32306
rect -17106 32254 -17054 32306
rect -17054 32254 -17052 32306
rect -17108 32252 -17052 32254
rect -16948 32306 -16892 32308
rect -16948 32254 -16946 32306
rect -16946 32254 -16894 32306
rect -16894 32254 -16892 32306
rect -16948 32252 -16892 32254
rect -16788 32306 -16732 32308
rect -16788 32254 -16786 32306
rect -16786 32254 -16734 32306
rect -16734 32254 -16732 32306
rect -16788 32252 -16732 32254
rect -16628 32306 -16572 32308
rect -16628 32254 -16626 32306
rect -16626 32254 -16574 32306
rect -16574 32254 -16572 32306
rect -16628 32252 -16572 32254
rect -16468 32306 -16412 32308
rect -16468 32254 -16466 32306
rect -16466 32254 -16414 32306
rect -16414 32254 -16412 32306
rect -16468 32252 -16412 32254
rect -16308 32306 -16252 32308
rect -16308 32254 -16306 32306
rect -16306 32254 -16254 32306
rect -16254 32254 -16252 32306
rect -16308 32252 -16252 32254
rect -16148 32306 -16092 32308
rect -16148 32254 -16146 32306
rect -16146 32254 -16094 32306
rect -16094 32254 -16092 32306
rect -16148 32252 -16092 32254
rect -15988 32306 -15932 32308
rect -15988 32254 -15986 32306
rect -15986 32254 -15934 32306
rect -15934 32254 -15932 32306
rect -15988 32252 -15932 32254
rect -15828 32306 -15772 32308
rect -15828 32254 -15826 32306
rect -15826 32254 -15774 32306
rect -15774 32254 -15772 32306
rect -15828 32252 -15772 32254
rect -15668 32306 -15612 32308
rect -15668 32254 -15666 32306
rect -15666 32254 -15614 32306
rect -15614 32254 -15612 32306
rect -15668 32252 -15612 32254
rect -15508 32306 -15452 32308
rect -15508 32254 -15506 32306
rect -15506 32254 -15454 32306
rect -15454 32254 -15452 32306
rect -15508 32252 -15452 32254
rect -15348 32306 -15292 32308
rect -15348 32254 -15346 32306
rect -15346 32254 -15294 32306
rect -15294 32254 -15292 32306
rect -15348 32252 -15292 32254
rect -15188 32306 -15132 32308
rect -15188 32254 -15186 32306
rect -15186 32254 -15134 32306
rect -15134 32254 -15132 32306
rect -15188 32252 -15132 32254
rect -15028 32306 -14972 32308
rect -15028 32254 -15026 32306
rect -15026 32254 -14974 32306
rect -14974 32254 -14972 32306
rect -15028 32252 -14972 32254
rect -14868 32306 -14812 32308
rect -14868 32254 -14866 32306
rect -14866 32254 -14814 32306
rect -14814 32254 -14812 32306
rect -14868 32252 -14812 32254
rect -14708 32306 -14652 32308
rect -14708 32254 -14706 32306
rect -14706 32254 -14654 32306
rect -14654 32254 -14652 32306
rect -14708 32252 -14652 32254
rect -14548 32306 -14492 32308
rect -14548 32254 -14546 32306
rect -14546 32254 -14494 32306
rect -14494 32254 -14492 32306
rect -14548 32252 -14492 32254
rect -14388 32306 -14332 32308
rect -14388 32254 -14386 32306
rect -14386 32254 -14334 32306
rect -14334 32254 -14332 32306
rect -14388 32252 -14332 32254
rect -14228 32306 -14172 32308
rect -14228 32254 -14226 32306
rect -14226 32254 -14174 32306
rect -14174 32254 -14172 32306
rect -14228 32252 -14172 32254
rect -14068 32306 -14012 32308
rect -14068 32254 -14066 32306
rect -14066 32254 -14014 32306
rect -14014 32254 -14012 32306
rect -14068 32252 -14012 32254
rect -13908 32306 -13852 32308
rect -13908 32254 -13906 32306
rect -13906 32254 -13854 32306
rect -13854 32254 -13852 32306
rect -13908 32252 -13852 32254
rect -13748 32306 -13692 32308
rect -13748 32254 -13746 32306
rect -13746 32254 -13694 32306
rect -13694 32254 -13692 32306
rect -13748 32252 -13692 32254
rect -13588 32306 -13532 32308
rect -13588 32254 -13586 32306
rect -13586 32254 -13534 32306
rect -13534 32254 -13532 32306
rect -13588 32252 -13532 32254
rect -13428 32306 -13372 32308
rect -13428 32254 -13426 32306
rect -13426 32254 -13374 32306
rect -13374 32254 -13372 32306
rect -13428 32252 -13372 32254
rect -13268 32306 -13212 32308
rect -13268 32254 -13266 32306
rect -13266 32254 -13214 32306
rect -13214 32254 -13212 32306
rect -13268 32252 -13212 32254
rect -13108 32306 -13052 32308
rect -13108 32254 -13106 32306
rect -13106 32254 -13054 32306
rect -13054 32254 -13052 32306
rect -13108 32252 -13052 32254
rect -12948 32306 -12892 32308
rect -12948 32254 -12946 32306
rect -12946 32254 -12894 32306
rect -12894 32254 -12892 32306
rect -12948 32252 -12892 32254
rect -12788 32306 -12732 32308
rect -12788 32254 -12786 32306
rect -12786 32254 -12734 32306
rect -12734 32254 -12732 32306
rect -12788 32252 -12732 32254
rect -12628 32306 -12572 32308
rect -12628 32254 -12626 32306
rect -12626 32254 -12574 32306
rect -12574 32254 -12572 32306
rect -12628 32252 -12572 32254
rect -12468 32306 -12412 32308
rect -12468 32254 -12466 32306
rect -12466 32254 -12414 32306
rect -12414 32254 -12412 32306
rect -12468 32252 -12412 32254
rect -12308 32306 -12252 32308
rect -12308 32254 -12306 32306
rect -12306 32254 -12254 32306
rect -12254 32254 -12252 32306
rect -12308 32252 -12252 32254
rect -12148 32306 -12092 32308
rect -12148 32254 -12146 32306
rect -12146 32254 -12094 32306
rect -12094 32254 -12092 32306
rect -12148 32252 -12092 32254
rect -11988 32306 -11932 32308
rect -11988 32254 -11986 32306
rect -11986 32254 -11934 32306
rect -11934 32254 -11932 32306
rect -11988 32252 -11932 32254
rect -11828 32306 -11772 32308
rect -11828 32254 -11826 32306
rect -11826 32254 -11774 32306
rect -11774 32254 -11772 32306
rect -11828 32252 -11772 32254
rect -11668 32306 -11612 32308
rect -11668 32254 -11666 32306
rect -11666 32254 -11614 32306
rect -11614 32254 -11612 32306
rect -11668 32252 -11612 32254
rect -11508 32306 -11452 32308
rect -11508 32254 -11506 32306
rect -11506 32254 -11454 32306
rect -11454 32254 -11452 32306
rect -11508 32252 -11452 32254
rect -11348 32306 -11292 32308
rect -11348 32254 -11346 32306
rect -11346 32254 -11294 32306
rect -11294 32254 -11292 32306
rect -11348 32252 -11292 32254
rect -11188 32306 -11132 32308
rect -11188 32254 -11186 32306
rect -11186 32254 -11134 32306
rect -11134 32254 -11132 32306
rect -11188 32252 -11132 32254
rect -10868 32306 -10812 32308
rect -10868 32254 -10866 32306
rect -10866 32254 -10814 32306
rect -10814 32254 -10812 32306
rect -10868 32252 -10812 32254
rect -10708 32306 -10652 32308
rect -10708 32254 -10706 32306
rect -10706 32254 -10654 32306
rect -10654 32254 -10652 32306
rect -10708 32252 -10652 32254
rect -10548 32306 -10492 32308
rect -10548 32254 -10546 32306
rect -10546 32254 -10494 32306
rect -10494 32254 -10492 32306
rect -10548 32252 -10492 32254
rect -10388 32306 -10332 32308
rect -10388 32254 -10386 32306
rect -10386 32254 -10334 32306
rect -10334 32254 -10332 32306
rect -10388 32252 -10332 32254
rect -10228 32306 -10172 32308
rect -10228 32254 -10226 32306
rect -10226 32254 -10174 32306
rect -10174 32254 -10172 32306
rect -10228 32252 -10172 32254
rect -10068 32306 -10012 32308
rect -10068 32254 -10066 32306
rect -10066 32254 -10014 32306
rect -10014 32254 -10012 32306
rect -10068 32252 -10012 32254
rect -9908 32306 -9852 32308
rect -9908 32254 -9906 32306
rect -9906 32254 -9854 32306
rect -9854 32254 -9852 32306
rect -9908 32252 -9852 32254
rect -9748 32306 -9692 32308
rect -9748 32254 -9746 32306
rect -9746 32254 -9694 32306
rect -9694 32254 -9692 32306
rect -9748 32252 -9692 32254
rect -9588 32306 -9532 32308
rect -9588 32254 -9586 32306
rect -9586 32254 -9534 32306
rect -9534 32254 -9532 32306
rect -9588 32252 -9532 32254
rect -9428 32306 -9372 32308
rect -9428 32254 -9426 32306
rect -9426 32254 -9374 32306
rect -9374 32254 -9372 32306
rect -9428 32252 -9372 32254
rect -9268 32306 -9212 32308
rect -9268 32254 -9266 32306
rect -9266 32254 -9214 32306
rect -9214 32254 -9212 32306
rect -9268 32252 -9212 32254
rect -9108 32306 -9052 32308
rect -9108 32254 -9106 32306
rect -9106 32254 -9054 32306
rect -9054 32254 -9052 32306
rect -9108 32252 -9052 32254
rect -8948 32306 -8892 32308
rect -8948 32254 -8946 32306
rect -8946 32254 -8894 32306
rect -8894 32254 -8892 32306
rect -8948 32252 -8892 32254
rect -8788 32306 -8732 32308
rect -8788 32254 -8786 32306
rect -8786 32254 -8734 32306
rect -8734 32254 -8732 32306
rect -8788 32252 -8732 32254
rect -8628 32306 -8572 32308
rect -8628 32254 -8626 32306
rect -8626 32254 -8574 32306
rect -8574 32254 -8572 32306
rect -8628 32252 -8572 32254
rect -8468 32306 -8412 32308
rect -8468 32254 -8466 32306
rect -8466 32254 -8414 32306
rect -8414 32254 -8412 32306
rect -8468 32252 -8412 32254
rect -8308 32306 -8252 32308
rect -8308 32254 -8306 32306
rect -8306 32254 -8254 32306
rect -8254 32254 -8252 32306
rect -8308 32252 -8252 32254
rect -8148 32306 -8092 32308
rect -8148 32254 -8146 32306
rect -8146 32254 -8094 32306
rect -8094 32254 -8092 32306
rect -8148 32252 -8092 32254
rect -7988 32306 -7932 32308
rect -7988 32254 -7986 32306
rect -7986 32254 -7934 32306
rect -7934 32254 -7932 32306
rect -7988 32252 -7932 32254
rect -7828 32306 -7772 32308
rect -7828 32254 -7826 32306
rect -7826 32254 -7774 32306
rect -7774 32254 -7772 32306
rect -7828 32252 -7772 32254
rect -7668 32306 -7612 32308
rect -7668 32254 -7666 32306
rect -7666 32254 -7614 32306
rect -7614 32254 -7612 32306
rect -7668 32252 -7612 32254
rect -7508 32306 -7452 32308
rect -7508 32254 -7506 32306
rect -7506 32254 -7454 32306
rect -7454 32254 -7452 32306
rect -7508 32252 -7452 32254
rect -7348 32306 -7292 32308
rect -7348 32254 -7346 32306
rect -7346 32254 -7294 32306
rect -7294 32254 -7292 32306
rect -7348 32252 -7292 32254
rect -7188 32306 -7132 32308
rect -7188 32254 -7186 32306
rect -7186 32254 -7134 32306
rect -7134 32254 -7132 32306
rect -7188 32252 -7132 32254
rect -7028 32306 -6972 32308
rect -7028 32254 -7026 32306
rect -7026 32254 -6974 32306
rect -6974 32254 -6972 32306
rect -7028 32252 -6972 32254
rect -6868 32306 -6812 32308
rect -6868 32254 -6866 32306
rect -6866 32254 -6814 32306
rect -6814 32254 -6812 32306
rect -6868 32252 -6812 32254
rect -6708 32306 -6652 32308
rect -6708 32254 -6706 32306
rect -6706 32254 -6654 32306
rect -6654 32254 -6652 32306
rect -6708 32252 -6652 32254
rect -6548 32306 -6492 32308
rect -6548 32254 -6546 32306
rect -6546 32254 -6494 32306
rect -6494 32254 -6492 32306
rect -6548 32252 -6492 32254
rect -6388 32306 -6332 32308
rect -6388 32254 -6386 32306
rect -6386 32254 -6334 32306
rect -6334 32254 -6332 32306
rect -6388 32252 -6332 32254
rect -6228 32306 -6172 32308
rect -6228 32254 -6226 32306
rect -6226 32254 -6174 32306
rect -6174 32254 -6172 32306
rect -6228 32252 -6172 32254
rect -6068 32306 -6012 32308
rect -6068 32254 -6066 32306
rect -6066 32254 -6014 32306
rect -6014 32254 -6012 32306
rect -6068 32252 -6012 32254
rect -5908 32306 -5852 32308
rect -5908 32254 -5906 32306
rect -5906 32254 -5854 32306
rect -5854 32254 -5852 32306
rect -5908 32252 -5852 32254
rect -5748 32306 -5692 32308
rect -5748 32254 -5746 32306
rect -5746 32254 -5694 32306
rect -5694 32254 -5692 32306
rect -5748 32252 -5692 32254
rect -5588 32306 -5532 32308
rect -5588 32254 -5586 32306
rect -5586 32254 -5534 32306
rect -5534 32254 -5532 32306
rect -5588 32252 -5532 32254
rect -5428 32306 -5372 32308
rect -5428 32254 -5426 32306
rect -5426 32254 -5374 32306
rect -5374 32254 -5372 32306
rect -5428 32252 -5372 32254
rect -5268 32306 -5212 32308
rect -5268 32254 -5266 32306
rect -5266 32254 -5214 32306
rect -5214 32254 -5212 32306
rect -5268 32252 -5212 32254
rect -5108 32306 -5052 32308
rect -5108 32254 -5106 32306
rect -5106 32254 -5054 32306
rect -5054 32254 -5052 32306
rect -5108 32252 -5052 32254
rect -4948 32306 -4892 32308
rect -4948 32254 -4946 32306
rect -4946 32254 -4894 32306
rect -4894 32254 -4892 32306
rect -4948 32252 -4892 32254
rect -4788 32306 -4732 32308
rect -4788 32254 -4786 32306
rect -4786 32254 -4734 32306
rect -4734 32254 -4732 32306
rect -4788 32252 -4732 32254
rect -4628 32306 -4572 32308
rect -4628 32254 -4626 32306
rect -4626 32254 -4574 32306
rect -4574 32254 -4572 32306
rect -4628 32252 -4572 32254
rect -4468 32306 -4412 32308
rect -4468 32254 -4466 32306
rect -4466 32254 -4414 32306
rect -4414 32254 -4412 32306
rect -4468 32252 -4412 32254
rect -4308 32306 -4252 32308
rect -4308 32254 -4306 32306
rect -4306 32254 -4254 32306
rect -4254 32254 -4252 32306
rect -4308 32252 -4252 32254
rect -4148 32306 -4092 32308
rect -4148 32254 -4146 32306
rect -4146 32254 -4094 32306
rect -4094 32254 -4092 32306
rect -4148 32252 -4092 32254
rect -3988 32306 -3932 32308
rect -3988 32254 -3986 32306
rect -3986 32254 -3934 32306
rect -3934 32254 -3932 32306
rect -3988 32252 -3932 32254
rect -3668 32306 -3612 32308
rect -3668 32254 -3666 32306
rect -3666 32254 -3614 32306
rect -3614 32254 -3612 32306
rect -3668 32252 -3612 32254
rect -3508 32306 -3452 32308
rect -3508 32254 -3506 32306
rect -3506 32254 -3454 32306
rect -3454 32254 -3452 32306
rect -3508 32252 -3452 32254
rect -3348 32306 -3292 32308
rect -3348 32254 -3346 32306
rect -3346 32254 -3294 32306
rect -3294 32254 -3292 32306
rect -3348 32252 -3292 32254
rect -3188 32306 -3132 32308
rect -3188 32254 -3186 32306
rect -3186 32254 -3134 32306
rect -3134 32254 -3132 32306
rect -3188 32252 -3132 32254
rect -3028 32306 -2972 32308
rect -3028 32254 -3026 32306
rect -3026 32254 -2974 32306
rect -2974 32254 -2972 32306
rect -3028 32252 -2972 32254
rect -2868 32306 -2812 32308
rect -2868 32254 -2866 32306
rect -2866 32254 -2814 32306
rect -2814 32254 -2812 32306
rect -2868 32252 -2812 32254
rect -2708 32306 -2652 32308
rect -2708 32254 -2706 32306
rect -2706 32254 -2654 32306
rect -2654 32254 -2652 32306
rect -2708 32252 -2652 32254
rect -2388 32306 -2332 32308
rect -2388 32254 -2386 32306
rect -2386 32254 -2334 32306
rect -2334 32254 -2332 32306
rect -2388 32252 -2332 32254
rect -2068 32306 -2012 32308
rect -2068 32254 -2066 32306
rect -2066 32254 -2014 32306
rect -2014 32254 -2012 32306
rect -2068 32252 -2012 32254
rect -1748 32306 -1692 32308
rect -1748 32254 -1746 32306
rect -1746 32254 -1694 32306
rect -1694 32254 -1692 32306
rect -1748 32252 -1692 32254
rect -1428 32306 -1372 32308
rect -1428 32254 -1426 32306
rect -1426 32254 -1374 32306
rect -1374 32254 -1372 32306
rect -1428 32252 -1372 32254
rect -1108 32306 -1052 32308
rect -1108 32254 -1106 32306
rect -1106 32254 -1054 32306
rect -1054 32254 -1052 32306
rect -1108 32252 -1052 32254
rect -31028 32092 -30972 32148
rect -30708 32092 -30652 32148
rect -30548 32092 -30492 32148
rect -11028 32092 -10972 32148
rect -2228 32092 -2172 32148
rect -31028 31932 -30972 31988
rect -30708 31932 -30652 31988
rect -30388 31932 -30332 31988
rect -30068 31932 -30012 31988
rect -29908 31986 -29852 31988
rect -29908 31934 -29906 31986
rect -29906 31934 -29854 31986
rect -29854 31934 -29852 31986
rect -29908 31932 -29852 31934
rect -29748 31986 -29692 31988
rect -29748 31934 -29746 31986
rect -29746 31934 -29694 31986
rect -29694 31934 -29692 31986
rect -29748 31932 -29692 31934
rect -29588 31986 -29532 31988
rect -29588 31934 -29586 31986
rect -29586 31934 -29534 31986
rect -29534 31934 -29532 31986
rect -29588 31932 -29532 31934
rect -29428 31986 -29372 31988
rect -29428 31934 -29426 31986
rect -29426 31934 -29374 31986
rect -29374 31934 -29372 31986
rect -29428 31932 -29372 31934
rect -29268 31986 -29212 31988
rect -29268 31934 -29266 31986
rect -29266 31934 -29214 31986
rect -29214 31934 -29212 31986
rect -29268 31932 -29212 31934
rect -29108 31986 -29052 31988
rect -29108 31934 -29106 31986
rect -29106 31934 -29054 31986
rect -29054 31934 -29052 31986
rect -29108 31932 -29052 31934
rect -28948 31986 -28892 31988
rect -28948 31934 -28946 31986
rect -28946 31934 -28894 31986
rect -28894 31934 -28892 31986
rect -28948 31932 -28892 31934
rect -28788 31986 -28732 31988
rect -28788 31934 -28786 31986
rect -28786 31934 -28734 31986
rect -28734 31934 -28732 31986
rect -28788 31932 -28732 31934
rect -28628 31986 -28572 31988
rect -28628 31934 -28626 31986
rect -28626 31934 -28574 31986
rect -28574 31934 -28572 31986
rect -28628 31932 -28572 31934
rect -28468 31986 -28412 31988
rect -28468 31934 -28466 31986
rect -28466 31934 -28414 31986
rect -28414 31934 -28412 31986
rect -28468 31932 -28412 31934
rect -28308 31986 -28252 31988
rect -28308 31934 -28306 31986
rect -28306 31934 -28254 31986
rect -28254 31934 -28252 31986
rect -28308 31932 -28252 31934
rect -28148 31986 -28092 31988
rect -28148 31934 -28146 31986
rect -28146 31934 -28094 31986
rect -28094 31934 -28092 31986
rect -28148 31932 -28092 31934
rect -27988 31986 -27932 31988
rect -27988 31934 -27986 31986
rect -27986 31934 -27934 31986
rect -27934 31934 -27932 31986
rect -27988 31932 -27932 31934
rect -27828 31986 -27772 31988
rect -27828 31934 -27826 31986
rect -27826 31934 -27774 31986
rect -27774 31934 -27772 31986
rect -27828 31932 -27772 31934
rect -27668 31986 -27612 31988
rect -27668 31934 -27666 31986
rect -27666 31934 -27614 31986
rect -27614 31934 -27612 31986
rect -27668 31932 -27612 31934
rect -27508 31986 -27452 31988
rect -27508 31934 -27506 31986
rect -27506 31934 -27454 31986
rect -27454 31934 -27452 31986
rect -27508 31932 -27452 31934
rect -27348 31986 -27292 31988
rect -27348 31934 -27346 31986
rect -27346 31934 -27294 31986
rect -27294 31934 -27292 31986
rect -27348 31932 -27292 31934
rect -27188 31986 -27132 31988
rect -27188 31934 -27186 31986
rect -27186 31934 -27134 31986
rect -27134 31934 -27132 31986
rect -27188 31932 -27132 31934
rect -27028 31986 -26972 31988
rect -27028 31934 -27026 31986
rect -27026 31934 -26974 31986
rect -26974 31934 -26972 31986
rect -27028 31932 -26972 31934
rect -26868 31986 -26812 31988
rect -26868 31934 -26866 31986
rect -26866 31934 -26814 31986
rect -26814 31934 -26812 31986
rect -26868 31932 -26812 31934
rect -26708 31986 -26652 31988
rect -26708 31934 -26706 31986
rect -26706 31934 -26654 31986
rect -26654 31934 -26652 31986
rect -26708 31932 -26652 31934
rect -26548 31986 -26492 31988
rect -26548 31934 -26546 31986
rect -26546 31934 -26494 31986
rect -26494 31934 -26492 31986
rect -26548 31932 -26492 31934
rect -26388 31986 -26332 31988
rect -26388 31934 -26386 31986
rect -26386 31934 -26334 31986
rect -26334 31934 -26332 31986
rect -26388 31932 -26332 31934
rect -26228 31986 -26172 31988
rect -26228 31934 -26226 31986
rect -26226 31934 -26174 31986
rect -26174 31934 -26172 31986
rect -26228 31932 -26172 31934
rect -26068 31986 -26012 31988
rect -26068 31934 -26066 31986
rect -26066 31934 -26014 31986
rect -26014 31934 -26012 31986
rect -26068 31932 -26012 31934
rect -25908 31986 -25852 31988
rect -25908 31934 -25906 31986
rect -25906 31934 -25854 31986
rect -25854 31934 -25852 31986
rect -25908 31932 -25852 31934
rect -25748 31986 -25692 31988
rect -25748 31934 -25746 31986
rect -25746 31934 -25694 31986
rect -25694 31934 -25692 31986
rect -25748 31932 -25692 31934
rect -25588 31986 -25532 31988
rect -25588 31934 -25586 31986
rect -25586 31934 -25534 31986
rect -25534 31934 -25532 31986
rect -25588 31932 -25532 31934
rect -25428 31986 -25372 31988
rect -25428 31934 -25426 31986
rect -25426 31934 -25374 31986
rect -25374 31934 -25372 31986
rect -25428 31932 -25372 31934
rect -25268 31986 -25212 31988
rect -25268 31934 -25266 31986
rect -25266 31934 -25214 31986
rect -25214 31934 -25212 31986
rect -25268 31932 -25212 31934
rect -25108 31986 -25052 31988
rect -25108 31934 -25106 31986
rect -25106 31934 -25054 31986
rect -25054 31934 -25052 31986
rect -25108 31932 -25052 31934
rect -24948 31986 -24892 31988
rect -24948 31934 -24946 31986
rect -24946 31934 -24894 31986
rect -24894 31934 -24892 31986
rect -24948 31932 -24892 31934
rect -24788 31986 -24732 31988
rect -24788 31934 -24786 31986
rect -24786 31934 -24734 31986
rect -24734 31934 -24732 31986
rect -24788 31932 -24732 31934
rect -24628 31986 -24572 31988
rect -24628 31934 -24626 31986
rect -24626 31934 -24574 31986
rect -24574 31934 -24572 31986
rect -24628 31932 -24572 31934
rect -24468 31986 -24412 31988
rect -24468 31934 -24466 31986
rect -24466 31934 -24414 31986
rect -24414 31934 -24412 31986
rect -24468 31932 -24412 31934
rect -24308 31986 -24252 31988
rect -24308 31934 -24306 31986
rect -24306 31934 -24254 31986
rect -24254 31934 -24252 31986
rect -24308 31932 -24252 31934
rect -24148 31986 -24092 31988
rect -24148 31934 -24146 31986
rect -24146 31934 -24094 31986
rect -24094 31934 -24092 31986
rect -24148 31932 -24092 31934
rect -23988 31986 -23932 31988
rect -23988 31934 -23986 31986
rect -23986 31934 -23934 31986
rect -23934 31934 -23932 31986
rect -23988 31932 -23932 31934
rect -23828 31986 -23772 31988
rect -23828 31934 -23826 31986
rect -23826 31934 -23774 31986
rect -23774 31934 -23772 31986
rect -23828 31932 -23772 31934
rect -23668 31986 -23612 31988
rect -23668 31934 -23666 31986
rect -23666 31934 -23614 31986
rect -23614 31934 -23612 31986
rect -23668 31932 -23612 31934
rect -23508 31986 -23452 31988
rect -23508 31934 -23506 31986
rect -23506 31934 -23454 31986
rect -23454 31934 -23452 31986
rect -23508 31932 -23452 31934
rect -23348 31986 -23292 31988
rect -23348 31934 -23346 31986
rect -23346 31934 -23294 31986
rect -23294 31934 -23292 31986
rect -23348 31932 -23292 31934
rect -23188 31986 -23132 31988
rect -23188 31934 -23186 31986
rect -23186 31934 -23134 31986
rect -23134 31934 -23132 31986
rect -23188 31932 -23132 31934
rect -23028 31986 -22972 31988
rect -23028 31934 -23026 31986
rect -23026 31934 -22974 31986
rect -22974 31934 -22972 31986
rect -23028 31932 -22972 31934
rect -22868 31986 -22812 31988
rect -22868 31934 -22866 31986
rect -22866 31934 -22814 31986
rect -22814 31934 -22812 31986
rect -22868 31932 -22812 31934
rect -22708 31986 -22652 31988
rect -22708 31934 -22706 31986
rect -22706 31934 -22654 31986
rect -22654 31934 -22652 31986
rect -22708 31932 -22652 31934
rect -22548 31986 -22492 31988
rect -22548 31934 -22546 31986
rect -22546 31934 -22494 31986
rect -22494 31934 -22492 31986
rect -22548 31932 -22492 31934
rect -22388 31986 -22332 31988
rect -22388 31934 -22386 31986
rect -22386 31934 -22334 31986
rect -22334 31934 -22332 31986
rect -22388 31932 -22332 31934
rect -22228 31986 -22172 31988
rect -22228 31934 -22226 31986
rect -22226 31934 -22174 31986
rect -22174 31934 -22172 31986
rect -22228 31932 -22172 31934
rect -22068 31986 -22012 31988
rect -22068 31934 -22066 31986
rect -22066 31934 -22014 31986
rect -22014 31934 -22012 31986
rect -22068 31932 -22012 31934
rect -21908 31986 -21852 31988
rect -21908 31934 -21906 31986
rect -21906 31934 -21854 31986
rect -21854 31934 -21852 31986
rect -21908 31932 -21852 31934
rect -21748 31986 -21692 31988
rect -21748 31934 -21746 31986
rect -21746 31934 -21694 31986
rect -21694 31934 -21692 31986
rect -21748 31932 -21692 31934
rect -21588 31986 -21532 31988
rect -21588 31934 -21586 31986
rect -21586 31934 -21534 31986
rect -21534 31934 -21532 31986
rect -21588 31932 -21532 31934
rect -21428 31986 -21372 31988
rect -21428 31934 -21426 31986
rect -21426 31934 -21374 31986
rect -21374 31934 -21372 31986
rect -21428 31932 -21372 31934
rect -21268 31986 -21212 31988
rect -21268 31934 -21266 31986
rect -21266 31934 -21214 31986
rect -21214 31934 -21212 31986
rect -21268 31932 -21212 31934
rect -21108 31986 -21052 31988
rect -21108 31934 -21106 31986
rect -21106 31934 -21054 31986
rect -21054 31934 -21052 31986
rect -21108 31932 -21052 31934
rect -20948 31986 -20892 31988
rect -20948 31934 -20946 31986
rect -20946 31934 -20894 31986
rect -20894 31934 -20892 31986
rect -20948 31932 -20892 31934
rect -20788 31986 -20732 31988
rect -20788 31934 -20786 31986
rect -20786 31934 -20734 31986
rect -20734 31934 -20732 31986
rect -20788 31932 -20732 31934
rect -20628 31986 -20572 31988
rect -20628 31934 -20626 31986
rect -20626 31934 -20574 31986
rect -20574 31934 -20572 31986
rect -20628 31932 -20572 31934
rect -20468 31986 -20412 31988
rect -20468 31934 -20466 31986
rect -20466 31934 -20414 31986
rect -20414 31934 -20412 31986
rect -20468 31932 -20412 31934
rect -20308 31986 -20252 31988
rect -20308 31934 -20306 31986
rect -20306 31934 -20254 31986
rect -20254 31934 -20252 31986
rect -20308 31932 -20252 31934
rect -20148 31986 -20092 31988
rect -20148 31934 -20146 31986
rect -20146 31934 -20094 31986
rect -20094 31934 -20092 31986
rect -20148 31932 -20092 31934
rect -19988 31986 -19932 31988
rect -19988 31934 -19986 31986
rect -19986 31934 -19934 31986
rect -19934 31934 -19932 31986
rect -19988 31932 -19932 31934
rect -19828 31986 -19772 31988
rect -19828 31934 -19826 31986
rect -19826 31934 -19774 31986
rect -19774 31934 -19772 31986
rect -19828 31932 -19772 31934
rect -19668 31986 -19612 31988
rect -19668 31934 -19666 31986
rect -19666 31934 -19614 31986
rect -19614 31934 -19612 31986
rect -19668 31932 -19612 31934
rect -19508 31986 -19452 31988
rect -19508 31934 -19506 31986
rect -19506 31934 -19454 31986
rect -19454 31934 -19452 31986
rect -19508 31932 -19452 31934
rect -19348 31986 -19292 31988
rect -19348 31934 -19346 31986
rect -19346 31934 -19294 31986
rect -19294 31934 -19292 31986
rect -19348 31932 -19292 31934
rect -19188 31986 -19132 31988
rect -19188 31934 -19186 31986
rect -19186 31934 -19134 31986
rect -19134 31934 -19132 31986
rect -19188 31932 -19132 31934
rect -19028 31986 -18972 31988
rect -19028 31934 -19026 31986
rect -19026 31934 -18974 31986
rect -18974 31934 -18972 31986
rect -19028 31932 -18972 31934
rect -18868 31986 -18812 31988
rect -18868 31934 -18866 31986
rect -18866 31934 -18814 31986
rect -18814 31934 -18812 31986
rect -18868 31932 -18812 31934
rect -18708 31986 -18652 31988
rect -18708 31934 -18706 31986
rect -18706 31934 -18654 31986
rect -18654 31934 -18652 31986
rect -18708 31932 -18652 31934
rect -18548 31986 -18492 31988
rect -18548 31934 -18546 31986
rect -18546 31934 -18494 31986
rect -18494 31934 -18492 31986
rect -18548 31932 -18492 31934
rect -18388 31986 -18332 31988
rect -18388 31934 -18386 31986
rect -18386 31934 -18334 31986
rect -18334 31934 -18332 31986
rect -18388 31932 -18332 31934
rect -18228 31986 -18172 31988
rect -18228 31934 -18226 31986
rect -18226 31934 -18174 31986
rect -18174 31934 -18172 31986
rect -18228 31932 -18172 31934
rect -18068 31986 -18012 31988
rect -18068 31934 -18066 31986
rect -18066 31934 -18014 31986
rect -18014 31934 -18012 31986
rect -18068 31932 -18012 31934
rect -17908 31986 -17852 31988
rect -17908 31934 -17906 31986
rect -17906 31934 -17854 31986
rect -17854 31934 -17852 31986
rect -17908 31932 -17852 31934
rect -17748 31986 -17692 31988
rect -17748 31934 -17746 31986
rect -17746 31934 -17694 31986
rect -17694 31934 -17692 31986
rect -17748 31932 -17692 31934
rect -17588 31986 -17532 31988
rect -17588 31934 -17586 31986
rect -17586 31934 -17534 31986
rect -17534 31934 -17532 31986
rect -17588 31932 -17532 31934
rect -17428 31986 -17372 31988
rect -17428 31934 -17426 31986
rect -17426 31934 -17374 31986
rect -17374 31934 -17372 31986
rect -17428 31932 -17372 31934
rect -17268 31986 -17212 31988
rect -17268 31934 -17266 31986
rect -17266 31934 -17214 31986
rect -17214 31934 -17212 31986
rect -17268 31932 -17212 31934
rect -17108 31986 -17052 31988
rect -17108 31934 -17106 31986
rect -17106 31934 -17054 31986
rect -17054 31934 -17052 31986
rect -17108 31932 -17052 31934
rect -16948 31986 -16892 31988
rect -16948 31934 -16946 31986
rect -16946 31934 -16894 31986
rect -16894 31934 -16892 31986
rect -16948 31932 -16892 31934
rect -16788 31986 -16732 31988
rect -16788 31934 -16786 31986
rect -16786 31934 -16734 31986
rect -16734 31934 -16732 31986
rect -16788 31932 -16732 31934
rect -16628 31986 -16572 31988
rect -16628 31934 -16626 31986
rect -16626 31934 -16574 31986
rect -16574 31934 -16572 31986
rect -16628 31932 -16572 31934
rect -16468 31986 -16412 31988
rect -16468 31934 -16466 31986
rect -16466 31934 -16414 31986
rect -16414 31934 -16412 31986
rect -16468 31932 -16412 31934
rect -16308 31986 -16252 31988
rect -16308 31934 -16306 31986
rect -16306 31934 -16254 31986
rect -16254 31934 -16252 31986
rect -16308 31932 -16252 31934
rect -16148 31986 -16092 31988
rect -16148 31934 -16146 31986
rect -16146 31934 -16094 31986
rect -16094 31934 -16092 31986
rect -16148 31932 -16092 31934
rect -15988 31986 -15932 31988
rect -15988 31934 -15986 31986
rect -15986 31934 -15934 31986
rect -15934 31934 -15932 31986
rect -15988 31932 -15932 31934
rect -15828 31986 -15772 31988
rect -15828 31934 -15826 31986
rect -15826 31934 -15774 31986
rect -15774 31934 -15772 31986
rect -15828 31932 -15772 31934
rect -15668 31986 -15612 31988
rect -15668 31934 -15666 31986
rect -15666 31934 -15614 31986
rect -15614 31934 -15612 31986
rect -15668 31932 -15612 31934
rect -15508 31986 -15452 31988
rect -15508 31934 -15506 31986
rect -15506 31934 -15454 31986
rect -15454 31934 -15452 31986
rect -15508 31932 -15452 31934
rect -15348 31986 -15292 31988
rect -15348 31934 -15346 31986
rect -15346 31934 -15294 31986
rect -15294 31934 -15292 31986
rect -15348 31932 -15292 31934
rect -15188 31986 -15132 31988
rect -15188 31934 -15186 31986
rect -15186 31934 -15134 31986
rect -15134 31934 -15132 31986
rect -15188 31932 -15132 31934
rect -15028 31986 -14972 31988
rect -15028 31934 -15026 31986
rect -15026 31934 -14974 31986
rect -14974 31934 -14972 31986
rect -15028 31932 -14972 31934
rect -14868 31986 -14812 31988
rect -14868 31934 -14866 31986
rect -14866 31934 -14814 31986
rect -14814 31934 -14812 31986
rect -14868 31932 -14812 31934
rect -14708 31986 -14652 31988
rect -14708 31934 -14706 31986
rect -14706 31934 -14654 31986
rect -14654 31934 -14652 31986
rect -14708 31932 -14652 31934
rect -14548 31986 -14492 31988
rect -14548 31934 -14546 31986
rect -14546 31934 -14494 31986
rect -14494 31934 -14492 31986
rect -14548 31932 -14492 31934
rect -14388 31986 -14332 31988
rect -14388 31934 -14386 31986
rect -14386 31934 -14334 31986
rect -14334 31934 -14332 31986
rect -14388 31932 -14332 31934
rect -14228 31986 -14172 31988
rect -14228 31934 -14226 31986
rect -14226 31934 -14174 31986
rect -14174 31934 -14172 31986
rect -14228 31932 -14172 31934
rect -14068 31986 -14012 31988
rect -14068 31934 -14066 31986
rect -14066 31934 -14014 31986
rect -14014 31934 -14012 31986
rect -14068 31932 -14012 31934
rect -13908 31986 -13852 31988
rect -13908 31934 -13906 31986
rect -13906 31934 -13854 31986
rect -13854 31934 -13852 31986
rect -13908 31932 -13852 31934
rect -13748 31986 -13692 31988
rect -13748 31934 -13746 31986
rect -13746 31934 -13694 31986
rect -13694 31934 -13692 31986
rect -13748 31932 -13692 31934
rect -13588 31986 -13532 31988
rect -13588 31934 -13586 31986
rect -13586 31934 -13534 31986
rect -13534 31934 -13532 31986
rect -13588 31932 -13532 31934
rect -13428 31986 -13372 31988
rect -13428 31934 -13426 31986
rect -13426 31934 -13374 31986
rect -13374 31934 -13372 31986
rect -13428 31932 -13372 31934
rect -13268 31986 -13212 31988
rect -13268 31934 -13266 31986
rect -13266 31934 -13214 31986
rect -13214 31934 -13212 31986
rect -13268 31932 -13212 31934
rect -13108 31986 -13052 31988
rect -13108 31934 -13106 31986
rect -13106 31934 -13054 31986
rect -13054 31934 -13052 31986
rect -13108 31932 -13052 31934
rect -12948 31986 -12892 31988
rect -12948 31934 -12946 31986
rect -12946 31934 -12894 31986
rect -12894 31934 -12892 31986
rect -12948 31932 -12892 31934
rect -12788 31986 -12732 31988
rect -12788 31934 -12786 31986
rect -12786 31934 -12734 31986
rect -12734 31934 -12732 31986
rect -12788 31932 -12732 31934
rect -12628 31986 -12572 31988
rect -12628 31934 -12626 31986
rect -12626 31934 -12574 31986
rect -12574 31934 -12572 31986
rect -12628 31932 -12572 31934
rect -12468 31986 -12412 31988
rect -12468 31934 -12466 31986
rect -12466 31934 -12414 31986
rect -12414 31934 -12412 31986
rect -12468 31932 -12412 31934
rect -12308 31986 -12252 31988
rect -12308 31934 -12306 31986
rect -12306 31934 -12254 31986
rect -12254 31934 -12252 31986
rect -12308 31932 -12252 31934
rect -12148 31986 -12092 31988
rect -12148 31934 -12146 31986
rect -12146 31934 -12094 31986
rect -12094 31934 -12092 31986
rect -12148 31932 -12092 31934
rect -11988 31986 -11932 31988
rect -11988 31934 -11986 31986
rect -11986 31934 -11934 31986
rect -11934 31934 -11932 31986
rect -11988 31932 -11932 31934
rect -11828 31986 -11772 31988
rect -11828 31934 -11826 31986
rect -11826 31934 -11774 31986
rect -11774 31934 -11772 31986
rect -11828 31932 -11772 31934
rect -11668 31986 -11612 31988
rect -11668 31934 -11666 31986
rect -11666 31934 -11614 31986
rect -11614 31934 -11612 31986
rect -11668 31932 -11612 31934
rect -11508 31986 -11452 31988
rect -11508 31934 -11506 31986
rect -11506 31934 -11454 31986
rect -11454 31934 -11452 31986
rect -11508 31932 -11452 31934
rect -11348 31986 -11292 31988
rect -11348 31934 -11346 31986
rect -11346 31934 -11294 31986
rect -11294 31934 -11292 31986
rect -11348 31932 -11292 31934
rect -11188 31986 -11132 31988
rect -11188 31934 -11186 31986
rect -11186 31934 -11134 31986
rect -11134 31934 -11132 31986
rect -11188 31932 -11132 31934
rect -10868 31986 -10812 31988
rect -10868 31934 -10866 31986
rect -10866 31934 -10814 31986
rect -10814 31934 -10812 31986
rect -10868 31932 -10812 31934
rect -10708 31986 -10652 31988
rect -10708 31934 -10706 31986
rect -10706 31934 -10654 31986
rect -10654 31934 -10652 31986
rect -10708 31932 -10652 31934
rect -10548 31986 -10492 31988
rect -10548 31934 -10546 31986
rect -10546 31934 -10494 31986
rect -10494 31934 -10492 31986
rect -10548 31932 -10492 31934
rect -10388 31986 -10332 31988
rect -10388 31934 -10386 31986
rect -10386 31934 -10334 31986
rect -10334 31934 -10332 31986
rect -10388 31932 -10332 31934
rect -10228 31986 -10172 31988
rect -10228 31934 -10226 31986
rect -10226 31934 -10174 31986
rect -10174 31934 -10172 31986
rect -10228 31932 -10172 31934
rect -10068 31986 -10012 31988
rect -10068 31934 -10066 31986
rect -10066 31934 -10014 31986
rect -10014 31934 -10012 31986
rect -10068 31932 -10012 31934
rect -9908 31986 -9852 31988
rect -9908 31934 -9906 31986
rect -9906 31934 -9854 31986
rect -9854 31934 -9852 31986
rect -9908 31932 -9852 31934
rect -9748 31986 -9692 31988
rect -9748 31934 -9746 31986
rect -9746 31934 -9694 31986
rect -9694 31934 -9692 31986
rect -9748 31932 -9692 31934
rect -9588 31986 -9532 31988
rect -9588 31934 -9586 31986
rect -9586 31934 -9534 31986
rect -9534 31934 -9532 31986
rect -9588 31932 -9532 31934
rect -9428 31986 -9372 31988
rect -9428 31934 -9426 31986
rect -9426 31934 -9374 31986
rect -9374 31934 -9372 31986
rect -9428 31932 -9372 31934
rect -9268 31986 -9212 31988
rect -9268 31934 -9266 31986
rect -9266 31934 -9214 31986
rect -9214 31934 -9212 31986
rect -9268 31932 -9212 31934
rect -9108 31986 -9052 31988
rect -9108 31934 -9106 31986
rect -9106 31934 -9054 31986
rect -9054 31934 -9052 31986
rect -9108 31932 -9052 31934
rect -8948 31986 -8892 31988
rect -8948 31934 -8946 31986
rect -8946 31934 -8894 31986
rect -8894 31934 -8892 31986
rect -8948 31932 -8892 31934
rect -8788 31986 -8732 31988
rect -8788 31934 -8786 31986
rect -8786 31934 -8734 31986
rect -8734 31934 -8732 31986
rect -8788 31932 -8732 31934
rect -8628 31986 -8572 31988
rect -8628 31934 -8626 31986
rect -8626 31934 -8574 31986
rect -8574 31934 -8572 31986
rect -8628 31932 -8572 31934
rect -8468 31986 -8412 31988
rect -8468 31934 -8466 31986
rect -8466 31934 -8414 31986
rect -8414 31934 -8412 31986
rect -8468 31932 -8412 31934
rect -8308 31986 -8252 31988
rect -8308 31934 -8306 31986
rect -8306 31934 -8254 31986
rect -8254 31934 -8252 31986
rect -8308 31932 -8252 31934
rect -8148 31986 -8092 31988
rect -8148 31934 -8146 31986
rect -8146 31934 -8094 31986
rect -8094 31934 -8092 31986
rect -8148 31932 -8092 31934
rect -7988 31986 -7932 31988
rect -7988 31934 -7986 31986
rect -7986 31934 -7934 31986
rect -7934 31934 -7932 31986
rect -7988 31932 -7932 31934
rect -7828 31986 -7772 31988
rect -7828 31934 -7826 31986
rect -7826 31934 -7774 31986
rect -7774 31934 -7772 31986
rect -7828 31932 -7772 31934
rect -7668 31986 -7612 31988
rect -7668 31934 -7666 31986
rect -7666 31934 -7614 31986
rect -7614 31934 -7612 31986
rect -7668 31932 -7612 31934
rect -7508 31986 -7452 31988
rect -7508 31934 -7506 31986
rect -7506 31934 -7454 31986
rect -7454 31934 -7452 31986
rect -7508 31932 -7452 31934
rect -7348 31986 -7292 31988
rect -7348 31934 -7346 31986
rect -7346 31934 -7294 31986
rect -7294 31934 -7292 31986
rect -7348 31932 -7292 31934
rect -7188 31986 -7132 31988
rect -7188 31934 -7186 31986
rect -7186 31934 -7134 31986
rect -7134 31934 -7132 31986
rect -7188 31932 -7132 31934
rect -7028 31986 -6972 31988
rect -7028 31934 -7026 31986
rect -7026 31934 -6974 31986
rect -6974 31934 -6972 31986
rect -7028 31932 -6972 31934
rect -6868 31986 -6812 31988
rect -6868 31934 -6866 31986
rect -6866 31934 -6814 31986
rect -6814 31934 -6812 31986
rect -6868 31932 -6812 31934
rect -6708 31986 -6652 31988
rect -6708 31934 -6706 31986
rect -6706 31934 -6654 31986
rect -6654 31934 -6652 31986
rect -6708 31932 -6652 31934
rect -6548 31986 -6492 31988
rect -6548 31934 -6546 31986
rect -6546 31934 -6494 31986
rect -6494 31934 -6492 31986
rect -6548 31932 -6492 31934
rect -6388 31986 -6332 31988
rect -6388 31934 -6386 31986
rect -6386 31934 -6334 31986
rect -6334 31934 -6332 31986
rect -6388 31932 -6332 31934
rect -6228 31986 -6172 31988
rect -6228 31934 -6226 31986
rect -6226 31934 -6174 31986
rect -6174 31934 -6172 31986
rect -6228 31932 -6172 31934
rect -6068 31986 -6012 31988
rect -6068 31934 -6066 31986
rect -6066 31934 -6014 31986
rect -6014 31934 -6012 31986
rect -6068 31932 -6012 31934
rect -5908 31986 -5852 31988
rect -5908 31934 -5906 31986
rect -5906 31934 -5854 31986
rect -5854 31934 -5852 31986
rect -5908 31932 -5852 31934
rect -5748 31986 -5692 31988
rect -5748 31934 -5746 31986
rect -5746 31934 -5694 31986
rect -5694 31934 -5692 31986
rect -5748 31932 -5692 31934
rect -5588 31986 -5532 31988
rect -5588 31934 -5586 31986
rect -5586 31934 -5534 31986
rect -5534 31934 -5532 31986
rect -5588 31932 -5532 31934
rect -5428 31986 -5372 31988
rect -5428 31934 -5426 31986
rect -5426 31934 -5374 31986
rect -5374 31934 -5372 31986
rect -5428 31932 -5372 31934
rect -5268 31986 -5212 31988
rect -5268 31934 -5266 31986
rect -5266 31934 -5214 31986
rect -5214 31934 -5212 31986
rect -5268 31932 -5212 31934
rect -5108 31986 -5052 31988
rect -5108 31934 -5106 31986
rect -5106 31934 -5054 31986
rect -5054 31934 -5052 31986
rect -5108 31932 -5052 31934
rect -4948 31986 -4892 31988
rect -4948 31934 -4946 31986
rect -4946 31934 -4894 31986
rect -4894 31934 -4892 31986
rect -4948 31932 -4892 31934
rect -4788 31986 -4732 31988
rect -4788 31934 -4786 31986
rect -4786 31934 -4734 31986
rect -4734 31934 -4732 31986
rect -4788 31932 -4732 31934
rect -4628 31986 -4572 31988
rect -4628 31934 -4626 31986
rect -4626 31934 -4574 31986
rect -4574 31934 -4572 31986
rect -4628 31932 -4572 31934
rect -4468 31986 -4412 31988
rect -4468 31934 -4466 31986
rect -4466 31934 -4414 31986
rect -4414 31934 -4412 31986
rect -4468 31932 -4412 31934
rect -4308 31986 -4252 31988
rect -4308 31934 -4306 31986
rect -4306 31934 -4254 31986
rect -4254 31934 -4252 31986
rect -4308 31932 -4252 31934
rect -4148 31986 -4092 31988
rect -4148 31934 -4146 31986
rect -4146 31934 -4094 31986
rect -4094 31934 -4092 31986
rect -4148 31932 -4092 31934
rect -3988 31986 -3932 31988
rect -3988 31934 -3986 31986
rect -3986 31934 -3934 31986
rect -3934 31934 -3932 31986
rect -3988 31932 -3932 31934
rect -3668 31986 -3612 31988
rect -3668 31934 -3666 31986
rect -3666 31934 -3614 31986
rect -3614 31934 -3612 31986
rect -3668 31932 -3612 31934
rect -3508 31986 -3452 31988
rect -3508 31934 -3506 31986
rect -3506 31934 -3454 31986
rect -3454 31934 -3452 31986
rect -3508 31932 -3452 31934
rect -3348 31986 -3292 31988
rect -3348 31934 -3346 31986
rect -3346 31934 -3294 31986
rect -3294 31934 -3292 31986
rect -3348 31932 -3292 31934
rect -3188 31986 -3132 31988
rect -3188 31934 -3186 31986
rect -3186 31934 -3134 31986
rect -3134 31934 -3132 31986
rect -3188 31932 -3132 31934
rect -3028 31986 -2972 31988
rect -3028 31934 -3026 31986
rect -3026 31934 -2974 31986
rect -2974 31934 -2972 31986
rect -3028 31932 -2972 31934
rect -2868 31986 -2812 31988
rect -2868 31934 -2866 31986
rect -2866 31934 -2814 31986
rect -2814 31934 -2812 31986
rect -2868 31932 -2812 31934
rect -2708 31986 -2652 31988
rect -2708 31934 -2706 31986
rect -2706 31934 -2654 31986
rect -2654 31934 -2652 31986
rect -2708 31932 -2652 31934
rect -2388 31986 -2332 31988
rect -2388 31934 -2386 31986
rect -2386 31934 -2334 31986
rect -2334 31934 -2332 31986
rect -2388 31932 -2332 31934
rect -2068 31986 -2012 31988
rect -2068 31934 -2066 31986
rect -2066 31934 -2014 31986
rect -2014 31934 -2012 31986
rect -2068 31932 -2012 31934
rect -1748 31986 -1692 31988
rect -1748 31934 -1746 31986
rect -1746 31934 -1694 31986
rect -1694 31934 -1692 31986
rect -1748 31932 -1692 31934
rect -1428 31986 -1372 31988
rect -1428 31934 -1426 31986
rect -1426 31934 -1374 31986
rect -1374 31934 -1372 31986
rect -1428 31932 -1372 31934
rect -1108 31986 -1052 31988
rect -1108 31934 -1106 31986
rect -1106 31934 -1054 31986
rect -1054 31934 -1052 31986
rect -1108 31932 -1052 31934
<< metal3 >>
rect -31040 42868 -30960 42960
rect -31040 42812 -31028 42868
rect -30972 42812 -30960 42868
rect -31040 42708 -30960 42812
rect -31040 42652 -31028 42708
rect -30972 42652 -30960 42708
rect -31040 42548 -30960 42652
rect -31040 42492 -31028 42548
rect -30972 42492 -30960 42548
rect -31040 42388 -30960 42492
rect -31040 42332 -31028 42388
rect -30972 42332 -30960 42388
rect -31040 42228 -30960 42332
rect -31040 42172 -31028 42228
rect -30972 42172 -30960 42228
rect -31040 42068 -30960 42172
rect -31040 42012 -31028 42068
rect -30972 42012 -30960 42068
rect -31040 41908 -30960 42012
rect -31040 41852 -31028 41908
rect -30972 41852 -30960 41908
rect -31040 41752 -30960 41852
rect -31040 41688 -31032 41752
rect -30968 41688 -30960 41752
rect -31040 41592 -30960 41688
rect -31040 41528 -31032 41592
rect -30968 41528 -30960 41592
rect -33120 41348 -33040 41360
rect -33120 41292 -33108 41348
rect -33052 41292 -33040 41348
rect -33120 41028 -33040 41292
rect -33120 40972 -33108 41028
rect -33052 40972 -33040 41028
rect -33120 40960 -33040 40972
rect -32960 41348 -32880 41360
rect -32960 41292 -32948 41348
rect -32892 41292 -32880 41348
rect -32960 41028 -32880 41292
rect -32960 40972 -32948 41028
rect -32892 40972 -32880 41028
rect -32960 40960 -32880 40972
rect -32800 41348 -32720 41360
rect -32800 41292 -32788 41348
rect -32732 41292 -32720 41348
rect -32800 41028 -32720 41292
rect -32800 40972 -32788 41028
rect -32732 40972 -32720 41028
rect -32800 40960 -32720 40972
rect -32640 41348 -32560 41360
rect -32640 41292 -32628 41348
rect -32572 41292 -32560 41348
rect -32640 41028 -32560 41292
rect -32640 40972 -32628 41028
rect -32572 40972 -32560 41028
rect -32640 40960 -32560 40972
rect -32480 41348 -32400 41360
rect -32480 41292 -32468 41348
rect -32412 41292 -32400 41348
rect -32480 41028 -32400 41292
rect -32480 40972 -32468 41028
rect -32412 40972 -32400 41028
rect -32480 40960 -32400 40972
rect -32320 41348 -32240 41360
rect -32320 41292 -32308 41348
rect -32252 41292 -32240 41348
rect -32320 41028 -32240 41292
rect -32320 40972 -32308 41028
rect -32252 40972 -32240 41028
rect -32320 40960 -32240 40972
rect -32160 41348 -32080 41360
rect -32160 41292 -32148 41348
rect -32092 41292 -32080 41348
rect -32160 41028 -32080 41292
rect -32160 40972 -32148 41028
rect -32092 40972 -32080 41028
rect -32160 40960 -32080 40972
rect -32000 41348 -31920 41360
rect -32000 41292 -31988 41348
rect -31932 41292 -31920 41348
rect -32000 41028 -31920 41292
rect -32000 40972 -31988 41028
rect -31932 40972 -31920 41028
rect -32000 40960 -31920 40972
rect -31840 41348 -31760 41360
rect -31840 41292 -31828 41348
rect -31772 41292 -31760 41348
rect -31840 41028 -31760 41292
rect -31840 40972 -31828 41028
rect -31772 40972 -31760 41028
rect -31840 40960 -31760 40972
rect -31680 41348 -31600 41360
rect -31680 41292 -31668 41348
rect -31612 41292 -31600 41348
rect -31680 41028 -31600 41292
rect -31680 40972 -31668 41028
rect -31612 40972 -31600 41028
rect -31680 40960 -31600 40972
rect -31520 41348 -31440 41360
rect -31520 41292 -31508 41348
rect -31452 41292 -31440 41348
rect -31520 41028 -31440 41292
rect -31520 40972 -31508 41028
rect -31452 40972 -31440 41028
rect -31520 40960 -31440 40972
rect -31360 41348 -31280 41360
rect -31360 41292 -31348 41348
rect -31292 41292 -31280 41348
rect -31360 41028 -31280 41292
rect -31360 40972 -31348 41028
rect -31292 40972 -31280 41028
rect -31360 40960 -31280 40972
rect -31200 41348 -31120 41360
rect -31200 41292 -31188 41348
rect -31132 41292 -31120 41348
rect -31200 41028 -31120 41292
rect -31200 40972 -31188 41028
rect -31132 40972 -31120 41028
rect -31200 40960 -31120 40972
rect -31040 40792 -30960 41528
rect -31040 40728 -31032 40792
rect -30968 40728 -30960 40792
rect -31040 40632 -30960 40728
rect -31040 40568 -31032 40632
rect -30968 40568 -30960 40632
rect -31040 40472 -30960 40568
rect -31040 40408 -31032 40472
rect -30968 40408 -30960 40472
rect -31040 40312 -30960 40408
rect -31040 40248 -31032 40312
rect -30968 40248 -30960 40312
rect -31040 40152 -30960 40248
rect -31040 40088 -31032 40152
rect -30968 40088 -30960 40152
rect -31040 39992 -30960 40088
rect -31040 39928 -31032 39992
rect -30968 39928 -30960 39992
rect -31040 39832 -30960 39928
rect -31040 39768 -31032 39832
rect -30968 39768 -30960 39832
rect -31040 39672 -30960 39768
rect -31040 39608 -31032 39672
rect -30968 39608 -30960 39672
rect -31040 39512 -30960 39608
rect -31040 39448 -31032 39512
rect -30968 39448 -30960 39512
rect -31040 39352 -30960 39448
rect -31040 39288 -31032 39352
rect -30968 39288 -30960 39352
rect -31040 39192 -30960 39288
rect -31040 39128 -31032 39192
rect -30968 39128 -30960 39192
rect -31040 39032 -30960 39128
rect -31040 38968 -31032 39032
rect -30968 38968 -30960 39032
rect -31040 38872 -30960 38968
rect -31040 38808 -31032 38872
rect -30968 38808 -30960 38872
rect -31040 38712 -30960 38808
rect -31040 38648 -31032 38712
rect -30968 38648 -30960 38712
rect -31040 38552 -30960 38648
rect -31040 38488 -31032 38552
rect -30968 38488 -30960 38552
rect -31040 38392 -30960 38488
rect -31040 38328 -31032 38392
rect -30968 38328 -30960 38392
rect -31040 38232 -30960 38328
rect -31040 38168 -31032 38232
rect -30968 38168 -30960 38232
rect -31040 38072 -30960 38168
rect -31040 38008 -31032 38072
rect -30968 38008 -30960 38072
rect -31040 37912 -30960 38008
rect -31040 37848 -31032 37912
rect -30968 37848 -30960 37912
rect -33120 37748 -33040 37760
rect -33120 37692 -33108 37748
rect -33052 37692 -33040 37748
rect -33120 37428 -33040 37692
rect -33120 37372 -33108 37428
rect -33052 37372 -33040 37428
rect -33120 37108 -33040 37372
rect -33120 37052 -33108 37108
rect -33052 37052 -33040 37108
rect -33120 37040 -33040 37052
rect -32960 37748 -32880 37760
rect -32960 37692 -32948 37748
rect -32892 37692 -32880 37748
rect -32960 37428 -32880 37692
rect -32960 37372 -32948 37428
rect -32892 37372 -32880 37428
rect -32960 37108 -32880 37372
rect -32960 37052 -32948 37108
rect -32892 37052 -32880 37108
rect -32960 37040 -32880 37052
rect -32800 37748 -32720 37760
rect -32800 37692 -32788 37748
rect -32732 37692 -32720 37748
rect -32800 37428 -32720 37692
rect -32800 37372 -32788 37428
rect -32732 37372 -32720 37428
rect -32800 37108 -32720 37372
rect -32800 37052 -32788 37108
rect -32732 37052 -32720 37108
rect -32800 37040 -32720 37052
rect -32640 37748 -32560 37760
rect -32640 37692 -32628 37748
rect -32572 37692 -32560 37748
rect -32640 37428 -32560 37692
rect -32640 37372 -32628 37428
rect -32572 37372 -32560 37428
rect -32640 37108 -32560 37372
rect -32640 37052 -32628 37108
rect -32572 37052 -32560 37108
rect -32640 37040 -32560 37052
rect -32480 37748 -32400 37760
rect -32480 37692 -32468 37748
rect -32412 37692 -32400 37748
rect -32480 37428 -32400 37692
rect -32480 37372 -32468 37428
rect -32412 37372 -32400 37428
rect -32480 37108 -32400 37372
rect -32480 37052 -32468 37108
rect -32412 37052 -32400 37108
rect -32480 37040 -32400 37052
rect -32320 37748 -32240 37760
rect -32320 37692 -32308 37748
rect -32252 37692 -32240 37748
rect -32320 37428 -32240 37692
rect -32320 37372 -32308 37428
rect -32252 37372 -32240 37428
rect -32320 37108 -32240 37372
rect -32320 37052 -32308 37108
rect -32252 37052 -32240 37108
rect -32320 37040 -32240 37052
rect -32160 37748 -32080 37760
rect -32160 37692 -32148 37748
rect -32092 37692 -32080 37748
rect -32160 37428 -32080 37692
rect -32160 37372 -32148 37428
rect -32092 37372 -32080 37428
rect -32160 37108 -32080 37372
rect -32160 37052 -32148 37108
rect -32092 37052 -32080 37108
rect -32160 37040 -32080 37052
rect -32000 37748 -31920 37760
rect -32000 37692 -31988 37748
rect -31932 37692 -31920 37748
rect -32000 37428 -31920 37692
rect -32000 37372 -31988 37428
rect -31932 37372 -31920 37428
rect -32000 37108 -31920 37372
rect -32000 37052 -31988 37108
rect -31932 37052 -31920 37108
rect -32000 37040 -31920 37052
rect -31840 37748 -31760 37760
rect -31840 37692 -31828 37748
rect -31772 37692 -31760 37748
rect -31840 37428 -31760 37692
rect -31840 37372 -31828 37428
rect -31772 37372 -31760 37428
rect -31840 37108 -31760 37372
rect -31840 37052 -31828 37108
rect -31772 37052 -31760 37108
rect -31840 37040 -31760 37052
rect -31680 37748 -31600 37760
rect -31680 37692 -31668 37748
rect -31612 37692 -31600 37748
rect -31680 37428 -31600 37692
rect -31680 37372 -31668 37428
rect -31612 37372 -31600 37428
rect -31680 37108 -31600 37372
rect -31680 37052 -31668 37108
rect -31612 37052 -31600 37108
rect -31680 37040 -31600 37052
rect -31520 37748 -31440 37760
rect -31520 37692 -31508 37748
rect -31452 37692 -31440 37748
rect -31520 37428 -31440 37692
rect -31520 37372 -31508 37428
rect -31452 37372 -31440 37428
rect -31520 37108 -31440 37372
rect -31520 37052 -31508 37108
rect -31452 37052 -31440 37108
rect -31520 37040 -31440 37052
rect -31360 37748 -31280 37760
rect -31360 37692 -31348 37748
rect -31292 37692 -31280 37748
rect -31360 37428 -31280 37692
rect -31360 37372 -31348 37428
rect -31292 37372 -31280 37428
rect -31360 37108 -31280 37372
rect -31360 37052 -31348 37108
rect -31292 37052 -31280 37108
rect -31360 37040 -31280 37052
rect -31200 37748 -31120 37760
rect -31200 37692 -31188 37748
rect -31132 37692 -31120 37748
rect -31200 37428 -31120 37692
rect -31200 37372 -31188 37428
rect -31132 37372 -31120 37428
rect -31200 37108 -31120 37372
rect -31200 37052 -31188 37108
rect -31132 37052 -31120 37108
rect -31200 37040 -31120 37052
rect -31040 37752 -30960 37848
rect -31040 37688 -31032 37752
rect -30968 37688 -30960 37752
rect -31040 37428 -30960 37688
rect -30880 37588 -30800 42960
rect -30880 37532 -30868 37588
rect -30812 37532 -30800 37588
rect -30880 37520 -30800 37532
rect -30720 42868 -30640 42960
rect -30720 42812 -30708 42868
rect -30652 42812 -30640 42868
rect -30720 42708 -30640 42812
rect -30720 42652 -30708 42708
rect -30652 42652 -30640 42708
rect -30720 42548 -30640 42652
rect -30720 42492 -30708 42548
rect -30652 42492 -30640 42548
rect -30720 42388 -30640 42492
rect -30720 42332 -30708 42388
rect -30652 42332 -30640 42388
rect -30720 42228 -30640 42332
rect -30560 42388 -30480 42960
rect -30560 42332 -30548 42388
rect -30492 42332 -30480 42388
rect -30560 42320 -30480 42332
rect -30400 42868 -30320 42960
rect -30400 42812 -30388 42868
rect -30332 42812 -30320 42868
rect -30400 42708 -30320 42812
rect -30400 42652 -30388 42708
rect -30332 42652 -30320 42708
rect -30400 42548 -30320 42652
rect -30240 42708 -30160 42960
rect -30240 42652 -30228 42708
rect -30172 42652 -30160 42708
rect -30240 42640 -30160 42652
rect -30080 42868 -30000 42960
rect -30080 42812 -30068 42868
rect -30012 42812 -30000 42868
rect -30400 42492 -30388 42548
rect -30332 42492 -30320 42548
rect -30720 42172 -30708 42228
rect -30652 42172 -30640 42228
rect -30720 42068 -30640 42172
rect -30720 42012 -30708 42068
rect -30652 42012 -30640 42068
rect -30720 41908 -30640 42012
rect -30720 41852 -30708 41908
rect -30652 41852 -30640 41908
rect -30720 41752 -30640 41852
rect -30720 41688 -30712 41752
rect -30648 41688 -30640 41752
rect -30720 41592 -30640 41688
rect -30720 41528 -30712 41592
rect -30648 41528 -30640 41592
rect -30720 40792 -30640 41528
rect -30720 40728 -30712 40792
rect -30648 40728 -30640 40792
rect -30720 40632 -30640 40728
rect -30720 40568 -30712 40632
rect -30648 40568 -30640 40632
rect -30720 40472 -30640 40568
rect -30720 40408 -30712 40472
rect -30648 40408 -30640 40472
rect -30720 40312 -30640 40408
rect -30720 40248 -30712 40312
rect -30648 40248 -30640 40312
rect -30720 40152 -30640 40248
rect -30720 40088 -30712 40152
rect -30648 40088 -30640 40152
rect -30720 39992 -30640 40088
rect -30720 39928 -30712 39992
rect -30648 39928 -30640 39992
rect -30720 39832 -30640 39928
rect -30720 39768 -30712 39832
rect -30648 39768 -30640 39832
rect -30720 39672 -30640 39768
rect -30720 39608 -30712 39672
rect -30648 39608 -30640 39672
rect -30720 39512 -30640 39608
rect -30720 39448 -30712 39512
rect -30648 39448 -30640 39512
rect -30720 39352 -30640 39448
rect -30720 39288 -30712 39352
rect -30648 39288 -30640 39352
rect -30720 39192 -30640 39288
rect -30720 39128 -30712 39192
rect -30648 39128 -30640 39192
rect -30720 39032 -30640 39128
rect -30720 38968 -30712 39032
rect -30648 38968 -30640 39032
rect -30720 38872 -30640 38968
rect -30720 38808 -30712 38872
rect -30648 38808 -30640 38872
rect -30720 38712 -30640 38808
rect -30720 38648 -30712 38712
rect -30648 38648 -30640 38712
rect -30720 38552 -30640 38648
rect -30720 38488 -30712 38552
rect -30648 38488 -30640 38552
rect -30720 38392 -30640 38488
rect -30720 38328 -30712 38392
rect -30648 38328 -30640 38392
rect -30720 38232 -30640 38328
rect -30720 38168 -30712 38232
rect -30648 38168 -30640 38232
rect -30720 38072 -30640 38168
rect -30720 38008 -30712 38072
rect -30648 38008 -30640 38072
rect -30720 37912 -30640 38008
rect -30720 37848 -30712 37912
rect -30648 37848 -30640 37912
rect -30720 37752 -30640 37848
rect -30720 37688 -30712 37752
rect -30648 37688 -30640 37752
rect -31040 37372 -31028 37428
rect -30972 37372 -30960 37428
rect -31040 37112 -30960 37372
rect -30720 37428 -30640 37688
rect -30400 42228 -30320 42492
rect -30400 42172 -30388 42228
rect -30332 42172 -30320 42228
rect -30400 42068 -30320 42172
rect -30080 42548 -30000 42812
rect -30080 42492 -30068 42548
rect -30012 42492 -30000 42548
rect -30080 42228 -30000 42492
rect -30080 42172 -30068 42228
rect -30012 42172 -30000 42228
rect -30400 42012 -30388 42068
rect -30332 42012 -30320 42068
rect -30400 41908 -30320 42012
rect -30400 41852 -30388 41908
rect -30332 41852 -30320 41908
rect -30400 41752 -30320 41852
rect -30400 41688 -30392 41752
rect -30328 41688 -30320 41752
rect -30400 41592 -30320 41688
rect -30400 41528 -30392 41592
rect -30328 41528 -30320 41592
rect -30400 40792 -30320 41528
rect -30400 40728 -30392 40792
rect -30328 40728 -30320 40792
rect -30400 40632 -30320 40728
rect -30400 40568 -30392 40632
rect -30328 40568 -30320 40632
rect -30400 40472 -30320 40568
rect -30400 40408 -30392 40472
rect -30328 40408 -30320 40472
rect -30400 40312 -30320 40408
rect -30400 40248 -30392 40312
rect -30328 40248 -30320 40312
rect -30400 40152 -30320 40248
rect -30400 40088 -30392 40152
rect -30328 40088 -30320 40152
rect -30400 39992 -30320 40088
rect -30400 39928 -30392 39992
rect -30328 39928 -30320 39992
rect -30400 39832 -30320 39928
rect -30400 39768 -30392 39832
rect -30328 39768 -30320 39832
rect -30400 39672 -30320 39768
rect -30400 39608 -30392 39672
rect -30328 39608 -30320 39672
rect -30400 39512 -30320 39608
rect -30400 39448 -30392 39512
rect -30328 39448 -30320 39512
rect -30400 39352 -30320 39448
rect -30400 39288 -30392 39352
rect -30328 39288 -30320 39352
rect -30400 39192 -30320 39288
rect -30400 39128 -30392 39192
rect -30328 39128 -30320 39192
rect -30400 39032 -30320 39128
rect -30400 38968 -30392 39032
rect -30328 38968 -30320 39032
rect -30400 38872 -30320 38968
rect -30400 38808 -30392 38872
rect -30328 38808 -30320 38872
rect -30400 38712 -30320 38808
rect -30400 38648 -30392 38712
rect -30328 38648 -30320 38712
rect -30400 38552 -30320 38648
rect -30400 38488 -30392 38552
rect -30328 38488 -30320 38552
rect -30400 38392 -30320 38488
rect -30400 38328 -30392 38392
rect -30328 38328 -30320 38392
rect -30400 38232 -30320 38328
rect -30400 38168 -30392 38232
rect -30328 38168 -30320 38232
rect -30400 38072 -30320 38168
rect -30400 38008 -30392 38072
rect -30328 38008 -30320 38072
rect -30400 37912 -30320 38008
rect -30400 37848 -30392 37912
rect -30328 37848 -30320 37912
rect -30400 37752 -30320 37848
rect -30400 37688 -30392 37752
rect -30328 37688 -30320 37752
rect -30720 37372 -30708 37428
rect -30652 37372 -30640 37428
rect -31040 37048 -31032 37112
rect -30968 37048 -30960 37112
rect -31040 36952 -30960 37048
rect -31040 36888 -31032 36952
rect -30968 36888 -30960 36952
rect -31040 36792 -30960 36888
rect -31040 36728 -31032 36792
rect -30968 36728 -30960 36792
rect -31040 36632 -30960 36728
rect -31040 36568 -31032 36632
rect -30968 36568 -30960 36632
rect -31040 36472 -30960 36568
rect -31040 36408 -31032 36472
rect -30968 36408 -30960 36472
rect -31040 36312 -30960 36408
rect -31040 36248 -31032 36312
rect -30968 36248 -30960 36312
rect -31040 36152 -30960 36248
rect -31040 36088 -31032 36152
rect -30968 36088 -30960 36152
rect -31040 35992 -30960 36088
rect -31040 35928 -31032 35992
rect -30968 35928 -30960 35992
rect -31040 35832 -30960 35928
rect -31040 35768 -31032 35832
rect -30968 35768 -30960 35832
rect -31040 35672 -30960 35768
rect -31040 35608 -31032 35672
rect -30968 35608 -30960 35672
rect -31040 35512 -30960 35608
rect -31040 35448 -31032 35512
rect -30968 35448 -30960 35512
rect -31040 35352 -30960 35448
rect -31040 35288 -31032 35352
rect -30968 35288 -30960 35352
rect -31040 35192 -30960 35288
rect -31040 35128 -31032 35192
rect -30968 35128 -30960 35192
rect -31040 35032 -30960 35128
rect -31040 34968 -31032 35032
rect -30968 34968 -30960 35032
rect -31040 34872 -30960 34968
rect -31040 34808 -31032 34872
rect -30968 34808 -30960 34872
rect -33120 34708 -33040 34720
rect -33120 34652 -33108 34708
rect -33052 34652 -33040 34708
rect -33120 34388 -33040 34652
rect -33120 34332 -33108 34388
rect -33052 34332 -33040 34388
rect -33120 34320 -33040 34332
rect -32960 34708 -32880 34720
rect -32960 34652 -32948 34708
rect -32892 34652 -32880 34708
rect -32960 34388 -32880 34652
rect -32960 34332 -32948 34388
rect -32892 34332 -32880 34388
rect -32960 34320 -32880 34332
rect -32800 34708 -32720 34720
rect -32800 34652 -32788 34708
rect -32732 34652 -32720 34708
rect -32800 34388 -32720 34652
rect -32800 34332 -32788 34388
rect -32732 34332 -32720 34388
rect -32800 34320 -32720 34332
rect -32640 34708 -32560 34720
rect -32640 34652 -32628 34708
rect -32572 34652 -32560 34708
rect -32640 34388 -32560 34652
rect -32640 34332 -32628 34388
rect -32572 34332 -32560 34388
rect -32640 34320 -32560 34332
rect -32480 34708 -32400 34720
rect -32480 34652 -32468 34708
rect -32412 34652 -32400 34708
rect -32480 34388 -32400 34652
rect -32480 34332 -32468 34388
rect -32412 34332 -32400 34388
rect -32480 34320 -32400 34332
rect -32320 34708 -32240 34720
rect -32320 34652 -32308 34708
rect -32252 34652 -32240 34708
rect -32320 34388 -32240 34652
rect -32320 34332 -32308 34388
rect -32252 34332 -32240 34388
rect -32320 34320 -32240 34332
rect -32160 34708 -32080 34720
rect -32160 34652 -32148 34708
rect -32092 34652 -32080 34708
rect -32160 34388 -32080 34652
rect -32160 34332 -32148 34388
rect -32092 34332 -32080 34388
rect -32160 34320 -32080 34332
rect -32000 34708 -31920 34720
rect -32000 34652 -31988 34708
rect -31932 34652 -31920 34708
rect -32000 34388 -31920 34652
rect -32000 34332 -31988 34388
rect -31932 34332 -31920 34388
rect -32000 34320 -31920 34332
rect -31840 34708 -31760 34720
rect -31840 34652 -31828 34708
rect -31772 34652 -31760 34708
rect -31840 34388 -31760 34652
rect -31840 34332 -31828 34388
rect -31772 34332 -31760 34388
rect -31840 34320 -31760 34332
rect -31680 34708 -31600 34720
rect -31680 34652 -31668 34708
rect -31612 34652 -31600 34708
rect -31680 34388 -31600 34652
rect -31680 34332 -31668 34388
rect -31612 34332 -31600 34388
rect -31680 34320 -31600 34332
rect -31520 34708 -31440 34720
rect -31520 34652 -31508 34708
rect -31452 34652 -31440 34708
rect -31520 34388 -31440 34652
rect -31520 34332 -31508 34388
rect -31452 34332 -31440 34388
rect -31520 34320 -31440 34332
rect -31360 34708 -31280 34720
rect -31360 34652 -31348 34708
rect -31292 34652 -31280 34708
rect -31360 34388 -31280 34652
rect -31360 34332 -31348 34388
rect -31292 34332 -31280 34388
rect -31360 34320 -31280 34332
rect -31200 34708 -31120 34720
rect -31200 34652 -31188 34708
rect -31132 34652 -31120 34708
rect -31200 34388 -31120 34652
rect -31200 34332 -31188 34388
rect -31132 34332 -31120 34388
rect -31200 34320 -31120 34332
rect -31040 34708 -30960 34808
rect -31040 34652 -31028 34708
rect -30972 34652 -30960 34708
rect -31040 34388 -30960 34652
rect -31040 34332 -31028 34388
rect -30972 34332 -30960 34388
rect -31040 34232 -30960 34332
rect -31040 34168 -31032 34232
rect -30968 34168 -30960 34232
rect -31040 34072 -30960 34168
rect -31040 34008 -31032 34072
rect -30968 34008 -30960 34072
rect -31040 33912 -30960 34008
rect -31040 33848 -31032 33912
rect -30968 33848 -30960 33912
rect -31040 33752 -30960 33848
rect -31040 33688 -31032 33752
rect -30968 33688 -30960 33752
rect -31040 33592 -30960 33688
rect -31040 33528 -31032 33592
rect -30968 33528 -30960 33592
rect -31040 33432 -30960 33528
rect -31040 33368 -31032 33432
rect -30968 33368 -30960 33432
rect -31040 33272 -30960 33368
rect -31040 33208 -31032 33272
rect -30968 33208 -30960 33272
rect -31040 33112 -30960 33208
rect -31040 33048 -31032 33112
rect -30968 33048 -30960 33112
rect -31040 32952 -30960 33048
rect -31040 32888 -31032 32952
rect -30968 32888 -30960 32952
rect -31040 32788 -30960 32888
rect -31040 32732 -31028 32788
rect -30972 32732 -30960 32788
rect -31040 32628 -30960 32732
rect -31040 32572 -31028 32628
rect -30972 32572 -30960 32628
rect -31040 32468 -30960 32572
rect -31040 32412 -31028 32468
rect -30972 32412 -30960 32468
rect -31040 32308 -30960 32412
rect -31040 32252 -31028 32308
rect -30972 32252 -30960 32308
rect -31040 32148 -30960 32252
rect -31040 32092 -31028 32148
rect -30972 32092 -30960 32148
rect -31040 31988 -30960 32092
rect -31040 31932 -31028 31988
rect -30972 31932 -30960 31988
rect -31040 31840 -30960 31932
rect -30880 37268 -30800 37280
rect -30880 37212 -30868 37268
rect -30812 37212 -30800 37268
rect -30880 31840 -30800 37212
rect -30720 37112 -30640 37372
rect -30720 37048 -30712 37112
rect -30648 37048 -30640 37112
rect -30720 36952 -30640 37048
rect -30720 36888 -30712 36952
rect -30648 36888 -30640 36952
rect -30720 36792 -30640 36888
rect -30720 36728 -30712 36792
rect -30648 36728 -30640 36792
rect -30720 36632 -30640 36728
rect -30720 36568 -30712 36632
rect -30648 36568 -30640 36632
rect -30720 36472 -30640 36568
rect -30720 36408 -30712 36472
rect -30648 36408 -30640 36472
rect -30720 36312 -30640 36408
rect -30720 36248 -30712 36312
rect -30648 36248 -30640 36312
rect -30720 36152 -30640 36248
rect -30720 36088 -30712 36152
rect -30648 36088 -30640 36152
rect -30720 35992 -30640 36088
rect -30720 35928 -30712 35992
rect -30648 35928 -30640 35992
rect -30720 35832 -30640 35928
rect -30720 35768 -30712 35832
rect -30648 35768 -30640 35832
rect -30720 35672 -30640 35768
rect -30720 35608 -30712 35672
rect -30648 35608 -30640 35672
rect -30720 35512 -30640 35608
rect -30720 35448 -30712 35512
rect -30648 35448 -30640 35512
rect -30720 35352 -30640 35448
rect -30720 35288 -30712 35352
rect -30648 35288 -30640 35352
rect -30720 35192 -30640 35288
rect -30720 35128 -30712 35192
rect -30648 35128 -30640 35192
rect -30720 35032 -30640 35128
rect -30720 34968 -30712 35032
rect -30648 34968 -30640 35032
rect -30720 34872 -30640 34968
rect -30720 34808 -30712 34872
rect -30648 34808 -30640 34872
rect -30720 34708 -30640 34808
rect -30720 34652 -30708 34708
rect -30652 34652 -30640 34708
rect -30720 34388 -30640 34652
rect -30720 34332 -30708 34388
rect -30652 34332 -30640 34388
rect -30720 34232 -30640 34332
rect -30720 34168 -30712 34232
rect -30648 34168 -30640 34232
rect -30720 34072 -30640 34168
rect -30720 34008 -30712 34072
rect -30648 34008 -30640 34072
rect -30720 33912 -30640 34008
rect -30720 33848 -30712 33912
rect -30648 33848 -30640 33912
rect -30720 33752 -30640 33848
rect -30720 33688 -30712 33752
rect -30648 33688 -30640 33752
rect -30720 33592 -30640 33688
rect -30720 33528 -30712 33592
rect -30648 33528 -30640 33592
rect -30720 33432 -30640 33528
rect -30720 33368 -30712 33432
rect -30648 33368 -30640 33432
rect -30720 33272 -30640 33368
rect -30720 33208 -30712 33272
rect -30648 33208 -30640 33272
rect -30720 33112 -30640 33208
rect -30720 33048 -30712 33112
rect -30648 33048 -30640 33112
rect -30720 32952 -30640 33048
rect -30720 32888 -30712 32952
rect -30648 32888 -30640 32952
rect -30720 32788 -30640 32888
rect -30720 32732 -30708 32788
rect -30652 32732 -30640 32788
rect -30720 32628 -30640 32732
rect -30560 37588 -30480 37600
rect -30560 37532 -30548 37588
rect -30492 37532 -30480 37588
rect -30560 32788 -30480 37532
rect -30560 32732 -30548 32788
rect -30492 32732 -30480 32788
rect -30560 32720 -30480 32732
rect -30400 37428 -30320 37688
rect -30400 37372 -30388 37428
rect -30332 37372 -30320 37428
rect -30400 37112 -30320 37372
rect -30240 42068 -30160 42080
rect -30240 42012 -30228 42068
rect -30172 42012 -30160 42068
rect -30240 37268 -30160 42012
rect -30240 37212 -30228 37268
rect -30172 37212 -30160 37268
rect -30240 37200 -30160 37212
rect -30080 41908 -30000 42172
rect -30080 41852 -30068 41908
rect -30012 41852 -30000 41908
rect -30080 41752 -30000 41852
rect -29920 42868 -29840 42880
rect -29920 42812 -29908 42868
rect -29852 42812 -29840 42868
rect -29920 42548 -29840 42812
rect -29920 42492 -29908 42548
rect -29852 42492 -29840 42548
rect -29920 42228 -29840 42492
rect -29920 42172 -29908 42228
rect -29852 42172 -29840 42228
rect -29920 41908 -29840 42172
rect -29920 41852 -29908 41908
rect -29852 41852 -29840 41908
rect -29920 41840 -29840 41852
rect -29760 42868 -29680 42880
rect -29760 42812 -29748 42868
rect -29692 42812 -29680 42868
rect -29760 42548 -29680 42812
rect -29760 42492 -29748 42548
rect -29692 42492 -29680 42548
rect -29760 42228 -29680 42492
rect -29760 42172 -29748 42228
rect -29692 42172 -29680 42228
rect -29760 41908 -29680 42172
rect -29760 41852 -29748 41908
rect -29692 41852 -29680 41908
rect -29760 41840 -29680 41852
rect -29600 42868 -29520 42880
rect -29600 42812 -29588 42868
rect -29532 42812 -29520 42868
rect -29600 42548 -29520 42812
rect -29600 42492 -29588 42548
rect -29532 42492 -29520 42548
rect -29600 42228 -29520 42492
rect -29600 42172 -29588 42228
rect -29532 42172 -29520 42228
rect -29600 41908 -29520 42172
rect -29600 41852 -29588 41908
rect -29532 41852 -29520 41908
rect -29600 41840 -29520 41852
rect -29440 42868 -29360 42880
rect -29440 42812 -29428 42868
rect -29372 42812 -29360 42868
rect -29440 42548 -29360 42812
rect -29440 42492 -29428 42548
rect -29372 42492 -29360 42548
rect -29440 42228 -29360 42492
rect -29440 42172 -29428 42228
rect -29372 42172 -29360 42228
rect -29440 41908 -29360 42172
rect -29440 41852 -29428 41908
rect -29372 41852 -29360 41908
rect -29440 41840 -29360 41852
rect -29280 42868 -29200 42880
rect -29280 42812 -29268 42868
rect -29212 42812 -29200 42868
rect -29280 42548 -29200 42812
rect -29280 42492 -29268 42548
rect -29212 42492 -29200 42548
rect -29280 42228 -29200 42492
rect -29280 42172 -29268 42228
rect -29212 42172 -29200 42228
rect -29280 41908 -29200 42172
rect -29280 41852 -29268 41908
rect -29212 41852 -29200 41908
rect -29280 41840 -29200 41852
rect -29120 42868 -29040 42880
rect -29120 42812 -29108 42868
rect -29052 42812 -29040 42868
rect -29120 42548 -29040 42812
rect -29120 42492 -29108 42548
rect -29052 42492 -29040 42548
rect -29120 42228 -29040 42492
rect -29120 42172 -29108 42228
rect -29052 42172 -29040 42228
rect -29120 41908 -29040 42172
rect -29120 41852 -29108 41908
rect -29052 41852 -29040 41908
rect -29120 41840 -29040 41852
rect -28960 42868 -28880 42880
rect -28960 42812 -28948 42868
rect -28892 42812 -28880 42868
rect -28960 42548 -28880 42812
rect -28960 42492 -28948 42548
rect -28892 42492 -28880 42548
rect -28960 42228 -28880 42492
rect -28960 42172 -28948 42228
rect -28892 42172 -28880 42228
rect -28960 41908 -28880 42172
rect -28960 41852 -28948 41908
rect -28892 41852 -28880 41908
rect -28960 41840 -28880 41852
rect -28800 42868 -28720 42880
rect -28800 42812 -28788 42868
rect -28732 42812 -28720 42868
rect -28800 42548 -28720 42812
rect -28800 42492 -28788 42548
rect -28732 42492 -28720 42548
rect -28800 42228 -28720 42492
rect -28800 42172 -28788 42228
rect -28732 42172 -28720 42228
rect -28800 41908 -28720 42172
rect -28800 41852 -28788 41908
rect -28732 41852 -28720 41908
rect -28800 41840 -28720 41852
rect -28640 42868 -28560 42880
rect -28640 42812 -28628 42868
rect -28572 42812 -28560 42868
rect -28640 42548 -28560 42812
rect -28640 42492 -28628 42548
rect -28572 42492 -28560 42548
rect -28640 42228 -28560 42492
rect -28640 42172 -28628 42228
rect -28572 42172 -28560 42228
rect -28640 41908 -28560 42172
rect -28640 41852 -28628 41908
rect -28572 41852 -28560 41908
rect -28640 41840 -28560 41852
rect -28480 42868 -28400 42880
rect -28480 42812 -28468 42868
rect -28412 42812 -28400 42868
rect -28480 42548 -28400 42812
rect -28480 42492 -28468 42548
rect -28412 42492 -28400 42548
rect -28480 42228 -28400 42492
rect -28480 42172 -28468 42228
rect -28412 42172 -28400 42228
rect -28480 41908 -28400 42172
rect -28480 41852 -28468 41908
rect -28412 41852 -28400 41908
rect -28480 41840 -28400 41852
rect -28320 42868 -28240 42880
rect -28320 42812 -28308 42868
rect -28252 42812 -28240 42868
rect -28320 42548 -28240 42812
rect -28320 42492 -28308 42548
rect -28252 42492 -28240 42548
rect -28320 42228 -28240 42492
rect -28320 42172 -28308 42228
rect -28252 42172 -28240 42228
rect -28320 41908 -28240 42172
rect -28320 41852 -28308 41908
rect -28252 41852 -28240 41908
rect -28320 41840 -28240 41852
rect -28160 42868 -28080 42880
rect -28160 42812 -28148 42868
rect -28092 42812 -28080 42868
rect -28160 42548 -28080 42812
rect -28160 42492 -28148 42548
rect -28092 42492 -28080 42548
rect -28160 42228 -28080 42492
rect -28160 42172 -28148 42228
rect -28092 42172 -28080 42228
rect -28160 41908 -28080 42172
rect -28160 41852 -28148 41908
rect -28092 41852 -28080 41908
rect -28160 41840 -28080 41852
rect -28000 42868 -27920 42880
rect -28000 42812 -27988 42868
rect -27932 42812 -27920 42868
rect -28000 42548 -27920 42812
rect -28000 42492 -27988 42548
rect -27932 42492 -27920 42548
rect -28000 42228 -27920 42492
rect -28000 42172 -27988 42228
rect -27932 42172 -27920 42228
rect -28000 41908 -27920 42172
rect -28000 41852 -27988 41908
rect -27932 41852 -27920 41908
rect -28000 41840 -27920 41852
rect -27840 42868 -27760 42880
rect -27840 42812 -27828 42868
rect -27772 42812 -27760 42868
rect -27840 42548 -27760 42812
rect -27840 42492 -27828 42548
rect -27772 42492 -27760 42548
rect -27840 42228 -27760 42492
rect -27840 42172 -27828 42228
rect -27772 42172 -27760 42228
rect -27840 41908 -27760 42172
rect -27840 41852 -27828 41908
rect -27772 41852 -27760 41908
rect -27840 41840 -27760 41852
rect -27680 42868 -27600 42880
rect -27680 42812 -27668 42868
rect -27612 42812 -27600 42868
rect -27680 42548 -27600 42812
rect -27680 42492 -27668 42548
rect -27612 42492 -27600 42548
rect -27680 42228 -27600 42492
rect -27680 42172 -27668 42228
rect -27612 42172 -27600 42228
rect -27680 41908 -27600 42172
rect -27680 41852 -27668 41908
rect -27612 41852 -27600 41908
rect -27680 41840 -27600 41852
rect -27520 42868 -27440 42880
rect -27520 42812 -27508 42868
rect -27452 42812 -27440 42868
rect -27520 42548 -27440 42812
rect -27520 42492 -27508 42548
rect -27452 42492 -27440 42548
rect -27520 42228 -27440 42492
rect -27520 42172 -27508 42228
rect -27452 42172 -27440 42228
rect -27520 41908 -27440 42172
rect -27520 41852 -27508 41908
rect -27452 41852 -27440 41908
rect -27520 41840 -27440 41852
rect -27360 42868 -27280 42880
rect -27360 42812 -27348 42868
rect -27292 42812 -27280 42868
rect -27360 42548 -27280 42812
rect -27360 42492 -27348 42548
rect -27292 42492 -27280 42548
rect -27360 42228 -27280 42492
rect -27360 42172 -27348 42228
rect -27292 42172 -27280 42228
rect -27360 41908 -27280 42172
rect -27360 41852 -27348 41908
rect -27292 41852 -27280 41908
rect -27360 41840 -27280 41852
rect -27200 42868 -27120 42880
rect -27200 42812 -27188 42868
rect -27132 42812 -27120 42868
rect -27200 42548 -27120 42812
rect -27200 42492 -27188 42548
rect -27132 42492 -27120 42548
rect -27200 42228 -27120 42492
rect -27200 42172 -27188 42228
rect -27132 42172 -27120 42228
rect -27200 41908 -27120 42172
rect -27200 41852 -27188 41908
rect -27132 41852 -27120 41908
rect -27200 41840 -27120 41852
rect -27040 42868 -26960 42880
rect -27040 42812 -27028 42868
rect -26972 42812 -26960 42868
rect -27040 42548 -26960 42812
rect -27040 42492 -27028 42548
rect -26972 42492 -26960 42548
rect -27040 42228 -26960 42492
rect -27040 42172 -27028 42228
rect -26972 42172 -26960 42228
rect -27040 41908 -26960 42172
rect -27040 41852 -27028 41908
rect -26972 41852 -26960 41908
rect -27040 41840 -26960 41852
rect -26880 42868 -26800 42880
rect -26880 42812 -26868 42868
rect -26812 42812 -26800 42868
rect -26880 42548 -26800 42812
rect -26880 42492 -26868 42548
rect -26812 42492 -26800 42548
rect -26880 42228 -26800 42492
rect -26880 42172 -26868 42228
rect -26812 42172 -26800 42228
rect -26880 41908 -26800 42172
rect -26880 41852 -26868 41908
rect -26812 41852 -26800 41908
rect -26880 41840 -26800 41852
rect -26720 42868 -26640 42880
rect -26720 42812 -26708 42868
rect -26652 42812 -26640 42868
rect -26720 42548 -26640 42812
rect -26720 42492 -26708 42548
rect -26652 42492 -26640 42548
rect -26720 42228 -26640 42492
rect -26720 42172 -26708 42228
rect -26652 42172 -26640 42228
rect -26720 41908 -26640 42172
rect -26720 41852 -26708 41908
rect -26652 41852 -26640 41908
rect -26720 41840 -26640 41852
rect -26560 42868 -26480 42880
rect -26560 42812 -26548 42868
rect -26492 42812 -26480 42868
rect -26560 42548 -26480 42812
rect -26560 42492 -26548 42548
rect -26492 42492 -26480 42548
rect -26560 42228 -26480 42492
rect -26560 42172 -26548 42228
rect -26492 42172 -26480 42228
rect -26560 41908 -26480 42172
rect -26560 41852 -26548 41908
rect -26492 41852 -26480 41908
rect -26560 41840 -26480 41852
rect -26400 42868 -26320 42880
rect -26400 42812 -26388 42868
rect -26332 42812 -26320 42868
rect -26400 42548 -26320 42812
rect -26400 42492 -26388 42548
rect -26332 42492 -26320 42548
rect -26400 42228 -26320 42492
rect -26400 42172 -26388 42228
rect -26332 42172 -26320 42228
rect -26400 41908 -26320 42172
rect -26400 41852 -26388 41908
rect -26332 41852 -26320 41908
rect -26400 41840 -26320 41852
rect -26240 42868 -26160 42880
rect -26240 42812 -26228 42868
rect -26172 42812 -26160 42868
rect -26240 42548 -26160 42812
rect -26240 42492 -26228 42548
rect -26172 42492 -26160 42548
rect -26240 42228 -26160 42492
rect -26240 42172 -26228 42228
rect -26172 42172 -26160 42228
rect -26240 41908 -26160 42172
rect -26240 41852 -26228 41908
rect -26172 41852 -26160 41908
rect -26240 41840 -26160 41852
rect -26080 42868 -26000 42880
rect -26080 42812 -26068 42868
rect -26012 42812 -26000 42868
rect -26080 42548 -26000 42812
rect -26080 42492 -26068 42548
rect -26012 42492 -26000 42548
rect -26080 42228 -26000 42492
rect -26080 42172 -26068 42228
rect -26012 42172 -26000 42228
rect -26080 41908 -26000 42172
rect -26080 41852 -26068 41908
rect -26012 41852 -26000 41908
rect -26080 41840 -26000 41852
rect -25920 42868 -25840 42880
rect -25920 42812 -25908 42868
rect -25852 42812 -25840 42868
rect -25920 42548 -25840 42812
rect -25920 42492 -25908 42548
rect -25852 42492 -25840 42548
rect -25920 42228 -25840 42492
rect -25920 42172 -25908 42228
rect -25852 42172 -25840 42228
rect -25920 41908 -25840 42172
rect -25920 41852 -25908 41908
rect -25852 41852 -25840 41908
rect -25920 41840 -25840 41852
rect -25760 42868 -25680 42880
rect -25760 42812 -25748 42868
rect -25692 42812 -25680 42868
rect -25760 42548 -25680 42812
rect -25760 42492 -25748 42548
rect -25692 42492 -25680 42548
rect -25760 42228 -25680 42492
rect -25760 42172 -25748 42228
rect -25692 42172 -25680 42228
rect -25760 41908 -25680 42172
rect -25760 41852 -25748 41908
rect -25692 41852 -25680 41908
rect -25760 41840 -25680 41852
rect -25600 42868 -25520 42880
rect -25600 42812 -25588 42868
rect -25532 42812 -25520 42868
rect -25600 42548 -25520 42812
rect -25600 42492 -25588 42548
rect -25532 42492 -25520 42548
rect -25600 42228 -25520 42492
rect -25600 42172 -25588 42228
rect -25532 42172 -25520 42228
rect -25600 41908 -25520 42172
rect -25600 41852 -25588 41908
rect -25532 41852 -25520 41908
rect -25600 41840 -25520 41852
rect -25440 42868 -25360 42880
rect -25440 42812 -25428 42868
rect -25372 42812 -25360 42868
rect -25440 42548 -25360 42812
rect -25440 42492 -25428 42548
rect -25372 42492 -25360 42548
rect -25440 42228 -25360 42492
rect -25440 42172 -25428 42228
rect -25372 42172 -25360 42228
rect -25440 41908 -25360 42172
rect -25440 41852 -25428 41908
rect -25372 41852 -25360 41908
rect -25440 41840 -25360 41852
rect -25280 42868 -25200 42880
rect -25280 42812 -25268 42868
rect -25212 42812 -25200 42868
rect -25280 42548 -25200 42812
rect -25280 42492 -25268 42548
rect -25212 42492 -25200 42548
rect -25280 42228 -25200 42492
rect -25280 42172 -25268 42228
rect -25212 42172 -25200 42228
rect -25280 41908 -25200 42172
rect -25280 41852 -25268 41908
rect -25212 41852 -25200 41908
rect -25280 41840 -25200 41852
rect -25120 42868 -25040 42880
rect -25120 42812 -25108 42868
rect -25052 42812 -25040 42868
rect -25120 42548 -25040 42812
rect -25120 42492 -25108 42548
rect -25052 42492 -25040 42548
rect -25120 42228 -25040 42492
rect -25120 42172 -25108 42228
rect -25052 42172 -25040 42228
rect -25120 41908 -25040 42172
rect -25120 41852 -25108 41908
rect -25052 41852 -25040 41908
rect -25120 41840 -25040 41852
rect -24960 42868 -24880 42880
rect -24960 42812 -24948 42868
rect -24892 42812 -24880 42868
rect -24960 42548 -24880 42812
rect -24960 42492 -24948 42548
rect -24892 42492 -24880 42548
rect -24960 42228 -24880 42492
rect -24960 42172 -24948 42228
rect -24892 42172 -24880 42228
rect -24960 41908 -24880 42172
rect -24960 41852 -24948 41908
rect -24892 41852 -24880 41908
rect -24960 41840 -24880 41852
rect -24800 42868 -24720 42880
rect -24800 42812 -24788 42868
rect -24732 42812 -24720 42868
rect -24800 42548 -24720 42812
rect -24800 42492 -24788 42548
rect -24732 42492 -24720 42548
rect -24800 42228 -24720 42492
rect -24800 42172 -24788 42228
rect -24732 42172 -24720 42228
rect -24800 41908 -24720 42172
rect -24800 41852 -24788 41908
rect -24732 41852 -24720 41908
rect -24800 41840 -24720 41852
rect -24640 42868 -24560 42880
rect -24640 42812 -24628 42868
rect -24572 42812 -24560 42868
rect -24640 42548 -24560 42812
rect -24640 42492 -24628 42548
rect -24572 42492 -24560 42548
rect -24640 42228 -24560 42492
rect -24640 42172 -24628 42228
rect -24572 42172 -24560 42228
rect -24640 41908 -24560 42172
rect -24640 41852 -24628 41908
rect -24572 41852 -24560 41908
rect -24640 41840 -24560 41852
rect -24480 42868 -24400 42880
rect -24480 42812 -24468 42868
rect -24412 42812 -24400 42868
rect -24480 42548 -24400 42812
rect -24480 42492 -24468 42548
rect -24412 42492 -24400 42548
rect -24480 42228 -24400 42492
rect -24480 42172 -24468 42228
rect -24412 42172 -24400 42228
rect -24480 41908 -24400 42172
rect -24480 41852 -24468 41908
rect -24412 41852 -24400 41908
rect -24480 41840 -24400 41852
rect -24320 42868 -24240 42880
rect -24320 42812 -24308 42868
rect -24252 42812 -24240 42868
rect -24320 42548 -24240 42812
rect -24320 42492 -24308 42548
rect -24252 42492 -24240 42548
rect -24320 42228 -24240 42492
rect -24320 42172 -24308 42228
rect -24252 42172 -24240 42228
rect -24320 41908 -24240 42172
rect -24320 41852 -24308 41908
rect -24252 41852 -24240 41908
rect -24320 41840 -24240 41852
rect -24160 42868 -24080 42880
rect -24160 42812 -24148 42868
rect -24092 42812 -24080 42868
rect -24160 42548 -24080 42812
rect -24160 42492 -24148 42548
rect -24092 42492 -24080 42548
rect -24160 42228 -24080 42492
rect -24160 42172 -24148 42228
rect -24092 42172 -24080 42228
rect -24160 41908 -24080 42172
rect -24160 41852 -24148 41908
rect -24092 41852 -24080 41908
rect -24160 41840 -24080 41852
rect -24000 42868 -23920 42880
rect -24000 42812 -23988 42868
rect -23932 42812 -23920 42868
rect -24000 42548 -23920 42812
rect -24000 42492 -23988 42548
rect -23932 42492 -23920 42548
rect -24000 42228 -23920 42492
rect -24000 42172 -23988 42228
rect -23932 42172 -23920 42228
rect -24000 41908 -23920 42172
rect -24000 41852 -23988 41908
rect -23932 41852 -23920 41908
rect -24000 41840 -23920 41852
rect -23840 42868 -23760 42880
rect -23840 42812 -23828 42868
rect -23772 42812 -23760 42868
rect -23840 42548 -23760 42812
rect -23840 42492 -23828 42548
rect -23772 42492 -23760 42548
rect -23840 42228 -23760 42492
rect -23840 42172 -23828 42228
rect -23772 42172 -23760 42228
rect -23840 41908 -23760 42172
rect -23840 41852 -23828 41908
rect -23772 41852 -23760 41908
rect -23840 41840 -23760 41852
rect -23680 42868 -23600 42880
rect -23680 42812 -23668 42868
rect -23612 42812 -23600 42868
rect -23680 42548 -23600 42812
rect -23680 42492 -23668 42548
rect -23612 42492 -23600 42548
rect -23680 42228 -23600 42492
rect -23680 42172 -23668 42228
rect -23612 42172 -23600 42228
rect -23680 41908 -23600 42172
rect -23680 41852 -23668 41908
rect -23612 41852 -23600 41908
rect -23680 41840 -23600 41852
rect -23520 42868 -23440 42880
rect -23520 42812 -23508 42868
rect -23452 42812 -23440 42868
rect -23520 42548 -23440 42812
rect -23520 42492 -23508 42548
rect -23452 42492 -23440 42548
rect -23520 42228 -23440 42492
rect -23520 42172 -23508 42228
rect -23452 42172 -23440 42228
rect -23520 41908 -23440 42172
rect -23520 41852 -23508 41908
rect -23452 41852 -23440 41908
rect -23520 41840 -23440 41852
rect -23360 42868 -23280 42880
rect -23360 42812 -23348 42868
rect -23292 42812 -23280 42868
rect -23360 42548 -23280 42812
rect -23360 42492 -23348 42548
rect -23292 42492 -23280 42548
rect -23360 42228 -23280 42492
rect -23360 42172 -23348 42228
rect -23292 42172 -23280 42228
rect -23360 41908 -23280 42172
rect -23360 41852 -23348 41908
rect -23292 41852 -23280 41908
rect -23360 41840 -23280 41852
rect -23200 42868 -23120 42880
rect -23200 42812 -23188 42868
rect -23132 42812 -23120 42868
rect -23200 42548 -23120 42812
rect -23200 42492 -23188 42548
rect -23132 42492 -23120 42548
rect -23200 42228 -23120 42492
rect -23200 42172 -23188 42228
rect -23132 42172 -23120 42228
rect -23200 41908 -23120 42172
rect -23200 41852 -23188 41908
rect -23132 41852 -23120 41908
rect -23200 41840 -23120 41852
rect -23040 42868 -22960 42880
rect -23040 42812 -23028 42868
rect -22972 42812 -22960 42868
rect -23040 42548 -22960 42812
rect -23040 42492 -23028 42548
rect -22972 42492 -22960 42548
rect -23040 42228 -22960 42492
rect -23040 42172 -23028 42228
rect -22972 42172 -22960 42228
rect -23040 41908 -22960 42172
rect -23040 41852 -23028 41908
rect -22972 41852 -22960 41908
rect -23040 41840 -22960 41852
rect -22880 42868 -22800 42880
rect -22880 42812 -22868 42868
rect -22812 42812 -22800 42868
rect -22880 42548 -22800 42812
rect -22880 42492 -22868 42548
rect -22812 42492 -22800 42548
rect -22880 42228 -22800 42492
rect -22880 42172 -22868 42228
rect -22812 42172 -22800 42228
rect -22880 41908 -22800 42172
rect -22880 41852 -22868 41908
rect -22812 41852 -22800 41908
rect -22880 41840 -22800 41852
rect -22720 42868 -22640 42880
rect -22720 42812 -22708 42868
rect -22652 42812 -22640 42868
rect -22720 42548 -22640 42812
rect -22720 42492 -22708 42548
rect -22652 42492 -22640 42548
rect -22720 42228 -22640 42492
rect -22720 42172 -22708 42228
rect -22652 42172 -22640 42228
rect -22720 41908 -22640 42172
rect -22720 41852 -22708 41908
rect -22652 41852 -22640 41908
rect -22720 41840 -22640 41852
rect -22560 42868 -22480 42880
rect -22560 42812 -22548 42868
rect -22492 42812 -22480 42868
rect -22560 42548 -22480 42812
rect -22560 42492 -22548 42548
rect -22492 42492 -22480 42548
rect -22560 42228 -22480 42492
rect -22560 42172 -22548 42228
rect -22492 42172 -22480 42228
rect -22560 41908 -22480 42172
rect -22560 41852 -22548 41908
rect -22492 41852 -22480 41908
rect -22560 41840 -22480 41852
rect -22400 42868 -22320 42880
rect -22400 42812 -22388 42868
rect -22332 42812 -22320 42868
rect -22400 42548 -22320 42812
rect -22400 42492 -22388 42548
rect -22332 42492 -22320 42548
rect -22400 42228 -22320 42492
rect -22400 42172 -22388 42228
rect -22332 42172 -22320 42228
rect -22400 41908 -22320 42172
rect -22400 41852 -22388 41908
rect -22332 41852 -22320 41908
rect -22400 41840 -22320 41852
rect -22240 42868 -22160 42880
rect -22240 42812 -22228 42868
rect -22172 42812 -22160 42868
rect -22240 42548 -22160 42812
rect -22240 42492 -22228 42548
rect -22172 42492 -22160 42548
rect -22240 42228 -22160 42492
rect -22240 42172 -22228 42228
rect -22172 42172 -22160 42228
rect -22240 41908 -22160 42172
rect -22240 41852 -22228 41908
rect -22172 41852 -22160 41908
rect -22240 41840 -22160 41852
rect -22080 42868 -22000 42880
rect -22080 42812 -22068 42868
rect -22012 42812 -22000 42868
rect -22080 42548 -22000 42812
rect -22080 42492 -22068 42548
rect -22012 42492 -22000 42548
rect -22080 42228 -22000 42492
rect -22080 42172 -22068 42228
rect -22012 42172 -22000 42228
rect -22080 41908 -22000 42172
rect -22080 41852 -22068 41908
rect -22012 41852 -22000 41908
rect -22080 41840 -22000 41852
rect -21920 42868 -21840 42880
rect -21920 42812 -21908 42868
rect -21852 42812 -21840 42868
rect -21920 42548 -21840 42812
rect -21920 42492 -21908 42548
rect -21852 42492 -21840 42548
rect -21920 42228 -21840 42492
rect -21920 42172 -21908 42228
rect -21852 42172 -21840 42228
rect -21920 41908 -21840 42172
rect -21920 41852 -21908 41908
rect -21852 41852 -21840 41908
rect -21920 41840 -21840 41852
rect -21760 42868 -21680 42880
rect -21760 42812 -21748 42868
rect -21692 42812 -21680 42868
rect -21760 42548 -21680 42812
rect -21760 42492 -21748 42548
rect -21692 42492 -21680 42548
rect -21760 42228 -21680 42492
rect -21760 42172 -21748 42228
rect -21692 42172 -21680 42228
rect -21760 41908 -21680 42172
rect -21760 41852 -21748 41908
rect -21692 41852 -21680 41908
rect -21760 41840 -21680 41852
rect -21600 42868 -21520 42880
rect -21600 42812 -21588 42868
rect -21532 42812 -21520 42868
rect -21600 42548 -21520 42812
rect -21600 42492 -21588 42548
rect -21532 42492 -21520 42548
rect -21600 42228 -21520 42492
rect -21600 42172 -21588 42228
rect -21532 42172 -21520 42228
rect -21600 41908 -21520 42172
rect -21600 41852 -21588 41908
rect -21532 41852 -21520 41908
rect -21600 41840 -21520 41852
rect -21440 42868 -21360 42880
rect -21440 42812 -21428 42868
rect -21372 42812 -21360 42868
rect -21440 42548 -21360 42812
rect -21440 42492 -21428 42548
rect -21372 42492 -21360 42548
rect -21440 42228 -21360 42492
rect -21440 42172 -21428 42228
rect -21372 42172 -21360 42228
rect -21440 41908 -21360 42172
rect -21440 41852 -21428 41908
rect -21372 41852 -21360 41908
rect -21440 41840 -21360 41852
rect -21280 42868 -21200 42880
rect -21280 42812 -21268 42868
rect -21212 42812 -21200 42868
rect -21280 42548 -21200 42812
rect -21280 42492 -21268 42548
rect -21212 42492 -21200 42548
rect -21280 42228 -21200 42492
rect -21280 42172 -21268 42228
rect -21212 42172 -21200 42228
rect -21280 41908 -21200 42172
rect -21280 41852 -21268 41908
rect -21212 41852 -21200 41908
rect -21280 41840 -21200 41852
rect -21120 42868 -21040 42880
rect -21120 42812 -21108 42868
rect -21052 42812 -21040 42868
rect -21120 42548 -21040 42812
rect -21120 42492 -21108 42548
rect -21052 42492 -21040 42548
rect -21120 42228 -21040 42492
rect -21120 42172 -21108 42228
rect -21052 42172 -21040 42228
rect -21120 41908 -21040 42172
rect -21120 41852 -21108 41908
rect -21052 41852 -21040 41908
rect -21120 41840 -21040 41852
rect -20960 42868 -20880 42880
rect -20960 42812 -20948 42868
rect -20892 42812 -20880 42868
rect -20960 42548 -20880 42812
rect -20960 42492 -20948 42548
rect -20892 42492 -20880 42548
rect -20960 42228 -20880 42492
rect -20960 42172 -20948 42228
rect -20892 42172 -20880 42228
rect -20960 41908 -20880 42172
rect -20960 41852 -20948 41908
rect -20892 41852 -20880 41908
rect -20960 41840 -20880 41852
rect -20800 42868 -20720 42880
rect -20800 42812 -20788 42868
rect -20732 42812 -20720 42868
rect -20800 42548 -20720 42812
rect -20800 42492 -20788 42548
rect -20732 42492 -20720 42548
rect -20800 42228 -20720 42492
rect -20800 42172 -20788 42228
rect -20732 42172 -20720 42228
rect -20800 41908 -20720 42172
rect -20800 41852 -20788 41908
rect -20732 41852 -20720 41908
rect -20800 41840 -20720 41852
rect -20640 42868 -20560 42880
rect -20640 42812 -20628 42868
rect -20572 42812 -20560 42868
rect -20640 42548 -20560 42812
rect -20640 42492 -20628 42548
rect -20572 42492 -20560 42548
rect -20640 42228 -20560 42492
rect -20640 42172 -20628 42228
rect -20572 42172 -20560 42228
rect -20640 41908 -20560 42172
rect -20640 41852 -20628 41908
rect -20572 41852 -20560 41908
rect -20640 41840 -20560 41852
rect -20480 42868 -20400 42880
rect -20480 42812 -20468 42868
rect -20412 42812 -20400 42868
rect -20480 42548 -20400 42812
rect -20480 42492 -20468 42548
rect -20412 42492 -20400 42548
rect -20480 42228 -20400 42492
rect -20480 42172 -20468 42228
rect -20412 42172 -20400 42228
rect -20480 41908 -20400 42172
rect -20480 41852 -20468 41908
rect -20412 41852 -20400 41908
rect -20480 41840 -20400 41852
rect -20320 42868 -20240 42880
rect -20320 42812 -20308 42868
rect -20252 42812 -20240 42868
rect -20320 42548 -20240 42812
rect -20320 42492 -20308 42548
rect -20252 42492 -20240 42548
rect -20320 42228 -20240 42492
rect -20320 42172 -20308 42228
rect -20252 42172 -20240 42228
rect -20320 41908 -20240 42172
rect -20320 41852 -20308 41908
rect -20252 41852 -20240 41908
rect -20320 41840 -20240 41852
rect -20160 42868 -20080 42880
rect -20160 42812 -20148 42868
rect -20092 42812 -20080 42868
rect -20160 42548 -20080 42812
rect -20160 42492 -20148 42548
rect -20092 42492 -20080 42548
rect -20160 42228 -20080 42492
rect -20160 42172 -20148 42228
rect -20092 42172 -20080 42228
rect -20160 41908 -20080 42172
rect -20160 41852 -20148 41908
rect -20092 41852 -20080 41908
rect -20160 41840 -20080 41852
rect -20000 42868 -19920 42880
rect -20000 42812 -19988 42868
rect -19932 42812 -19920 42868
rect -20000 42548 -19920 42812
rect -20000 42492 -19988 42548
rect -19932 42492 -19920 42548
rect -20000 42228 -19920 42492
rect -20000 42172 -19988 42228
rect -19932 42172 -19920 42228
rect -20000 41908 -19920 42172
rect -20000 41852 -19988 41908
rect -19932 41852 -19920 41908
rect -20000 41840 -19920 41852
rect -19840 42868 -19760 42880
rect -19840 42812 -19828 42868
rect -19772 42812 -19760 42868
rect -19840 42548 -19760 42812
rect -19840 42492 -19828 42548
rect -19772 42492 -19760 42548
rect -19840 42228 -19760 42492
rect -19840 42172 -19828 42228
rect -19772 42172 -19760 42228
rect -19840 41908 -19760 42172
rect -19840 41852 -19828 41908
rect -19772 41852 -19760 41908
rect -19840 41840 -19760 41852
rect -19680 42868 -19600 42880
rect -19680 42812 -19668 42868
rect -19612 42812 -19600 42868
rect -19680 42548 -19600 42812
rect -19680 42492 -19668 42548
rect -19612 42492 -19600 42548
rect -19680 42228 -19600 42492
rect -19680 42172 -19668 42228
rect -19612 42172 -19600 42228
rect -19680 41908 -19600 42172
rect -19680 41852 -19668 41908
rect -19612 41852 -19600 41908
rect -19680 41840 -19600 41852
rect -19520 42868 -19440 42880
rect -19520 42812 -19508 42868
rect -19452 42812 -19440 42868
rect -19520 42548 -19440 42812
rect -19520 42492 -19508 42548
rect -19452 42492 -19440 42548
rect -19520 42228 -19440 42492
rect -19520 42172 -19508 42228
rect -19452 42172 -19440 42228
rect -19520 41908 -19440 42172
rect -19520 41852 -19508 41908
rect -19452 41852 -19440 41908
rect -19520 41840 -19440 41852
rect -19360 42868 -19280 42880
rect -19360 42812 -19348 42868
rect -19292 42812 -19280 42868
rect -19360 42548 -19280 42812
rect -19360 42492 -19348 42548
rect -19292 42492 -19280 42548
rect -19360 42228 -19280 42492
rect -19360 42172 -19348 42228
rect -19292 42172 -19280 42228
rect -19360 41908 -19280 42172
rect -19360 41852 -19348 41908
rect -19292 41852 -19280 41908
rect -19360 41840 -19280 41852
rect -19200 42868 -19120 42880
rect -19200 42812 -19188 42868
rect -19132 42812 -19120 42868
rect -19200 42548 -19120 42812
rect -19200 42492 -19188 42548
rect -19132 42492 -19120 42548
rect -19200 42228 -19120 42492
rect -19200 42172 -19188 42228
rect -19132 42172 -19120 42228
rect -19200 41908 -19120 42172
rect -19200 41852 -19188 41908
rect -19132 41852 -19120 41908
rect -19200 41840 -19120 41852
rect -19040 42868 -18960 42880
rect -19040 42812 -19028 42868
rect -18972 42812 -18960 42868
rect -19040 42548 -18960 42812
rect -19040 42492 -19028 42548
rect -18972 42492 -18960 42548
rect -19040 42228 -18960 42492
rect -19040 42172 -19028 42228
rect -18972 42172 -18960 42228
rect -19040 41908 -18960 42172
rect -19040 41852 -19028 41908
rect -18972 41852 -18960 41908
rect -19040 41840 -18960 41852
rect -18880 42868 -18800 42880
rect -18880 42812 -18868 42868
rect -18812 42812 -18800 42868
rect -18880 42548 -18800 42812
rect -18880 42492 -18868 42548
rect -18812 42492 -18800 42548
rect -18880 42228 -18800 42492
rect -18880 42172 -18868 42228
rect -18812 42172 -18800 42228
rect -18880 41908 -18800 42172
rect -18880 41852 -18868 41908
rect -18812 41852 -18800 41908
rect -18880 41840 -18800 41852
rect -18720 42868 -18640 42880
rect -18720 42812 -18708 42868
rect -18652 42812 -18640 42868
rect -18720 42548 -18640 42812
rect -18720 42492 -18708 42548
rect -18652 42492 -18640 42548
rect -18720 42228 -18640 42492
rect -18720 42172 -18708 42228
rect -18652 42172 -18640 42228
rect -18720 41908 -18640 42172
rect -18720 41852 -18708 41908
rect -18652 41852 -18640 41908
rect -18720 41840 -18640 41852
rect -18560 42868 -18480 42880
rect -18560 42812 -18548 42868
rect -18492 42812 -18480 42868
rect -18560 42548 -18480 42812
rect -18560 42492 -18548 42548
rect -18492 42492 -18480 42548
rect -18560 42228 -18480 42492
rect -18560 42172 -18548 42228
rect -18492 42172 -18480 42228
rect -18560 41908 -18480 42172
rect -18560 41852 -18548 41908
rect -18492 41852 -18480 41908
rect -18560 41840 -18480 41852
rect -18400 42868 -18320 42880
rect -18400 42812 -18388 42868
rect -18332 42812 -18320 42868
rect -18400 42548 -18320 42812
rect -18400 42492 -18388 42548
rect -18332 42492 -18320 42548
rect -18400 42228 -18320 42492
rect -18400 42172 -18388 42228
rect -18332 42172 -18320 42228
rect -18400 41908 -18320 42172
rect -18400 41852 -18388 41908
rect -18332 41852 -18320 41908
rect -18400 41840 -18320 41852
rect -18240 42868 -18160 42880
rect -18240 42812 -18228 42868
rect -18172 42812 -18160 42868
rect -18240 42548 -18160 42812
rect -18240 42492 -18228 42548
rect -18172 42492 -18160 42548
rect -18240 42228 -18160 42492
rect -18240 42172 -18228 42228
rect -18172 42172 -18160 42228
rect -18240 41908 -18160 42172
rect -18240 41852 -18228 41908
rect -18172 41852 -18160 41908
rect -18240 41840 -18160 41852
rect -18080 42868 -18000 42880
rect -18080 42812 -18068 42868
rect -18012 42812 -18000 42868
rect -18080 42548 -18000 42812
rect -18080 42492 -18068 42548
rect -18012 42492 -18000 42548
rect -18080 42228 -18000 42492
rect -18080 42172 -18068 42228
rect -18012 42172 -18000 42228
rect -18080 41908 -18000 42172
rect -18080 41852 -18068 41908
rect -18012 41852 -18000 41908
rect -18080 41840 -18000 41852
rect -17920 42868 -17840 42880
rect -17920 42812 -17908 42868
rect -17852 42812 -17840 42868
rect -17920 42548 -17840 42812
rect -17920 42492 -17908 42548
rect -17852 42492 -17840 42548
rect -17920 42228 -17840 42492
rect -17920 42172 -17908 42228
rect -17852 42172 -17840 42228
rect -17920 41908 -17840 42172
rect -17920 41852 -17908 41908
rect -17852 41852 -17840 41908
rect -17920 41840 -17840 41852
rect -17760 42868 -17680 42880
rect -17760 42812 -17748 42868
rect -17692 42812 -17680 42868
rect -17760 42548 -17680 42812
rect -17760 42492 -17748 42548
rect -17692 42492 -17680 42548
rect -17760 42228 -17680 42492
rect -17760 42172 -17748 42228
rect -17692 42172 -17680 42228
rect -17760 41908 -17680 42172
rect -17760 41852 -17748 41908
rect -17692 41852 -17680 41908
rect -17760 41840 -17680 41852
rect -17600 42868 -17520 42880
rect -17600 42812 -17588 42868
rect -17532 42812 -17520 42868
rect -17600 42548 -17520 42812
rect -17600 42492 -17588 42548
rect -17532 42492 -17520 42548
rect -17600 42228 -17520 42492
rect -17600 42172 -17588 42228
rect -17532 42172 -17520 42228
rect -17600 41908 -17520 42172
rect -17600 41852 -17588 41908
rect -17532 41852 -17520 41908
rect -17600 41840 -17520 41852
rect -17440 42868 -17360 42880
rect -17440 42812 -17428 42868
rect -17372 42812 -17360 42868
rect -17440 42548 -17360 42812
rect -17440 42492 -17428 42548
rect -17372 42492 -17360 42548
rect -17440 42228 -17360 42492
rect -17440 42172 -17428 42228
rect -17372 42172 -17360 42228
rect -17440 41908 -17360 42172
rect -17440 41852 -17428 41908
rect -17372 41852 -17360 41908
rect -17440 41840 -17360 41852
rect -17280 42868 -17200 42880
rect -17280 42812 -17268 42868
rect -17212 42812 -17200 42868
rect -17280 42548 -17200 42812
rect -17280 42492 -17268 42548
rect -17212 42492 -17200 42548
rect -17280 42228 -17200 42492
rect -17280 42172 -17268 42228
rect -17212 42172 -17200 42228
rect -17280 41908 -17200 42172
rect -17280 41852 -17268 41908
rect -17212 41852 -17200 41908
rect -17280 41840 -17200 41852
rect -17120 42868 -17040 42880
rect -17120 42812 -17108 42868
rect -17052 42812 -17040 42868
rect -17120 42548 -17040 42812
rect -17120 42492 -17108 42548
rect -17052 42492 -17040 42548
rect -17120 42228 -17040 42492
rect -17120 42172 -17108 42228
rect -17052 42172 -17040 42228
rect -17120 41908 -17040 42172
rect -17120 41852 -17108 41908
rect -17052 41852 -17040 41908
rect -17120 41840 -17040 41852
rect -16960 42868 -16880 42880
rect -16960 42812 -16948 42868
rect -16892 42812 -16880 42868
rect -16960 42548 -16880 42812
rect -16960 42492 -16948 42548
rect -16892 42492 -16880 42548
rect -16960 42228 -16880 42492
rect -16960 42172 -16948 42228
rect -16892 42172 -16880 42228
rect -16960 41908 -16880 42172
rect -16960 41852 -16948 41908
rect -16892 41852 -16880 41908
rect -16960 41840 -16880 41852
rect -16800 42868 -16720 42880
rect -16800 42812 -16788 42868
rect -16732 42812 -16720 42868
rect -16800 42548 -16720 42812
rect -16800 42492 -16788 42548
rect -16732 42492 -16720 42548
rect -16800 42228 -16720 42492
rect -16800 42172 -16788 42228
rect -16732 42172 -16720 42228
rect -16800 41908 -16720 42172
rect -16800 41852 -16788 41908
rect -16732 41852 -16720 41908
rect -16800 41840 -16720 41852
rect -16640 42868 -16560 42880
rect -16640 42812 -16628 42868
rect -16572 42812 -16560 42868
rect -16640 42548 -16560 42812
rect -16640 42492 -16628 42548
rect -16572 42492 -16560 42548
rect -16640 42228 -16560 42492
rect -16640 42172 -16628 42228
rect -16572 42172 -16560 42228
rect -16640 41908 -16560 42172
rect -16640 41852 -16628 41908
rect -16572 41852 -16560 41908
rect -16640 41840 -16560 41852
rect -16480 42868 -16400 42880
rect -16480 42812 -16468 42868
rect -16412 42812 -16400 42868
rect -16480 42548 -16400 42812
rect -16480 42492 -16468 42548
rect -16412 42492 -16400 42548
rect -16480 42228 -16400 42492
rect -16480 42172 -16468 42228
rect -16412 42172 -16400 42228
rect -16480 41908 -16400 42172
rect -16480 41852 -16468 41908
rect -16412 41852 -16400 41908
rect -16480 41840 -16400 41852
rect -16320 42868 -16240 42880
rect -16320 42812 -16308 42868
rect -16252 42812 -16240 42868
rect -16320 42548 -16240 42812
rect -16320 42492 -16308 42548
rect -16252 42492 -16240 42548
rect -16320 42228 -16240 42492
rect -16320 42172 -16308 42228
rect -16252 42172 -16240 42228
rect -16320 41908 -16240 42172
rect -16320 41852 -16308 41908
rect -16252 41852 -16240 41908
rect -16320 41840 -16240 41852
rect -16160 42868 -16080 42880
rect -16160 42812 -16148 42868
rect -16092 42812 -16080 42868
rect -16160 42548 -16080 42812
rect -16160 42492 -16148 42548
rect -16092 42492 -16080 42548
rect -16160 42228 -16080 42492
rect -16160 42172 -16148 42228
rect -16092 42172 -16080 42228
rect -16160 41908 -16080 42172
rect -16160 41852 -16148 41908
rect -16092 41852 -16080 41908
rect -16160 41840 -16080 41852
rect -16000 42868 -15920 42880
rect -16000 42812 -15988 42868
rect -15932 42812 -15920 42868
rect -16000 42548 -15920 42812
rect -16000 42492 -15988 42548
rect -15932 42492 -15920 42548
rect -16000 42228 -15920 42492
rect -16000 42172 -15988 42228
rect -15932 42172 -15920 42228
rect -16000 41908 -15920 42172
rect -16000 41852 -15988 41908
rect -15932 41852 -15920 41908
rect -16000 41840 -15920 41852
rect -15840 42868 -15760 42880
rect -15840 42812 -15828 42868
rect -15772 42812 -15760 42868
rect -15840 42548 -15760 42812
rect -15840 42492 -15828 42548
rect -15772 42492 -15760 42548
rect -15840 42228 -15760 42492
rect -15840 42172 -15828 42228
rect -15772 42172 -15760 42228
rect -15840 41908 -15760 42172
rect -15840 41852 -15828 41908
rect -15772 41852 -15760 41908
rect -15840 41840 -15760 41852
rect -15680 42868 -15600 42880
rect -15680 42812 -15668 42868
rect -15612 42812 -15600 42868
rect -15680 42548 -15600 42812
rect -15680 42492 -15668 42548
rect -15612 42492 -15600 42548
rect -15680 42228 -15600 42492
rect -15680 42172 -15668 42228
rect -15612 42172 -15600 42228
rect -15680 41908 -15600 42172
rect -15680 41852 -15668 41908
rect -15612 41852 -15600 41908
rect -15680 41840 -15600 41852
rect -15520 42868 -15440 42880
rect -15520 42812 -15508 42868
rect -15452 42812 -15440 42868
rect -15520 42548 -15440 42812
rect -15520 42492 -15508 42548
rect -15452 42492 -15440 42548
rect -15520 42228 -15440 42492
rect -15520 42172 -15508 42228
rect -15452 42172 -15440 42228
rect -15520 41908 -15440 42172
rect -15520 41852 -15508 41908
rect -15452 41852 -15440 41908
rect -15520 41840 -15440 41852
rect -15360 42868 -15280 42880
rect -15360 42812 -15348 42868
rect -15292 42812 -15280 42868
rect -15360 42548 -15280 42812
rect -15360 42492 -15348 42548
rect -15292 42492 -15280 42548
rect -15360 42228 -15280 42492
rect -15360 42172 -15348 42228
rect -15292 42172 -15280 42228
rect -15360 41908 -15280 42172
rect -15360 41852 -15348 41908
rect -15292 41852 -15280 41908
rect -15360 41840 -15280 41852
rect -15200 42868 -15120 42880
rect -15200 42812 -15188 42868
rect -15132 42812 -15120 42868
rect -15200 42548 -15120 42812
rect -15200 42492 -15188 42548
rect -15132 42492 -15120 42548
rect -15200 42228 -15120 42492
rect -15200 42172 -15188 42228
rect -15132 42172 -15120 42228
rect -15200 41908 -15120 42172
rect -15200 41852 -15188 41908
rect -15132 41852 -15120 41908
rect -15200 41840 -15120 41852
rect -15040 42868 -14960 42880
rect -15040 42812 -15028 42868
rect -14972 42812 -14960 42868
rect -15040 42548 -14960 42812
rect -15040 42492 -15028 42548
rect -14972 42492 -14960 42548
rect -15040 42228 -14960 42492
rect -15040 42172 -15028 42228
rect -14972 42172 -14960 42228
rect -15040 41908 -14960 42172
rect -15040 41852 -15028 41908
rect -14972 41852 -14960 41908
rect -15040 41840 -14960 41852
rect -14880 42868 -14800 42880
rect -14880 42812 -14868 42868
rect -14812 42812 -14800 42868
rect -14880 42548 -14800 42812
rect -14880 42492 -14868 42548
rect -14812 42492 -14800 42548
rect -14880 42228 -14800 42492
rect -14880 42172 -14868 42228
rect -14812 42172 -14800 42228
rect -14880 41908 -14800 42172
rect -14880 41852 -14868 41908
rect -14812 41852 -14800 41908
rect -14880 41840 -14800 41852
rect -14720 42868 -14640 42880
rect -14720 42812 -14708 42868
rect -14652 42812 -14640 42868
rect -14720 42548 -14640 42812
rect -14720 42492 -14708 42548
rect -14652 42492 -14640 42548
rect -14720 42228 -14640 42492
rect -14720 42172 -14708 42228
rect -14652 42172 -14640 42228
rect -14720 41908 -14640 42172
rect -14720 41852 -14708 41908
rect -14652 41852 -14640 41908
rect -14720 41840 -14640 41852
rect -14560 42868 -14480 42880
rect -14560 42812 -14548 42868
rect -14492 42812 -14480 42868
rect -14560 42548 -14480 42812
rect -14560 42492 -14548 42548
rect -14492 42492 -14480 42548
rect -14560 42228 -14480 42492
rect -14560 42172 -14548 42228
rect -14492 42172 -14480 42228
rect -14560 41908 -14480 42172
rect -14560 41852 -14548 41908
rect -14492 41852 -14480 41908
rect -14560 41840 -14480 41852
rect -14400 42868 -14320 42880
rect -14400 42812 -14388 42868
rect -14332 42812 -14320 42868
rect -14400 42548 -14320 42812
rect -14400 42492 -14388 42548
rect -14332 42492 -14320 42548
rect -14400 42228 -14320 42492
rect -14400 42172 -14388 42228
rect -14332 42172 -14320 42228
rect -14400 41908 -14320 42172
rect -14400 41852 -14388 41908
rect -14332 41852 -14320 41908
rect -14400 41840 -14320 41852
rect -14240 42868 -14160 42880
rect -14240 42812 -14228 42868
rect -14172 42812 -14160 42868
rect -14240 42548 -14160 42812
rect -14240 42492 -14228 42548
rect -14172 42492 -14160 42548
rect -14240 42228 -14160 42492
rect -14240 42172 -14228 42228
rect -14172 42172 -14160 42228
rect -14240 41908 -14160 42172
rect -14240 41852 -14228 41908
rect -14172 41852 -14160 41908
rect -14240 41840 -14160 41852
rect -14080 42868 -14000 42880
rect -14080 42812 -14068 42868
rect -14012 42812 -14000 42868
rect -14080 42548 -14000 42812
rect -14080 42492 -14068 42548
rect -14012 42492 -14000 42548
rect -14080 42228 -14000 42492
rect -14080 42172 -14068 42228
rect -14012 42172 -14000 42228
rect -14080 41908 -14000 42172
rect -14080 41852 -14068 41908
rect -14012 41852 -14000 41908
rect -14080 41840 -14000 41852
rect -13920 42868 -13840 42880
rect -13920 42812 -13908 42868
rect -13852 42812 -13840 42868
rect -13920 42548 -13840 42812
rect -13920 42492 -13908 42548
rect -13852 42492 -13840 42548
rect -13920 42228 -13840 42492
rect -13920 42172 -13908 42228
rect -13852 42172 -13840 42228
rect -13920 41908 -13840 42172
rect -13920 41852 -13908 41908
rect -13852 41852 -13840 41908
rect -13920 41840 -13840 41852
rect -13760 42868 -13680 42880
rect -13760 42812 -13748 42868
rect -13692 42812 -13680 42868
rect -13760 42548 -13680 42812
rect -13760 42492 -13748 42548
rect -13692 42492 -13680 42548
rect -13760 42228 -13680 42492
rect -13760 42172 -13748 42228
rect -13692 42172 -13680 42228
rect -13760 41908 -13680 42172
rect -13760 41852 -13748 41908
rect -13692 41852 -13680 41908
rect -13760 41840 -13680 41852
rect -13600 42868 -13520 42880
rect -13600 42812 -13588 42868
rect -13532 42812 -13520 42868
rect -13600 42548 -13520 42812
rect -13600 42492 -13588 42548
rect -13532 42492 -13520 42548
rect -13600 42228 -13520 42492
rect -13600 42172 -13588 42228
rect -13532 42172 -13520 42228
rect -13600 41908 -13520 42172
rect -13600 41852 -13588 41908
rect -13532 41852 -13520 41908
rect -13600 41840 -13520 41852
rect -13440 42868 -13360 42880
rect -13440 42812 -13428 42868
rect -13372 42812 -13360 42868
rect -13440 42548 -13360 42812
rect -13440 42492 -13428 42548
rect -13372 42492 -13360 42548
rect -13440 42228 -13360 42492
rect -13440 42172 -13428 42228
rect -13372 42172 -13360 42228
rect -13440 41908 -13360 42172
rect -13440 41852 -13428 41908
rect -13372 41852 -13360 41908
rect -13440 41840 -13360 41852
rect -13280 42868 -13200 42880
rect -13280 42812 -13268 42868
rect -13212 42812 -13200 42868
rect -13280 42548 -13200 42812
rect -13280 42492 -13268 42548
rect -13212 42492 -13200 42548
rect -13280 42228 -13200 42492
rect -13280 42172 -13268 42228
rect -13212 42172 -13200 42228
rect -13280 41908 -13200 42172
rect -13280 41852 -13268 41908
rect -13212 41852 -13200 41908
rect -13280 41840 -13200 41852
rect -13120 42868 -13040 42880
rect -13120 42812 -13108 42868
rect -13052 42812 -13040 42868
rect -13120 42548 -13040 42812
rect -13120 42492 -13108 42548
rect -13052 42492 -13040 42548
rect -13120 42228 -13040 42492
rect -13120 42172 -13108 42228
rect -13052 42172 -13040 42228
rect -13120 41908 -13040 42172
rect -13120 41852 -13108 41908
rect -13052 41852 -13040 41908
rect -13120 41840 -13040 41852
rect -12960 42868 -12880 42880
rect -12960 42812 -12948 42868
rect -12892 42812 -12880 42868
rect -12960 42548 -12880 42812
rect -12960 42492 -12948 42548
rect -12892 42492 -12880 42548
rect -12960 42228 -12880 42492
rect -12960 42172 -12948 42228
rect -12892 42172 -12880 42228
rect -12960 41908 -12880 42172
rect -12960 41852 -12948 41908
rect -12892 41852 -12880 41908
rect -12960 41840 -12880 41852
rect -12800 42868 -12720 42880
rect -12800 42812 -12788 42868
rect -12732 42812 -12720 42868
rect -12800 42548 -12720 42812
rect -12800 42492 -12788 42548
rect -12732 42492 -12720 42548
rect -12800 42228 -12720 42492
rect -12800 42172 -12788 42228
rect -12732 42172 -12720 42228
rect -12800 41908 -12720 42172
rect -12800 41852 -12788 41908
rect -12732 41852 -12720 41908
rect -12800 41840 -12720 41852
rect -12640 42868 -12560 42880
rect -12640 42812 -12628 42868
rect -12572 42812 -12560 42868
rect -12640 42548 -12560 42812
rect -12640 42492 -12628 42548
rect -12572 42492 -12560 42548
rect -12640 42228 -12560 42492
rect -12640 42172 -12628 42228
rect -12572 42172 -12560 42228
rect -12640 41908 -12560 42172
rect -12640 41852 -12628 41908
rect -12572 41852 -12560 41908
rect -12640 41840 -12560 41852
rect -12480 42868 -12400 42880
rect -12480 42812 -12468 42868
rect -12412 42812 -12400 42868
rect -12480 42548 -12400 42812
rect -12480 42492 -12468 42548
rect -12412 42492 -12400 42548
rect -12480 42228 -12400 42492
rect -12480 42172 -12468 42228
rect -12412 42172 -12400 42228
rect -12480 41908 -12400 42172
rect -12480 41852 -12468 41908
rect -12412 41852 -12400 41908
rect -12480 41840 -12400 41852
rect -12320 42868 -12240 42880
rect -12320 42812 -12308 42868
rect -12252 42812 -12240 42868
rect -12320 42548 -12240 42812
rect -12320 42492 -12308 42548
rect -12252 42492 -12240 42548
rect -12320 42228 -12240 42492
rect -12320 42172 -12308 42228
rect -12252 42172 -12240 42228
rect -12320 41908 -12240 42172
rect -12320 41852 -12308 41908
rect -12252 41852 -12240 41908
rect -12320 41840 -12240 41852
rect -12160 42868 -12080 42880
rect -12160 42812 -12148 42868
rect -12092 42812 -12080 42868
rect -12160 42548 -12080 42812
rect -11840 42868 -11760 42880
rect -11840 42812 -11828 42868
rect -11772 42812 -11760 42868
rect -12160 42492 -12148 42548
rect -12092 42492 -12080 42548
rect -12160 42228 -12080 42492
rect -12160 42172 -12148 42228
rect -12092 42172 -12080 42228
rect -12160 41908 -12080 42172
rect -12160 41852 -12148 41908
rect -12092 41852 -12080 41908
rect -30080 41688 -30072 41752
rect -30008 41688 -30000 41752
rect -30080 41592 -30000 41688
rect -30080 41528 -30072 41592
rect -30008 41528 -30000 41592
rect -30080 40792 -30000 41528
rect -12160 41748 -12080 41852
rect -12160 41692 -12148 41748
rect -12092 41692 -12080 41748
rect -12160 41588 -12080 41692
rect -12160 41532 -12148 41588
rect -12092 41532 -12080 41588
rect -29920 41348 -29840 41360
rect -29920 41292 -29908 41348
rect -29852 41292 -29840 41348
rect -29920 41028 -29840 41292
rect -29920 40972 -29908 41028
rect -29852 40972 -29840 41028
rect -29920 40960 -29840 40972
rect -29760 41348 -29680 41360
rect -29760 41292 -29748 41348
rect -29692 41292 -29680 41348
rect -29760 41028 -29680 41292
rect -29760 40972 -29748 41028
rect -29692 40972 -29680 41028
rect -29760 40960 -29680 40972
rect -29600 41348 -29520 41360
rect -29600 41292 -29588 41348
rect -29532 41292 -29520 41348
rect -29600 41028 -29520 41292
rect -29600 40972 -29588 41028
rect -29532 40972 -29520 41028
rect -29600 40960 -29520 40972
rect -29440 41348 -29360 41360
rect -29440 41292 -29428 41348
rect -29372 41292 -29360 41348
rect -29440 41028 -29360 41292
rect -29440 40972 -29428 41028
rect -29372 40972 -29360 41028
rect -29440 40960 -29360 40972
rect -29280 41348 -29200 41360
rect -29280 41292 -29268 41348
rect -29212 41292 -29200 41348
rect -29280 41028 -29200 41292
rect -29280 40972 -29268 41028
rect -29212 40972 -29200 41028
rect -29280 40960 -29200 40972
rect -29120 41348 -29040 41360
rect -29120 41292 -29108 41348
rect -29052 41292 -29040 41348
rect -29120 41028 -29040 41292
rect -29120 40972 -29108 41028
rect -29052 40972 -29040 41028
rect -29120 40960 -29040 40972
rect -28960 41348 -28880 41360
rect -28960 41292 -28948 41348
rect -28892 41292 -28880 41348
rect -28960 41028 -28880 41292
rect -28960 40972 -28948 41028
rect -28892 40972 -28880 41028
rect -28960 40960 -28880 40972
rect -28800 41348 -28720 41360
rect -28800 41292 -28788 41348
rect -28732 41292 -28720 41348
rect -28800 41028 -28720 41292
rect -28800 40972 -28788 41028
rect -28732 40972 -28720 41028
rect -28800 40960 -28720 40972
rect -28640 41348 -28560 41360
rect -28640 41292 -28628 41348
rect -28572 41292 -28560 41348
rect -28640 41028 -28560 41292
rect -28640 40972 -28628 41028
rect -28572 40972 -28560 41028
rect -28640 40960 -28560 40972
rect -28480 41348 -28400 41360
rect -28480 41292 -28468 41348
rect -28412 41292 -28400 41348
rect -28480 41028 -28400 41292
rect -28480 40972 -28468 41028
rect -28412 40972 -28400 41028
rect -28480 40960 -28400 40972
rect -28320 41348 -28240 41360
rect -28320 41292 -28308 41348
rect -28252 41292 -28240 41348
rect -28320 41028 -28240 41292
rect -28320 40972 -28308 41028
rect -28252 40972 -28240 41028
rect -28320 40960 -28240 40972
rect -28160 41348 -28080 41360
rect -28160 41292 -28148 41348
rect -28092 41292 -28080 41348
rect -28160 41028 -28080 41292
rect -28160 40972 -28148 41028
rect -28092 40972 -28080 41028
rect -28160 40960 -28080 40972
rect -28000 41348 -27920 41360
rect -28000 41292 -27988 41348
rect -27932 41292 -27920 41348
rect -28000 41028 -27920 41292
rect -28000 40972 -27988 41028
rect -27932 40972 -27920 41028
rect -28000 40960 -27920 40972
rect -27840 41348 -27760 41360
rect -27840 41292 -27828 41348
rect -27772 41292 -27760 41348
rect -27840 41028 -27760 41292
rect -27840 40972 -27828 41028
rect -27772 40972 -27760 41028
rect -27840 40960 -27760 40972
rect -27680 41348 -27600 41360
rect -27680 41292 -27668 41348
rect -27612 41292 -27600 41348
rect -27680 41028 -27600 41292
rect -27680 40972 -27668 41028
rect -27612 40972 -27600 41028
rect -27680 40960 -27600 40972
rect -27520 41348 -27440 41360
rect -27520 41292 -27508 41348
rect -27452 41292 -27440 41348
rect -27520 41028 -27440 41292
rect -27520 40972 -27508 41028
rect -27452 40972 -27440 41028
rect -27520 40960 -27440 40972
rect -27360 41348 -27280 41360
rect -27360 41292 -27348 41348
rect -27292 41292 -27280 41348
rect -27360 41028 -27280 41292
rect -27360 40972 -27348 41028
rect -27292 40972 -27280 41028
rect -27360 40960 -27280 40972
rect -27200 41348 -27120 41360
rect -27200 41292 -27188 41348
rect -27132 41292 -27120 41348
rect -27200 41028 -27120 41292
rect -27200 40972 -27188 41028
rect -27132 40972 -27120 41028
rect -27200 40960 -27120 40972
rect -27040 41348 -26960 41360
rect -27040 41292 -27028 41348
rect -26972 41292 -26960 41348
rect -27040 41028 -26960 41292
rect -27040 40972 -27028 41028
rect -26972 40972 -26960 41028
rect -27040 40960 -26960 40972
rect -26880 41348 -26800 41360
rect -26880 41292 -26868 41348
rect -26812 41292 -26800 41348
rect -26880 41028 -26800 41292
rect -26880 40972 -26868 41028
rect -26812 40972 -26800 41028
rect -26880 40960 -26800 40972
rect -26720 41348 -26640 41360
rect -26720 41292 -26708 41348
rect -26652 41292 -26640 41348
rect -26720 41028 -26640 41292
rect -26720 40972 -26708 41028
rect -26652 40972 -26640 41028
rect -26720 40960 -26640 40972
rect -26560 41348 -26480 41360
rect -26560 41292 -26548 41348
rect -26492 41292 -26480 41348
rect -26560 41028 -26480 41292
rect -26560 40972 -26548 41028
rect -26492 40972 -26480 41028
rect -26560 40960 -26480 40972
rect -26400 41348 -26320 41360
rect -26400 41292 -26388 41348
rect -26332 41292 -26320 41348
rect -26400 41028 -26320 41292
rect -26400 40972 -26388 41028
rect -26332 40972 -26320 41028
rect -26400 40960 -26320 40972
rect -26240 41348 -26160 41360
rect -26240 41292 -26228 41348
rect -26172 41292 -26160 41348
rect -26240 41028 -26160 41292
rect -26240 40972 -26228 41028
rect -26172 40972 -26160 41028
rect -26240 40960 -26160 40972
rect -26080 41348 -26000 41360
rect -26080 41292 -26068 41348
rect -26012 41292 -26000 41348
rect -26080 41028 -26000 41292
rect -26080 40972 -26068 41028
rect -26012 40972 -26000 41028
rect -26080 40960 -26000 40972
rect -25920 41348 -25840 41360
rect -25920 41292 -25908 41348
rect -25852 41292 -25840 41348
rect -25920 41028 -25840 41292
rect -25920 40972 -25908 41028
rect -25852 40972 -25840 41028
rect -25920 40960 -25840 40972
rect -25760 41348 -25680 41360
rect -25760 41292 -25748 41348
rect -25692 41292 -25680 41348
rect -25760 41028 -25680 41292
rect -25760 40972 -25748 41028
rect -25692 40972 -25680 41028
rect -25760 40960 -25680 40972
rect -25600 41348 -25520 41360
rect -25600 41292 -25588 41348
rect -25532 41292 -25520 41348
rect -25600 41028 -25520 41292
rect -25600 40972 -25588 41028
rect -25532 40972 -25520 41028
rect -25600 40960 -25520 40972
rect -25440 41348 -25360 41360
rect -25440 41292 -25428 41348
rect -25372 41292 -25360 41348
rect -25440 41028 -25360 41292
rect -25440 40972 -25428 41028
rect -25372 40972 -25360 41028
rect -25440 40960 -25360 40972
rect -25280 41348 -25200 41360
rect -25280 41292 -25268 41348
rect -25212 41292 -25200 41348
rect -25280 41028 -25200 41292
rect -25280 40972 -25268 41028
rect -25212 40972 -25200 41028
rect -25280 40960 -25200 40972
rect -25120 41348 -25040 41360
rect -25120 41292 -25108 41348
rect -25052 41292 -25040 41348
rect -25120 41028 -25040 41292
rect -25120 40972 -25108 41028
rect -25052 40972 -25040 41028
rect -25120 40960 -25040 40972
rect -24960 41348 -24880 41360
rect -24960 41292 -24948 41348
rect -24892 41292 -24880 41348
rect -24960 41028 -24880 41292
rect -24960 40972 -24948 41028
rect -24892 40972 -24880 41028
rect -24960 40960 -24880 40972
rect -24800 41348 -24720 41360
rect -24800 41292 -24788 41348
rect -24732 41292 -24720 41348
rect -24800 41028 -24720 41292
rect -24800 40972 -24788 41028
rect -24732 40972 -24720 41028
rect -24800 40960 -24720 40972
rect -24640 41348 -24560 41360
rect -24640 41292 -24628 41348
rect -24572 41292 -24560 41348
rect -24640 41028 -24560 41292
rect -24640 40972 -24628 41028
rect -24572 40972 -24560 41028
rect -24640 40960 -24560 40972
rect -24480 41348 -24400 41360
rect -24480 41292 -24468 41348
rect -24412 41292 -24400 41348
rect -24480 41028 -24400 41292
rect -24480 40972 -24468 41028
rect -24412 40972 -24400 41028
rect -24480 40960 -24400 40972
rect -24320 41348 -24240 41360
rect -24320 41292 -24308 41348
rect -24252 41292 -24240 41348
rect -24320 41028 -24240 41292
rect -24320 40972 -24308 41028
rect -24252 40972 -24240 41028
rect -24320 40960 -24240 40972
rect -24160 41348 -24080 41360
rect -24160 41292 -24148 41348
rect -24092 41292 -24080 41348
rect -24160 41028 -24080 41292
rect -24160 40972 -24148 41028
rect -24092 40972 -24080 41028
rect -24160 40960 -24080 40972
rect -24000 41348 -23920 41360
rect -24000 41292 -23988 41348
rect -23932 41292 -23920 41348
rect -24000 41028 -23920 41292
rect -24000 40972 -23988 41028
rect -23932 40972 -23920 41028
rect -24000 40960 -23920 40972
rect -23840 41348 -23760 41360
rect -23840 41292 -23828 41348
rect -23772 41292 -23760 41348
rect -23840 41028 -23760 41292
rect -23840 40972 -23828 41028
rect -23772 40972 -23760 41028
rect -23840 40960 -23760 40972
rect -23680 41348 -23600 41360
rect -23680 41292 -23668 41348
rect -23612 41292 -23600 41348
rect -23680 41028 -23600 41292
rect -23680 40972 -23668 41028
rect -23612 40972 -23600 41028
rect -23680 40960 -23600 40972
rect -23520 41348 -23440 41360
rect -23520 41292 -23508 41348
rect -23452 41292 -23440 41348
rect -23520 41028 -23440 41292
rect -23520 40972 -23508 41028
rect -23452 40972 -23440 41028
rect -23520 40960 -23440 40972
rect -23360 41348 -23280 41360
rect -23360 41292 -23348 41348
rect -23292 41292 -23280 41348
rect -23360 41028 -23280 41292
rect -23360 40972 -23348 41028
rect -23292 40972 -23280 41028
rect -23360 40960 -23280 40972
rect -23200 41348 -23120 41360
rect -23200 41292 -23188 41348
rect -23132 41292 -23120 41348
rect -23200 41028 -23120 41292
rect -23200 40972 -23188 41028
rect -23132 40972 -23120 41028
rect -23200 40960 -23120 40972
rect -23040 41348 -22960 41360
rect -23040 41292 -23028 41348
rect -22972 41292 -22960 41348
rect -23040 41028 -22960 41292
rect -23040 40972 -23028 41028
rect -22972 40972 -22960 41028
rect -23040 40960 -22960 40972
rect -22880 41348 -22800 41360
rect -22880 41292 -22868 41348
rect -22812 41292 -22800 41348
rect -22880 41028 -22800 41292
rect -22880 40972 -22868 41028
rect -22812 40972 -22800 41028
rect -22880 40960 -22800 40972
rect -22720 41348 -22640 41360
rect -22720 41292 -22708 41348
rect -22652 41292 -22640 41348
rect -22720 41028 -22640 41292
rect -22720 40972 -22708 41028
rect -22652 40972 -22640 41028
rect -22720 40960 -22640 40972
rect -22560 41348 -22480 41360
rect -22560 41292 -22548 41348
rect -22492 41292 -22480 41348
rect -22560 41028 -22480 41292
rect -22560 40972 -22548 41028
rect -22492 40972 -22480 41028
rect -22560 40960 -22480 40972
rect -22400 41348 -22320 41360
rect -22400 41292 -22388 41348
rect -22332 41292 -22320 41348
rect -22400 41028 -22320 41292
rect -22400 40972 -22388 41028
rect -22332 40972 -22320 41028
rect -22400 40960 -22320 40972
rect -22240 41348 -22160 41360
rect -22240 41292 -22228 41348
rect -22172 41292 -22160 41348
rect -22240 41028 -22160 41292
rect -22240 40972 -22228 41028
rect -22172 40972 -22160 41028
rect -22240 40960 -22160 40972
rect -22080 41348 -22000 41360
rect -22080 41292 -22068 41348
rect -22012 41292 -22000 41348
rect -22080 41028 -22000 41292
rect -22080 40972 -22068 41028
rect -22012 40972 -22000 41028
rect -22080 40960 -22000 40972
rect -21920 41348 -21840 41360
rect -21920 41292 -21908 41348
rect -21852 41292 -21840 41348
rect -21920 41028 -21840 41292
rect -21920 40972 -21908 41028
rect -21852 40972 -21840 41028
rect -21920 40960 -21840 40972
rect -21760 41348 -21680 41360
rect -21760 41292 -21748 41348
rect -21692 41292 -21680 41348
rect -21760 41028 -21680 41292
rect -21760 40972 -21748 41028
rect -21692 40972 -21680 41028
rect -21760 40960 -21680 40972
rect -21600 41348 -21520 41360
rect -21600 41292 -21588 41348
rect -21532 41292 -21520 41348
rect -21600 41028 -21520 41292
rect -21600 40972 -21588 41028
rect -21532 40972 -21520 41028
rect -21600 40960 -21520 40972
rect -21440 41348 -21360 41360
rect -21440 41292 -21428 41348
rect -21372 41292 -21360 41348
rect -21440 41028 -21360 41292
rect -21440 40972 -21428 41028
rect -21372 40972 -21360 41028
rect -21440 40960 -21360 40972
rect -21280 41348 -21200 41360
rect -21280 41292 -21268 41348
rect -21212 41292 -21200 41348
rect -21280 41028 -21200 41292
rect -21280 40972 -21268 41028
rect -21212 40972 -21200 41028
rect -21280 40960 -21200 40972
rect -21120 41348 -21040 41360
rect -21120 41292 -21108 41348
rect -21052 41292 -21040 41348
rect -21120 41028 -21040 41292
rect -21120 40972 -21108 41028
rect -21052 40972 -21040 41028
rect -21120 40960 -21040 40972
rect -20960 41348 -20880 41360
rect -20960 41292 -20948 41348
rect -20892 41292 -20880 41348
rect -20960 41028 -20880 41292
rect -20960 40972 -20948 41028
rect -20892 40972 -20880 41028
rect -20960 40960 -20880 40972
rect -20800 41348 -20720 41360
rect -20800 41292 -20788 41348
rect -20732 41292 -20720 41348
rect -20800 41028 -20720 41292
rect -20800 40972 -20788 41028
rect -20732 40972 -20720 41028
rect -20800 40960 -20720 40972
rect -20640 41348 -20560 41360
rect -20640 41292 -20628 41348
rect -20572 41292 -20560 41348
rect -20640 41028 -20560 41292
rect -20640 40972 -20628 41028
rect -20572 40972 -20560 41028
rect -20640 40960 -20560 40972
rect -20480 41348 -20400 41360
rect -20480 41292 -20468 41348
rect -20412 41292 -20400 41348
rect -20480 41028 -20400 41292
rect -20480 40972 -20468 41028
rect -20412 40972 -20400 41028
rect -20480 40960 -20400 40972
rect -20320 41348 -20240 41360
rect -20320 41292 -20308 41348
rect -20252 41292 -20240 41348
rect -20320 41028 -20240 41292
rect -20320 40972 -20308 41028
rect -20252 40972 -20240 41028
rect -20320 40960 -20240 40972
rect -20160 41348 -20080 41360
rect -20160 41292 -20148 41348
rect -20092 41292 -20080 41348
rect -20160 41028 -20080 41292
rect -20160 40972 -20148 41028
rect -20092 40972 -20080 41028
rect -20160 40960 -20080 40972
rect -20000 41348 -19920 41360
rect -20000 41292 -19988 41348
rect -19932 41292 -19920 41348
rect -20000 41028 -19920 41292
rect -20000 40972 -19988 41028
rect -19932 40972 -19920 41028
rect -20000 40960 -19920 40972
rect -19840 41348 -19760 41360
rect -19840 41292 -19828 41348
rect -19772 41292 -19760 41348
rect -19840 41028 -19760 41292
rect -19840 40972 -19828 41028
rect -19772 40972 -19760 41028
rect -19840 40960 -19760 40972
rect -19680 41348 -19600 41360
rect -19680 41292 -19668 41348
rect -19612 41292 -19600 41348
rect -19680 41028 -19600 41292
rect -19680 40972 -19668 41028
rect -19612 40972 -19600 41028
rect -19680 40960 -19600 40972
rect -19520 41348 -19440 41360
rect -19520 41292 -19508 41348
rect -19452 41292 -19440 41348
rect -19520 41028 -19440 41292
rect -19520 40972 -19508 41028
rect -19452 40972 -19440 41028
rect -19520 40960 -19440 40972
rect -19360 41348 -19280 41360
rect -19360 41292 -19348 41348
rect -19292 41292 -19280 41348
rect -19360 41028 -19280 41292
rect -19360 40972 -19348 41028
rect -19292 40972 -19280 41028
rect -19360 40960 -19280 40972
rect -19200 41348 -19120 41360
rect -19200 41292 -19188 41348
rect -19132 41292 -19120 41348
rect -19200 41028 -19120 41292
rect -19200 40972 -19188 41028
rect -19132 40972 -19120 41028
rect -19200 40960 -19120 40972
rect -19040 41348 -18960 41360
rect -19040 41292 -19028 41348
rect -18972 41292 -18960 41348
rect -19040 41028 -18960 41292
rect -19040 40972 -19028 41028
rect -18972 40972 -18960 41028
rect -19040 40960 -18960 40972
rect -18880 41348 -18800 41360
rect -18880 41292 -18868 41348
rect -18812 41292 -18800 41348
rect -18880 41028 -18800 41292
rect -18880 40972 -18868 41028
rect -18812 40972 -18800 41028
rect -18880 40960 -18800 40972
rect -18720 41348 -18640 41360
rect -18720 41292 -18708 41348
rect -18652 41292 -18640 41348
rect -18720 41028 -18640 41292
rect -18720 40972 -18708 41028
rect -18652 40972 -18640 41028
rect -18720 40960 -18640 40972
rect -18560 41348 -18480 41360
rect -18560 41292 -18548 41348
rect -18492 41292 -18480 41348
rect -18560 41028 -18480 41292
rect -18560 40972 -18548 41028
rect -18492 40972 -18480 41028
rect -18560 40960 -18480 40972
rect -18400 41348 -18320 41360
rect -18400 41292 -18388 41348
rect -18332 41292 -18320 41348
rect -18400 41028 -18320 41292
rect -18400 40972 -18388 41028
rect -18332 40972 -18320 41028
rect -18400 40960 -18320 40972
rect -18240 41348 -18160 41360
rect -18240 41292 -18228 41348
rect -18172 41292 -18160 41348
rect -18240 41028 -18160 41292
rect -18240 40972 -18228 41028
rect -18172 40972 -18160 41028
rect -18240 40960 -18160 40972
rect -18080 41348 -18000 41360
rect -18080 41292 -18068 41348
rect -18012 41292 -18000 41348
rect -18080 41028 -18000 41292
rect -18080 40972 -18068 41028
rect -18012 40972 -18000 41028
rect -18080 40960 -18000 40972
rect -17920 41348 -17840 41360
rect -17920 41292 -17908 41348
rect -17852 41292 -17840 41348
rect -17920 41028 -17840 41292
rect -17920 40972 -17908 41028
rect -17852 40972 -17840 41028
rect -17920 40960 -17840 40972
rect -17760 41348 -17680 41360
rect -17760 41292 -17748 41348
rect -17692 41292 -17680 41348
rect -17760 41028 -17680 41292
rect -17760 40972 -17748 41028
rect -17692 40972 -17680 41028
rect -17760 40960 -17680 40972
rect -17600 41348 -17520 41360
rect -17600 41292 -17588 41348
rect -17532 41292 -17520 41348
rect -17600 41028 -17520 41292
rect -17600 40972 -17588 41028
rect -17532 40972 -17520 41028
rect -17600 40960 -17520 40972
rect -17440 41348 -17360 41360
rect -17440 41292 -17428 41348
rect -17372 41292 -17360 41348
rect -17440 41028 -17360 41292
rect -17440 40972 -17428 41028
rect -17372 40972 -17360 41028
rect -17440 40960 -17360 40972
rect -17280 41348 -17200 41360
rect -17280 41292 -17268 41348
rect -17212 41292 -17200 41348
rect -17280 41028 -17200 41292
rect -17280 40972 -17268 41028
rect -17212 40972 -17200 41028
rect -17280 40960 -17200 40972
rect -17120 41348 -17040 41360
rect -17120 41292 -17108 41348
rect -17052 41292 -17040 41348
rect -17120 41028 -17040 41292
rect -17120 40972 -17108 41028
rect -17052 40972 -17040 41028
rect -17120 40960 -17040 40972
rect -16960 41348 -16880 41360
rect -16960 41292 -16948 41348
rect -16892 41292 -16880 41348
rect -16960 41028 -16880 41292
rect -16960 40972 -16948 41028
rect -16892 40972 -16880 41028
rect -16960 40960 -16880 40972
rect -16800 41348 -16720 41360
rect -16800 41292 -16788 41348
rect -16732 41292 -16720 41348
rect -16800 41028 -16720 41292
rect -16800 40972 -16788 41028
rect -16732 40972 -16720 41028
rect -16800 40960 -16720 40972
rect -16640 41348 -16560 41360
rect -16640 41292 -16628 41348
rect -16572 41292 -16560 41348
rect -16640 41028 -16560 41292
rect -16640 40972 -16628 41028
rect -16572 40972 -16560 41028
rect -16640 40960 -16560 40972
rect -16480 41348 -16400 41360
rect -16480 41292 -16468 41348
rect -16412 41292 -16400 41348
rect -16480 41028 -16400 41292
rect -16480 40972 -16468 41028
rect -16412 40972 -16400 41028
rect -16480 40960 -16400 40972
rect -16320 41348 -16240 41360
rect -16320 41292 -16308 41348
rect -16252 41292 -16240 41348
rect -16320 41028 -16240 41292
rect -16320 40972 -16308 41028
rect -16252 40972 -16240 41028
rect -16320 40960 -16240 40972
rect -16160 41348 -16080 41360
rect -16160 41292 -16148 41348
rect -16092 41292 -16080 41348
rect -16160 41028 -16080 41292
rect -16160 40972 -16148 41028
rect -16092 40972 -16080 41028
rect -16160 40960 -16080 40972
rect -16000 41348 -15920 41360
rect -16000 41292 -15988 41348
rect -15932 41292 -15920 41348
rect -16000 41028 -15920 41292
rect -16000 40972 -15988 41028
rect -15932 40972 -15920 41028
rect -16000 40960 -15920 40972
rect -15840 41348 -15760 41360
rect -15840 41292 -15828 41348
rect -15772 41292 -15760 41348
rect -15840 41028 -15760 41292
rect -15840 40972 -15828 41028
rect -15772 40972 -15760 41028
rect -15840 40960 -15760 40972
rect -15680 41348 -15600 41360
rect -15680 41292 -15668 41348
rect -15612 41292 -15600 41348
rect -15680 41028 -15600 41292
rect -15680 40972 -15668 41028
rect -15612 40972 -15600 41028
rect -15680 40960 -15600 40972
rect -15520 41348 -15440 41360
rect -15520 41292 -15508 41348
rect -15452 41292 -15440 41348
rect -15520 41028 -15440 41292
rect -15520 40972 -15508 41028
rect -15452 40972 -15440 41028
rect -15520 40960 -15440 40972
rect -15360 41348 -15280 41360
rect -15360 41292 -15348 41348
rect -15292 41292 -15280 41348
rect -15360 41028 -15280 41292
rect -15360 40972 -15348 41028
rect -15292 40972 -15280 41028
rect -15360 40960 -15280 40972
rect -15200 41348 -15120 41360
rect -15200 41292 -15188 41348
rect -15132 41292 -15120 41348
rect -15200 41028 -15120 41292
rect -15200 40972 -15188 41028
rect -15132 40972 -15120 41028
rect -15200 40960 -15120 40972
rect -15040 41348 -14960 41360
rect -15040 41292 -15028 41348
rect -14972 41292 -14960 41348
rect -15040 41028 -14960 41292
rect -15040 40972 -15028 41028
rect -14972 40972 -14960 41028
rect -15040 40960 -14960 40972
rect -14880 41348 -14800 41360
rect -14880 41292 -14868 41348
rect -14812 41292 -14800 41348
rect -14880 41028 -14800 41292
rect -14880 40972 -14868 41028
rect -14812 40972 -14800 41028
rect -14880 40960 -14800 40972
rect -14720 41348 -14640 41360
rect -14720 41292 -14708 41348
rect -14652 41292 -14640 41348
rect -14720 41028 -14640 41292
rect -14720 40972 -14708 41028
rect -14652 40972 -14640 41028
rect -14720 40960 -14640 40972
rect -14560 41348 -14480 41360
rect -14560 41292 -14548 41348
rect -14492 41292 -14480 41348
rect -14560 41028 -14480 41292
rect -14560 40972 -14548 41028
rect -14492 40972 -14480 41028
rect -14560 40960 -14480 40972
rect -14400 41348 -14320 41360
rect -14400 41292 -14388 41348
rect -14332 41292 -14320 41348
rect -14400 41028 -14320 41292
rect -14400 40972 -14388 41028
rect -14332 40972 -14320 41028
rect -14400 40960 -14320 40972
rect -14240 41348 -14160 41360
rect -14240 41292 -14228 41348
rect -14172 41292 -14160 41348
rect -14240 41028 -14160 41292
rect -14240 40972 -14228 41028
rect -14172 40972 -14160 41028
rect -14240 40960 -14160 40972
rect -14080 41348 -14000 41360
rect -14080 41292 -14068 41348
rect -14012 41292 -14000 41348
rect -14080 41028 -14000 41292
rect -14080 40972 -14068 41028
rect -14012 40972 -14000 41028
rect -14080 40960 -14000 40972
rect -13920 41348 -13840 41360
rect -13920 41292 -13908 41348
rect -13852 41292 -13840 41348
rect -13920 41028 -13840 41292
rect -13920 40972 -13908 41028
rect -13852 40972 -13840 41028
rect -13920 40960 -13840 40972
rect -13760 41348 -13680 41360
rect -13760 41292 -13748 41348
rect -13692 41292 -13680 41348
rect -13760 41028 -13680 41292
rect -13760 40972 -13748 41028
rect -13692 40972 -13680 41028
rect -13760 40960 -13680 40972
rect -13600 41348 -13520 41360
rect -13600 41292 -13588 41348
rect -13532 41292 -13520 41348
rect -13600 41028 -13520 41292
rect -13600 40972 -13588 41028
rect -13532 40972 -13520 41028
rect -13600 40960 -13520 40972
rect -13440 41348 -13360 41360
rect -13440 41292 -13428 41348
rect -13372 41292 -13360 41348
rect -13440 41028 -13360 41292
rect -13440 40972 -13428 41028
rect -13372 40972 -13360 41028
rect -13440 40960 -13360 40972
rect -13280 41348 -13200 41360
rect -13280 41292 -13268 41348
rect -13212 41292 -13200 41348
rect -13280 41028 -13200 41292
rect -13280 40972 -13268 41028
rect -13212 40972 -13200 41028
rect -13280 40960 -13200 40972
rect -13120 41348 -13040 41360
rect -13120 41292 -13108 41348
rect -13052 41292 -13040 41348
rect -13120 41028 -13040 41292
rect -13120 40972 -13108 41028
rect -13052 40972 -13040 41028
rect -13120 40960 -13040 40972
rect -12960 41348 -12880 41360
rect -12960 41292 -12948 41348
rect -12892 41292 -12880 41348
rect -12960 41028 -12880 41292
rect -12960 40972 -12948 41028
rect -12892 40972 -12880 41028
rect -12960 40960 -12880 40972
rect -12800 41348 -12720 41360
rect -12800 41292 -12788 41348
rect -12732 41292 -12720 41348
rect -12800 41028 -12720 41292
rect -12800 40972 -12788 41028
rect -12732 40972 -12720 41028
rect -12800 40960 -12720 40972
rect -12640 41348 -12560 41360
rect -12640 41292 -12628 41348
rect -12572 41292 -12560 41348
rect -12640 41028 -12560 41292
rect -12640 40972 -12628 41028
rect -12572 40972 -12560 41028
rect -12640 40960 -12560 40972
rect -12480 41348 -12400 41360
rect -12480 41292 -12468 41348
rect -12412 41292 -12400 41348
rect -12480 41028 -12400 41292
rect -12480 40972 -12468 41028
rect -12412 40972 -12400 41028
rect -12480 40960 -12400 40972
rect -12320 41348 -12240 41360
rect -12320 41292 -12308 41348
rect -12252 41292 -12240 41348
rect -12320 41028 -12240 41292
rect -12320 40972 -12308 41028
rect -12252 40972 -12240 41028
rect -12320 40960 -12240 40972
rect -30080 40728 -30072 40792
rect -30008 40728 -30000 40792
rect -30080 40632 -30000 40728
rect -30080 40568 -30072 40632
rect -30008 40568 -30000 40632
rect -30080 40472 -30000 40568
rect -30080 40408 -30072 40472
rect -30008 40408 -30000 40472
rect -30080 40312 -30000 40408
rect -12160 40868 -12080 41532
rect -12160 40812 -12148 40868
rect -12092 40812 -12080 40868
rect -12160 40708 -12080 40812
rect -12160 40652 -12148 40708
rect -12092 40652 -12080 40708
rect -12160 40388 -12080 40652
rect -12160 40332 -12148 40388
rect -12092 40332 -12080 40388
rect -12160 40320 -12080 40332
rect -12000 42708 -11920 42720
rect -12000 42652 -11988 42708
rect -11932 42652 -11920 42708
rect -30080 40248 -30072 40312
rect -30008 40248 -30000 40312
rect -30080 40152 -30000 40248
rect -30080 40088 -30072 40152
rect -30008 40088 -30000 40152
rect -30080 39992 -30000 40088
rect -30080 39928 -30072 39992
rect -30008 39928 -30000 39992
rect -30080 39832 -30000 39928
rect -12000 39920 -11920 42652
rect -11840 42548 -11760 42812
rect -11840 42492 -11828 42548
rect -11772 42492 -11760 42548
rect -11840 42228 -11760 42492
rect -11520 42868 -11440 42880
rect -11520 42812 -11508 42868
rect -11452 42812 -11440 42868
rect -11520 42548 -11440 42812
rect -11520 42492 -11508 42548
rect -11452 42492 -11440 42548
rect -11840 42172 -11828 42228
rect -11772 42172 -11760 42228
rect -11840 41908 -11760 42172
rect -11840 41852 -11828 41908
rect -11772 41852 -11760 41908
rect -11840 41748 -11760 41852
rect -11840 41692 -11828 41748
rect -11772 41692 -11760 41748
rect -11840 41588 -11760 41692
rect -11840 41532 -11828 41588
rect -11772 41532 -11760 41588
rect -11840 40868 -11760 41532
rect -11840 40812 -11828 40868
rect -11772 40812 -11760 40868
rect -11840 40708 -11760 40812
rect -11840 40652 -11828 40708
rect -11772 40652 -11760 40708
rect -11840 40388 -11760 40652
rect -11840 40332 -11828 40388
rect -11772 40332 -11760 40388
rect -11840 40320 -11760 40332
rect -11680 42388 -11600 42400
rect -11680 42332 -11668 42388
rect -11612 42332 -11600 42388
rect -11680 39920 -11600 42332
rect -11520 42228 -11440 42492
rect -11520 42172 -11508 42228
rect -11452 42172 -11440 42228
rect -11520 41908 -11440 42172
rect -11520 41852 -11508 41908
rect -11452 41852 -11440 41908
rect -11520 41748 -11440 41852
rect -11360 42868 -11280 42880
rect -11360 42812 -11348 42868
rect -11292 42812 -11280 42868
rect -11360 42548 -11280 42812
rect -11360 42492 -11348 42548
rect -11292 42492 -11280 42548
rect -11360 42228 -11280 42492
rect -11360 42172 -11348 42228
rect -11292 42172 -11280 42228
rect -11360 41908 -11280 42172
rect -11360 41852 -11348 41908
rect -11292 41852 -11280 41908
rect -11360 41840 -11280 41852
rect -11200 42868 -11120 42880
rect -11200 42812 -11188 42868
rect -11132 42812 -11120 42868
rect -11200 42548 -11120 42812
rect -11200 42492 -11188 42548
rect -11132 42492 -11120 42548
rect -11200 42228 -11120 42492
rect -11200 42172 -11188 42228
rect -11132 42172 -11120 42228
rect -11200 41908 -11120 42172
rect -11200 41852 -11188 41908
rect -11132 41852 -11120 41908
rect -11200 41840 -11120 41852
rect -11040 42868 -10960 42880
rect -11040 42812 -11028 42868
rect -10972 42812 -10960 42868
rect -11040 42548 -10960 42812
rect -11040 42492 -11028 42548
rect -10972 42492 -10960 42548
rect -11040 42228 -10960 42492
rect -11040 42172 -11028 42228
rect -10972 42172 -10960 42228
rect -11040 41908 -10960 42172
rect -11040 41852 -11028 41908
rect -10972 41852 -10960 41908
rect -11040 41840 -10960 41852
rect -10880 42868 -10800 42880
rect -10880 42812 -10868 42868
rect -10812 42812 -10800 42868
rect -10880 42548 -10800 42812
rect -10880 42492 -10868 42548
rect -10812 42492 -10800 42548
rect -10880 42228 -10800 42492
rect -10880 42172 -10868 42228
rect -10812 42172 -10800 42228
rect -10880 41908 -10800 42172
rect -10880 41852 -10868 41908
rect -10812 41852 -10800 41908
rect -10880 41840 -10800 41852
rect -10720 42868 -10640 42880
rect -10720 42812 -10708 42868
rect -10652 42812 -10640 42868
rect -10720 42548 -10640 42812
rect -10720 42492 -10708 42548
rect -10652 42492 -10640 42548
rect -10720 42228 -10640 42492
rect -10720 42172 -10708 42228
rect -10652 42172 -10640 42228
rect -10720 41908 -10640 42172
rect -10720 41852 -10708 41908
rect -10652 41852 -10640 41908
rect -10720 41840 -10640 41852
rect -10560 42868 -10480 42880
rect -10560 42812 -10548 42868
rect -10492 42812 -10480 42868
rect -10560 42548 -10480 42812
rect -10560 42492 -10548 42548
rect -10492 42492 -10480 42548
rect -10560 42228 -10480 42492
rect -10560 42172 -10548 42228
rect -10492 42172 -10480 42228
rect -10560 41908 -10480 42172
rect -10560 41852 -10548 41908
rect -10492 41852 -10480 41908
rect -10560 41840 -10480 41852
rect -10400 42868 -10320 42880
rect -10400 42812 -10388 42868
rect -10332 42812 -10320 42868
rect -10400 42548 -10320 42812
rect -10400 42492 -10388 42548
rect -10332 42492 -10320 42548
rect -10400 42228 -10320 42492
rect -10400 42172 -10388 42228
rect -10332 42172 -10320 42228
rect -10400 41908 -10320 42172
rect -10400 41852 -10388 41908
rect -10332 41852 -10320 41908
rect -10400 41840 -10320 41852
rect -10240 42868 -10160 42880
rect -10240 42812 -10228 42868
rect -10172 42812 -10160 42868
rect -10240 42548 -10160 42812
rect -10240 42492 -10228 42548
rect -10172 42492 -10160 42548
rect -10240 42228 -10160 42492
rect -10240 42172 -10228 42228
rect -10172 42172 -10160 42228
rect -10240 41908 -10160 42172
rect -10240 41852 -10228 41908
rect -10172 41852 -10160 41908
rect -10240 41840 -10160 41852
rect -10080 42868 -10000 42880
rect -10080 42812 -10068 42868
rect -10012 42812 -10000 42868
rect -10080 42548 -10000 42812
rect -10080 42492 -10068 42548
rect -10012 42492 -10000 42548
rect -10080 42228 -10000 42492
rect -10080 42172 -10068 42228
rect -10012 42172 -10000 42228
rect -10080 41908 -10000 42172
rect -10080 41852 -10068 41908
rect -10012 41852 -10000 41908
rect -10080 41840 -10000 41852
rect -9920 42868 -9840 42880
rect -9920 42812 -9908 42868
rect -9852 42812 -9840 42868
rect -9920 42548 -9840 42812
rect -9920 42492 -9908 42548
rect -9852 42492 -9840 42548
rect -9920 42228 -9840 42492
rect -9920 42172 -9908 42228
rect -9852 42172 -9840 42228
rect -9920 41908 -9840 42172
rect -9920 41852 -9908 41908
rect -9852 41852 -9840 41908
rect -9920 41840 -9840 41852
rect -9760 42868 -9680 42880
rect -9760 42812 -9748 42868
rect -9692 42812 -9680 42868
rect -9760 42548 -9680 42812
rect -9760 42492 -9748 42548
rect -9692 42492 -9680 42548
rect -9760 42228 -9680 42492
rect -9760 42172 -9748 42228
rect -9692 42172 -9680 42228
rect -9760 41908 -9680 42172
rect -9760 41852 -9748 41908
rect -9692 41852 -9680 41908
rect -9760 41840 -9680 41852
rect -9600 42868 -9520 42880
rect -9600 42812 -9588 42868
rect -9532 42812 -9520 42868
rect -9600 42548 -9520 42812
rect -9600 42492 -9588 42548
rect -9532 42492 -9520 42548
rect -9600 42228 -9520 42492
rect -9600 42172 -9588 42228
rect -9532 42172 -9520 42228
rect -9600 41908 -9520 42172
rect -9600 41852 -9588 41908
rect -9532 41852 -9520 41908
rect -9600 41840 -9520 41852
rect -9440 42868 -9360 42880
rect -9440 42812 -9428 42868
rect -9372 42812 -9360 42868
rect -9440 42548 -9360 42812
rect -9440 42492 -9428 42548
rect -9372 42492 -9360 42548
rect -9440 42228 -9360 42492
rect -9440 42172 -9428 42228
rect -9372 42172 -9360 42228
rect -9440 41908 -9360 42172
rect -9440 41852 -9428 41908
rect -9372 41852 -9360 41908
rect -9440 41840 -9360 41852
rect -9280 42868 -9200 42880
rect -9280 42812 -9268 42868
rect -9212 42812 -9200 42868
rect -9280 42548 -9200 42812
rect -9280 42492 -9268 42548
rect -9212 42492 -9200 42548
rect -9280 42228 -9200 42492
rect -9280 42172 -9268 42228
rect -9212 42172 -9200 42228
rect -9280 41908 -9200 42172
rect -9280 41852 -9268 41908
rect -9212 41852 -9200 41908
rect -9280 41840 -9200 41852
rect -9120 42868 -9040 42880
rect -9120 42812 -9108 42868
rect -9052 42812 -9040 42868
rect -9120 42548 -9040 42812
rect -9120 42492 -9108 42548
rect -9052 42492 -9040 42548
rect -9120 42228 -9040 42492
rect -9120 42172 -9108 42228
rect -9052 42172 -9040 42228
rect -9120 41908 -9040 42172
rect -9120 41852 -9108 41908
rect -9052 41852 -9040 41908
rect -9120 41840 -9040 41852
rect -8960 42868 -8880 42880
rect -8960 42812 -8948 42868
rect -8892 42812 -8880 42868
rect -8960 42548 -8880 42812
rect -8960 42492 -8948 42548
rect -8892 42492 -8880 42548
rect -8960 42228 -8880 42492
rect -8960 42172 -8948 42228
rect -8892 42172 -8880 42228
rect -8960 41908 -8880 42172
rect -8960 41852 -8948 41908
rect -8892 41852 -8880 41908
rect -8960 41840 -8880 41852
rect -8800 42868 -8720 42880
rect -8800 42812 -8788 42868
rect -8732 42812 -8720 42868
rect -8800 42548 -8720 42812
rect -8800 42492 -8788 42548
rect -8732 42492 -8720 42548
rect -8800 42228 -8720 42492
rect -8800 42172 -8788 42228
rect -8732 42172 -8720 42228
rect -8800 41908 -8720 42172
rect -8800 41852 -8788 41908
rect -8732 41852 -8720 41908
rect -8800 41840 -8720 41852
rect -8640 42868 -8560 42880
rect -8640 42812 -8628 42868
rect -8572 42812 -8560 42868
rect -8640 42548 -8560 42812
rect -8640 42492 -8628 42548
rect -8572 42492 -8560 42548
rect -8640 42228 -8560 42492
rect -8640 42172 -8628 42228
rect -8572 42172 -8560 42228
rect -8640 41908 -8560 42172
rect -8640 41852 -8628 41908
rect -8572 41852 -8560 41908
rect -8640 41840 -8560 41852
rect -8480 42868 -8400 42880
rect -8480 42812 -8468 42868
rect -8412 42812 -8400 42868
rect -8480 42548 -8400 42812
rect -8480 42492 -8468 42548
rect -8412 42492 -8400 42548
rect -8480 42228 -8400 42492
rect -8480 42172 -8468 42228
rect -8412 42172 -8400 42228
rect -8480 41908 -8400 42172
rect -8480 41852 -8468 41908
rect -8412 41852 -8400 41908
rect -8480 41840 -8400 41852
rect -8320 42868 -8240 42880
rect -8320 42812 -8308 42868
rect -8252 42812 -8240 42868
rect -8320 42548 -8240 42812
rect -8320 42492 -8308 42548
rect -8252 42492 -8240 42548
rect -8320 42228 -8240 42492
rect -8320 42172 -8308 42228
rect -8252 42172 -8240 42228
rect -8320 41908 -8240 42172
rect -8320 41852 -8308 41908
rect -8252 41852 -8240 41908
rect -8320 41840 -8240 41852
rect -8160 42868 -8080 42880
rect -8160 42812 -8148 42868
rect -8092 42812 -8080 42868
rect -8160 42548 -8080 42812
rect -8160 42492 -8148 42548
rect -8092 42492 -8080 42548
rect -8160 42228 -8080 42492
rect -8160 42172 -8148 42228
rect -8092 42172 -8080 42228
rect -8160 41908 -8080 42172
rect -8160 41852 -8148 41908
rect -8092 41852 -8080 41908
rect -8160 41840 -8080 41852
rect -8000 42868 -7920 42880
rect -8000 42812 -7988 42868
rect -7932 42812 -7920 42868
rect -8000 42548 -7920 42812
rect -8000 42492 -7988 42548
rect -7932 42492 -7920 42548
rect -8000 42228 -7920 42492
rect -8000 42172 -7988 42228
rect -7932 42172 -7920 42228
rect -8000 41908 -7920 42172
rect -8000 41852 -7988 41908
rect -7932 41852 -7920 41908
rect -8000 41840 -7920 41852
rect -7840 42868 -7760 42880
rect -7840 42812 -7828 42868
rect -7772 42812 -7760 42868
rect -7840 42548 -7760 42812
rect -7840 42492 -7828 42548
rect -7772 42492 -7760 42548
rect -7840 42228 -7760 42492
rect -7840 42172 -7828 42228
rect -7772 42172 -7760 42228
rect -7840 41908 -7760 42172
rect -7840 41852 -7828 41908
rect -7772 41852 -7760 41908
rect -7840 41840 -7760 41852
rect -7680 42868 -7600 42880
rect -7680 42812 -7668 42868
rect -7612 42812 -7600 42868
rect -7680 42548 -7600 42812
rect -7680 42492 -7668 42548
rect -7612 42492 -7600 42548
rect -7680 42228 -7600 42492
rect -7680 42172 -7668 42228
rect -7612 42172 -7600 42228
rect -7680 41908 -7600 42172
rect -7680 41852 -7668 41908
rect -7612 41852 -7600 41908
rect -7680 41840 -7600 41852
rect -7520 42868 -7440 42880
rect -7520 42812 -7508 42868
rect -7452 42812 -7440 42868
rect -7520 42548 -7440 42812
rect -7520 42492 -7508 42548
rect -7452 42492 -7440 42548
rect -7520 42228 -7440 42492
rect -7520 42172 -7508 42228
rect -7452 42172 -7440 42228
rect -7520 41908 -7440 42172
rect -7520 41852 -7508 41908
rect -7452 41852 -7440 41908
rect -7520 41840 -7440 41852
rect -7360 42868 -7280 42880
rect -7360 42812 -7348 42868
rect -7292 42812 -7280 42868
rect -7360 42548 -7280 42812
rect -7360 42492 -7348 42548
rect -7292 42492 -7280 42548
rect -7360 42228 -7280 42492
rect -7360 42172 -7348 42228
rect -7292 42172 -7280 42228
rect -7360 41908 -7280 42172
rect -7360 41852 -7348 41908
rect -7292 41852 -7280 41908
rect -7360 41840 -7280 41852
rect -7200 42868 -7120 42880
rect -7200 42812 -7188 42868
rect -7132 42812 -7120 42868
rect -7200 42548 -7120 42812
rect -7200 42492 -7188 42548
rect -7132 42492 -7120 42548
rect -7200 42228 -7120 42492
rect -7200 42172 -7188 42228
rect -7132 42172 -7120 42228
rect -7200 41908 -7120 42172
rect -7200 41852 -7188 41908
rect -7132 41852 -7120 41908
rect -7200 41840 -7120 41852
rect -7040 42868 -6960 42880
rect -7040 42812 -7028 42868
rect -6972 42812 -6960 42868
rect -7040 42548 -6960 42812
rect -7040 42492 -7028 42548
rect -6972 42492 -6960 42548
rect -7040 42228 -6960 42492
rect -7040 42172 -7028 42228
rect -6972 42172 -6960 42228
rect -7040 41908 -6960 42172
rect -7040 41852 -7028 41908
rect -6972 41852 -6960 41908
rect -7040 41840 -6960 41852
rect -6880 42868 -6800 42880
rect -6880 42812 -6868 42868
rect -6812 42812 -6800 42868
rect -6880 42548 -6800 42812
rect -6880 42492 -6868 42548
rect -6812 42492 -6800 42548
rect -6880 42228 -6800 42492
rect -6880 42172 -6868 42228
rect -6812 42172 -6800 42228
rect -6880 41908 -6800 42172
rect -6880 41852 -6868 41908
rect -6812 41852 -6800 41908
rect -6880 41840 -6800 41852
rect -6720 42868 -6640 42880
rect -6720 42812 -6708 42868
rect -6652 42812 -6640 42868
rect -6720 42548 -6640 42812
rect -6720 42492 -6708 42548
rect -6652 42492 -6640 42548
rect -6720 42228 -6640 42492
rect -6720 42172 -6708 42228
rect -6652 42172 -6640 42228
rect -6720 41908 -6640 42172
rect -6720 41852 -6708 41908
rect -6652 41852 -6640 41908
rect -6720 41840 -6640 41852
rect -6560 42868 -6480 42880
rect -6560 42812 -6548 42868
rect -6492 42812 -6480 42868
rect -6560 42548 -6480 42812
rect -6560 42492 -6548 42548
rect -6492 42492 -6480 42548
rect -6560 42228 -6480 42492
rect -6560 42172 -6548 42228
rect -6492 42172 -6480 42228
rect -6560 41908 -6480 42172
rect -6560 41852 -6548 41908
rect -6492 41852 -6480 41908
rect -6560 41840 -6480 41852
rect -6400 42868 -6320 42880
rect -6400 42812 -6388 42868
rect -6332 42812 -6320 42868
rect -6400 42548 -6320 42812
rect -6400 42492 -6388 42548
rect -6332 42492 -6320 42548
rect -6400 42228 -6320 42492
rect -6400 42172 -6388 42228
rect -6332 42172 -6320 42228
rect -6400 41908 -6320 42172
rect -6400 41852 -6388 41908
rect -6332 41852 -6320 41908
rect -6400 41840 -6320 41852
rect -6240 42868 -6160 42880
rect -6240 42812 -6228 42868
rect -6172 42812 -6160 42868
rect -6240 42548 -6160 42812
rect -6240 42492 -6228 42548
rect -6172 42492 -6160 42548
rect -6240 42228 -6160 42492
rect -6240 42172 -6228 42228
rect -6172 42172 -6160 42228
rect -6240 41908 -6160 42172
rect -6240 41852 -6228 41908
rect -6172 41852 -6160 41908
rect -6240 41840 -6160 41852
rect -6080 42868 -6000 42880
rect -6080 42812 -6068 42868
rect -6012 42812 -6000 42868
rect -6080 42548 -6000 42812
rect -6080 42492 -6068 42548
rect -6012 42492 -6000 42548
rect -6080 42228 -6000 42492
rect -6080 42172 -6068 42228
rect -6012 42172 -6000 42228
rect -6080 41908 -6000 42172
rect -6080 41852 -6068 41908
rect -6012 41852 -6000 41908
rect -6080 41840 -6000 41852
rect -5920 42868 -5840 42880
rect -5920 42812 -5908 42868
rect -5852 42812 -5840 42868
rect -5920 42548 -5840 42812
rect -5920 42492 -5908 42548
rect -5852 42492 -5840 42548
rect -5920 42228 -5840 42492
rect -5920 42172 -5908 42228
rect -5852 42172 -5840 42228
rect -5920 41908 -5840 42172
rect -5920 41852 -5908 41908
rect -5852 41852 -5840 41908
rect -5920 41840 -5840 41852
rect -5760 42868 -5680 42880
rect -5760 42812 -5748 42868
rect -5692 42812 -5680 42868
rect -5760 42548 -5680 42812
rect -5760 42492 -5748 42548
rect -5692 42492 -5680 42548
rect -5760 42228 -5680 42492
rect -5760 42172 -5748 42228
rect -5692 42172 -5680 42228
rect -5760 41908 -5680 42172
rect -5760 41852 -5748 41908
rect -5692 41852 -5680 41908
rect -5760 41840 -5680 41852
rect -5600 42868 -5520 42880
rect -5600 42812 -5588 42868
rect -5532 42812 -5520 42868
rect -5600 42548 -5520 42812
rect -5600 42492 -5588 42548
rect -5532 42492 -5520 42548
rect -5600 42228 -5520 42492
rect -5600 42172 -5588 42228
rect -5532 42172 -5520 42228
rect -5600 41908 -5520 42172
rect -5600 41852 -5588 41908
rect -5532 41852 -5520 41908
rect -5600 41840 -5520 41852
rect -5440 42868 -5360 42880
rect -5440 42812 -5428 42868
rect -5372 42812 -5360 42868
rect -5440 42548 -5360 42812
rect -5440 42492 -5428 42548
rect -5372 42492 -5360 42548
rect -5440 42228 -5360 42492
rect -5440 42172 -5428 42228
rect -5372 42172 -5360 42228
rect -5440 41908 -5360 42172
rect -5440 41852 -5428 41908
rect -5372 41852 -5360 41908
rect -5440 41840 -5360 41852
rect -5280 42868 -5200 42880
rect -5280 42812 -5268 42868
rect -5212 42812 -5200 42868
rect -5280 42548 -5200 42812
rect -5280 42492 -5268 42548
rect -5212 42492 -5200 42548
rect -5280 42228 -5200 42492
rect -5280 42172 -5268 42228
rect -5212 42172 -5200 42228
rect -5280 41908 -5200 42172
rect -5280 41852 -5268 41908
rect -5212 41852 -5200 41908
rect -5280 41840 -5200 41852
rect -5120 42868 -5040 42880
rect -5120 42812 -5108 42868
rect -5052 42812 -5040 42868
rect -5120 42548 -5040 42812
rect -5120 42492 -5108 42548
rect -5052 42492 -5040 42548
rect -5120 42228 -5040 42492
rect -5120 42172 -5108 42228
rect -5052 42172 -5040 42228
rect -5120 41908 -5040 42172
rect -5120 41852 -5108 41908
rect -5052 41852 -5040 41908
rect -5120 41840 -5040 41852
rect -4960 42868 -4880 42880
rect -4960 42812 -4948 42868
rect -4892 42812 -4880 42868
rect -4960 42548 -4880 42812
rect -4960 42492 -4948 42548
rect -4892 42492 -4880 42548
rect -4960 42228 -4880 42492
rect -4960 42172 -4948 42228
rect -4892 42172 -4880 42228
rect -4960 41908 -4880 42172
rect -4960 41852 -4948 41908
rect -4892 41852 -4880 41908
rect -4960 41840 -4880 41852
rect -4800 42868 -4720 42880
rect -4800 42812 -4788 42868
rect -4732 42812 -4720 42868
rect -4800 42548 -4720 42812
rect -4800 42492 -4788 42548
rect -4732 42492 -4720 42548
rect -4800 42228 -4720 42492
rect -4800 42172 -4788 42228
rect -4732 42172 -4720 42228
rect -4800 41908 -4720 42172
rect -4800 41852 -4788 41908
rect -4732 41852 -4720 41908
rect -4800 41840 -4720 41852
rect -4640 42868 -4560 42880
rect -4640 42812 -4628 42868
rect -4572 42812 -4560 42868
rect -4640 42548 -4560 42812
rect -4640 42492 -4628 42548
rect -4572 42492 -4560 42548
rect -4640 42228 -4560 42492
rect -4640 42172 -4628 42228
rect -4572 42172 -4560 42228
rect -4640 41908 -4560 42172
rect -4640 41852 -4628 41908
rect -4572 41852 -4560 41908
rect -4640 41840 -4560 41852
rect -4480 42868 -4400 42880
rect -4480 42812 -4468 42868
rect -4412 42812 -4400 42868
rect -4480 42548 -4400 42812
rect -4480 42492 -4468 42548
rect -4412 42492 -4400 42548
rect -4480 42228 -4400 42492
rect -4480 42172 -4468 42228
rect -4412 42172 -4400 42228
rect -4480 41908 -4400 42172
rect -4480 41852 -4468 41908
rect -4412 41852 -4400 41908
rect -4480 41840 -4400 41852
rect -4320 42868 -4240 42880
rect -4320 42812 -4308 42868
rect -4252 42812 -4240 42868
rect -4320 42548 -4240 42812
rect -4320 42492 -4308 42548
rect -4252 42492 -4240 42548
rect -4320 42228 -4240 42492
rect -4320 42172 -4308 42228
rect -4252 42172 -4240 42228
rect -4320 41908 -4240 42172
rect -4320 41852 -4308 41908
rect -4252 41852 -4240 41908
rect -4320 41840 -4240 41852
rect -4160 42868 -4080 42880
rect -4160 42812 -4148 42868
rect -4092 42812 -4080 42868
rect -4160 42548 -4080 42812
rect -4160 42492 -4148 42548
rect -4092 42492 -4080 42548
rect -4160 42228 -4080 42492
rect -4160 42172 -4148 42228
rect -4092 42172 -4080 42228
rect -4160 41908 -4080 42172
rect -4160 41852 -4148 41908
rect -4092 41852 -4080 41908
rect -4160 41840 -4080 41852
rect -4000 42868 -3920 42880
rect -4000 42812 -3988 42868
rect -3932 42812 -3920 42868
rect -4000 42548 -3920 42812
rect -4000 42492 -3988 42548
rect -3932 42492 -3920 42548
rect -4000 42228 -3920 42492
rect -4000 42172 -3988 42228
rect -3932 42172 -3920 42228
rect -4000 41908 -3920 42172
rect -4000 41852 -3988 41908
rect -3932 41852 -3920 41908
rect -4000 41840 -3920 41852
rect -3680 42868 -3600 42880
rect -3680 42812 -3668 42868
rect -3612 42812 -3600 42868
rect -3680 42548 -3600 42812
rect -3680 42492 -3668 42548
rect -3612 42492 -3600 42548
rect -3680 42228 -3600 42492
rect -3680 42172 -3668 42228
rect -3612 42172 -3600 42228
rect -3680 41908 -3600 42172
rect -3680 41852 -3668 41908
rect -3612 41852 -3600 41908
rect -3680 41840 -3600 41852
rect -3520 42868 -3440 42880
rect -3520 42812 -3508 42868
rect -3452 42812 -3440 42868
rect -3520 42548 -3440 42812
rect -3520 42492 -3508 42548
rect -3452 42492 -3440 42548
rect -3520 42228 -3440 42492
rect -3520 42172 -3508 42228
rect -3452 42172 -3440 42228
rect -3520 41908 -3440 42172
rect -3520 41852 -3508 41908
rect -3452 41852 -3440 41908
rect -3520 41840 -3440 41852
rect -3360 42868 -3280 42880
rect -3360 42812 -3348 42868
rect -3292 42812 -3280 42868
rect -3360 42548 -3280 42812
rect -3360 42492 -3348 42548
rect -3292 42492 -3280 42548
rect -3360 42228 -3280 42492
rect -3200 42868 -3120 42880
rect -3200 42812 -3188 42868
rect -3132 42812 -3120 42868
rect -3200 42548 -3120 42812
rect -3200 42492 -3188 42548
rect -3132 42492 -3120 42548
rect -3200 42480 -3120 42492
rect -3040 42868 -2960 42880
rect -3040 42812 -3028 42868
rect -2972 42812 -2960 42868
rect -3040 42548 -2960 42812
rect -2720 42868 -2640 42880
rect -2720 42812 -2708 42868
rect -2652 42812 -2640 42868
rect -3040 42492 -3028 42548
rect -2972 42492 -2960 42548
rect -3360 42172 -3348 42228
rect -3292 42172 -3280 42228
rect -3360 41908 -3280 42172
rect -3360 41852 -3348 41908
rect -3292 41852 -3280 41908
rect -11520 41692 -11508 41748
rect -11452 41692 -11440 41748
rect -11520 41588 -11440 41692
rect -11520 41532 -11508 41588
rect -11452 41532 -11440 41588
rect -11520 40868 -11440 41532
rect -3360 41748 -3280 41852
rect -3360 41692 -3348 41748
rect -3292 41692 -3280 41748
rect -3360 41588 -3280 41692
rect -3360 41532 -3348 41588
rect -3292 41532 -3280 41588
rect -11360 41348 -11280 41360
rect -11360 41292 -11348 41348
rect -11292 41292 -11280 41348
rect -11360 41028 -11280 41292
rect -11360 40972 -11348 41028
rect -11292 40972 -11280 41028
rect -11360 40960 -11280 40972
rect -11200 41348 -11120 41360
rect -11200 41292 -11188 41348
rect -11132 41292 -11120 41348
rect -11200 41028 -11120 41292
rect -11200 40972 -11188 41028
rect -11132 40972 -11120 41028
rect -11200 40960 -11120 40972
rect -11040 41348 -10960 41360
rect -11040 41292 -11028 41348
rect -10972 41292 -10960 41348
rect -11040 41028 -10960 41292
rect -11040 40972 -11028 41028
rect -10972 40972 -10960 41028
rect -11040 40960 -10960 40972
rect -10880 41348 -10800 41360
rect -10880 41292 -10868 41348
rect -10812 41292 -10800 41348
rect -10880 41028 -10800 41292
rect -10880 40972 -10868 41028
rect -10812 40972 -10800 41028
rect -10880 40960 -10800 40972
rect -10720 41348 -10640 41360
rect -10720 41292 -10708 41348
rect -10652 41292 -10640 41348
rect -10720 41028 -10640 41292
rect -10720 40972 -10708 41028
rect -10652 40972 -10640 41028
rect -10720 40960 -10640 40972
rect -10560 41348 -10480 41360
rect -10560 41292 -10548 41348
rect -10492 41292 -10480 41348
rect -10560 41028 -10480 41292
rect -10560 40972 -10548 41028
rect -10492 40972 -10480 41028
rect -10560 40960 -10480 40972
rect -10400 41348 -10320 41360
rect -10400 41292 -10388 41348
rect -10332 41292 -10320 41348
rect -10400 41028 -10320 41292
rect -10400 40972 -10388 41028
rect -10332 40972 -10320 41028
rect -10400 40960 -10320 40972
rect -10240 41348 -10160 41360
rect -10240 41292 -10228 41348
rect -10172 41292 -10160 41348
rect -10240 41028 -10160 41292
rect -10240 40972 -10228 41028
rect -10172 40972 -10160 41028
rect -10240 40960 -10160 40972
rect -10080 41348 -10000 41360
rect -10080 41292 -10068 41348
rect -10012 41292 -10000 41348
rect -10080 41028 -10000 41292
rect -10080 40972 -10068 41028
rect -10012 40972 -10000 41028
rect -10080 40960 -10000 40972
rect -9920 41348 -9840 41360
rect -9920 41292 -9908 41348
rect -9852 41292 -9840 41348
rect -9920 41028 -9840 41292
rect -9920 40972 -9908 41028
rect -9852 40972 -9840 41028
rect -9920 40960 -9840 40972
rect -9760 41348 -9680 41360
rect -9760 41292 -9748 41348
rect -9692 41292 -9680 41348
rect -9760 41028 -9680 41292
rect -9760 40972 -9748 41028
rect -9692 40972 -9680 41028
rect -9760 40960 -9680 40972
rect -9600 41348 -9520 41360
rect -9600 41292 -9588 41348
rect -9532 41292 -9520 41348
rect -9600 41028 -9520 41292
rect -9600 40972 -9588 41028
rect -9532 40972 -9520 41028
rect -9600 40960 -9520 40972
rect -9440 41348 -9360 41360
rect -9440 41292 -9428 41348
rect -9372 41292 -9360 41348
rect -9440 41028 -9360 41292
rect -9440 40972 -9428 41028
rect -9372 40972 -9360 41028
rect -9440 40960 -9360 40972
rect -9280 41348 -9200 41360
rect -9280 41292 -9268 41348
rect -9212 41292 -9200 41348
rect -9280 41028 -9200 41292
rect -9280 40972 -9268 41028
rect -9212 40972 -9200 41028
rect -9280 40960 -9200 40972
rect -9120 41348 -9040 41360
rect -9120 41292 -9108 41348
rect -9052 41292 -9040 41348
rect -9120 41028 -9040 41292
rect -9120 40972 -9108 41028
rect -9052 40972 -9040 41028
rect -9120 40960 -9040 40972
rect -8960 41348 -8880 41360
rect -8960 41292 -8948 41348
rect -8892 41292 -8880 41348
rect -8960 41028 -8880 41292
rect -8960 40972 -8948 41028
rect -8892 40972 -8880 41028
rect -8960 40960 -8880 40972
rect -8800 41348 -8720 41360
rect -8800 41292 -8788 41348
rect -8732 41292 -8720 41348
rect -8800 41028 -8720 41292
rect -8800 40972 -8788 41028
rect -8732 40972 -8720 41028
rect -8800 40960 -8720 40972
rect -8640 41348 -8560 41360
rect -8640 41292 -8628 41348
rect -8572 41292 -8560 41348
rect -8640 41028 -8560 41292
rect -8640 40972 -8628 41028
rect -8572 40972 -8560 41028
rect -8640 40960 -8560 40972
rect -8480 41348 -8400 41360
rect -8480 41292 -8468 41348
rect -8412 41292 -8400 41348
rect -8480 41028 -8400 41292
rect -8480 40972 -8468 41028
rect -8412 40972 -8400 41028
rect -8480 40960 -8400 40972
rect -8320 41348 -8240 41360
rect -8320 41292 -8308 41348
rect -8252 41292 -8240 41348
rect -8320 41028 -8240 41292
rect -8320 40972 -8308 41028
rect -8252 40972 -8240 41028
rect -8320 40960 -8240 40972
rect -8160 41348 -8080 41360
rect -8160 41292 -8148 41348
rect -8092 41292 -8080 41348
rect -8160 41028 -8080 41292
rect -8160 40972 -8148 41028
rect -8092 40972 -8080 41028
rect -8160 40960 -8080 40972
rect -8000 41348 -7920 41360
rect -8000 41292 -7988 41348
rect -7932 41292 -7920 41348
rect -8000 41028 -7920 41292
rect -8000 40972 -7988 41028
rect -7932 40972 -7920 41028
rect -8000 40960 -7920 40972
rect -7840 41348 -7760 41360
rect -7840 41292 -7828 41348
rect -7772 41292 -7760 41348
rect -7840 41028 -7760 41292
rect -7840 40972 -7828 41028
rect -7772 40972 -7760 41028
rect -7840 40960 -7760 40972
rect -7680 41348 -7600 41360
rect -7680 41292 -7668 41348
rect -7612 41292 -7600 41348
rect -7680 41028 -7600 41292
rect -7680 40972 -7668 41028
rect -7612 40972 -7600 41028
rect -7680 40960 -7600 40972
rect -7520 41348 -7440 41360
rect -7520 41292 -7508 41348
rect -7452 41292 -7440 41348
rect -7520 41028 -7440 41292
rect -7520 40972 -7508 41028
rect -7452 40972 -7440 41028
rect -7520 40960 -7440 40972
rect -7360 41348 -7280 41360
rect -7360 41292 -7348 41348
rect -7292 41292 -7280 41348
rect -7360 41028 -7280 41292
rect -7360 40972 -7348 41028
rect -7292 40972 -7280 41028
rect -7360 40960 -7280 40972
rect -7200 41348 -7120 41360
rect -7200 41292 -7188 41348
rect -7132 41292 -7120 41348
rect -7200 41028 -7120 41292
rect -7200 40972 -7188 41028
rect -7132 40972 -7120 41028
rect -7200 40960 -7120 40972
rect -7040 41348 -6960 41360
rect -7040 41292 -7028 41348
rect -6972 41292 -6960 41348
rect -7040 41028 -6960 41292
rect -7040 40972 -7028 41028
rect -6972 40972 -6960 41028
rect -7040 40960 -6960 40972
rect -6880 41348 -6800 41360
rect -6880 41292 -6868 41348
rect -6812 41292 -6800 41348
rect -6880 41028 -6800 41292
rect -6880 40972 -6868 41028
rect -6812 40972 -6800 41028
rect -6880 40960 -6800 40972
rect -6720 41348 -6640 41360
rect -6720 41292 -6708 41348
rect -6652 41292 -6640 41348
rect -6720 41028 -6640 41292
rect -6720 40972 -6708 41028
rect -6652 40972 -6640 41028
rect -6720 40960 -6640 40972
rect -6560 41348 -6480 41360
rect -6560 41292 -6548 41348
rect -6492 41292 -6480 41348
rect -6560 41028 -6480 41292
rect -6560 40972 -6548 41028
rect -6492 40972 -6480 41028
rect -6560 40960 -6480 40972
rect -6400 41348 -6320 41360
rect -6400 41292 -6388 41348
rect -6332 41292 -6320 41348
rect -6400 41028 -6320 41292
rect -6400 40972 -6388 41028
rect -6332 40972 -6320 41028
rect -6400 40960 -6320 40972
rect -6240 41348 -6160 41360
rect -6240 41292 -6228 41348
rect -6172 41292 -6160 41348
rect -6240 41028 -6160 41292
rect -6240 40972 -6228 41028
rect -6172 40972 -6160 41028
rect -6240 40960 -6160 40972
rect -6080 41348 -6000 41360
rect -6080 41292 -6068 41348
rect -6012 41292 -6000 41348
rect -6080 41028 -6000 41292
rect -6080 40972 -6068 41028
rect -6012 40972 -6000 41028
rect -6080 40960 -6000 40972
rect -5920 41348 -5840 41360
rect -5920 41292 -5908 41348
rect -5852 41292 -5840 41348
rect -5920 41028 -5840 41292
rect -5920 40972 -5908 41028
rect -5852 40972 -5840 41028
rect -5920 40960 -5840 40972
rect -5760 41348 -5680 41360
rect -5760 41292 -5748 41348
rect -5692 41292 -5680 41348
rect -5760 41028 -5680 41292
rect -5760 40972 -5748 41028
rect -5692 40972 -5680 41028
rect -5760 40960 -5680 40972
rect -5600 41348 -5520 41360
rect -5600 41292 -5588 41348
rect -5532 41292 -5520 41348
rect -5600 41028 -5520 41292
rect -5600 40972 -5588 41028
rect -5532 40972 -5520 41028
rect -5600 40960 -5520 40972
rect -5440 41348 -5360 41360
rect -5440 41292 -5428 41348
rect -5372 41292 -5360 41348
rect -5440 41028 -5360 41292
rect -5440 40972 -5428 41028
rect -5372 40972 -5360 41028
rect -5440 40960 -5360 40972
rect -5280 41348 -5200 41360
rect -5280 41292 -5268 41348
rect -5212 41292 -5200 41348
rect -5280 41028 -5200 41292
rect -5280 40972 -5268 41028
rect -5212 40972 -5200 41028
rect -5280 40960 -5200 40972
rect -5120 41348 -5040 41360
rect -5120 41292 -5108 41348
rect -5052 41292 -5040 41348
rect -5120 41028 -5040 41292
rect -5120 40972 -5108 41028
rect -5052 40972 -5040 41028
rect -5120 40960 -5040 40972
rect -4960 41348 -4880 41360
rect -4960 41292 -4948 41348
rect -4892 41292 -4880 41348
rect -4960 41028 -4880 41292
rect -4960 40972 -4948 41028
rect -4892 40972 -4880 41028
rect -4960 40960 -4880 40972
rect -4800 41348 -4720 41360
rect -4800 41292 -4788 41348
rect -4732 41292 -4720 41348
rect -4800 41028 -4720 41292
rect -4800 40972 -4788 41028
rect -4732 40972 -4720 41028
rect -4800 40960 -4720 40972
rect -4640 41348 -4560 41360
rect -4640 41292 -4628 41348
rect -4572 41292 -4560 41348
rect -4640 41028 -4560 41292
rect -4640 40972 -4628 41028
rect -4572 40972 -4560 41028
rect -4640 40960 -4560 40972
rect -4480 41348 -4400 41360
rect -4480 41292 -4468 41348
rect -4412 41292 -4400 41348
rect -4480 41028 -4400 41292
rect -4480 40972 -4468 41028
rect -4412 40972 -4400 41028
rect -4480 40960 -4400 40972
rect -4320 41348 -4240 41360
rect -4320 41292 -4308 41348
rect -4252 41292 -4240 41348
rect -4320 41028 -4240 41292
rect -4320 40972 -4308 41028
rect -4252 40972 -4240 41028
rect -4320 40960 -4240 40972
rect -4160 41348 -4080 41360
rect -4160 41292 -4148 41348
rect -4092 41292 -4080 41348
rect -4160 41028 -4080 41292
rect -4160 40972 -4148 41028
rect -4092 40972 -4080 41028
rect -4160 40960 -4080 40972
rect -4000 41348 -3920 41360
rect -4000 41292 -3988 41348
rect -3932 41292 -3920 41348
rect -4000 41028 -3920 41292
rect -4000 40972 -3988 41028
rect -3932 40972 -3920 41028
rect -4000 40960 -3920 40972
rect -3840 41348 -3760 41360
rect -3840 41292 -3828 41348
rect -3772 41292 -3760 41348
rect -3840 41028 -3760 41292
rect -3840 40972 -3828 41028
rect -3772 40972 -3760 41028
rect -3840 40960 -3760 40972
rect -3680 41348 -3600 41360
rect -3680 41292 -3668 41348
rect -3612 41292 -3600 41348
rect -3680 41028 -3600 41292
rect -3680 40972 -3668 41028
rect -3612 40972 -3600 41028
rect -3680 40960 -3600 40972
rect -3520 41348 -3440 41360
rect -3520 41292 -3508 41348
rect -3452 41292 -3440 41348
rect -3520 41028 -3440 41292
rect -3520 40972 -3508 41028
rect -3452 40972 -3440 41028
rect -3520 40960 -3440 40972
rect -11520 40812 -11508 40868
rect -11452 40812 -11440 40868
rect -11520 40708 -11440 40812
rect -3360 40868 -3280 41532
rect -3360 40812 -3348 40868
rect -3292 40812 -3280 40868
rect -11520 40652 -11508 40708
rect -11452 40652 -11440 40708
rect -11520 40388 -11440 40652
rect -11520 40332 -11508 40388
rect -11452 40332 -11440 40388
rect -11520 40320 -11440 40332
rect -10560 40708 -10480 40720
rect -10560 40652 -10548 40708
rect -10492 40652 -10480 40708
rect -10560 40388 -10480 40652
rect -10240 40708 -10160 40720
rect -10240 40652 -10228 40708
rect -10172 40652 -10160 40708
rect -10560 40332 -10548 40388
rect -10492 40332 -10480 40388
rect -10560 40320 -10480 40332
rect -10400 40548 -10320 40560
rect -10400 40492 -10388 40548
rect -10332 40492 -10320 40548
rect -10400 39920 -10320 40492
rect -10240 40388 -10160 40652
rect -10240 40332 -10228 40388
rect -10172 40332 -10160 40388
rect -10240 40320 -10160 40332
rect -10080 40708 -10000 40720
rect -10080 40652 -10068 40708
rect -10012 40652 -10000 40708
rect -10080 40388 -10000 40652
rect -10080 40332 -10068 40388
rect -10012 40332 -10000 40388
rect -10080 40320 -10000 40332
rect -9920 40708 -9840 40720
rect -9920 40652 -9908 40708
rect -9852 40652 -9840 40708
rect -9920 40388 -9840 40652
rect -9920 40332 -9908 40388
rect -9852 40332 -9840 40388
rect -9920 40320 -9840 40332
rect -9760 40708 -9680 40720
rect -9760 40652 -9748 40708
rect -9692 40652 -9680 40708
rect -9760 40388 -9680 40652
rect -9760 40332 -9748 40388
rect -9692 40332 -9680 40388
rect -9760 40320 -9680 40332
rect -9600 40708 -9520 40720
rect -9600 40652 -9588 40708
rect -9532 40652 -9520 40708
rect -9600 40388 -9520 40652
rect -9600 40332 -9588 40388
rect -9532 40332 -9520 40388
rect -9600 40320 -9520 40332
rect -9440 40708 -9360 40720
rect -9440 40652 -9428 40708
rect -9372 40652 -9360 40708
rect -9440 40388 -9360 40652
rect -9440 40332 -9428 40388
rect -9372 40332 -9360 40388
rect -9440 40320 -9360 40332
rect -9280 40708 -9200 40720
rect -9280 40652 -9268 40708
rect -9212 40652 -9200 40708
rect -9280 40388 -9200 40652
rect -9280 40332 -9268 40388
rect -9212 40332 -9200 40388
rect -9280 40320 -9200 40332
rect -9120 40708 -9040 40720
rect -9120 40652 -9108 40708
rect -9052 40652 -9040 40708
rect -9120 40388 -9040 40652
rect -9120 40332 -9108 40388
rect -9052 40332 -9040 40388
rect -9120 40320 -9040 40332
rect -8960 40708 -8880 40720
rect -8960 40652 -8948 40708
rect -8892 40652 -8880 40708
rect -8960 40388 -8880 40652
rect -8960 40332 -8948 40388
rect -8892 40332 -8880 40388
rect -8960 40320 -8880 40332
rect -8800 40708 -8720 40720
rect -8800 40652 -8788 40708
rect -8732 40652 -8720 40708
rect -8800 40388 -8720 40652
rect -8800 40332 -8788 40388
rect -8732 40332 -8720 40388
rect -8800 40320 -8720 40332
rect -8640 40708 -8560 40720
rect -8640 40652 -8628 40708
rect -8572 40652 -8560 40708
rect -8640 40388 -8560 40652
rect -8640 40332 -8628 40388
rect -8572 40332 -8560 40388
rect -8640 40320 -8560 40332
rect -8480 40708 -8400 40720
rect -8480 40652 -8468 40708
rect -8412 40652 -8400 40708
rect -8480 40388 -8400 40652
rect -8480 40332 -8468 40388
rect -8412 40332 -8400 40388
rect -8480 40320 -8400 40332
rect -8320 40708 -8240 40720
rect -8320 40652 -8308 40708
rect -8252 40652 -8240 40708
rect -8320 40388 -8240 40652
rect -8320 40332 -8308 40388
rect -8252 40332 -8240 40388
rect -8320 40320 -8240 40332
rect -8160 40708 -8080 40720
rect -8160 40652 -8148 40708
rect -8092 40652 -8080 40708
rect -8160 40388 -8080 40652
rect -8160 40332 -8148 40388
rect -8092 40332 -8080 40388
rect -8160 40320 -8080 40332
rect -8000 40708 -7920 40720
rect -8000 40652 -7988 40708
rect -7932 40652 -7920 40708
rect -8000 40388 -7920 40652
rect -8000 40332 -7988 40388
rect -7932 40332 -7920 40388
rect -8000 40320 -7920 40332
rect -7840 40708 -7760 40720
rect -7840 40652 -7828 40708
rect -7772 40652 -7760 40708
rect -7840 40388 -7760 40652
rect -7840 40332 -7828 40388
rect -7772 40332 -7760 40388
rect -7840 40320 -7760 40332
rect -7680 40708 -7600 40720
rect -7680 40652 -7668 40708
rect -7612 40652 -7600 40708
rect -7680 40388 -7600 40652
rect -7680 40332 -7668 40388
rect -7612 40332 -7600 40388
rect -7680 40320 -7600 40332
rect -7520 40708 -7440 40720
rect -7520 40652 -7508 40708
rect -7452 40652 -7440 40708
rect -7520 40388 -7440 40652
rect -7520 40332 -7508 40388
rect -7452 40332 -7440 40388
rect -7520 40320 -7440 40332
rect -7360 40708 -7280 40720
rect -7360 40652 -7348 40708
rect -7292 40652 -7280 40708
rect -7360 40388 -7280 40652
rect -7360 40332 -7348 40388
rect -7292 40332 -7280 40388
rect -7360 40320 -7280 40332
rect -7200 40708 -7120 40720
rect -7200 40652 -7188 40708
rect -7132 40652 -7120 40708
rect -7200 40388 -7120 40652
rect -7200 40332 -7188 40388
rect -7132 40332 -7120 40388
rect -7200 40320 -7120 40332
rect -7040 40708 -6960 40720
rect -7040 40652 -7028 40708
rect -6972 40652 -6960 40708
rect -7040 40388 -6960 40652
rect -7040 40332 -7028 40388
rect -6972 40332 -6960 40388
rect -7040 40320 -6960 40332
rect -6880 40708 -6800 40720
rect -6880 40652 -6868 40708
rect -6812 40652 -6800 40708
rect -6880 40388 -6800 40652
rect -6880 40332 -6868 40388
rect -6812 40332 -6800 40388
rect -6880 40320 -6800 40332
rect -6720 40708 -6640 40720
rect -6720 40652 -6708 40708
rect -6652 40652 -6640 40708
rect -6720 40388 -6640 40652
rect -6720 40332 -6708 40388
rect -6652 40332 -6640 40388
rect -6720 40320 -6640 40332
rect -6560 40708 -6480 40720
rect -6560 40652 -6548 40708
rect -6492 40652 -6480 40708
rect -6560 40388 -6480 40652
rect -6560 40332 -6548 40388
rect -6492 40332 -6480 40388
rect -6560 40320 -6480 40332
rect -6400 40708 -6320 40720
rect -6400 40652 -6388 40708
rect -6332 40652 -6320 40708
rect -6400 40388 -6320 40652
rect -6400 40332 -6388 40388
rect -6332 40332 -6320 40388
rect -6400 40320 -6320 40332
rect -6240 40708 -6160 40720
rect -6240 40652 -6228 40708
rect -6172 40652 -6160 40708
rect -6240 40388 -6160 40652
rect -6240 40332 -6228 40388
rect -6172 40332 -6160 40388
rect -6240 40320 -6160 40332
rect -6080 40708 -6000 40720
rect -6080 40652 -6068 40708
rect -6012 40652 -6000 40708
rect -6080 40388 -6000 40652
rect -6080 40332 -6068 40388
rect -6012 40332 -6000 40388
rect -6080 40320 -6000 40332
rect -5920 40708 -5840 40720
rect -5920 40652 -5908 40708
rect -5852 40652 -5840 40708
rect -5920 40388 -5840 40652
rect -5920 40332 -5908 40388
rect -5852 40332 -5840 40388
rect -5920 40320 -5840 40332
rect -5760 40708 -5680 40720
rect -5760 40652 -5748 40708
rect -5692 40652 -5680 40708
rect -5760 40388 -5680 40652
rect -5760 40332 -5748 40388
rect -5692 40332 -5680 40388
rect -5760 40320 -5680 40332
rect -5600 40708 -5520 40720
rect -5600 40652 -5588 40708
rect -5532 40652 -5520 40708
rect -5600 40388 -5520 40652
rect -5600 40332 -5588 40388
rect -5532 40332 -5520 40388
rect -5600 40320 -5520 40332
rect -5440 40708 -5360 40720
rect -5440 40652 -5428 40708
rect -5372 40652 -5360 40708
rect -5440 40388 -5360 40652
rect -5440 40332 -5428 40388
rect -5372 40332 -5360 40388
rect -5440 40320 -5360 40332
rect -5280 40708 -5200 40720
rect -5280 40652 -5268 40708
rect -5212 40652 -5200 40708
rect -5280 40388 -5200 40652
rect -5280 40332 -5268 40388
rect -5212 40332 -5200 40388
rect -5280 40320 -5200 40332
rect -5120 40708 -5040 40720
rect -5120 40652 -5108 40708
rect -5052 40652 -5040 40708
rect -5120 40388 -5040 40652
rect -5120 40332 -5108 40388
rect -5052 40332 -5040 40388
rect -5120 40320 -5040 40332
rect -4960 40708 -4880 40720
rect -4960 40652 -4948 40708
rect -4892 40652 -4880 40708
rect -4960 40388 -4880 40652
rect -4960 40332 -4948 40388
rect -4892 40332 -4880 40388
rect -4960 40320 -4880 40332
rect -4800 40708 -4720 40720
rect -4800 40652 -4788 40708
rect -4732 40652 -4720 40708
rect -4800 40388 -4720 40652
rect -4800 40332 -4788 40388
rect -4732 40332 -4720 40388
rect -4800 40320 -4720 40332
rect -4640 40708 -4560 40720
rect -4640 40652 -4628 40708
rect -4572 40652 -4560 40708
rect -4640 40388 -4560 40652
rect -4640 40332 -4628 40388
rect -4572 40332 -4560 40388
rect -4640 40320 -4560 40332
rect -4480 40708 -4400 40720
rect -4480 40652 -4468 40708
rect -4412 40652 -4400 40708
rect -4480 40388 -4400 40652
rect -4480 40332 -4468 40388
rect -4412 40332 -4400 40388
rect -4480 40320 -4400 40332
rect -4320 40708 -4240 40720
rect -4320 40652 -4308 40708
rect -4252 40652 -4240 40708
rect -4320 40388 -4240 40652
rect -4320 40332 -4308 40388
rect -4252 40332 -4240 40388
rect -4320 40320 -4240 40332
rect -4160 40708 -4080 40720
rect -4160 40652 -4148 40708
rect -4092 40652 -4080 40708
rect -4160 40388 -4080 40652
rect -4160 40332 -4148 40388
rect -4092 40332 -4080 40388
rect -4160 40320 -4080 40332
rect -4000 40708 -3920 40720
rect -4000 40652 -3988 40708
rect -3932 40652 -3920 40708
rect -4000 40388 -3920 40652
rect -4000 40332 -3988 40388
rect -3932 40332 -3920 40388
rect -4000 40320 -3920 40332
rect -3680 40708 -3600 40720
rect -3680 40652 -3668 40708
rect -3612 40652 -3600 40708
rect -3680 40388 -3600 40652
rect -3680 40332 -3668 40388
rect -3612 40332 -3600 40388
rect -3680 40320 -3600 40332
rect -3520 40708 -3440 40720
rect -3520 40652 -3508 40708
rect -3452 40652 -3440 40708
rect -3520 40388 -3440 40652
rect -3520 40332 -3508 40388
rect -3452 40332 -3440 40388
rect -3520 40320 -3440 40332
rect -3360 40708 -3280 40812
rect -3360 40652 -3348 40708
rect -3292 40652 -3280 40708
rect -3360 40388 -3280 40652
rect -3360 40332 -3348 40388
rect -3292 40332 -3280 40388
rect -3360 40228 -3280 40332
rect -3360 40172 -3348 40228
rect -3292 40172 -3280 40228
rect -3360 40068 -3280 40172
rect -3360 40012 -3348 40068
rect -3292 40012 -3280 40068
rect -30080 39768 -30072 39832
rect -30008 39768 -30000 39832
rect -30080 39672 -30000 39768
rect -30080 39608 -30072 39672
rect -30008 39608 -30000 39672
rect -30080 39512 -30000 39608
rect -30080 39448 -30072 39512
rect -30008 39448 -30000 39512
rect -30080 39352 -30000 39448
rect -30080 39288 -30072 39352
rect -30008 39288 -30000 39352
rect -30080 39192 -30000 39288
rect -30080 39128 -30072 39192
rect -30008 39128 -30000 39192
rect -30080 39032 -30000 39128
rect -30080 38968 -30072 39032
rect -30008 38968 -30000 39032
rect -30080 38872 -30000 38968
rect -30080 38808 -30072 38872
rect -30008 38808 -30000 38872
rect -30080 38712 -30000 38808
rect -30080 38648 -30072 38712
rect -30008 38648 -30000 38712
rect -30080 38552 -30000 38648
rect -30080 38488 -30072 38552
rect -30008 38488 -30000 38552
rect -30080 38392 -30000 38488
rect -30080 38328 -30072 38392
rect -30008 38328 -30000 38392
rect -30080 38232 -30000 38328
rect -30080 38168 -30072 38232
rect -30008 38168 -30000 38232
rect -30080 38072 -30000 38168
rect -30080 38008 -30072 38072
rect -30008 38008 -30000 38072
rect -30080 37912 -30000 38008
rect -30080 37848 -30072 37912
rect -30008 37848 -30000 37912
rect -30080 37752 -30000 37848
rect -30080 37688 -30072 37752
rect -30008 37688 -30000 37752
rect -30080 37428 -30000 37688
rect -30080 37372 -30068 37428
rect -30012 37372 -30000 37428
rect -30400 37048 -30392 37112
rect -30328 37048 -30320 37112
rect -30400 36952 -30320 37048
rect -30400 36888 -30392 36952
rect -30328 36888 -30320 36952
rect -30400 36792 -30320 36888
rect -30400 36728 -30392 36792
rect -30328 36728 -30320 36792
rect -30400 36632 -30320 36728
rect -30400 36568 -30392 36632
rect -30328 36568 -30320 36632
rect -30400 36472 -30320 36568
rect -30400 36408 -30392 36472
rect -30328 36408 -30320 36472
rect -30400 36312 -30320 36408
rect -30400 36248 -30392 36312
rect -30328 36248 -30320 36312
rect -30400 36152 -30320 36248
rect -30400 36088 -30392 36152
rect -30328 36088 -30320 36152
rect -30400 35992 -30320 36088
rect -30400 35928 -30392 35992
rect -30328 35928 -30320 35992
rect -30400 35832 -30320 35928
rect -30400 35768 -30392 35832
rect -30328 35768 -30320 35832
rect -30400 35672 -30320 35768
rect -30240 35760 -30160 37120
rect -30080 37112 -30000 37372
rect -30080 37048 -30072 37112
rect -30008 37048 -30000 37112
rect -30080 36952 -30000 37048
rect -30080 36888 -30072 36952
rect -30008 36888 -30000 36952
rect -30080 36792 -30000 36888
rect -30080 36728 -30072 36792
rect -30008 36728 -30000 36792
rect -30080 36632 -30000 36728
rect -30080 36568 -30072 36632
rect -30008 36568 -30000 36632
rect -30080 36472 -30000 36568
rect -30080 36408 -30072 36472
rect -30008 36408 -30000 36472
rect -30080 36312 -30000 36408
rect -30080 36248 -30072 36312
rect -30008 36248 -30000 36312
rect -30080 36152 -30000 36248
rect -30080 36088 -30072 36152
rect -30008 36088 -30000 36152
rect -30080 35992 -30000 36088
rect -30080 35928 -30072 35992
rect -30008 35928 -30000 35992
rect -30080 35832 -30000 35928
rect -30080 35768 -30072 35832
rect -30008 35768 -30000 35832
rect -30400 35608 -30392 35672
rect -30328 35608 -30320 35672
rect -30400 35512 -30320 35608
rect -30400 35448 -30392 35512
rect -30328 35448 -30320 35512
rect -30400 35352 -30320 35448
rect -30400 35288 -30392 35352
rect -30328 35288 -30320 35352
rect -30400 35192 -30320 35288
rect -30400 35128 -30392 35192
rect -30328 35128 -30320 35192
rect -30400 35032 -30320 35128
rect -30400 34968 -30392 35032
rect -30328 34968 -30320 35032
rect -30400 34872 -30320 34968
rect -30400 34808 -30392 34872
rect -30328 34808 -30320 34872
rect -30400 34708 -30320 34808
rect -30240 34800 -30160 35680
rect -30080 35672 -30000 35768
rect -30080 35608 -30072 35672
rect -30008 35608 -30000 35672
rect -30080 35512 -30000 35608
rect -30080 35448 -30072 35512
rect -30008 35448 -30000 35512
rect -30080 35352 -30000 35448
rect -30080 35288 -30072 35352
rect -30008 35288 -30000 35352
rect -30080 35192 -30000 35288
rect -30080 35128 -30072 35192
rect -30008 35128 -30000 35192
rect -30080 35032 -30000 35128
rect -30080 34968 -30072 35032
rect -30008 34968 -30000 35032
rect -30080 34872 -30000 34968
rect -3360 39908 -3280 40012
rect -3360 39852 -3348 39908
rect -3292 39852 -3280 39908
rect -3360 39752 -3280 39852
rect -3360 39688 -3352 39752
rect -3288 39688 -3280 39752
rect -3360 39592 -3280 39688
rect -3360 39528 -3352 39592
rect -3288 39528 -3280 39592
rect -3360 39432 -3280 39528
rect -3360 39368 -3352 39432
rect -3288 39368 -3280 39432
rect -3360 39272 -3280 39368
rect -3360 39208 -3352 39272
rect -3288 39208 -3280 39272
rect -3360 39112 -3280 39208
rect -3360 39048 -3352 39112
rect -3288 39048 -3280 39112
rect -3360 38952 -3280 39048
rect -3360 38888 -3352 38952
rect -3288 38888 -3280 38952
rect -3360 38792 -3280 38888
rect -3360 38728 -3352 38792
rect -3288 38728 -3280 38792
rect -3360 38632 -3280 38728
rect -3360 38568 -3352 38632
rect -3288 38568 -3280 38632
rect -3360 38472 -3280 38568
rect -3360 38408 -3352 38472
rect -3288 38408 -3280 38472
rect -3360 38312 -3280 38408
rect -3360 38248 -3352 38312
rect -3288 38248 -3280 38312
rect -3360 38152 -3280 38248
rect -3360 38088 -3352 38152
rect -3288 38088 -3280 38152
rect -3360 37992 -3280 38088
rect -3360 37928 -3352 37992
rect -3288 37928 -3280 37992
rect -3360 37832 -3280 37928
rect -3360 37768 -3352 37832
rect -3288 37768 -3280 37832
rect -3360 37668 -3280 37768
rect -3360 37612 -3348 37668
rect -3292 37612 -3280 37668
rect -3360 37512 -3280 37612
rect -3360 37448 -3352 37512
rect -3288 37448 -3280 37512
rect -3360 37352 -3280 37448
rect -3360 37288 -3352 37352
rect -3288 37288 -3280 37352
rect -3360 37192 -3280 37288
rect -3360 37128 -3352 37192
rect -3288 37128 -3280 37192
rect -3360 37032 -3280 37128
rect -3360 36968 -3352 37032
rect -3288 36968 -3280 37032
rect -3360 36872 -3280 36968
rect -3360 36808 -3352 36872
rect -3288 36808 -3280 36872
rect -3360 36712 -3280 36808
rect -3360 36648 -3352 36712
rect -3288 36648 -3280 36712
rect -3360 36552 -3280 36648
rect -3360 36488 -3352 36552
rect -3288 36488 -3280 36552
rect -3360 36392 -3280 36488
rect -3360 36328 -3352 36392
rect -3288 36328 -3280 36392
rect -3360 36228 -3280 36328
rect -3360 36172 -3348 36228
rect -3292 36172 -3280 36228
rect -3360 36068 -3280 36172
rect -3360 36012 -3348 36068
rect -3292 36012 -3280 36068
rect -3360 35752 -3280 36012
rect -3200 42388 -3120 42400
rect -3200 42332 -3188 42388
rect -3132 42332 -3120 42388
rect -3200 35908 -3120 42332
rect -3200 35852 -3188 35908
rect -3132 35852 -3120 35908
rect -3200 35840 -3120 35852
rect -3040 42228 -2960 42492
rect -3040 42172 -3028 42228
rect -2972 42172 -2960 42228
rect -3040 41908 -2960 42172
rect -3040 41852 -3028 41908
rect -2972 41852 -2960 41908
rect -3040 41748 -2960 41852
rect -3040 41692 -3028 41748
rect -2972 41692 -2960 41748
rect -3040 41588 -2960 41692
rect -3040 41532 -3028 41588
rect -2972 41532 -2960 41588
rect -3040 40868 -2960 41532
rect -3040 40812 -3028 40868
rect -2972 40812 -2960 40868
rect -3040 40708 -2960 40812
rect -3040 40652 -3028 40708
rect -2972 40652 -2960 40708
rect -3040 40388 -2960 40652
rect -3040 40332 -3028 40388
rect -2972 40332 -2960 40388
rect -3040 40228 -2960 40332
rect -3040 40172 -3028 40228
rect -2972 40172 -2960 40228
rect -3040 40068 -2960 40172
rect -3040 40012 -3028 40068
rect -2972 40012 -2960 40068
rect -3040 39908 -2960 40012
rect -3040 39852 -3028 39908
rect -2972 39852 -2960 39908
rect -3040 39752 -2960 39852
rect -3040 39688 -3032 39752
rect -2968 39688 -2960 39752
rect -3040 39592 -2960 39688
rect -3040 39528 -3032 39592
rect -2968 39528 -2960 39592
rect -3040 39432 -2960 39528
rect -3040 39368 -3032 39432
rect -2968 39368 -2960 39432
rect -3040 39272 -2960 39368
rect -3040 39208 -3032 39272
rect -2968 39208 -2960 39272
rect -3040 39112 -2960 39208
rect -3040 39048 -3032 39112
rect -2968 39048 -2960 39112
rect -3040 38952 -2960 39048
rect -3040 38888 -3032 38952
rect -2968 38888 -2960 38952
rect -3040 38792 -2960 38888
rect -3040 38728 -3032 38792
rect -2968 38728 -2960 38792
rect -3040 38632 -2960 38728
rect -3040 38568 -3032 38632
rect -2968 38568 -2960 38632
rect -3040 38472 -2960 38568
rect -3040 38408 -3032 38472
rect -2968 38408 -2960 38472
rect -3040 38312 -2960 38408
rect -3040 38248 -3032 38312
rect -2968 38248 -2960 38312
rect -3040 38152 -2960 38248
rect -3040 38088 -3032 38152
rect -2968 38088 -2960 38152
rect -3040 37992 -2960 38088
rect -3040 37928 -3032 37992
rect -2968 37928 -2960 37992
rect -3040 37832 -2960 37928
rect -3040 37768 -3032 37832
rect -2968 37768 -2960 37832
rect -3040 37668 -2960 37768
rect -3040 37612 -3028 37668
rect -2972 37612 -2960 37668
rect -3040 37512 -2960 37612
rect -3040 37448 -3032 37512
rect -2968 37448 -2960 37512
rect -3040 37352 -2960 37448
rect -3040 37288 -3032 37352
rect -2968 37288 -2960 37352
rect -3040 37192 -2960 37288
rect -3040 37128 -3032 37192
rect -2968 37128 -2960 37192
rect -3040 37032 -2960 37128
rect -3040 36968 -3032 37032
rect -2968 36968 -2960 37032
rect -3040 36872 -2960 36968
rect -3040 36808 -3032 36872
rect -2968 36808 -2960 36872
rect -3040 36712 -2960 36808
rect -3040 36648 -3032 36712
rect -2968 36648 -2960 36712
rect -3040 36552 -2960 36648
rect -3040 36488 -3032 36552
rect -2968 36488 -2960 36552
rect -3040 36392 -2960 36488
rect -3040 36328 -3032 36392
rect -2968 36328 -2960 36392
rect -3040 36228 -2960 36328
rect -3040 36172 -3028 36228
rect -2972 36172 -2960 36228
rect -3040 36068 -2960 36172
rect -2880 42708 -2800 42720
rect -2880 42652 -2868 42708
rect -2812 42652 -2800 42708
rect -2880 36228 -2800 42652
rect -2880 36172 -2868 36228
rect -2812 36172 -2800 36228
rect -2880 36160 -2800 36172
rect -2720 42548 -2640 42812
rect -2720 42492 -2708 42548
rect -2652 42492 -2640 42548
rect -2720 42228 -2640 42492
rect -2720 42172 -2708 42228
rect -2652 42172 -2640 42228
rect -2720 41908 -2640 42172
rect -2720 41852 -2708 41908
rect -2652 41852 -2640 41908
rect -2720 41748 -2640 41852
rect -2560 42868 -2480 42880
rect -2560 42812 -2548 42868
rect -2492 42812 -2480 42868
rect -2560 42548 -2480 42812
rect -2560 42492 -2548 42548
rect -2492 42492 -2480 42548
rect -2560 42228 -2480 42492
rect -2560 42172 -2548 42228
rect -2492 42172 -2480 42228
rect -2560 41908 -2480 42172
rect -2560 41852 -2548 41908
rect -2492 41852 -2480 41908
rect -2560 41840 -2480 41852
rect -2400 42868 -2320 42880
rect -2400 42812 -2388 42868
rect -2332 42812 -2320 42868
rect -2400 42548 -2320 42812
rect -2400 42492 -2388 42548
rect -2332 42492 -2320 42548
rect -2400 42228 -2320 42492
rect -2400 42172 -2388 42228
rect -2332 42172 -2320 42228
rect -2400 41908 -2320 42172
rect -2400 41852 -2388 41908
rect -2332 41852 -2320 41908
rect -2720 41692 -2708 41748
rect -2652 41692 -2640 41748
rect -2720 41588 -2640 41692
rect -2720 41532 -2708 41588
rect -2652 41532 -2640 41588
rect -2720 40868 -2640 41532
rect -2720 40812 -2708 40868
rect -2652 40812 -2640 40868
rect -2720 40708 -2640 40812
rect -2720 40652 -2708 40708
rect -2652 40652 -2640 40708
rect -2720 40388 -2640 40652
rect -2720 40332 -2708 40388
rect -2652 40332 -2640 40388
rect -2720 40228 -2640 40332
rect -2400 41748 -2320 41852
rect -2240 42868 -2160 42880
rect -2240 42812 -2228 42868
rect -2172 42812 -2160 42868
rect -2240 42548 -2160 42812
rect -2240 42492 -2228 42548
rect -2172 42492 -2160 42548
rect -2240 42228 -2160 42492
rect -2240 42172 -2228 42228
rect -2172 42172 -2160 42228
rect -2240 41908 -2160 42172
rect -2240 41852 -2228 41908
rect -2172 41852 -2160 41908
rect -2240 41840 -2160 41852
rect -2080 42868 -2000 42960
rect -2080 42812 -2068 42868
rect -2012 42812 -2000 42868
rect -2080 42548 -2000 42812
rect -2080 42492 -2068 42548
rect -2012 42492 -2000 42548
rect -2080 42228 -2000 42492
rect -2080 42172 -2068 42228
rect -2012 42172 -2000 42228
rect -2080 41908 -2000 42172
rect -2080 41852 -2068 41908
rect -2012 41852 -2000 41908
rect -2400 41692 -2388 41748
rect -2332 41692 -2320 41748
rect -2400 41588 -2320 41692
rect -2400 41532 -2388 41588
rect -2332 41532 -2320 41588
rect -2400 40868 -2320 41532
rect -2400 40812 -2388 40868
rect -2332 40812 -2320 40868
rect -2400 40708 -2320 40812
rect -2400 40652 -2388 40708
rect -2332 40652 -2320 40708
rect -2400 40388 -2320 40652
rect -2400 40332 -2388 40388
rect -2332 40332 -2320 40388
rect -2720 40172 -2708 40228
rect -2652 40172 -2640 40228
rect -2720 40068 -2640 40172
rect -2720 40012 -2708 40068
rect -2652 40012 -2640 40068
rect -2720 39908 -2640 40012
rect -2720 39852 -2708 39908
rect -2652 39852 -2640 39908
rect -2720 39752 -2640 39852
rect -2720 39688 -2712 39752
rect -2648 39688 -2640 39752
rect -2720 39592 -2640 39688
rect -2720 39528 -2712 39592
rect -2648 39528 -2640 39592
rect -2720 39432 -2640 39528
rect -2720 39368 -2712 39432
rect -2648 39368 -2640 39432
rect -2720 39272 -2640 39368
rect -2720 39208 -2712 39272
rect -2648 39208 -2640 39272
rect -2720 39112 -2640 39208
rect -2720 39048 -2712 39112
rect -2648 39048 -2640 39112
rect -2720 38952 -2640 39048
rect -2720 38888 -2712 38952
rect -2648 38888 -2640 38952
rect -2720 38792 -2640 38888
rect -2720 38728 -2712 38792
rect -2648 38728 -2640 38792
rect -2720 38632 -2640 38728
rect -2720 38568 -2712 38632
rect -2648 38568 -2640 38632
rect -2720 38472 -2640 38568
rect -2720 38408 -2712 38472
rect -2648 38408 -2640 38472
rect -2720 38312 -2640 38408
rect -2720 38248 -2712 38312
rect -2648 38248 -2640 38312
rect -2720 38152 -2640 38248
rect -2720 38088 -2712 38152
rect -2648 38088 -2640 38152
rect -2720 37992 -2640 38088
rect -2720 37928 -2712 37992
rect -2648 37928 -2640 37992
rect -2720 37832 -2640 37928
rect -2720 37768 -2712 37832
rect -2648 37768 -2640 37832
rect -2720 37668 -2640 37768
rect -2720 37612 -2708 37668
rect -2652 37612 -2640 37668
rect -2720 37512 -2640 37612
rect -2720 37448 -2712 37512
rect -2648 37448 -2640 37512
rect -2720 37352 -2640 37448
rect -2720 37288 -2712 37352
rect -2648 37288 -2640 37352
rect -2720 37192 -2640 37288
rect -2720 37128 -2712 37192
rect -2648 37128 -2640 37192
rect -2720 37032 -2640 37128
rect -2720 36968 -2712 37032
rect -2648 36968 -2640 37032
rect -2720 36872 -2640 36968
rect -2720 36808 -2712 36872
rect -2648 36808 -2640 36872
rect -2720 36712 -2640 36808
rect -2720 36648 -2712 36712
rect -2648 36648 -2640 36712
rect -2720 36552 -2640 36648
rect -2720 36488 -2712 36552
rect -2648 36488 -2640 36552
rect -2720 36392 -2640 36488
rect -2720 36328 -2712 36392
rect -2648 36328 -2640 36392
rect -3040 36012 -3028 36068
rect -2972 36012 -2960 36068
rect -3360 35688 -3352 35752
rect -3288 35688 -3280 35752
rect -3360 35592 -3280 35688
rect -3360 35528 -3352 35592
rect -3288 35528 -3280 35592
rect -3360 35432 -3280 35528
rect -3360 35368 -3352 35432
rect -3288 35368 -3280 35432
rect -3360 35272 -3280 35368
rect -3360 35208 -3352 35272
rect -3288 35208 -3280 35272
rect -3360 35112 -3280 35208
rect -3360 35048 -3352 35112
rect -3288 35048 -3280 35112
rect -3360 34952 -3280 35048
rect -3360 34888 -3352 34952
rect -3288 34888 -3280 34952
rect -30080 34808 -30072 34872
rect -30008 34808 -30000 34872
rect -30400 34652 -30388 34708
rect -30332 34652 -30320 34708
rect -30400 34388 -30320 34652
rect -30400 34332 -30388 34388
rect -30332 34332 -30320 34388
rect -30400 34232 -30320 34332
rect -30080 34708 -30000 34808
rect -30080 34652 -30068 34708
rect -30012 34652 -30000 34708
rect -30080 34388 -30000 34652
rect -30080 34332 -30068 34388
rect -30012 34332 -30000 34388
rect -30400 34168 -30392 34232
rect -30328 34168 -30320 34232
rect -30400 34072 -30320 34168
rect -30400 34008 -30392 34072
rect -30328 34008 -30320 34072
rect -30400 33912 -30320 34008
rect -30400 33848 -30392 33912
rect -30328 33848 -30320 33912
rect -30400 33752 -30320 33848
rect -30400 33688 -30392 33752
rect -30328 33688 -30320 33752
rect -30400 33592 -30320 33688
rect -30400 33528 -30392 33592
rect -30328 33528 -30320 33592
rect -30400 33432 -30320 33528
rect -30400 33368 -30392 33432
rect -30328 33368 -30320 33432
rect -30400 33272 -30320 33368
rect -30400 33208 -30392 33272
rect -30328 33208 -30320 33272
rect -30400 33112 -30320 33208
rect -30400 33048 -30392 33112
rect -30328 33048 -30320 33112
rect -30400 32952 -30320 33048
rect -30400 32888 -30392 32952
rect -30328 32888 -30320 32952
rect -30720 32572 -30708 32628
rect -30652 32572 -30640 32628
rect -30720 32468 -30640 32572
rect -30720 32412 -30708 32468
rect -30652 32412 -30640 32468
rect -30720 32308 -30640 32412
rect -30720 32252 -30708 32308
rect -30652 32252 -30640 32308
rect -30720 32148 -30640 32252
rect -30400 32628 -30320 32888
rect -30240 32880 -30160 34240
rect -30080 34232 -30000 34332
rect -29920 34708 -29840 34720
rect -29920 34652 -29908 34708
rect -29852 34652 -29840 34708
rect -29920 34388 -29840 34652
rect -29920 34332 -29908 34388
rect -29852 34332 -29840 34388
rect -29920 34320 -29840 34332
rect -29760 34708 -29680 34720
rect -29760 34652 -29748 34708
rect -29692 34652 -29680 34708
rect -29760 34388 -29680 34652
rect -29760 34332 -29748 34388
rect -29692 34332 -29680 34388
rect -29760 34320 -29680 34332
rect -29600 34708 -29520 34720
rect -29600 34652 -29588 34708
rect -29532 34652 -29520 34708
rect -29600 34388 -29520 34652
rect -29600 34332 -29588 34388
rect -29532 34332 -29520 34388
rect -29600 34320 -29520 34332
rect -29440 34708 -29360 34720
rect -29440 34652 -29428 34708
rect -29372 34652 -29360 34708
rect -29440 34388 -29360 34652
rect -29440 34332 -29428 34388
rect -29372 34332 -29360 34388
rect -29440 34320 -29360 34332
rect -29280 34708 -29200 34720
rect -29280 34652 -29268 34708
rect -29212 34652 -29200 34708
rect -29280 34388 -29200 34652
rect -29280 34332 -29268 34388
rect -29212 34332 -29200 34388
rect -29280 34320 -29200 34332
rect -29120 34708 -29040 34720
rect -29120 34652 -29108 34708
rect -29052 34652 -29040 34708
rect -29120 34388 -29040 34652
rect -29120 34332 -29108 34388
rect -29052 34332 -29040 34388
rect -29120 34320 -29040 34332
rect -28960 34708 -28880 34720
rect -28960 34652 -28948 34708
rect -28892 34652 -28880 34708
rect -28960 34388 -28880 34652
rect -28960 34332 -28948 34388
rect -28892 34332 -28880 34388
rect -28960 34320 -28880 34332
rect -28800 34708 -28720 34720
rect -28800 34652 -28788 34708
rect -28732 34652 -28720 34708
rect -28800 34388 -28720 34652
rect -28800 34332 -28788 34388
rect -28732 34332 -28720 34388
rect -28800 34320 -28720 34332
rect -28640 34708 -28560 34720
rect -28640 34652 -28628 34708
rect -28572 34652 -28560 34708
rect -28640 34388 -28560 34652
rect -28640 34332 -28628 34388
rect -28572 34332 -28560 34388
rect -28640 34320 -28560 34332
rect -28480 34708 -28400 34720
rect -28480 34652 -28468 34708
rect -28412 34652 -28400 34708
rect -28480 34388 -28400 34652
rect -28480 34332 -28468 34388
rect -28412 34332 -28400 34388
rect -28480 34320 -28400 34332
rect -28320 34708 -28240 34720
rect -28320 34652 -28308 34708
rect -28252 34652 -28240 34708
rect -28320 34388 -28240 34652
rect -28320 34332 -28308 34388
rect -28252 34332 -28240 34388
rect -28320 34320 -28240 34332
rect -28160 34708 -28080 34720
rect -28160 34652 -28148 34708
rect -28092 34652 -28080 34708
rect -28160 34388 -28080 34652
rect -28160 34332 -28148 34388
rect -28092 34332 -28080 34388
rect -28160 34320 -28080 34332
rect -28000 34708 -27920 34720
rect -28000 34652 -27988 34708
rect -27932 34652 -27920 34708
rect -28000 34388 -27920 34652
rect -28000 34332 -27988 34388
rect -27932 34332 -27920 34388
rect -28000 34320 -27920 34332
rect -27840 34708 -27760 34720
rect -27840 34652 -27828 34708
rect -27772 34652 -27760 34708
rect -27840 34388 -27760 34652
rect -27840 34332 -27828 34388
rect -27772 34332 -27760 34388
rect -27840 34320 -27760 34332
rect -27680 34708 -27600 34720
rect -27680 34652 -27668 34708
rect -27612 34652 -27600 34708
rect -27680 34388 -27600 34652
rect -27680 34332 -27668 34388
rect -27612 34332 -27600 34388
rect -27680 34320 -27600 34332
rect -27520 34708 -27440 34720
rect -27520 34652 -27508 34708
rect -27452 34652 -27440 34708
rect -27520 34388 -27440 34652
rect -27520 34332 -27508 34388
rect -27452 34332 -27440 34388
rect -27520 34320 -27440 34332
rect -27360 34708 -27280 34720
rect -27360 34652 -27348 34708
rect -27292 34652 -27280 34708
rect -27360 34388 -27280 34652
rect -27360 34332 -27348 34388
rect -27292 34332 -27280 34388
rect -27360 34320 -27280 34332
rect -27200 34708 -27120 34720
rect -27200 34652 -27188 34708
rect -27132 34652 -27120 34708
rect -27200 34388 -27120 34652
rect -27200 34332 -27188 34388
rect -27132 34332 -27120 34388
rect -27200 34320 -27120 34332
rect -27040 34708 -26960 34720
rect -27040 34652 -27028 34708
rect -26972 34652 -26960 34708
rect -27040 34388 -26960 34652
rect -27040 34332 -27028 34388
rect -26972 34332 -26960 34388
rect -27040 34320 -26960 34332
rect -26880 34708 -26800 34720
rect -26880 34652 -26868 34708
rect -26812 34652 -26800 34708
rect -26880 34388 -26800 34652
rect -26880 34332 -26868 34388
rect -26812 34332 -26800 34388
rect -26880 34320 -26800 34332
rect -26720 34708 -26640 34720
rect -26720 34652 -26708 34708
rect -26652 34652 -26640 34708
rect -26720 34388 -26640 34652
rect -26720 34332 -26708 34388
rect -26652 34332 -26640 34388
rect -26720 34320 -26640 34332
rect -26560 34708 -26480 34720
rect -26560 34652 -26548 34708
rect -26492 34652 -26480 34708
rect -26560 34388 -26480 34652
rect -26560 34332 -26548 34388
rect -26492 34332 -26480 34388
rect -26560 34320 -26480 34332
rect -26400 34708 -26320 34720
rect -26400 34652 -26388 34708
rect -26332 34652 -26320 34708
rect -26400 34388 -26320 34652
rect -26400 34332 -26388 34388
rect -26332 34332 -26320 34388
rect -26400 34320 -26320 34332
rect -26240 34708 -26160 34720
rect -26240 34652 -26228 34708
rect -26172 34652 -26160 34708
rect -26240 34388 -26160 34652
rect -26240 34332 -26228 34388
rect -26172 34332 -26160 34388
rect -26240 34320 -26160 34332
rect -26080 34708 -26000 34720
rect -26080 34652 -26068 34708
rect -26012 34652 -26000 34708
rect -26080 34388 -26000 34652
rect -26080 34332 -26068 34388
rect -26012 34332 -26000 34388
rect -26080 34320 -26000 34332
rect -25920 34708 -25840 34720
rect -25920 34652 -25908 34708
rect -25852 34652 -25840 34708
rect -25920 34388 -25840 34652
rect -25920 34332 -25908 34388
rect -25852 34332 -25840 34388
rect -25920 34320 -25840 34332
rect -25760 34708 -25680 34720
rect -25760 34652 -25748 34708
rect -25692 34652 -25680 34708
rect -25760 34388 -25680 34652
rect -25760 34332 -25748 34388
rect -25692 34332 -25680 34388
rect -25760 34320 -25680 34332
rect -25600 34708 -25520 34720
rect -25600 34652 -25588 34708
rect -25532 34652 -25520 34708
rect -25600 34388 -25520 34652
rect -25600 34332 -25588 34388
rect -25532 34332 -25520 34388
rect -25600 34320 -25520 34332
rect -25440 34708 -25360 34720
rect -25440 34652 -25428 34708
rect -25372 34652 -25360 34708
rect -25440 34388 -25360 34652
rect -25440 34332 -25428 34388
rect -25372 34332 -25360 34388
rect -25440 34320 -25360 34332
rect -25280 34708 -25200 34720
rect -25280 34652 -25268 34708
rect -25212 34652 -25200 34708
rect -25280 34388 -25200 34652
rect -25280 34332 -25268 34388
rect -25212 34332 -25200 34388
rect -25280 34320 -25200 34332
rect -25120 34708 -25040 34720
rect -25120 34652 -25108 34708
rect -25052 34652 -25040 34708
rect -25120 34388 -25040 34652
rect -25120 34332 -25108 34388
rect -25052 34332 -25040 34388
rect -25120 34320 -25040 34332
rect -24960 34708 -24880 34720
rect -24960 34652 -24948 34708
rect -24892 34652 -24880 34708
rect -24960 34388 -24880 34652
rect -24960 34332 -24948 34388
rect -24892 34332 -24880 34388
rect -24960 34320 -24880 34332
rect -24800 34708 -24720 34720
rect -24800 34652 -24788 34708
rect -24732 34652 -24720 34708
rect -24800 34388 -24720 34652
rect -24800 34332 -24788 34388
rect -24732 34332 -24720 34388
rect -24800 34320 -24720 34332
rect -24640 34708 -24560 34720
rect -24640 34652 -24628 34708
rect -24572 34652 -24560 34708
rect -24640 34388 -24560 34652
rect -24640 34332 -24628 34388
rect -24572 34332 -24560 34388
rect -24640 34320 -24560 34332
rect -24480 34708 -24400 34720
rect -24480 34652 -24468 34708
rect -24412 34652 -24400 34708
rect -24480 34388 -24400 34652
rect -24480 34332 -24468 34388
rect -24412 34332 -24400 34388
rect -24480 34320 -24400 34332
rect -24320 34708 -24240 34720
rect -24320 34652 -24308 34708
rect -24252 34652 -24240 34708
rect -24320 34388 -24240 34652
rect -24320 34332 -24308 34388
rect -24252 34332 -24240 34388
rect -24320 34320 -24240 34332
rect -24160 34708 -24080 34720
rect -24160 34652 -24148 34708
rect -24092 34652 -24080 34708
rect -24160 34388 -24080 34652
rect -24160 34332 -24148 34388
rect -24092 34332 -24080 34388
rect -24160 34320 -24080 34332
rect -24000 34708 -23920 34720
rect -24000 34652 -23988 34708
rect -23932 34652 -23920 34708
rect -24000 34388 -23920 34652
rect -24000 34332 -23988 34388
rect -23932 34332 -23920 34388
rect -24000 34320 -23920 34332
rect -23840 34708 -23760 34720
rect -23840 34652 -23828 34708
rect -23772 34652 -23760 34708
rect -23840 34388 -23760 34652
rect -23840 34332 -23828 34388
rect -23772 34332 -23760 34388
rect -23840 34320 -23760 34332
rect -23680 34708 -23600 34720
rect -23680 34652 -23668 34708
rect -23612 34652 -23600 34708
rect -23680 34388 -23600 34652
rect -23680 34332 -23668 34388
rect -23612 34332 -23600 34388
rect -23680 34320 -23600 34332
rect -23520 34708 -23440 34720
rect -23520 34652 -23508 34708
rect -23452 34652 -23440 34708
rect -23520 34388 -23440 34652
rect -23520 34332 -23508 34388
rect -23452 34332 -23440 34388
rect -23520 34320 -23440 34332
rect -23360 34708 -23280 34720
rect -23360 34652 -23348 34708
rect -23292 34652 -23280 34708
rect -23360 34388 -23280 34652
rect -23360 34332 -23348 34388
rect -23292 34332 -23280 34388
rect -23360 34320 -23280 34332
rect -23200 34708 -23120 34720
rect -23200 34652 -23188 34708
rect -23132 34652 -23120 34708
rect -23200 34388 -23120 34652
rect -23200 34332 -23188 34388
rect -23132 34332 -23120 34388
rect -23200 34320 -23120 34332
rect -23040 34708 -22960 34720
rect -23040 34652 -23028 34708
rect -22972 34652 -22960 34708
rect -23040 34388 -22960 34652
rect -23040 34332 -23028 34388
rect -22972 34332 -22960 34388
rect -23040 34320 -22960 34332
rect -22880 34708 -22800 34720
rect -22880 34652 -22868 34708
rect -22812 34652 -22800 34708
rect -22880 34388 -22800 34652
rect -22880 34332 -22868 34388
rect -22812 34332 -22800 34388
rect -22880 34320 -22800 34332
rect -22720 34708 -22640 34720
rect -22720 34652 -22708 34708
rect -22652 34652 -22640 34708
rect -22720 34388 -22640 34652
rect -22720 34332 -22708 34388
rect -22652 34332 -22640 34388
rect -22720 34320 -22640 34332
rect -22560 34708 -22480 34720
rect -22560 34652 -22548 34708
rect -22492 34652 -22480 34708
rect -22560 34388 -22480 34652
rect -22560 34332 -22548 34388
rect -22492 34332 -22480 34388
rect -22560 34320 -22480 34332
rect -22400 34708 -22320 34720
rect -22400 34652 -22388 34708
rect -22332 34652 -22320 34708
rect -22400 34388 -22320 34652
rect -22400 34332 -22388 34388
rect -22332 34332 -22320 34388
rect -22400 34320 -22320 34332
rect -22240 34708 -22160 34720
rect -22240 34652 -22228 34708
rect -22172 34652 -22160 34708
rect -22240 34388 -22160 34652
rect -22240 34332 -22228 34388
rect -22172 34332 -22160 34388
rect -22240 34320 -22160 34332
rect -22080 34708 -22000 34720
rect -22080 34652 -22068 34708
rect -22012 34652 -22000 34708
rect -22080 34388 -22000 34652
rect -22080 34332 -22068 34388
rect -22012 34332 -22000 34388
rect -22080 34320 -22000 34332
rect -21920 34708 -21840 34720
rect -21920 34652 -21908 34708
rect -21852 34652 -21840 34708
rect -21920 34388 -21840 34652
rect -21920 34332 -21908 34388
rect -21852 34332 -21840 34388
rect -21920 34320 -21840 34332
rect -21760 34708 -21680 34720
rect -21760 34652 -21748 34708
rect -21692 34652 -21680 34708
rect -21760 34388 -21680 34652
rect -21760 34332 -21748 34388
rect -21692 34332 -21680 34388
rect -21760 34320 -21680 34332
rect -21600 34708 -21520 34720
rect -21600 34652 -21588 34708
rect -21532 34652 -21520 34708
rect -21600 34388 -21520 34652
rect -21600 34332 -21588 34388
rect -21532 34332 -21520 34388
rect -21600 34320 -21520 34332
rect -21440 34708 -21360 34720
rect -21440 34652 -21428 34708
rect -21372 34652 -21360 34708
rect -21440 34388 -21360 34652
rect -21440 34332 -21428 34388
rect -21372 34332 -21360 34388
rect -21440 34320 -21360 34332
rect -21280 34708 -21200 34720
rect -21280 34652 -21268 34708
rect -21212 34652 -21200 34708
rect -21280 34388 -21200 34652
rect -21280 34332 -21268 34388
rect -21212 34332 -21200 34388
rect -21280 34320 -21200 34332
rect -21120 34708 -21040 34720
rect -21120 34652 -21108 34708
rect -21052 34652 -21040 34708
rect -21120 34388 -21040 34652
rect -21120 34332 -21108 34388
rect -21052 34332 -21040 34388
rect -21120 34320 -21040 34332
rect -20960 34708 -20880 34720
rect -20960 34652 -20948 34708
rect -20892 34652 -20880 34708
rect -20960 34388 -20880 34652
rect -20960 34332 -20948 34388
rect -20892 34332 -20880 34388
rect -20960 34320 -20880 34332
rect -20800 34708 -20720 34720
rect -20800 34652 -20788 34708
rect -20732 34652 -20720 34708
rect -20800 34388 -20720 34652
rect -20800 34332 -20788 34388
rect -20732 34332 -20720 34388
rect -20800 34320 -20720 34332
rect -20640 34708 -20560 34720
rect -20640 34652 -20628 34708
rect -20572 34652 -20560 34708
rect -20640 34388 -20560 34652
rect -20640 34332 -20628 34388
rect -20572 34332 -20560 34388
rect -20640 34320 -20560 34332
rect -20480 34708 -20400 34720
rect -20480 34652 -20468 34708
rect -20412 34652 -20400 34708
rect -20480 34388 -20400 34652
rect -20480 34332 -20468 34388
rect -20412 34332 -20400 34388
rect -20480 34320 -20400 34332
rect -20320 34708 -20240 34720
rect -20320 34652 -20308 34708
rect -20252 34652 -20240 34708
rect -20320 34388 -20240 34652
rect -20320 34332 -20308 34388
rect -20252 34332 -20240 34388
rect -20320 34320 -20240 34332
rect -20160 34708 -20080 34720
rect -20160 34652 -20148 34708
rect -20092 34652 -20080 34708
rect -20160 34388 -20080 34652
rect -20160 34332 -20148 34388
rect -20092 34332 -20080 34388
rect -20160 34320 -20080 34332
rect -20000 34708 -19920 34720
rect -20000 34652 -19988 34708
rect -19932 34652 -19920 34708
rect -20000 34388 -19920 34652
rect -20000 34332 -19988 34388
rect -19932 34332 -19920 34388
rect -20000 34320 -19920 34332
rect -19840 34708 -19760 34720
rect -19840 34652 -19828 34708
rect -19772 34652 -19760 34708
rect -19840 34388 -19760 34652
rect -19840 34332 -19828 34388
rect -19772 34332 -19760 34388
rect -19840 34320 -19760 34332
rect -19680 34708 -19600 34720
rect -19680 34652 -19668 34708
rect -19612 34652 -19600 34708
rect -19680 34388 -19600 34652
rect -19680 34332 -19668 34388
rect -19612 34332 -19600 34388
rect -19680 34320 -19600 34332
rect -19520 34708 -19440 34720
rect -19520 34652 -19508 34708
rect -19452 34652 -19440 34708
rect -19520 34388 -19440 34652
rect -19520 34332 -19508 34388
rect -19452 34332 -19440 34388
rect -19520 34320 -19440 34332
rect -19360 34708 -19280 34720
rect -19360 34652 -19348 34708
rect -19292 34652 -19280 34708
rect -19360 34388 -19280 34652
rect -19360 34332 -19348 34388
rect -19292 34332 -19280 34388
rect -19360 34320 -19280 34332
rect -19200 34708 -19120 34720
rect -19200 34652 -19188 34708
rect -19132 34652 -19120 34708
rect -19200 34388 -19120 34652
rect -19200 34332 -19188 34388
rect -19132 34332 -19120 34388
rect -19200 34320 -19120 34332
rect -19040 34708 -18960 34720
rect -19040 34652 -19028 34708
rect -18972 34652 -18960 34708
rect -19040 34388 -18960 34652
rect -19040 34332 -19028 34388
rect -18972 34332 -18960 34388
rect -19040 34320 -18960 34332
rect -18880 34708 -18800 34720
rect -18880 34652 -18868 34708
rect -18812 34652 -18800 34708
rect -18880 34388 -18800 34652
rect -18880 34332 -18868 34388
rect -18812 34332 -18800 34388
rect -18880 34320 -18800 34332
rect -18720 34708 -18640 34720
rect -18720 34652 -18708 34708
rect -18652 34652 -18640 34708
rect -18720 34388 -18640 34652
rect -18720 34332 -18708 34388
rect -18652 34332 -18640 34388
rect -18720 34320 -18640 34332
rect -18560 34708 -18480 34720
rect -18560 34652 -18548 34708
rect -18492 34652 -18480 34708
rect -18560 34388 -18480 34652
rect -18560 34332 -18548 34388
rect -18492 34332 -18480 34388
rect -18560 34320 -18480 34332
rect -18400 34708 -18320 34720
rect -18400 34652 -18388 34708
rect -18332 34652 -18320 34708
rect -18400 34388 -18320 34652
rect -18400 34332 -18388 34388
rect -18332 34332 -18320 34388
rect -18400 34320 -18320 34332
rect -18240 34708 -18160 34720
rect -18240 34652 -18228 34708
rect -18172 34652 -18160 34708
rect -18240 34388 -18160 34652
rect -18240 34332 -18228 34388
rect -18172 34332 -18160 34388
rect -18240 34320 -18160 34332
rect -18080 34708 -18000 34720
rect -18080 34652 -18068 34708
rect -18012 34652 -18000 34708
rect -18080 34388 -18000 34652
rect -18080 34332 -18068 34388
rect -18012 34332 -18000 34388
rect -18080 34320 -18000 34332
rect -17920 34708 -17840 34720
rect -17920 34652 -17908 34708
rect -17852 34652 -17840 34708
rect -17920 34388 -17840 34652
rect -17920 34332 -17908 34388
rect -17852 34332 -17840 34388
rect -17920 34320 -17840 34332
rect -17760 34708 -17680 34720
rect -17760 34652 -17748 34708
rect -17692 34652 -17680 34708
rect -17760 34388 -17680 34652
rect -17760 34332 -17748 34388
rect -17692 34332 -17680 34388
rect -17760 34320 -17680 34332
rect -17600 34708 -17520 34720
rect -17600 34652 -17588 34708
rect -17532 34652 -17520 34708
rect -17600 34388 -17520 34652
rect -17600 34332 -17588 34388
rect -17532 34332 -17520 34388
rect -17600 34320 -17520 34332
rect -17440 34708 -17360 34720
rect -17440 34652 -17428 34708
rect -17372 34652 -17360 34708
rect -17440 34388 -17360 34652
rect -17440 34332 -17428 34388
rect -17372 34332 -17360 34388
rect -17440 34320 -17360 34332
rect -17280 34708 -17200 34720
rect -17280 34652 -17268 34708
rect -17212 34652 -17200 34708
rect -17280 34388 -17200 34652
rect -17280 34332 -17268 34388
rect -17212 34332 -17200 34388
rect -17280 34320 -17200 34332
rect -17120 34708 -17040 34720
rect -17120 34652 -17108 34708
rect -17052 34652 -17040 34708
rect -17120 34388 -17040 34652
rect -17120 34332 -17108 34388
rect -17052 34332 -17040 34388
rect -17120 34320 -17040 34332
rect -16960 34708 -16880 34720
rect -16960 34652 -16948 34708
rect -16892 34652 -16880 34708
rect -16960 34388 -16880 34652
rect -16960 34332 -16948 34388
rect -16892 34332 -16880 34388
rect -16960 34320 -16880 34332
rect -16800 34708 -16720 34720
rect -16800 34652 -16788 34708
rect -16732 34652 -16720 34708
rect -16800 34388 -16720 34652
rect -16800 34332 -16788 34388
rect -16732 34332 -16720 34388
rect -16800 34320 -16720 34332
rect -16640 34708 -16560 34720
rect -16640 34652 -16628 34708
rect -16572 34652 -16560 34708
rect -16640 34388 -16560 34652
rect -16640 34332 -16628 34388
rect -16572 34332 -16560 34388
rect -16640 34320 -16560 34332
rect -16480 34708 -16400 34720
rect -16480 34652 -16468 34708
rect -16412 34652 -16400 34708
rect -16480 34388 -16400 34652
rect -16480 34332 -16468 34388
rect -16412 34332 -16400 34388
rect -16480 34320 -16400 34332
rect -16320 34708 -16240 34720
rect -16320 34652 -16308 34708
rect -16252 34652 -16240 34708
rect -16320 34388 -16240 34652
rect -16320 34332 -16308 34388
rect -16252 34332 -16240 34388
rect -16320 34320 -16240 34332
rect -16160 34708 -16080 34720
rect -16160 34652 -16148 34708
rect -16092 34652 -16080 34708
rect -16160 34388 -16080 34652
rect -16160 34332 -16148 34388
rect -16092 34332 -16080 34388
rect -16160 34320 -16080 34332
rect -16000 34708 -15920 34720
rect -16000 34652 -15988 34708
rect -15932 34652 -15920 34708
rect -16000 34388 -15920 34652
rect -16000 34332 -15988 34388
rect -15932 34332 -15920 34388
rect -16000 34320 -15920 34332
rect -15840 34708 -15760 34720
rect -15840 34652 -15828 34708
rect -15772 34652 -15760 34708
rect -15840 34388 -15760 34652
rect -15840 34332 -15828 34388
rect -15772 34332 -15760 34388
rect -15840 34320 -15760 34332
rect -15680 34708 -15600 34720
rect -15680 34652 -15668 34708
rect -15612 34652 -15600 34708
rect -15680 34388 -15600 34652
rect -15680 34332 -15668 34388
rect -15612 34332 -15600 34388
rect -15680 34320 -15600 34332
rect -15520 34708 -15440 34720
rect -15520 34652 -15508 34708
rect -15452 34652 -15440 34708
rect -15520 34388 -15440 34652
rect -15520 34332 -15508 34388
rect -15452 34332 -15440 34388
rect -15520 34320 -15440 34332
rect -15360 34708 -15280 34720
rect -15360 34652 -15348 34708
rect -15292 34652 -15280 34708
rect -15360 34388 -15280 34652
rect -15360 34332 -15348 34388
rect -15292 34332 -15280 34388
rect -15360 34320 -15280 34332
rect -15200 34708 -15120 34720
rect -15200 34652 -15188 34708
rect -15132 34652 -15120 34708
rect -15200 34388 -15120 34652
rect -15200 34332 -15188 34388
rect -15132 34332 -15120 34388
rect -15200 34320 -15120 34332
rect -15040 34708 -14960 34720
rect -15040 34652 -15028 34708
rect -14972 34652 -14960 34708
rect -15040 34388 -14960 34652
rect -15040 34332 -15028 34388
rect -14972 34332 -14960 34388
rect -15040 34320 -14960 34332
rect -14880 34708 -14800 34720
rect -14880 34652 -14868 34708
rect -14812 34652 -14800 34708
rect -14880 34388 -14800 34652
rect -14880 34332 -14868 34388
rect -14812 34332 -14800 34388
rect -14880 34320 -14800 34332
rect -14720 34708 -14640 34720
rect -14720 34652 -14708 34708
rect -14652 34652 -14640 34708
rect -14720 34388 -14640 34652
rect -14720 34332 -14708 34388
rect -14652 34332 -14640 34388
rect -14720 34320 -14640 34332
rect -14560 34708 -14480 34720
rect -14560 34652 -14548 34708
rect -14492 34652 -14480 34708
rect -14560 34388 -14480 34652
rect -14560 34332 -14548 34388
rect -14492 34332 -14480 34388
rect -14560 34320 -14480 34332
rect -14400 34708 -14320 34720
rect -14400 34652 -14388 34708
rect -14332 34652 -14320 34708
rect -14400 34388 -14320 34652
rect -14400 34332 -14388 34388
rect -14332 34332 -14320 34388
rect -14400 34320 -14320 34332
rect -14240 34708 -14160 34720
rect -14240 34652 -14228 34708
rect -14172 34652 -14160 34708
rect -14240 34388 -14160 34652
rect -14240 34332 -14228 34388
rect -14172 34332 -14160 34388
rect -14240 34320 -14160 34332
rect -14080 34708 -14000 34720
rect -14080 34652 -14068 34708
rect -14012 34652 -14000 34708
rect -14080 34388 -14000 34652
rect -14080 34332 -14068 34388
rect -14012 34332 -14000 34388
rect -14080 34320 -14000 34332
rect -13920 34708 -13840 34720
rect -13920 34652 -13908 34708
rect -13852 34652 -13840 34708
rect -13920 34388 -13840 34652
rect -13920 34332 -13908 34388
rect -13852 34332 -13840 34388
rect -13920 34320 -13840 34332
rect -13760 34708 -13680 34720
rect -13760 34652 -13748 34708
rect -13692 34652 -13680 34708
rect -13760 34388 -13680 34652
rect -13760 34332 -13748 34388
rect -13692 34332 -13680 34388
rect -13760 34320 -13680 34332
rect -13600 34708 -13520 34720
rect -13600 34652 -13588 34708
rect -13532 34652 -13520 34708
rect -13600 34388 -13520 34652
rect -13600 34332 -13588 34388
rect -13532 34332 -13520 34388
rect -13600 34320 -13520 34332
rect -13440 34708 -13360 34720
rect -13440 34652 -13428 34708
rect -13372 34652 -13360 34708
rect -13440 34388 -13360 34652
rect -13440 34332 -13428 34388
rect -13372 34332 -13360 34388
rect -13440 34320 -13360 34332
rect -13280 34708 -13200 34720
rect -13280 34652 -13268 34708
rect -13212 34652 -13200 34708
rect -13280 34388 -13200 34652
rect -13280 34332 -13268 34388
rect -13212 34332 -13200 34388
rect -13280 34320 -13200 34332
rect -13120 34708 -13040 34720
rect -13120 34652 -13108 34708
rect -13052 34652 -13040 34708
rect -13120 34388 -13040 34652
rect -13120 34332 -13108 34388
rect -13052 34332 -13040 34388
rect -13120 34320 -13040 34332
rect -12960 34708 -12880 34720
rect -12960 34652 -12948 34708
rect -12892 34652 -12880 34708
rect -12960 34388 -12880 34652
rect -12960 34332 -12948 34388
rect -12892 34332 -12880 34388
rect -12960 34320 -12880 34332
rect -12800 34708 -12720 34720
rect -12800 34652 -12788 34708
rect -12732 34652 -12720 34708
rect -12800 34388 -12720 34652
rect -12800 34332 -12788 34388
rect -12732 34332 -12720 34388
rect -12800 34320 -12720 34332
rect -12640 34708 -12560 34720
rect -12640 34652 -12628 34708
rect -12572 34652 -12560 34708
rect -12640 34388 -12560 34652
rect -12640 34332 -12628 34388
rect -12572 34332 -12560 34388
rect -12640 34320 -12560 34332
rect -12480 34708 -12400 34720
rect -12480 34652 -12468 34708
rect -12412 34652 -12400 34708
rect -12480 34388 -12400 34652
rect -12480 34332 -12468 34388
rect -12412 34332 -12400 34388
rect -12480 34320 -12400 34332
rect -12320 34708 -12240 34720
rect -12320 34652 -12308 34708
rect -12252 34652 -12240 34708
rect -12320 34388 -12240 34652
rect -12320 34332 -12308 34388
rect -12252 34332 -12240 34388
rect -12320 34320 -12240 34332
rect -12160 34708 -12080 34880
rect -12160 34652 -12148 34708
rect -12092 34652 -12080 34708
rect -12160 34388 -12080 34652
rect -12160 34332 -12148 34388
rect -12092 34332 -12080 34388
rect -12160 34320 -12080 34332
rect -12000 34708 -11920 34720
rect -12000 34652 -11988 34708
rect -11932 34652 -11920 34708
rect -12000 34388 -11920 34652
rect -12000 34332 -11988 34388
rect -11932 34332 -11920 34388
rect -12000 34320 -11920 34332
rect -11840 34708 -11760 34880
rect -11840 34652 -11828 34708
rect -11772 34652 -11760 34708
rect -11840 34388 -11760 34652
rect -11840 34332 -11828 34388
rect -11772 34332 -11760 34388
rect -11840 34320 -11760 34332
rect -11680 34708 -11600 34720
rect -11680 34652 -11668 34708
rect -11612 34652 -11600 34708
rect -11680 34388 -11600 34652
rect -11680 34332 -11668 34388
rect -11612 34332 -11600 34388
rect -11680 34320 -11600 34332
rect -11520 34708 -11440 34880
rect -11520 34652 -11508 34708
rect -11452 34652 -11440 34708
rect -11520 34388 -11440 34652
rect -11520 34332 -11508 34388
rect -11452 34332 -11440 34388
rect -11520 34320 -11440 34332
rect -30080 34168 -30072 34232
rect -30008 34168 -30000 34232
rect -30080 34072 -30000 34168
rect -30080 34008 -30072 34072
rect -30008 34008 -30000 34072
rect -30080 33912 -30000 34008
rect -30080 33848 -30072 33912
rect -30008 33848 -30000 33912
rect -30080 33752 -30000 33848
rect -30080 33688 -30072 33752
rect -30008 33688 -30000 33752
rect -30080 33592 -30000 33688
rect -30080 33528 -30072 33592
rect -30008 33528 -30000 33592
rect -30080 33432 -30000 33528
rect -30080 33368 -30072 33432
rect -30008 33368 -30000 33432
rect -30080 33272 -30000 33368
rect -30080 33208 -30072 33272
rect -30008 33208 -30000 33272
rect -30080 33112 -30000 33208
rect -30080 33048 -30072 33112
rect -30008 33048 -30000 33112
rect -30080 32952 -30000 33048
rect -30080 32888 -30072 32952
rect -30008 32888 -30000 32952
rect -30400 32572 -30388 32628
rect -30332 32572 -30320 32628
rect -30400 32308 -30320 32572
rect -30080 32628 -30000 32888
rect -30080 32572 -30068 32628
rect -30012 32572 -30000 32628
rect -30400 32252 -30388 32308
rect -30332 32252 -30320 32308
rect -30720 32092 -30708 32148
rect -30652 32092 -30640 32148
rect -30720 31988 -30640 32092
rect -30720 31932 -30708 31988
rect -30652 31932 -30640 31988
rect -30720 31840 -30640 31932
rect -30560 32148 -30480 32160
rect -30560 32092 -30548 32148
rect -30492 32092 -30480 32148
rect -30560 31840 -30480 32092
rect -30400 31988 -30320 32252
rect -30400 31932 -30388 31988
rect -30332 31932 -30320 31988
rect -30400 31840 -30320 31932
rect -30240 32468 -30160 32480
rect -30240 32412 -30228 32468
rect -30172 32412 -30160 32468
rect -30240 31840 -30160 32412
rect -30080 32308 -30000 32572
rect -30080 32252 -30068 32308
rect -30012 32252 -30000 32308
rect -30080 31988 -30000 32252
rect -30080 31932 -30068 31988
rect -30012 31932 -30000 31988
rect -30080 31840 -30000 31932
rect -29920 32948 -29840 32960
rect -29920 32892 -29908 32948
rect -29852 32892 -29840 32948
rect -29920 32628 -29840 32892
rect -29920 32572 -29908 32628
rect -29852 32572 -29840 32628
rect -29920 32308 -29840 32572
rect -29920 32252 -29908 32308
rect -29852 32252 -29840 32308
rect -29920 31988 -29840 32252
rect -29920 31932 -29908 31988
rect -29852 31932 -29840 31988
rect -29920 31920 -29840 31932
rect -29760 32948 -29680 32960
rect -29760 32892 -29748 32948
rect -29692 32892 -29680 32948
rect -29760 32628 -29680 32892
rect -29760 32572 -29748 32628
rect -29692 32572 -29680 32628
rect -29760 32308 -29680 32572
rect -29760 32252 -29748 32308
rect -29692 32252 -29680 32308
rect -29760 31988 -29680 32252
rect -29760 31932 -29748 31988
rect -29692 31932 -29680 31988
rect -29760 31920 -29680 31932
rect -29600 32948 -29520 32960
rect -29600 32892 -29588 32948
rect -29532 32892 -29520 32948
rect -29600 32628 -29520 32892
rect -29600 32572 -29588 32628
rect -29532 32572 -29520 32628
rect -29600 32308 -29520 32572
rect -29600 32252 -29588 32308
rect -29532 32252 -29520 32308
rect -29600 31988 -29520 32252
rect -29600 31932 -29588 31988
rect -29532 31932 -29520 31988
rect -29600 31920 -29520 31932
rect -29440 32948 -29360 32960
rect -29440 32892 -29428 32948
rect -29372 32892 -29360 32948
rect -29440 32628 -29360 32892
rect -29440 32572 -29428 32628
rect -29372 32572 -29360 32628
rect -29440 32308 -29360 32572
rect -29440 32252 -29428 32308
rect -29372 32252 -29360 32308
rect -29440 31988 -29360 32252
rect -29440 31932 -29428 31988
rect -29372 31932 -29360 31988
rect -29440 31920 -29360 31932
rect -29280 32948 -29200 32960
rect -29280 32892 -29268 32948
rect -29212 32892 -29200 32948
rect -29280 32628 -29200 32892
rect -29280 32572 -29268 32628
rect -29212 32572 -29200 32628
rect -29280 32308 -29200 32572
rect -29280 32252 -29268 32308
rect -29212 32252 -29200 32308
rect -29280 31988 -29200 32252
rect -29280 31932 -29268 31988
rect -29212 31932 -29200 31988
rect -29280 31920 -29200 31932
rect -29120 32948 -29040 32960
rect -29120 32892 -29108 32948
rect -29052 32892 -29040 32948
rect -29120 32628 -29040 32892
rect -29120 32572 -29108 32628
rect -29052 32572 -29040 32628
rect -29120 32308 -29040 32572
rect -29120 32252 -29108 32308
rect -29052 32252 -29040 32308
rect -29120 31988 -29040 32252
rect -29120 31932 -29108 31988
rect -29052 31932 -29040 31988
rect -29120 31920 -29040 31932
rect -28960 32948 -28880 32960
rect -28960 32892 -28948 32948
rect -28892 32892 -28880 32948
rect -28960 32628 -28880 32892
rect -28960 32572 -28948 32628
rect -28892 32572 -28880 32628
rect -28960 32308 -28880 32572
rect -28960 32252 -28948 32308
rect -28892 32252 -28880 32308
rect -28960 31988 -28880 32252
rect -28960 31932 -28948 31988
rect -28892 31932 -28880 31988
rect -28960 31920 -28880 31932
rect -28800 32948 -28720 32960
rect -28800 32892 -28788 32948
rect -28732 32892 -28720 32948
rect -28800 32628 -28720 32892
rect -28800 32572 -28788 32628
rect -28732 32572 -28720 32628
rect -28800 32308 -28720 32572
rect -28800 32252 -28788 32308
rect -28732 32252 -28720 32308
rect -28800 31988 -28720 32252
rect -28800 31932 -28788 31988
rect -28732 31932 -28720 31988
rect -28800 31920 -28720 31932
rect -28640 32948 -28560 32960
rect -28640 32892 -28628 32948
rect -28572 32892 -28560 32948
rect -28640 32628 -28560 32892
rect -28640 32572 -28628 32628
rect -28572 32572 -28560 32628
rect -28640 32308 -28560 32572
rect -28640 32252 -28628 32308
rect -28572 32252 -28560 32308
rect -28640 31988 -28560 32252
rect -28640 31932 -28628 31988
rect -28572 31932 -28560 31988
rect -28640 31920 -28560 31932
rect -28480 32948 -28400 32960
rect -28480 32892 -28468 32948
rect -28412 32892 -28400 32948
rect -28480 32628 -28400 32892
rect -28480 32572 -28468 32628
rect -28412 32572 -28400 32628
rect -28480 32308 -28400 32572
rect -28480 32252 -28468 32308
rect -28412 32252 -28400 32308
rect -28480 31988 -28400 32252
rect -28480 31932 -28468 31988
rect -28412 31932 -28400 31988
rect -28480 31920 -28400 31932
rect -28320 32948 -28240 32960
rect -28320 32892 -28308 32948
rect -28252 32892 -28240 32948
rect -28320 32628 -28240 32892
rect -28320 32572 -28308 32628
rect -28252 32572 -28240 32628
rect -28320 32308 -28240 32572
rect -28320 32252 -28308 32308
rect -28252 32252 -28240 32308
rect -28320 31988 -28240 32252
rect -28320 31932 -28308 31988
rect -28252 31932 -28240 31988
rect -28320 31920 -28240 31932
rect -28160 32948 -28080 32960
rect -28160 32892 -28148 32948
rect -28092 32892 -28080 32948
rect -28160 32628 -28080 32892
rect -28160 32572 -28148 32628
rect -28092 32572 -28080 32628
rect -28160 32308 -28080 32572
rect -28160 32252 -28148 32308
rect -28092 32252 -28080 32308
rect -28160 31988 -28080 32252
rect -28160 31932 -28148 31988
rect -28092 31932 -28080 31988
rect -28160 31920 -28080 31932
rect -28000 32948 -27920 32960
rect -28000 32892 -27988 32948
rect -27932 32892 -27920 32948
rect -28000 32628 -27920 32892
rect -28000 32572 -27988 32628
rect -27932 32572 -27920 32628
rect -28000 32308 -27920 32572
rect -28000 32252 -27988 32308
rect -27932 32252 -27920 32308
rect -28000 31988 -27920 32252
rect -28000 31932 -27988 31988
rect -27932 31932 -27920 31988
rect -28000 31920 -27920 31932
rect -27840 32948 -27760 32960
rect -27840 32892 -27828 32948
rect -27772 32892 -27760 32948
rect -27840 32628 -27760 32892
rect -27840 32572 -27828 32628
rect -27772 32572 -27760 32628
rect -27840 32308 -27760 32572
rect -27840 32252 -27828 32308
rect -27772 32252 -27760 32308
rect -27840 31988 -27760 32252
rect -27840 31932 -27828 31988
rect -27772 31932 -27760 31988
rect -27840 31920 -27760 31932
rect -27680 32948 -27600 32960
rect -27680 32892 -27668 32948
rect -27612 32892 -27600 32948
rect -27680 32628 -27600 32892
rect -27680 32572 -27668 32628
rect -27612 32572 -27600 32628
rect -27680 32308 -27600 32572
rect -27680 32252 -27668 32308
rect -27612 32252 -27600 32308
rect -27680 31988 -27600 32252
rect -27680 31932 -27668 31988
rect -27612 31932 -27600 31988
rect -27680 31920 -27600 31932
rect -27520 32948 -27440 32960
rect -27520 32892 -27508 32948
rect -27452 32892 -27440 32948
rect -27520 32628 -27440 32892
rect -27520 32572 -27508 32628
rect -27452 32572 -27440 32628
rect -27520 32308 -27440 32572
rect -27520 32252 -27508 32308
rect -27452 32252 -27440 32308
rect -27520 31988 -27440 32252
rect -27520 31932 -27508 31988
rect -27452 31932 -27440 31988
rect -27520 31920 -27440 31932
rect -27360 32948 -27280 32960
rect -27360 32892 -27348 32948
rect -27292 32892 -27280 32948
rect -27360 32628 -27280 32892
rect -27360 32572 -27348 32628
rect -27292 32572 -27280 32628
rect -27360 32308 -27280 32572
rect -27360 32252 -27348 32308
rect -27292 32252 -27280 32308
rect -27360 31988 -27280 32252
rect -27360 31932 -27348 31988
rect -27292 31932 -27280 31988
rect -27360 31920 -27280 31932
rect -27200 32948 -27120 32960
rect -27200 32892 -27188 32948
rect -27132 32892 -27120 32948
rect -27200 32628 -27120 32892
rect -27200 32572 -27188 32628
rect -27132 32572 -27120 32628
rect -27200 32308 -27120 32572
rect -27200 32252 -27188 32308
rect -27132 32252 -27120 32308
rect -27200 31988 -27120 32252
rect -27200 31932 -27188 31988
rect -27132 31932 -27120 31988
rect -27200 31920 -27120 31932
rect -27040 32948 -26960 32960
rect -27040 32892 -27028 32948
rect -26972 32892 -26960 32948
rect -27040 32628 -26960 32892
rect -27040 32572 -27028 32628
rect -26972 32572 -26960 32628
rect -27040 32308 -26960 32572
rect -27040 32252 -27028 32308
rect -26972 32252 -26960 32308
rect -27040 31988 -26960 32252
rect -27040 31932 -27028 31988
rect -26972 31932 -26960 31988
rect -27040 31920 -26960 31932
rect -26880 32948 -26800 32960
rect -26880 32892 -26868 32948
rect -26812 32892 -26800 32948
rect -26880 32628 -26800 32892
rect -26880 32572 -26868 32628
rect -26812 32572 -26800 32628
rect -26880 32308 -26800 32572
rect -26880 32252 -26868 32308
rect -26812 32252 -26800 32308
rect -26880 31988 -26800 32252
rect -26880 31932 -26868 31988
rect -26812 31932 -26800 31988
rect -26880 31920 -26800 31932
rect -26720 32948 -26640 32960
rect -26720 32892 -26708 32948
rect -26652 32892 -26640 32948
rect -26720 32628 -26640 32892
rect -26720 32572 -26708 32628
rect -26652 32572 -26640 32628
rect -26720 32308 -26640 32572
rect -26720 32252 -26708 32308
rect -26652 32252 -26640 32308
rect -26720 31988 -26640 32252
rect -26720 31932 -26708 31988
rect -26652 31932 -26640 31988
rect -26720 31920 -26640 31932
rect -26560 32948 -26480 32960
rect -26560 32892 -26548 32948
rect -26492 32892 -26480 32948
rect -26560 32628 -26480 32892
rect -26560 32572 -26548 32628
rect -26492 32572 -26480 32628
rect -26560 32308 -26480 32572
rect -26560 32252 -26548 32308
rect -26492 32252 -26480 32308
rect -26560 31988 -26480 32252
rect -26560 31932 -26548 31988
rect -26492 31932 -26480 31988
rect -26560 31920 -26480 31932
rect -26400 32948 -26320 32960
rect -26400 32892 -26388 32948
rect -26332 32892 -26320 32948
rect -26400 32628 -26320 32892
rect -26400 32572 -26388 32628
rect -26332 32572 -26320 32628
rect -26400 32308 -26320 32572
rect -26400 32252 -26388 32308
rect -26332 32252 -26320 32308
rect -26400 31988 -26320 32252
rect -26400 31932 -26388 31988
rect -26332 31932 -26320 31988
rect -26400 31920 -26320 31932
rect -26240 32948 -26160 32960
rect -26240 32892 -26228 32948
rect -26172 32892 -26160 32948
rect -26240 32628 -26160 32892
rect -26240 32572 -26228 32628
rect -26172 32572 -26160 32628
rect -26240 32308 -26160 32572
rect -26240 32252 -26228 32308
rect -26172 32252 -26160 32308
rect -26240 31988 -26160 32252
rect -26240 31932 -26228 31988
rect -26172 31932 -26160 31988
rect -26240 31920 -26160 31932
rect -26080 32948 -26000 32960
rect -26080 32892 -26068 32948
rect -26012 32892 -26000 32948
rect -26080 32628 -26000 32892
rect -26080 32572 -26068 32628
rect -26012 32572 -26000 32628
rect -26080 32308 -26000 32572
rect -26080 32252 -26068 32308
rect -26012 32252 -26000 32308
rect -26080 31988 -26000 32252
rect -26080 31932 -26068 31988
rect -26012 31932 -26000 31988
rect -26080 31920 -26000 31932
rect -25920 32948 -25840 32960
rect -25920 32892 -25908 32948
rect -25852 32892 -25840 32948
rect -25920 32628 -25840 32892
rect -25920 32572 -25908 32628
rect -25852 32572 -25840 32628
rect -25920 32308 -25840 32572
rect -25920 32252 -25908 32308
rect -25852 32252 -25840 32308
rect -25920 31988 -25840 32252
rect -25920 31932 -25908 31988
rect -25852 31932 -25840 31988
rect -25920 31920 -25840 31932
rect -25760 32948 -25680 32960
rect -25760 32892 -25748 32948
rect -25692 32892 -25680 32948
rect -25760 32628 -25680 32892
rect -25760 32572 -25748 32628
rect -25692 32572 -25680 32628
rect -25760 32308 -25680 32572
rect -25760 32252 -25748 32308
rect -25692 32252 -25680 32308
rect -25760 31988 -25680 32252
rect -25760 31932 -25748 31988
rect -25692 31932 -25680 31988
rect -25760 31920 -25680 31932
rect -25600 32948 -25520 32960
rect -25600 32892 -25588 32948
rect -25532 32892 -25520 32948
rect -25600 32628 -25520 32892
rect -25600 32572 -25588 32628
rect -25532 32572 -25520 32628
rect -25600 32308 -25520 32572
rect -25600 32252 -25588 32308
rect -25532 32252 -25520 32308
rect -25600 31988 -25520 32252
rect -25600 31932 -25588 31988
rect -25532 31932 -25520 31988
rect -25600 31920 -25520 31932
rect -25440 32948 -25360 32960
rect -25440 32892 -25428 32948
rect -25372 32892 -25360 32948
rect -25440 32628 -25360 32892
rect -25440 32572 -25428 32628
rect -25372 32572 -25360 32628
rect -25440 32308 -25360 32572
rect -25440 32252 -25428 32308
rect -25372 32252 -25360 32308
rect -25440 31988 -25360 32252
rect -25440 31932 -25428 31988
rect -25372 31932 -25360 31988
rect -25440 31920 -25360 31932
rect -25280 32948 -25200 32960
rect -25280 32892 -25268 32948
rect -25212 32892 -25200 32948
rect -25280 32628 -25200 32892
rect -25280 32572 -25268 32628
rect -25212 32572 -25200 32628
rect -25280 32308 -25200 32572
rect -25280 32252 -25268 32308
rect -25212 32252 -25200 32308
rect -25280 31988 -25200 32252
rect -25280 31932 -25268 31988
rect -25212 31932 -25200 31988
rect -25280 31920 -25200 31932
rect -25120 32948 -25040 32960
rect -25120 32892 -25108 32948
rect -25052 32892 -25040 32948
rect -25120 32628 -25040 32892
rect -25120 32572 -25108 32628
rect -25052 32572 -25040 32628
rect -25120 32308 -25040 32572
rect -25120 32252 -25108 32308
rect -25052 32252 -25040 32308
rect -25120 31988 -25040 32252
rect -25120 31932 -25108 31988
rect -25052 31932 -25040 31988
rect -25120 31920 -25040 31932
rect -24960 32948 -24880 32960
rect -24960 32892 -24948 32948
rect -24892 32892 -24880 32948
rect -24960 32628 -24880 32892
rect -24960 32572 -24948 32628
rect -24892 32572 -24880 32628
rect -24960 32308 -24880 32572
rect -24960 32252 -24948 32308
rect -24892 32252 -24880 32308
rect -24960 31988 -24880 32252
rect -24960 31932 -24948 31988
rect -24892 31932 -24880 31988
rect -24960 31920 -24880 31932
rect -24800 32948 -24720 32960
rect -24800 32892 -24788 32948
rect -24732 32892 -24720 32948
rect -24800 32628 -24720 32892
rect -24800 32572 -24788 32628
rect -24732 32572 -24720 32628
rect -24800 32308 -24720 32572
rect -24800 32252 -24788 32308
rect -24732 32252 -24720 32308
rect -24800 31988 -24720 32252
rect -24800 31932 -24788 31988
rect -24732 31932 -24720 31988
rect -24800 31920 -24720 31932
rect -24640 32948 -24560 32960
rect -24640 32892 -24628 32948
rect -24572 32892 -24560 32948
rect -24640 32628 -24560 32892
rect -24640 32572 -24628 32628
rect -24572 32572 -24560 32628
rect -24640 32308 -24560 32572
rect -24640 32252 -24628 32308
rect -24572 32252 -24560 32308
rect -24640 31988 -24560 32252
rect -24640 31932 -24628 31988
rect -24572 31932 -24560 31988
rect -24640 31920 -24560 31932
rect -24480 32948 -24400 32960
rect -24480 32892 -24468 32948
rect -24412 32892 -24400 32948
rect -24480 32628 -24400 32892
rect -24480 32572 -24468 32628
rect -24412 32572 -24400 32628
rect -24480 32308 -24400 32572
rect -24480 32252 -24468 32308
rect -24412 32252 -24400 32308
rect -24480 31988 -24400 32252
rect -24480 31932 -24468 31988
rect -24412 31932 -24400 31988
rect -24480 31920 -24400 31932
rect -24320 32948 -24240 32960
rect -24320 32892 -24308 32948
rect -24252 32892 -24240 32948
rect -24320 32628 -24240 32892
rect -24320 32572 -24308 32628
rect -24252 32572 -24240 32628
rect -24320 32308 -24240 32572
rect -24320 32252 -24308 32308
rect -24252 32252 -24240 32308
rect -24320 31988 -24240 32252
rect -24320 31932 -24308 31988
rect -24252 31932 -24240 31988
rect -24320 31920 -24240 31932
rect -24160 32948 -24080 32960
rect -24160 32892 -24148 32948
rect -24092 32892 -24080 32948
rect -24160 32628 -24080 32892
rect -24160 32572 -24148 32628
rect -24092 32572 -24080 32628
rect -24160 32308 -24080 32572
rect -24160 32252 -24148 32308
rect -24092 32252 -24080 32308
rect -24160 31988 -24080 32252
rect -24160 31932 -24148 31988
rect -24092 31932 -24080 31988
rect -24160 31920 -24080 31932
rect -24000 32948 -23920 32960
rect -24000 32892 -23988 32948
rect -23932 32892 -23920 32948
rect -24000 32628 -23920 32892
rect -24000 32572 -23988 32628
rect -23932 32572 -23920 32628
rect -24000 32308 -23920 32572
rect -24000 32252 -23988 32308
rect -23932 32252 -23920 32308
rect -24000 31988 -23920 32252
rect -24000 31932 -23988 31988
rect -23932 31932 -23920 31988
rect -24000 31920 -23920 31932
rect -23840 32948 -23760 32960
rect -23840 32892 -23828 32948
rect -23772 32892 -23760 32948
rect -23840 32628 -23760 32892
rect -23840 32572 -23828 32628
rect -23772 32572 -23760 32628
rect -23840 32308 -23760 32572
rect -23840 32252 -23828 32308
rect -23772 32252 -23760 32308
rect -23840 31988 -23760 32252
rect -23840 31932 -23828 31988
rect -23772 31932 -23760 31988
rect -23840 31920 -23760 31932
rect -23680 32948 -23600 32960
rect -23680 32892 -23668 32948
rect -23612 32892 -23600 32948
rect -23680 32628 -23600 32892
rect -23680 32572 -23668 32628
rect -23612 32572 -23600 32628
rect -23680 32308 -23600 32572
rect -23680 32252 -23668 32308
rect -23612 32252 -23600 32308
rect -23680 31988 -23600 32252
rect -23680 31932 -23668 31988
rect -23612 31932 -23600 31988
rect -23680 31920 -23600 31932
rect -23520 32948 -23440 32960
rect -23520 32892 -23508 32948
rect -23452 32892 -23440 32948
rect -23520 32628 -23440 32892
rect -23520 32572 -23508 32628
rect -23452 32572 -23440 32628
rect -23520 32308 -23440 32572
rect -23520 32252 -23508 32308
rect -23452 32252 -23440 32308
rect -23520 31988 -23440 32252
rect -23520 31932 -23508 31988
rect -23452 31932 -23440 31988
rect -23520 31920 -23440 31932
rect -23360 32948 -23280 32960
rect -23360 32892 -23348 32948
rect -23292 32892 -23280 32948
rect -23360 32628 -23280 32892
rect -23360 32572 -23348 32628
rect -23292 32572 -23280 32628
rect -23360 32308 -23280 32572
rect -23360 32252 -23348 32308
rect -23292 32252 -23280 32308
rect -23360 31988 -23280 32252
rect -23360 31932 -23348 31988
rect -23292 31932 -23280 31988
rect -23360 31920 -23280 31932
rect -23200 32948 -23120 32960
rect -23200 32892 -23188 32948
rect -23132 32892 -23120 32948
rect -23200 32628 -23120 32892
rect -23200 32572 -23188 32628
rect -23132 32572 -23120 32628
rect -23200 32308 -23120 32572
rect -23200 32252 -23188 32308
rect -23132 32252 -23120 32308
rect -23200 31988 -23120 32252
rect -23200 31932 -23188 31988
rect -23132 31932 -23120 31988
rect -23200 31920 -23120 31932
rect -23040 32948 -22960 32960
rect -23040 32892 -23028 32948
rect -22972 32892 -22960 32948
rect -23040 32628 -22960 32892
rect -23040 32572 -23028 32628
rect -22972 32572 -22960 32628
rect -23040 32308 -22960 32572
rect -23040 32252 -23028 32308
rect -22972 32252 -22960 32308
rect -23040 31988 -22960 32252
rect -23040 31932 -23028 31988
rect -22972 31932 -22960 31988
rect -23040 31920 -22960 31932
rect -22880 32948 -22800 32960
rect -22880 32892 -22868 32948
rect -22812 32892 -22800 32948
rect -22880 32628 -22800 32892
rect -22880 32572 -22868 32628
rect -22812 32572 -22800 32628
rect -22880 32308 -22800 32572
rect -22880 32252 -22868 32308
rect -22812 32252 -22800 32308
rect -22880 31988 -22800 32252
rect -22880 31932 -22868 31988
rect -22812 31932 -22800 31988
rect -22880 31920 -22800 31932
rect -22720 32948 -22640 32960
rect -22720 32892 -22708 32948
rect -22652 32892 -22640 32948
rect -22720 32628 -22640 32892
rect -22720 32572 -22708 32628
rect -22652 32572 -22640 32628
rect -22720 32308 -22640 32572
rect -22720 32252 -22708 32308
rect -22652 32252 -22640 32308
rect -22720 31988 -22640 32252
rect -22720 31932 -22708 31988
rect -22652 31932 -22640 31988
rect -22720 31920 -22640 31932
rect -22560 32948 -22480 32960
rect -22560 32892 -22548 32948
rect -22492 32892 -22480 32948
rect -22560 32628 -22480 32892
rect -22560 32572 -22548 32628
rect -22492 32572 -22480 32628
rect -22560 32308 -22480 32572
rect -22560 32252 -22548 32308
rect -22492 32252 -22480 32308
rect -22560 31988 -22480 32252
rect -22560 31932 -22548 31988
rect -22492 31932 -22480 31988
rect -22560 31920 -22480 31932
rect -22400 32948 -22320 32960
rect -22400 32892 -22388 32948
rect -22332 32892 -22320 32948
rect -22400 32628 -22320 32892
rect -22400 32572 -22388 32628
rect -22332 32572 -22320 32628
rect -22400 32308 -22320 32572
rect -22400 32252 -22388 32308
rect -22332 32252 -22320 32308
rect -22400 31988 -22320 32252
rect -22400 31932 -22388 31988
rect -22332 31932 -22320 31988
rect -22400 31920 -22320 31932
rect -22240 32948 -22160 32960
rect -22240 32892 -22228 32948
rect -22172 32892 -22160 32948
rect -22240 32628 -22160 32892
rect -22240 32572 -22228 32628
rect -22172 32572 -22160 32628
rect -22240 32308 -22160 32572
rect -22240 32252 -22228 32308
rect -22172 32252 -22160 32308
rect -22240 31988 -22160 32252
rect -22240 31932 -22228 31988
rect -22172 31932 -22160 31988
rect -22240 31920 -22160 31932
rect -22080 32948 -22000 32960
rect -22080 32892 -22068 32948
rect -22012 32892 -22000 32948
rect -22080 32628 -22000 32892
rect -22080 32572 -22068 32628
rect -22012 32572 -22000 32628
rect -22080 32308 -22000 32572
rect -22080 32252 -22068 32308
rect -22012 32252 -22000 32308
rect -22080 31988 -22000 32252
rect -22080 31932 -22068 31988
rect -22012 31932 -22000 31988
rect -22080 31920 -22000 31932
rect -21920 32948 -21840 32960
rect -21920 32892 -21908 32948
rect -21852 32892 -21840 32948
rect -21920 32628 -21840 32892
rect -21920 32572 -21908 32628
rect -21852 32572 -21840 32628
rect -21920 32308 -21840 32572
rect -21920 32252 -21908 32308
rect -21852 32252 -21840 32308
rect -21920 31988 -21840 32252
rect -21920 31932 -21908 31988
rect -21852 31932 -21840 31988
rect -21920 31920 -21840 31932
rect -21760 32948 -21680 32960
rect -21760 32892 -21748 32948
rect -21692 32892 -21680 32948
rect -21760 32628 -21680 32892
rect -21760 32572 -21748 32628
rect -21692 32572 -21680 32628
rect -21760 32308 -21680 32572
rect -21760 32252 -21748 32308
rect -21692 32252 -21680 32308
rect -21760 31988 -21680 32252
rect -21760 31932 -21748 31988
rect -21692 31932 -21680 31988
rect -21760 31920 -21680 31932
rect -21600 32948 -21520 32960
rect -21600 32892 -21588 32948
rect -21532 32892 -21520 32948
rect -21600 32628 -21520 32892
rect -21600 32572 -21588 32628
rect -21532 32572 -21520 32628
rect -21600 32308 -21520 32572
rect -21600 32252 -21588 32308
rect -21532 32252 -21520 32308
rect -21600 31988 -21520 32252
rect -21600 31932 -21588 31988
rect -21532 31932 -21520 31988
rect -21600 31920 -21520 31932
rect -21440 32948 -21360 32960
rect -21440 32892 -21428 32948
rect -21372 32892 -21360 32948
rect -21440 32628 -21360 32892
rect -21440 32572 -21428 32628
rect -21372 32572 -21360 32628
rect -21440 32308 -21360 32572
rect -21440 32252 -21428 32308
rect -21372 32252 -21360 32308
rect -21440 31988 -21360 32252
rect -21440 31932 -21428 31988
rect -21372 31932 -21360 31988
rect -21440 31920 -21360 31932
rect -21280 32948 -21200 32960
rect -21280 32892 -21268 32948
rect -21212 32892 -21200 32948
rect -21280 32628 -21200 32892
rect -21280 32572 -21268 32628
rect -21212 32572 -21200 32628
rect -21280 32308 -21200 32572
rect -21280 32252 -21268 32308
rect -21212 32252 -21200 32308
rect -21280 31988 -21200 32252
rect -21280 31932 -21268 31988
rect -21212 31932 -21200 31988
rect -21280 31920 -21200 31932
rect -21120 32948 -21040 32960
rect -21120 32892 -21108 32948
rect -21052 32892 -21040 32948
rect -21120 32628 -21040 32892
rect -21120 32572 -21108 32628
rect -21052 32572 -21040 32628
rect -21120 32308 -21040 32572
rect -21120 32252 -21108 32308
rect -21052 32252 -21040 32308
rect -21120 31988 -21040 32252
rect -21120 31932 -21108 31988
rect -21052 31932 -21040 31988
rect -21120 31920 -21040 31932
rect -20960 32948 -20880 32960
rect -20960 32892 -20948 32948
rect -20892 32892 -20880 32948
rect -20960 32628 -20880 32892
rect -20960 32572 -20948 32628
rect -20892 32572 -20880 32628
rect -20960 32308 -20880 32572
rect -20960 32252 -20948 32308
rect -20892 32252 -20880 32308
rect -20960 31988 -20880 32252
rect -20960 31932 -20948 31988
rect -20892 31932 -20880 31988
rect -20960 31920 -20880 31932
rect -20800 32948 -20720 32960
rect -20800 32892 -20788 32948
rect -20732 32892 -20720 32948
rect -20800 32628 -20720 32892
rect -20800 32572 -20788 32628
rect -20732 32572 -20720 32628
rect -20800 32308 -20720 32572
rect -20800 32252 -20788 32308
rect -20732 32252 -20720 32308
rect -20800 31988 -20720 32252
rect -20800 31932 -20788 31988
rect -20732 31932 -20720 31988
rect -20800 31920 -20720 31932
rect -20640 32948 -20560 32960
rect -20640 32892 -20628 32948
rect -20572 32892 -20560 32948
rect -20640 32628 -20560 32892
rect -20640 32572 -20628 32628
rect -20572 32572 -20560 32628
rect -20640 32308 -20560 32572
rect -20640 32252 -20628 32308
rect -20572 32252 -20560 32308
rect -20640 31988 -20560 32252
rect -20640 31932 -20628 31988
rect -20572 31932 -20560 31988
rect -20640 31920 -20560 31932
rect -20480 32948 -20400 32960
rect -20480 32892 -20468 32948
rect -20412 32892 -20400 32948
rect -20480 32628 -20400 32892
rect -20480 32572 -20468 32628
rect -20412 32572 -20400 32628
rect -20480 32308 -20400 32572
rect -20480 32252 -20468 32308
rect -20412 32252 -20400 32308
rect -20480 31988 -20400 32252
rect -20480 31932 -20468 31988
rect -20412 31932 -20400 31988
rect -20480 31920 -20400 31932
rect -20320 32948 -20240 32960
rect -20320 32892 -20308 32948
rect -20252 32892 -20240 32948
rect -20320 32628 -20240 32892
rect -20320 32572 -20308 32628
rect -20252 32572 -20240 32628
rect -20320 32308 -20240 32572
rect -20320 32252 -20308 32308
rect -20252 32252 -20240 32308
rect -20320 31988 -20240 32252
rect -20320 31932 -20308 31988
rect -20252 31932 -20240 31988
rect -20320 31920 -20240 31932
rect -20160 32948 -20080 32960
rect -20160 32892 -20148 32948
rect -20092 32892 -20080 32948
rect -20160 32628 -20080 32892
rect -20160 32572 -20148 32628
rect -20092 32572 -20080 32628
rect -20160 32308 -20080 32572
rect -20160 32252 -20148 32308
rect -20092 32252 -20080 32308
rect -20160 31988 -20080 32252
rect -20160 31932 -20148 31988
rect -20092 31932 -20080 31988
rect -20160 31920 -20080 31932
rect -20000 32948 -19920 32960
rect -20000 32892 -19988 32948
rect -19932 32892 -19920 32948
rect -20000 32628 -19920 32892
rect -20000 32572 -19988 32628
rect -19932 32572 -19920 32628
rect -20000 32308 -19920 32572
rect -20000 32252 -19988 32308
rect -19932 32252 -19920 32308
rect -20000 31988 -19920 32252
rect -20000 31932 -19988 31988
rect -19932 31932 -19920 31988
rect -20000 31920 -19920 31932
rect -19840 32948 -19760 32960
rect -19840 32892 -19828 32948
rect -19772 32892 -19760 32948
rect -19840 32628 -19760 32892
rect -19840 32572 -19828 32628
rect -19772 32572 -19760 32628
rect -19840 32308 -19760 32572
rect -19840 32252 -19828 32308
rect -19772 32252 -19760 32308
rect -19840 31988 -19760 32252
rect -19840 31932 -19828 31988
rect -19772 31932 -19760 31988
rect -19840 31920 -19760 31932
rect -19680 32948 -19600 32960
rect -19680 32892 -19668 32948
rect -19612 32892 -19600 32948
rect -19680 32628 -19600 32892
rect -19680 32572 -19668 32628
rect -19612 32572 -19600 32628
rect -19680 32308 -19600 32572
rect -19680 32252 -19668 32308
rect -19612 32252 -19600 32308
rect -19680 31988 -19600 32252
rect -19680 31932 -19668 31988
rect -19612 31932 -19600 31988
rect -19680 31920 -19600 31932
rect -19520 32948 -19440 32960
rect -19520 32892 -19508 32948
rect -19452 32892 -19440 32948
rect -19520 32628 -19440 32892
rect -19520 32572 -19508 32628
rect -19452 32572 -19440 32628
rect -19520 32308 -19440 32572
rect -19520 32252 -19508 32308
rect -19452 32252 -19440 32308
rect -19520 31988 -19440 32252
rect -19520 31932 -19508 31988
rect -19452 31932 -19440 31988
rect -19520 31920 -19440 31932
rect -19360 32948 -19280 32960
rect -19360 32892 -19348 32948
rect -19292 32892 -19280 32948
rect -19360 32628 -19280 32892
rect -19360 32572 -19348 32628
rect -19292 32572 -19280 32628
rect -19360 32308 -19280 32572
rect -19360 32252 -19348 32308
rect -19292 32252 -19280 32308
rect -19360 31988 -19280 32252
rect -19360 31932 -19348 31988
rect -19292 31932 -19280 31988
rect -19360 31920 -19280 31932
rect -19200 32948 -19120 32960
rect -19200 32892 -19188 32948
rect -19132 32892 -19120 32948
rect -19200 32628 -19120 32892
rect -19200 32572 -19188 32628
rect -19132 32572 -19120 32628
rect -19200 32308 -19120 32572
rect -19200 32252 -19188 32308
rect -19132 32252 -19120 32308
rect -19200 31988 -19120 32252
rect -19200 31932 -19188 31988
rect -19132 31932 -19120 31988
rect -19200 31920 -19120 31932
rect -19040 32948 -18960 32960
rect -19040 32892 -19028 32948
rect -18972 32892 -18960 32948
rect -19040 32628 -18960 32892
rect -19040 32572 -19028 32628
rect -18972 32572 -18960 32628
rect -19040 32308 -18960 32572
rect -19040 32252 -19028 32308
rect -18972 32252 -18960 32308
rect -19040 31988 -18960 32252
rect -19040 31932 -19028 31988
rect -18972 31932 -18960 31988
rect -19040 31920 -18960 31932
rect -18880 32948 -18800 32960
rect -18880 32892 -18868 32948
rect -18812 32892 -18800 32948
rect -18880 32628 -18800 32892
rect -18880 32572 -18868 32628
rect -18812 32572 -18800 32628
rect -18880 32308 -18800 32572
rect -18880 32252 -18868 32308
rect -18812 32252 -18800 32308
rect -18880 31988 -18800 32252
rect -18880 31932 -18868 31988
rect -18812 31932 -18800 31988
rect -18880 31920 -18800 31932
rect -18720 32948 -18640 32960
rect -18720 32892 -18708 32948
rect -18652 32892 -18640 32948
rect -18720 32628 -18640 32892
rect -18720 32572 -18708 32628
rect -18652 32572 -18640 32628
rect -18720 32308 -18640 32572
rect -18720 32252 -18708 32308
rect -18652 32252 -18640 32308
rect -18720 31988 -18640 32252
rect -18720 31932 -18708 31988
rect -18652 31932 -18640 31988
rect -18720 31920 -18640 31932
rect -18560 32948 -18480 32960
rect -18560 32892 -18548 32948
rect -18492 32892 -18480 32948
rect -18560 32628 -18480 32892
rect -18560 32572 -18548 32628
rect -18492 32572 -18480 32628
rect -18560 32308 -18480 32572
rect -18560 32252 -18548 32308
rect -18492 32252 -18480 32308
rect -18560 31988 -18480 32252
rect -18560 31932 -18548 31988
rect -18492 31932 -18480 31988
rect -18560 31920 -18480 31932
rect -18400 32948 -18320 32960
rect -18400 32892 -18388 32948
rect -18332 32892 -18320 32948
rect -18400 32628 -18320 32892
rect -18400 32572 -18388 32628
rect -18332 32572 -18320 32628
rect -18400 32308 -18320 32572
rect -18400 32252 -18388 32308
rect -18332 32252 -18320 32308
rect -18400 31988 -18320 32252
rect -18400 31932 -18388 31988
rect -18332 31932 -18320 31988
rect -18400 31920 -18320 31932
rect -18240 32948 -18160 32960
rect -18240 32892 -18228 32948
rect -18172 32892 -18160 32948
rect -18240 32628 -18160 32892
rect -18240 32572 -18228 32628
rect -18172 32572 -18160 32628
rect -18240 32308 -18160 32572
rect -18240 32252 -18228 32308
rect -18172 32252 -18160 32308
rect -18240 31988 -18160 32252
rect -18240 31932 -18228 31988
rect -18172 31932 -18160 31988
rect -18240 31920 -18160 31932
rect -18080 32948 -18000 32960
rect -18080 32892 -18068 32948
rect -18012 32892 -18000 32948
rect -18080 32628 -18000 32892
rect -18080 32572 -18068 32628
rect -18012 32572 -18000 32628
rect -18080 32308 -18000 32572
rect -18080 32252 -18068 32308
rect -18012 32252 -18000 32308
rect -18080 31988 -18000 32252
rect -18080 31932 -18068 31988
rect -18012 31932 -18000 31988
rect -18080 31920 -18000 31932
rect -17920 32948 -17840 32960
rect -17920 32892 -17908 32948
rect -17852 32892 -17840 32948
rect -17920 32628 -17840 32892
rect -17920 32572 -17908 32628
rect -17852 32572 -17840 32628
rect -17920 32308 -17840 32572
rect -17920 32252 -17908 32308
rect -17852 32252 -17840 32308
rect -17920 31988 -17840 32252
rect -17920 31932 -17908 31988
rect -17852 31932 -17840 31988
rect -17920 31920 -17840 31932
rect -17760 32948 -17680 32960
rect -17760 32892 -17748 32948
rect -17692 32892 -17680 32948
rect -17760 32628 -17680 32892
rect -17760 32572 -17748 32628
rect -17692 32572 -17680 32628
rect -17760 32308 -17680 32572
rect -17760 32252 -17748 32308
rect -17692 32252 -17680 32308
rect -17760 31988 -17680 32252
rect -17760 31932 -17748 31988
rect -17692 31932 -17680 31988
rect -17760 31920 -17680 31932
rect -17600 32948 -17520 32960
rect -17600 32892 -17588 32948
rect -17532 32892 -17520 32948
rect -17600 32628 -17520 32892
rect -17600 32572 -17588 32628
rect -17532 32572 -17520 32628
rect -17600 32308 -17520 32572
rect -17600 32252 -17588 32308
rect -17532 32252 -17520 32308
rect -17600 31988 -17520 32252
rect -17600 31932 -17588 31988
rect -17532 31932 -17520 31988
rect -17600 31920 -17520 31932
rect -17440 32948 -17360 32960
rect -17440 32892 -17428 32948
rect -17372 32892 -17360 32948
rect -17440 32628 -17360 32892
rect -17440 32572 -17428 32628
rect -17372 32572 -17360 32628
rect -17440 32308 -17360 32572
rect -17440 32252 -17428 32308
rect -17372 32252 -17360 32308
rect -17440 31988 -17360 32252
rect -17440 31932 -17428 31988
rect -17372 31932 -17360 31988
rect -17440 31920 -17360 31932
rect -17280 32948 -17200 32960
rect -17280 32892 -17268 32948
rect -17212 32892 -17200 32948
rect -17280 32628 -17200 32892
rect -17280 32572 -17268 32628
rect -17212 32572 -17200 32628
rect -17280 32308 -17200 32572
rect -17280 32252 -17268 32308
rect -17212 32252 -17200 32308
rect -17280 31988 -17200 32252
rect -17280 31932 -17268 31988
rect -17212 31932 -17200 31988
rect -17280 31920 -17200 31932
rect -17120 32948 -17040 32960
rect -17120 32892 -17108 32948
rect -17052 32892 -17040 32948
rect -17120 32628 -17040 32892
rect -17120 32572 -17108 32628
rect -17052 32572 -17040 32628
rect -17120 32308 -17040 32572
rect -17120 32252 -17108 32308
rect -17052 32252 -17040 32308
rect -17120 31988 -17040 32252
rect -17120 31932 -17108 31988
rect -17052 31932 -17040 31988
rect -17120 31920 -17040 31932
rect -16960 32948 -16880 32960
rect -16960 32892 -16948 32948
rect -16892 32892 -16880 32948
rect -16960 32628 -16880 32892
rect -16960 32572 -16948 32628
rect -16892 32572 -16880 32628
rect -16960 32308 -16880 32572
rect -16960 32252 -16948 32308
rect -16892 32252 -16880 32308
rect -16960 31988 -16880 32252
rect -16960 31932 -16948 31988
rect -16892 31932 -16880 31988
rect -16960 31920 -16880 31932
rect -16800 32948 -16720 32960
rect -16800 32892 -16788 32948
rect -16732 32892 -16720 32948
rect -16800 32628 -16720 32892
rect -16800 32572 -16788 32628
rect -16732 32572 -16720 32628
rect -16800 32308 -16720 32572
rect -16800 32252 -16788 32308
rect -16732 32252 -16720 32308
rect -16800 31988 -16720 32252
rect -16800 31932 -16788 31988
rect -16732 31932 -16720 31988
rect -16800 31920 -16720 31932
rect -16640 32948 -16560 32960
rect -16640 32892 -16628 32948
rect -16572 32892 -16560 32948
rect -16640 32628 -16560 32892
rect -16640 32572 -16628 32628
rect -16572 32572 -16560 32628
rect -16640 32308 -16560 32572
rect -16640 32252 -16628 32308
rect -16572 32252 -16560 32308
rect -16640 31988 -16560 32252
rect -16640 31932 -16628 31988
rect -16572 31932 -16560 31988
rect -16640 31920 -16560 31932
rect -16480 32948 -16400 32960
rect -16480 32892 -16468 32948
rect -16412 32892 -16400 32948
rect -16480 32628 -16400 32892
rect -16480 32572 -16468 32628
rect -16412 32572 -16400 32628
rect -16480 32308 -16400 32572
rect -16480 32252 -16468 32308
rect -16412 32252 -16400 32308
rect -16480 31988 -16400 32252
rect -16480 31932 -16468 31988
rect -16412 31932 -16400 31988
rect -16480 31920 -16400 31932
rect -16320 32948 -16240 32960
rect -16320 32892 -16308 32948
rect -16252 32892 -16240 32948
rect -16320 32628 -16240 32892
rect -16320 32572 -16308 32628
rect -16252 32572 -16240 32628
rect -16320 32308 -16240 32572
rect -16320 32252 -16308 32308
rect -16252 32252 -16240 32308
rect -16320 31988 -16240 32252
rect -16320 31932 -16308 31988
rect -16252 31932 -16240 31988
rect -16320 31920 -16240 31932
rect -16160 32948 -16080 32960
rect -16160 32892 -16148 32948
rect -16092 32892 -16080 32948
rect -16160 32628 -16080 32892
rect -16160 32572 -16148 32628
rect -16092 32572 -16080 32628
rect -16160 32308 -16080 32572
rect -16160 32252 -16148 32308
rect -16092 32252 -16080 32308
rect -16160 31988 -16080 32252
rect -16160 31932 -16148 31988
rect -16092 31932 -16080 31988
rect -16160 31920 -16080 31932
rect -16000 32948 -15920 32960
rect -16000 32892 -15988 32948
rect -15932 32892 -15920 32948
rect -16000 32628 -15920 32892
rect -16000 32572 -15988 32628
rect -15932 32572 -15920 32628
rect -16000 32308 -15920 32572
rect -16000 32252 -15988 32308
rect -15932 32252 -15920 32308
rect -16000 31988 -15920 32252
rect -16000 31932 -15988 31988
rect -15932 31932 -15920 31988
rect -16000 31920 -15920 31932
rect -15840 32948 -15760 32960
rect -15840 32892 -15828 32948
rect -15772 32892 -15760 32948
rect -15840 32628 -15760 32892
rect -15840 32572 -15828 32628
rect -15772 32572 -15760 32628
rect -15840 32308 -15760 32572
rect -15840 32252 -15828 32308
rect -15772 32252 -15760 32308
rect -15840 31988 -15760 32252
rect -15840 31932 -15828 31988
rect -15772 31932 -15760 31988
rect -15840 31920 -15760 31932
rect -15680 32948 -15600 32960
rect -15680 32892 -15668 32948
rect -15612 32892 -15600 32948
rect -15680 32628 -15600 32892
rect -15680 32572 -15668 32628
rect -15612 32572 -15600 32628
rect -15680 32308 -15600 32572
rect -15680 32252 -15668 32308
rect -15612 32252 -15600 32308
rect -15680 31988 -15600 32252
rect -15680 31932 -15668 31988
rect -15612 31932 -15600 31988
rect -15680 31920 -15600 31932
rect -15520 32948 -15440 32960
rect -15520 32892 -15508 32948
rect -15452 32892 -15440 32948
rect -15520 32628 -15440 32892
rect -15520 32572 -15508 32628
rect -15452 32572 -15440 32628
rect -15520 32308 -15440 32572
rect -15520 32252 -15508 32308
rect -15452 32252 -15440 32308
rect -15520 31988 -15440 32252
rect -15520 31932 -15508 31988
rect -15452 31932 -15440 31988
rect -15520 31920 -15440 31932
rect -15360 32948 -15280 32960
rect -15360 32892 -15348 32948
rect -15292 32892 -15280 32948
rect -15360 32628 -15280 32892
rect -15360 32572 -15348 32628
rect -15292 32572 -15280 32628
rect -15360 32308 -15280 32572
rect -15360 32252 -15348 32308
rect -15292 32252 -15280 32308
rect -15360 31988 -15280 32252
rect -15360 31932 -15348 31988
rect -15292 31932 -15280 31988
rect -15360 31920 -15280 31932
rect -15200 32948 -15120 32960
rect -15200 32892 -15188 32948
rect -15132 32892 -15120 32948
rect -15200 32628 -15120 32892
rect -15200 32572 -15188 32628
rect -15132 32572 -15120 32628
rect -15200 32308 -15120 32572
rect -15200 32252 -15188 32308
rect -15132 32252 -15120 32308
rect -15200 31988 -15120 32252
rect -15200 31932 -15188 31988
rect -15132 31932 -15120 31988
rect -15200 31920 -15120 31932
rect -15040 32948 -14960 32960
rect -15040 32892 -15028 32948
rect -14972 32892 -14960 32948
rect -15040 32628 -14960 32892
rect -15040 32572 -15028 32628
rect -14972 32572 -14960 32628
rect -15040 32308 -14960 32572
rect -15040 32252 -15028 32308
rect -14972 32252 -14960 32308
rect -15040 31988 -14960 32252
rect -15040 31932 -15028 31988
rect -14972 31932 -14960 31988
rect -15040 31920 -14960 31932
rect -14880 32948 -14800 32960
rect -14880 32892 -14868 32948
rect -14812 32892 -14800 32948
rect -14880 32628 -14800 32892
rect -14880 32572 -14868 32628
rect -14812 32572 -14800 32628
rect -14880 32308 -14800 32572
rect -14880 32252 -14868 32308
rect -14812 32252 -14800 32308
rect -14880 31988 -14800 32252
rect -14880 31932 -14868 31988
rect -14812 31932 -14800 31988
rect -14880 31920 -14800 31932
rect -14720 32948 -14640 32960
rect -14720 32892 -14708 32948
rect -14652 32892 -14640 32948
rect -14720 32628 -14640 32892
rect -14720 32572 -14708 32628
rect -14652 32572 -14640 32628
rect -14720 32308 -14640 32572
rect -14720 32252 -14708 32308
rect -14652 32252 -14640 32308
rect -14720 31988 -14640 32252
rect -14720 31932 -14708 31988
rect -14652 31932 -14640 31988
rect -14720 31920 -14640 31932
rect -14560 32948 -14480 32960
rect -14560 32892 -14548 32948
rect -14492 32892 -14480 32948
rect -14560 32628 -14480 32892
rect -14560 32572 -14548 32628
rect -14492 32572 -14480 32628
rect -14560 32308 -14480 32572
rect -14560 32252 -14548 32308
rect -14492 32252 -14480 32308
rect -14560 31988 -14480 32252
rect -14560 31932 -14548 31988
rect -14492 31932 -14480 31988
rect -14560 31920 -14480 31932
rect -14400 32948 -14320 32960
rect -14400 32892 -14388 32948
rect -14332 32892 -14320 32948
rect -14400 32628 -14320 32892
rect -14400 32572 -14388 32628
rect -14332 32572 -14320 32628
rect -14400 32308 -14320 32572
rect -14400 32252 -14388 32308
rect -14332 32252 -14320 32308
rect -14400 31988 -14320 32252
rect -14400 31932 -14388 31988
rect -14332 31932 -14320 31988
rect -14400 31920 -14320 31932
rect -14240 32948 -14160 32960
rect -14240 32892 -14228 32948
rect -14172 32892 -14160 32948
rect -14240 32628 -14160 32892
rect -14240 32572 -14228 32628
rect -14172 32572 -14160 32628
rect -14240 32308 -14160 32572
rect -14240 32252 -14228 32308
rect -14172 32252 -14160 32308
rect -14240 31988 -14160 32252
rect -14240 31932 -14228 31988
rect -14172 31932 -14160 31988
rect -14240 31920 -14160 31932
rect -14080 32948 -14000 32960
rect -14080 32892 -14068 32948
rect -14012 32892 -14000 32948
rect -14080 32628 -14000 32892
rect -14080 32572 -14068 32628
rect -14012 32572 -14000 32628
rect -14080 32308 -14000 32572
rect -14080 32252 -14068 32308
rect -14012 32252 -14000 32308
rect -14080 31988 -14000 32252
rect -14080 31932 -14068 31988
rect -14012 31932 -14000 31988
rect -14080 31920 -14000 31932
rect -13920 32948 -13840 32960
rect -13920 32892 -13908 32948
rect -13852 32892 -13840 32948
rect -13920 32628 -13840 32892
rect -13920 32572 -13908 32628
rect -13852 32572 -13840 32628
rect -13920 32308 -13840 32572
rect -13920 32252 -13908 32308
rect -13852 32252 -13840 32308
rect -13920 31988 -13840 32252
rect -13920 31932 -13908 31988
rect -13852 31932 -13840 31988
rect -13920 31920 -13840 31932
rect -13760 32948 -13680 32960
rect -13760 32892 -13748 32948
rect -13692 32892 -13680 32948
rect -13760 32628 -13680 32892
rect -13760 32572 -13748 32628
rect -13692 32572 -13680 32628
rect -13760 32308 -13680 32572
rect -13760 32252 -13748 32308
rect -13692 32252 -13680 32308
rect -13760 31988 -13680 32252
rect -13760 31932 -13748 31988
rect -13692 31932 -13680 31988
rect -13760 31920 -13680 31932
rect -13600 32948 -13520 32960
rect -13600 32892 -13588 32948
rect -13532 32892 -13520 32948
rect -13600 32628 -13520 32892
rect -13600 32572 -13588 32628
rect -13532 32572 -13520 32628
rect -13600 32308 -13520 32572
rect -13600 32252 -13588 32308
rect -13532 32252 -13520 32308
rect -13600 31988 -13520 32252
rect -13600 31932 -13588 31988
rect -13532 31932 -13520 31988
rect -13600 31920 -13520 31932
rect -13440 32948 -13360 32960
rect -13440 32892 -13428 32948
rect -13372 32892 -13360 32948
rect -13440 32628 -13360 32892
rect -13440 32572 -13428 32628
rect -13372 32572 -13360 32628
rect -13440 32308 -13360 32572
rect -13440 32252 -13428 32308
rect -13372 32252 -13360 32308
rect -13440 31988 -13360 32252
rect -13440 31932 -13428 31988
rect -13372 31932 -13360 31988
rect -13440 31920 -13360 31932
rect -13280 32948 -13200 32960
rect -13280 32892 -13268 32948
rect -13212 32892 -13200 32948
rect -13280 32628 -13200 32892
rect -13280 32572 -13268 32628
rect -13212 32572 -13200 32628
rect -13280 32308 -13200 32572
rect -13280 32252 -13268 32308
rect -13212 32252 -13200 32308
rect -13280 31988 -13200 32252
rect -13280 31932 -13268 31988
rect -13212 31932 -13200 31988
rect -13280 31920 -13200 31932
rect -13120 32948 -13040 32960
rect -13120 32892 -13108 32948
rect -13052 32892 -13040 32948
rect -13120 32628 -13040 32892
rect -13120 32572 -13108 32628
rect -13052 32572 -13040 32628
rect -13120 32308 -13040 32572
rect -13120 32252 -13108 32308
rect -13052 32252 -13040 32308
rect -13120 31988 -13040 32252
rect -13120 31932 -13108 31988
rect -13052 31932 -13040 31988
rect -13120 31920 -13040 31932
rect -12960 32948 -12880 32960
rect -12960 32892 -12948 32948
rect -12892 32892 -12880 32948
rect -12960 32628 -12880 32892
rect -12960 32572 -12948 32628
rect -12892 32572 -12880 32628
rect -12960 32308 -12880 32572
rect -12960 32252 -12948 32308
rect -12892 32252 -12880 32308
rect -12960 31988 -12880 32252
rect -12960 31932 -12948 31988
rect -12892 31932 -12880 31988
rect -12960 31920 -12880 31932
rect -12800 32948 -12720 32960
rect -12800 32892 -12788 32948
rect -12732 32892 -12720 32948
rect -12800 32628 -12720 32892
rect -12800 32572 -12788 32628
rect -12732 32572 -12720 32628
rect -12800 32308 -12720 32572
rect -12800 32252 -12788 32308
rect -12732 32252 -12720 32308
rect -12800 31988 -12720 32252
rect -12800 31932 -12788 31988
rect -12732 31932 -12720 31988
rect -12800 31920 -12720 31932
rect -12640 32948 -12560 32960
rect -12640 32892 -12628 32948
rect -12572 32892 -12560 32948
rect -12640 32628 -12560 32892
rect -12640 32572 -12628 32628
rect -12572 32572 -12560 32628
rect -12640 32308 -12560 32572
rect -12640 32252 -12628 32308
rect -12572 32252 -12560 32308
rect -12640 31988 -12560 32252
rect -12640 31932 -12628 31988
rect -12572 31932 -12560 31988
rect -12640 31920 -12560 31932
rect -12480 32948 -12400 32960
rect -12480 32892 -12468 32948
rect -12412 32892 -12400 32948
rect -12480 32628 -12400 32892
rect -12480 32572 -12468 32628
rect -12412 32572 -12400 32628
rect -12480 32308 -12400 32572
rect -12480 32252 -12468 32308
rect -12412 32252 -12400 32308
rect -12480 31988 -12400 32252
rect -12480 31932 -12468 31988
rect -12412 31932 -12400 31988
rect -12480 31920 -12400 31932
rect -12320 32948 -12240 32960
rect -12320 32892 -12308 32948
rect -12252 32892 -12240 32948
rect -12320 32628 -12240 32892
rect -12320 32572 -12308 32628
rect -12252 32572 -12240 32628
rect -12320 32308 -12240 32572
rect -12320 32252 -12308 32308
rect -12252 32252 -12240 32308
rect -12320 31988 -12240 32252
rect -12320 31932 -12308 31988
rect -12252 31932 -12240 31988
rect -12320 31920 -12240 31932
rect -12160 32948 -12080 32960
rect -12160 32892 -12148 32948
rect -12092 32892 -12080 32948
rect -12160 32628 -12080 32892
rect -12160 32572 -12148 32628
rect -12092 32572 -12080 32628
rect -12160 32308 -12080 32572
rect -12160 32252 -12148 32308
rect -12092 32252 -12080 32308
rect -12160 31988 -12080 32252
rect -12160 31932 -12148 31988
rect -12092 31932 -12080 31988
rect -12160 31920 -12080 31932
rect -12000 32948 -11920 32960
rect -12000 32892 -11988 32948
rect -11932 32892 -11920 32948
rect -12000 32628 -11920 32892
rect -12000 32572 -11988 32628
rect -11932 32572 -11920 32628
rect -12000 32308 -11920 32572
rect -12000 32252 -11988 32308
rect -11932 32252 -11920 32308
rect -12000 31988 -11920 32252
rect -12000 31932 -11988 31988
rect -11932 31932 -11920 31988
rect -12000 31920 -11920 31932
rect -11840 32948 -11760 32960
rect -11840 32892 -11828 32948
rect -11772 32892 -11760 32948
rect -11840 32628 -11760 32892
rect -11840 32572 -11828 32628
rect -11772 32572 -11760 32628
rect -11840 32308 -11760 32572
rect -11840 32252 -11828 32308
rect -11772 32252 -11760 32308
rect -11840 31988 -11760 32252
rect -11840 31932 -11828 31988
rect -11772 31932 -11760 31988
rect -11840 31920 -11760 31932
rect -11680 32948 -11600 32960
rect -11680 32892 -11668 32948
rect -11612 32892 -11600 32948
rect -11680 32628 -11600 32892
rect -11680 32572 -11668 32628
rect -11612 32572 -11600 32628
rect -11680 32308 -11600 32572
rect -11680 32252 -11668 32308
rect -11612 32252 -11600 32308
rect -11680 31988 -11600 32252
rect -11680 31932 -11668 31988
rect -11612 31932 -11600 31988
rect -11680 31920 -11600 31932
rect -11520 32948 -11440 32960
rect -11520 32892 -11508 32948
rect -11452 32892 -11440 32948
rect -11520 32628 -11440 32892
rect -11520 32572 -11508 32628
rect -11452 32572 -11440 32628
rect -11520 32308 -11440 32572
rect -11360 32468 -11280 34880
rect -11360 32412 -11348 32468
rect -11292 32412 -11280 32468
rect -11360 32400 -11280 32412
rect -11200 34708 -11120 34880
rect -11200 34652 -11188 34708
rect -11132 34652 -11120 34708
rect -11200 34388 -11120 34652
rect -11200 34332 -11188 34388
rect -11132 34332 -11120 34388
rect -11200 32948 -11120 34332
rect -11200 32892 -11188 32948
rect -11132 32892 -11120 32948
rect -11200 32628 -11120 32892
rect -11200 32572 -11188 32628
rect -11132 32572 -11120 32628
rect -11520 32252 -11508 32308
rect -11452 32252 -11440 32308
rect -11520 31988 -11440 32252
rect -11520 31932 -11508 31988
rect -11452 31932 -11440 31988
rect -11520 31920 -11440 31932
rect -11360 32308 -11280 32320
rect -11360 32252 -11348 32308
rect -11292 32252 -11280 32308
rect -11360 31988 -11280 32252
rect -11360 31932 -11348 31988
rect -11292 31932 -11280 31988
rect -11360 31920 -11280 31932
rect -11200 32308 -11120 32572
rect -11200 32252 -11188 32308
rect -11132 32252 -11120 32308
rect -11200 31988 -11120 32252
rect -11040 32148 -10960 34880
rect -10880 34708 -10800 34880
rect -10880 34652 -10868 34708
rect -10812 34652 -10800 34708
rect -10880 34388 -10800 34652
rect -10720 34548 -10640 34880
rect -10720 34492 -10708 34548
rect -10652 34492 -10640 34548
rect -10720 34480 -10640 34492
rect -10560 34708 -10480 34880
rect -10560 34652 -10548 34708
rect -10492 34652 -10480 34708
rect -10880 34332 -10868 34388
rect -10812 34332 -10800 34388
rect -10880 34320 -10800 34332
rect -10560 34388 -10480 34652
rect -10560 34332 -10548 34388
rect -10492 34332 -10480 34388
rect -10560 34320 -10480 34332
rect -3360 34792 -3280 34888
rect -3360 34728 -3352 34792
rect -3288 34728 -3280 34792
rect -3360 34632 -3280 34728
rect -3360 34568 -3352 34632
rect -3288 34568 -3280 34632
rect -3360 34472 -3280 34568
rect -3360 34408 -3352 34472
rect -3288 34408 -3280 34472
rect -3360 34312 -3280 34408
rect -3360 34248 -3352 34312
rect -3288 34248 -3280 34312
rect -3360 34152 -3280 34248
rect -3360 34088 -3352 34152
rect -3288 34088 -3280 34152
rect -3360 33992 -3280 34088
rect -3360 33928 -3352 33992
rect -3288 33928 -3280 33992
rect -3360 33832 -3280 33928
rect -3360 33768 -3352 33832
rect -3288 33768 -3280 33832
rect -3360 33672 -3280 33768
rect -3360 33608 -3352 33672
rect -3288 33608 -3280 33672
rect -3360 33512 -3280 33608
rect -3360 33448 -3352 33512
rect -3288 33448 -3280 33512
rect -3360 33272 -3280 33448
rect -3360 33208 -3352 33272
rect -3288 33208 -3280 33272
rect -3360 33112 -3280 33208
rect -3360 33048 -3352 33112
rect -3288 33048 -3280 33112
rect -11040 32092 -11028 32148
rect -10972 32092 -10960 32148
rect -11040 32080 -10960 32092
rect -10880 32948 -10800 32960
rect -10880 32892 -10868 32948
rect -10812 32892 -10800 32948
rect -10880 32628 -10800 32892
rect -10880 32572 -10868 32628
rect -10812 32572 -10800 32628
rect -10880 32308 -10800 32572
rect -10880 32252 -10868 32308
rect -10812 32252 -10800 32308
rect -11200 31932 -11188 31988
rect -11132 31932 -11120 31988
rect -11200 31920 -11120 31932
rect -10880 31988 -10800 32252
rect -10880 31932 -10868 31988
rect -10812 31932 -10800 31988
rect -10880 31920 -10800 31932
rect -10720 32948 -10640 32960
rect -10720 32892 -10708 32948
rect -10652 32892 -10640 32948
rect -10720 32628 -10640 32892
rect -10720 32572 -10708 32628
rect -10652 32572 -10640 32628
rect -10720 32308 -10640 32572
rect -10720 32252 -10708 32308
rect -10652 32252 -10640 32308
rect -10720 31988 -10640 32252
rect -10720 31932 -10708 31988
rect -10652 31932 -10640 31988
rect -10720 31920 -10640 31932
rect -10560 32948 -10480 32960
rect -10560 32892 -10548 32948
rect -10492 32892 -10480 32948
rect -10560 32628 -10480 32892
rect -10560 32572 -10548 32628
rect -10492 32572 -10480 32628
rect -10560 32308 -10480 32572
rect -10560 32252 -10548 32308
rect -10492 32252 -10480 32308
rect -10560 31988 -10480 32252
rect -10560 31932 -10548 31988
rect -10492 31932 -10480 31988
rect -10560 31920 -10480 31932
rect -10400 32948 -10320 32960
rect -10400 32892 -10388 32948
rect -10332 32892 -10320 32948
rect -10400 32628 -10320 32892
rect -10400 32572 -10388 32628
rect -10332 32572 -10320 32628
rect -10400 32308 -10320 32572
rect -10400 32252 -10388 32308
rect -10332 32252 -10320 32308
rect -10400 31988 -10320 32252
rect -10400 31932 -10388 31988
rect -10332 31932 -10320 31988
rect -10400 31920 -10320 31932
rect -10240 32948 -10160 32960
rect -10240 32892 -10228 32948
rect -10172 32892 -10160 32948
rect -10240 32628 -10160 32892
rect -10240 32572 -10228 32628
rect -10172 32572 -10160 32628
rect -10240 32308 -10160 32572
rect -10240 32252 -10228 32308
rect -10172 32252 -10160 32308
rect -10240 31988 -10160 32252
rect -10240 31932 -10228 31988
rect -10172 31932 -10160 31988
rect -10240 31920 -10160 31932
rect -10080 32948 -10000 32960
rect -10080 32892 -10068 32948
rect -10012 32892 -10000 32948
rect -10080 32628 -10000 32892
rect -10080 32572 -10068 32628
rect -10012 32572 -10000 32628
rect -10080 32308 -10000 32572
rect -10080 32252 -10068 32308
rect -10012 32252 -10000 32308
rect -10080 31988 -10000 32252
rect -10080 31932 -10068 31988
rect -10012 31932 -10000 31988
rect -10080 31920 -10000 31932
rect -9920 32948 -9840 32960
rect -9920 32892 -9908 32948
rect -9852 32892 -9840 32948
rect -9920 32628 -9840 32892
rect -9920 32572 -9908 32628
rect -9852 32572 -9840 32628
rect -9920 32308 -9840 32572
rect -9920 32252 -9908 32308
rect -9852 32252 -9840 32308
rect -9920 31988 -9840 32252
rect -9920 31932 -9908 31988
rect -9852 31932 -9840 31988
rect -9920 31920 -9840 31932
rect -9760 32948 -9680 32960
rect -9760 32892 -9748 32948
rect -9692 32892 -9680 32948
rect -9760 32628 -9680 32892
rect -9760 32572 -9748 32628
rect -9692 32572 -9680 32628
rect -9760 32308 -9680 32572
rect -9760 32252 -9748 32308
rect -9692 32252 -9680 32308
rect -9760 31988 -9680 32252
rect -9760 31932 -9748 31988
rect -9692 31932 -9680 31988
rect -9760 31920 -9680 31932
rect -9600 32948 -9520 32960
rect -9600 32892 -9588 32948
rect -9532 32892 -9520 32948
rect -9600 32628 -9520 32892
rect -9600 32572 -9588 32628
rect -9532 32572 -9520 32628
rect -9600 32308 -9520 32572
rect -9600 32252 -9588 32308
rect -9532 32252 -9520 32308
rect -9600 31988 -9520 32252
rect -9600 31932 -9588 31988
rect -9532 31932 -9520 31988
rect -9600 31920 -9520 31932
rect -9440 32948 -9360 32960
rect -9440 32892 -9428 32948
rect -9372 32892 -9360 32948
rect -9440 32628 -9360 32892
rect -9440 32572 -9428 32628
rect -9372 32572 -9360 32628
rect -9440 32308 -9360 32572
rect -9440 32252 -9428 32308
rect -9372 32252 -9360 32308
rect -9440 31988 -9360 32252
rect -9440 31932 -9428 31988
rect -9372 31932 -9360 31988
rect -9440 31920 -9360 31932
rect -9280 32948 -9200 32960
rect -9280 32892 -9268 32948
rect -9212 32892 -9200 32948
rect -9280 32628 -9200 32892
rect -9280 32572 -9268 32628
rect -9212 32572 -9200 32628
rect -9280 32308 -9200 32572
rect -9280 32252 -9268 32308
rect -9212 32252 -9200 32308
rect -9280 31988 -9200 32252
rect -9280 31932 -9268 31988
rect -9212 31932 -9200 31988
rect -9280 31920 -9200 31932
rect -9120 32948 -9040 32960
rect -9120 32892 -9108 32948
rect -9052 32892 -9040 32948
rect -9120 32628 -9040 32892
rect -9120 32572 -9108 32628
rect -9052 32572 -9040 32628
rect -9120 32308 -9040 32572
rect -9120 32252 -9108 32308
rect -9052 32252 -9040 32308
rect -9120 31988 -9040 32252
rect -9120 31932 -9108 31988
rect -9052 31932 -9040 31988
rect -9120 31920 -9040 31932
rect -8960 32948 -8880 32960
rect -8960 32892 -8948 32948
rect -8892 32892 -8880 32948
rect -8960 32628 -8880 32892
rect -8960 32572 -8948 32628
rect -8892 32572 -8880 32628
rect -8960 32308 -8880 32572
rect -8960 32252 -8948 32308
rect -8892 32252 -8880 32308
rect -8960 31988 -8880 32252
rect -8960 31932 -8948 31988
rect -8892 31932 -8880 31988
rect -8960 31920 -8880 31932
rect -8800 32948 -8720 32960
rect -8800 32892 -8788 32948
rect -8732 32892 -8720 32948
rect -8800 32628 -8720 32892
rect -8800 32572 -8788 32628
rect -8732 32572 -8720 32628
rect -8800 32308 -8720 32572
rect -8800 32252 -8788 32308
rect -8732 32252 -8720 32308
rect -8800 31988 -8720 32252
rect -8800 31932 -8788 31988
rect -8732 31932 -8720 31988
rect -8800 31920 -8720 31932
rect -8640 32948 -8560 32960
rect -8640 32892 -8628 32948
rect -8572 32892 -8560 32948
rect -8640 32628 -8560 32892
rect -8640 32572 -8628 32628
rect -8572 32572 -8560 32628
rect -8640 32308 -8560 32572
rect -8640 32252 -8628 32308
rect -8572 32252 -8560 32308
rect -8640 31988 -8560 32252
rect -8640 31932 -8628 31988
rect -8572 31932 -8560 31988
rect -8640 31920 -8560 31932
rect -8480 32948 -8400 32960
rect -8480 32892 -8468 32948
rect -8412 32892 -8400 32948
rect -8480 32628 -8400 32892
rect -8480 32572 -8468 32628
rect -8412 32572 -8400 32628
rect -8480 32308 -8400 32572
rect -8480 32252 -8468 32308
rect -8412 32252 -8400 32308
rect -8480 31988 -8400 32252
rect -8480 31932 -8468 31988
rect -8412 31932 -8400 31988
rect -8480 31920 -8400 31932
rect -8320 32948 -8240 32960
rect -8320 32892 -8308 32948
rect -8252 32892 -8240 32948
rect -8320 32628 -8240 32892
rect -8320 32572 -8308 32628
rect -8252 32572 -8240 32628
rect -8320 32308 -8240 32572
rect -8320 32252 -8308 32308
rect -8252 32252 -8240 32308
rect -8320 31988 -8240 32252
rect -8320 31932 -8308 31988
rect -8252 31932 -8240 31988
rect -8320 31920 -8240 31932
rect -8160 32948 -8080 32960
rect -8160 32892 -8148 32948
rect -8092 32892 -8080 32948
rect -8160 32628 -8080 32892
rect -8160 32572 -8148 32628
rect -8092 32572 -8080 32628
rect -8160 32308 -8080 32572
rect -8160 32252 -8148 32308
rect -8092 32252 -8080 32308
rect -8160 31988 -8080 32252
rect -8160 31932 -8148 31988
rect -8092 31932 -8080 31988
rect -8160 31920 -8080 31932
rect -8000 32948 -7920 32960
rect -8000 32892 -7988 32948
rect -7932 32892 -7920 32948
rect -8000 32628 -7920 32892
rect -8000 32572 -7988 32628
rect -7932 32572 -7920 32628
rect -8000 32308 -7920 32572
rect -8000 32252 -7988 32308
rect -7932 32252 -7920 32308
rect -8000 31988 -7920 32252
rect -8000 31932 -7988 31988
rect -7932 31932 -7920 31988
rect -8000 31920 -7920 31932
rect -7840 32948 -7760 32960
rect -7840 32892 -7828 32948
rect -7772 32892 -7760 32948
rect -7840 32628 -7760 32892
rect -7840 32572 -7828 32628
rect -7772 32572 -7760 32628
rect -7840 32308 -7760 32572
rect -7840 32252 -7828 32308
rect -7772 32252 -7760 32308
rect -7840 31988 -7760 32252
rect -7840 31932 -7828 31988
rect -7772 31932 -7760 31988
rect -7840 31920 -7760 31932
rect -7680 32948 -7600 32960
rect -7680 32892 -7668 32948
rect -7612 32892 -7600 32948
rect -7680 32628 -7600 32892
rect -7680 32572 -7668 32628
rect -7612 32572 -7600 32628
rect -7680 32308 -7600 32572
rect -7680 32252 -7668 32308
rect -7612 32252 -7600 32308
rect -7680 31988 -7600 32252
rect -7680 31932 -7668 31988
rect -7612 31932 -7600 31988
rect -7680 31920 -7600 31932
rect -7520 32948 -7440 32960
rect -7520 32892 -7508 32948
rect -7452 32892 -7440 32948
rect -7520 32628 -7440 32892
rect -7520 32572 -7508 32628
rect -7452 32572 -7440 32628
rect -7520 32308 -7440 32572
rect -7520 32252 -7508 32308
rect -7452 32252 -7440 32308
rect -7520 31988 -7440 32252
rect -7520 31932 -7508 31988
rect -7452 31932 -7440 31988
rect -7520 31920 -7440 31932
rect -7360 32948 -7280 32960
rect -7360 32892 -7348 32948
rect -7292 32892 -7280 32948
rect -7360 32628 -7280 32892
rect -7360 32572 -7348 32628
rect -7292 32572 -7280 32628
rect -7360 32308 -7280 32572
rect -7360 32252 -7348 32308
rect -7292 32252 -7280 32308
rect -7360 31988 -7280 32252
rect -7360 31932 -7348 31988
rect -7292 31932 -7280 31988
rect -7360 31920 -7280 31932
rect -7200 32948 -7120 32960
rect -7200 32892 -7188 32948
rect -7132 32892 -7120 32948
rect -7200 32628 -7120 32892
rect -7200 32572 -7188 32628
rect -7132 32572 -7120 32628
rect -7200 32308 -7120 32572
rect -7200 32252 -7188 32308
rect -7132 32252 -7120 32308
rect -7200 31988 -7120 32252
rect -7200 31932 -7188 31988
rect -7132 31932 -7120 31988
rect -7200 31920 -7120 31932
rect -7040 32948 -6960 32960
rect -7040 32892 -7028 32948
rect -6972 32892 -6960 32948
rect -7040 32628 -6960 32892
rect -7040 32572 -7028 32628
rect -6972 32572 -6960 32628
rect -7040 32308 -6960 32572
rect -7040 32252 -7028 32308
rect -6972 32252 -6960 32308
rect -7040 31988 -6960 32252
rect -7040 31932 -7028 31988
rect -6972 31932 -6960 31988
rect -7040 31920 -6960 31932
rect -6880 32948 -6800 32960
rect -6880 32892 -6868 32948
rect -6812 32892 -6800 32948
rect -6880 32628 -6800 32892
rect -6880 32572 -6868 32628
rect -6812 32572 -6800 32628
rect -6880 32308 -6800 32572
rect -6880 32252 -6868 32308
rect -6812 32252 -6800 32308
rect -6880 31988 -6800 32252
rect -6880 31932 -6868 31988
rect -6812 31932 -6800 31988
rect -6880 31920 -6800 31932
rect -6720 32948 -6640 32960
rect -6720 32892 -6708 32948
rect -6652 32892 -6640 32948
rect -6720 32628 -6640 32892
rect -6720 32572 -6708 32628
rect -6652 32572 -6640 32628
rect -6720 32308 -6640 32572
rect -6720 32252 -6708 32308
rect -6652 32252 -6640 32308
rect -6720 31988 -6640 32252
rect -6720 31932 -6708 31988
rect -6652 31932 -6640 31988
rect -6720 31920 -6640 31932
rect -6560 32948 -6480 32960
rect -6560 32892 -6548 32948
rect -6492 32892 -6480 32948
rect -6560 32628 -6480 32892
rect -6560 32572 -6548 32628
rect -6492 32572 -6480 32628
rect -6560 32308 -6480 32572
rect -6560 32252 -6548 32308
rect -6492 32252 -6480 32308
rect -6560 31988 -6480 32252
rect -6560 31932 -6548 31988
rect -6492 31932 -6480 31988
rect -6560 31920 -6480 31932
rect -6400 32948 -6320 32960
rect -6400 32892 -6388 32948
rect -6332 32892 -6320 32948
rect -6400 32628 -6320 32892
rect -6400 32572 -6388 32628
rect -6332 32572 -6320 32628
rect -6400 32308 -6320 32572
rect -6400 32252 -6388 32308
rect -6332 32252 -6320 32308
rect -6400 31988 -6320 32252
rect -6400 31932 -6388 31988
rect -6332 31932 -6320 31988
rect -6400 31920 -6320 31932
rect -6240 32948 -6160 32960
rect -6240 32892 -6228 32948
rect -6172 32892 -6160 32948
rect -6240 32628 -6160 32892
rect -6240 32572 -6228 32628
rect -6172 32572 -6160 32628
rect -6240 32308 -6160 32572
rect -6240 32252 -6228 32308
rect -6172 32252 -6160 32308
rect -6240 31988 -6160 32252
rect -6240 31932 -6228 31988
rect -6172 31932 -6160 31988
rect -6240 31920 -6160 31932
rect -6080 32948 -6000 32960
rect -6080 32892 -6068 32948
rect -6012 32892 -6000 32948
rect -6080 32628 -6000 32892
rect -6080 32572 -6068 32628
rect -6012 32572 -6000 32628
rect -6080 32308 -6000 32572
rect -6080 32252 -6068 32308
rect -6012 32252 -6000 32308
rect -6080 31988 -6000 32252
rect -6080 31932 -6068 31988
rect -6012 31932 -6000 31988
rect -6080 31920 -6000 31932
rect -5920 32948 -5840 32960
rect -5920 32892 -5908 32948
rect -5852 32892 -5840 32948
rect -5920 32628 -5840 32892
rect -5920 32572 -5908 32628
rect -5852 32572 -5840 32628
rect -5920 32308 -5840 32572
rect -5920 32252 -5908 32308
rect -5852 32252 -5840 32308
rect -5920 31988 -5840 32252
rect -5920 31932 -5908 31988
rect -5852 31932 -5840 31988
rect -5920 31920 -5840 31932
rect -5760 32948 -5680 32960
rect -5760 32892 -5748 32948
rect -5692 32892 -5680 32948
rect -5760 32628 -5680 32892
rect -5760 32572 -5748 32628
rect -5692 32572 -5680 32628
rect -5760 32308 -5680 32572
rect -5760 32252 -5748 32308
rect -5692 32252 -5680 32308
rect -5760 31988 -5680 32252
rect -5760 31932 -5748 31988
rect -5692 31932 -5680 31988
rect -5760 31920 -5680 31932
rect -5600 32948 -5520 32960
rect -5600 32892 -5588 32948
rect -5532 32892 -5520 32948
rect -5600 32628 -5520 32892
rect -5600 32572 -5588 32628
rect -5532 32572 -5520 32628
rect -5600 32308 -5520 32572
rect -5600 32252 -5588 32308
rect -5532 32252 -5520 32308
rect -5600 31988 -5520 32252
rect -5600 31932 -5588 31988
rect -5532 31932 -5520 31988
rect -5600 31920 -5520 31932
rect -5440 32948 -5360 32960
rect -5440 32892 -5428 32948
rect -5372 32892 -5360 32948
rect -5440 32628 -5360 32892
rect -5440 32572 -5428 32628
rect -5372 32572 -5360 32628
rect -5440 32308 -5360 32572
rect -5440 32252 -5428 32308
rect -5372 32252 -5360 32308
rect -5440 31988 -5360 32252
rect -5440 31932 -5428 31988
rect -5372 31932 -5360 31988
rect -5440 31920 -5360 31932
rect -5280 32948 -5200 32960
rect -5280 32892 -5268 32948
rect -5212 32892 -5200 32948
rect -5280 32628 -5200 32892
rect -5280 32572 -5268 32628
rect -5212 32572 -5200 32628
rect -5280 32308 -5200 32572
rect -5280 32252 -5268 32308
rect -5212 32252 -5200 32308
rect -5280 31988 -5200 32252
rect -5280 31932 -5268 31988
rect -5212 31932 -5200 31988
rect -5280 31920 -5200 31932
rect -5120 32948 -5040 32960
rect -5120 32892 -5108 32948
rect -5052 32892 -5040 32948
rect -5120 32628 -5040 32892
rect -5120 32572 -5108 32628
rect -5052 32572 -5040 32628
rect -5120 32308 -5040 32572
rect -5120 32252 -5108 32308
rect -5052 32252 -5040 32308
rect -5120 31988 -5040 32252
rect -5120 31932 -5108 31988
rect -5052 31932 -5040 31988
rect -5120 31920 -5040 31932
rect -4960 32948 -4880 32960
rect -4960 32892 -4948 32948
rect -4892 32892 -4880 32948
rect -4960 32628 -4880 32892
rect -4960 32572 -4948 32628
rect -4892 32572 -4880 32628
rect -4960 32308 -4880 32572
rect -4960 32252 -4948 32308
rect -4892 32252 -4880 32308
rect -4960 31988 -4880 32252
rect -4960 31932 -4948 31988
rect -4892 31932 -4880 31988
rect -4960 31920 -4880 31932
rect -4800 32948 -4720 32960
rect -4800 32892 -4788 32948
rect -4732 32892 -4720 32948
rect -4800 32628 -4720 32892
rect -4800 32572 -4788 32628
rect -4732 32572 -4720 32628
rect -4800 32308 -4720 32572
rect -4800 32252 -4788 32308
rect -4732 32252 -4720 32308
rect -4800 31988 -4720 32252
rect -4800 31932 -4788 31988
rect -4732 31932 -4720 31988
rect -4800 31920 -4720 31932
rect -4640 32948 -4560 32960
rect -4640 32892 -4628 32948
rect -4572 32892 -4560 32948
rect -4640 32628 -4560 32892
rect -4640 32572 -4628 32628
rect -4572 32572 -4560 32628
rect -4640 32308 -4560 32572
rect -4640 32252 -4628 32308
rect -4572 32252 -4560 32308
rect -4640 31988 -4560 32252
rect -4640 31932 -4628 31988
rect -4572 31932 -4560 31988
rect -4640 31920 -4560 31932
rect -4480 32948 -4400 32960
rect -4480 32892 -4468 32948
rect -4412 32892 -4400 32948
rect -4480 32628 -4400 32892
rect -4480 32572 -4468 32628
rect -4412 32572 -4400 32628
rect -4480 32308 -4400 32572
rect -4480 32252 -4468 32308
rect -4412 32252 -4400 32308
rect -4480 31988 -4400 32252
rect -4480 31932 -4468 31988
rect -4412 31932 -4400 31988
rect -4480 31920 -4400 31932
rect -4320 32948 -4240 32960
rect -4320 32892 -4308 32948
rect -4252 32892 -4240 32948
rect -4320 32628 -4240 32892
rect -4320 32572 -4308 32628
rect -4252 32572 -4240 32628
rect -4320 32308 -4240 32572
rect -4320 32252 -4308 32308
rect -4252 32252 -4240 32308
rect -4320 31988 -4240 32252
rect -4320 31932 -4308 31988
rect -4252 31932 -4240 31988
rect -4320 31920 -4240 31932
rect -4160 32948 -4080 32960
rect -4160 32892 -4148 32948
rect -4092 32892 -4080 32948
rect -4160 32628 -4080 32892
rect -4160 32572 -4148 32628
rect -4092 32572 -4080 32628
rect -4160 32308 -4080 32572
rect -4160 32252 -4148 32308
rect -4092 32252 -4080 32308
rect -4160 31988 -4080 32252
rect -4160 31932 -4148 31988
rect -4092 31932 -4080 31988
rect -4160 31920 -4080 31932
rect -4000 32948 -3920 32960
rect -4000 32892 -3988 32948
rect -3932 32892 -3920 32948
rect -4000 32628 -3920 32892
rect -4000 32572 -3988 32628
rect -3932 32572 -3920 32628
rect -4000 32308 -3920 32572
rect -4000 32252 -3988 32308
rect -3932 32252 -3920 32308
rect -4000 31988 -3920 32252
rect -4000 31932 -3988 31988
rect -3932 31932 -3920 31988
rect -4000 31920 -3920 31932
rect -3680 32948 -3600 32960
rect -3680 32892 -3668 32948
rect -3612 32892 -3600 32948
rect -3680 32628 -3600 32892
rect -3680 32572 -3668 32628
rect -3612 32572 -3600 32628
rect -3680 32308 -3600 32572
rect -3680 32252 -3668 32308
rect -3612 32252 -3600 32308
rect -3680 31988 -3600 32252
rect -3680 31932 -3668 31988
rect -3612 31932 -3600 31988
rect -3680 31920 -3600 31932
rect -3520 32948 -3440 32960
rect -3520 32892 -3508 32948
rect -3452 32892 -3440 32948
rect -3520 32628 -3440 32892
rect -3520 32572 -3508 32628
rect -3452 32572 -3440 32628
rect -3520 32308 -3440 32572
rect -3520 32252 -3508 32308
rect -3452 32252 -3440 32308
rect -3520 31988 -3440 32252
rect -3520 31932 -3508 31988
rect -3452 31932 -3440 31988
rect -3520 31920 -3440 31932
rect -3360 32948 -3280 33048
rect -3040 35752 -2960 36012
rect -3040 35688 -3032 35752
rect -2968 35688 -2960 35752
rect -3040 35592 -2960 35688
rect -3040 35528 -3032 35592
rect -2968 35528 -2960 35592
rect -3040 35432 -2960 35528
rect -3040 35368 -3032 35432
rect -2968 35368 -2960 35432
rect -3040 35272 -2960 35368
rect -3040 35208 -3032 35272
rect -2968 35208 -2960 35272
rect -3040 35112 -2960 35208
rect -3040 35048 -3032 35112
rect -2968 35048 -2960 35112
rect -3040 34952 -2960 35048
rect -3040 34888 -3032 34952
rect -2968 34888 -2960 34952
rect -3040 34792 -2960 34888
rect -3040 34728 -3032 34792
rect -2968 34728 -2960 34792
rect -3040 34632 -2960 34728
rect -3040 34568 -3032 34632
rect -2968 34568 -2960 34632
rect -3040 34472 -2960 34568
rect -3040 34408 -3032 34472
rect -2968 34408 -2960 34472
rect -3040 34312 -2960 34408
rect -3040 34248 -3032 34312
rect -2968 34248 -2960 34312
rect -3040 34152 -2960 34248
rect -3040 34088 -3032 34152
rect -2968 34088 -2960 34152
rect -3040 33992 -2960 34088
rect -3040 33928 -3032 33992
rect -2968 33928 -2960 33992
rect -3040 33832 -2960 33928
rect -3040 33768 -3032 33832
rect -2968 33768 -2960 33832
rect -3040 33672 -2960 33768
rect -3040 33608 -3032 33672
rect -2968 33608 -2960 33672
rect -3040 33512 -2960 33608
rect -3040 33448 -3032 33512
rect -2968 33448 -2960 33512
rect -3040 33272 -2960 33448
rect -3040 33208 -3032 33272
rect -2968 33208 -2960 33272
rect -3040 33112 -2960 33208
rect -3040 33048 -3032 33112
rect -2968 33048 -2960 33112
rect -3360 32892 -3348 32948
rect -3292 32892 -3280 32948
rect -3360 32628 -3280 32892
rect -3360 32572 -3348 32628
rect -3292 32572 -3280 32628
rect -3360 32308 -3280 32572
rect -3360 32252 -3348 32308
rect -3292 32252 -3280 32308
rect -3360 31988 -3280 32252
rect -3360 31932 -3348 31988
rect -3292 31932 -3280 31988
rect -3360 31920 -3280 31932
rect -3200 32948 -3120 32960
rect -3200 32892 -3188 32948
rect -3132 32892 -3120 32948
rect -3200 32628 -3120 32892
rect -3200 32572 -3188 32628
rect -3132 32572 -3120 32628
rect -3200 32308 -3120 32572
rect -3200 32252 -3188 32308
rect -3132 32252 -3120 32308
rect -3200 31988 -3120 32252
rect -3200 31932 -3188 31988
rect -3132 31932 -3120 31988
rect -3200 31920 -3120 31932
rect -3040 32948 -2960 33048
rect -2720 36068 -2640 36328
rect -2720 36012 -2708 36068
rect -2652 36012 -2640 36068
rect -2720 35752 -2640 36012
rect -2720 35688 -2712 35752
rect -2648 35688 -2640 35752
rect -2720 35592 -2640 35688
rect -2720 35528 -2712 35592
rect -2648 35528 -2640 35592
rect -2720 35432 -2640 35528
rect -2720 35368 -2712 35432
rect -2648 35368 -2640 35432
rect -2720 35272 -2640 35368
rect -2720 35208 -2712 35272
rect -2648 35208 -2640 35272
rect -2720 35112 -2640 35208
rect -2720 35048 -2712 35112
rect -2648 35048 -2640 35112
rect -2720 34952 -2640 35048
rect -2720 34888 -2712 34952
rect -2648 34888 -2640 34952
rect -2720 34792 -2640 34888
rect -2720 34728 -2712 34792
rect -2648 34728 -2640 34792
rect -2720 34632 -2640 34728
rect -2720 34568 -2712 34632
rect -2648 34568 -2640 34632
rect -2720 34472 -2640 34568
rect -2720 34408 -2712 34472
rect -2648 34408 -2640 34472
rect -2720 34312 -2640 34408
rect -2720 34248 -2712 34312
rect -2648 34248 -2640 34312
rect -2720 34152 -2640 34248
rect -2720 34088 -2712 34152
rect -2648 34088 -2640 34152
rect -2720 33992 -2640 34088
rect -2720 33928 -2712 33992
rect -2648 33928 -2640 33992
rect -2720 33832 -2640 33928
rect -2720 33768 -2712 33832
rect -2648 33768 -2640 33832
rect -2720 33672 -2640 33768
rect -2720 33608 -2712 33672
rect -2648 33608 -2640 33672
rect -2720 33512 -2640 33608
rect -2720 33448 -2712 33512
rect -2648 33448 -2640 33512
rect -2720 33272 -2640 33448
rect -2720 33208 -2712 33272
rect -2648 33208 -2640 33272
rect -2720 33112 -2640 33208
rect -2720 33048 -2712 33112
rect -2648 33048 -2640 33112
rect -3040 32892 -3028 32948
rect -2972 32892 -2960 32948
rect -3040 32628 -2960 32892
rect -3040 32572 -3028 32628
rect -2972 32572 -2960 32628
rect -3040 32308 -2960 32572
rect -3040 32252 -3028 32308
rect -2972 32252 -2960 32308
rect -3040 31988 -2960 32252
rect -3040 31932 -3028 31988
rect -2972 31932 -2960 31988
rect -3040 31920 -2960 31932
rect -2880 32948 -2800 32960
rect -2880 32892 -2868 32948
rect -2812 32892 -2800 32948
rect -2880 32628 -2800 32892
rect -2880 32572 -2868 32628
rect -2812 32572 -2800 32628
rect -2880 32308 -2800 32572
rect -2880 32252 -2868 32308
rect -2812 32252 -2800 32308
rect -2880 31988 -2800 32252
rect -2880 31932 -2868 31988
rect -2812 31932 -2800 31988
rect -2880 31920 -2800 31932
rect -2720 32948 -2640 33048
rect -2720 32892 -2708 32948
rect -2652 32892 -2640 32948
rect -2720 32628 -2640 32892
rect -2720 32572 -2708 32628
rect -2652 32572 -2640 32628
rect -2720 32308 -2640 32572
rect -2560 40228 -2480 40240
rect -2560 40172 -2548 40228
rect -2492 40172 -2480 40228
rect -2560 32468 -2480 40172
rect -2400 40068 -2320 40332
rect -2400 40012 -2388 40068
rect -2332 40012 -2320 40068
rect -2400 39908 -2320 40012
rect -2080 41748 -2000 41852
rect -2080 41692 -2068 41748
rect -2012 41692 -2000 41748
rect -2080 41588 -2000 41692
rect -2080 41532 -2068 41588
rect -2012 41532 -2000 41588
rect -2080 40868 -2000 41532
rect -2080 40812 -2068 40868
rect -2012 40812 -2000 40868
rect -2080 40708 -2000 40812
rect -2080 40652 -2068 40708
rect -2012 40652 -2000 40708
rect -2080 40388 -2000 40652
rect -2080 40332 -2068 40388
rect -2012 40332 -2000 40388
rect -2080 40068 -2000 40332
rect -1920 40228 -1840 42960
rect -1920 40172 -1908 40228
rect -1852 40172 -1840 40228
rect -1920 40160 -1840 40172
rect -1760 42868 -1680 42960
rect -1760 42812 -1748 42868
rect -1692 42812 -1680 42868
rect -1760 42548 -1680 42812
rect -1760 42492 -1748 42548
rect -1692 42492 -1680 42548
rect -1760 42228 -1680 42492
rect -1760 42172 -1748 42228
rect -1692 42172 -1680 42228
rect -1760 41908 -1680 42172
rect -1760 41852 -1748 41908
rect -1692 41852 -1680 41908
rect -1760 41748 -1680 41852
rect -1760 41692 -1748 41748
rect -1692 41692 -1680 41748
rect -1760 41588 -1680 41692
rect -1760 41532 -1748 41588
rect -1692 41532 -1680 41588
rect -1760 40868 -1680 41532
rect -1760 40812 -1748 40868
rect -1692 40812 -1680 40868
rect -1760 40708 -1680 40812
rect -1760 40652 -1748 40708
rect -1692 40652 -1680 40708
rect -1760 40388 -1680 40652
rect -1760 40332 -1748 40388
rect -1692 40332 -1680 40388
rect -2080 40012 -2068 40068
rect -2012 40012 -2000 40068
rect -2400 39852 -2388 39908
rect -2332 39852 -2320 39908
rect -2400 39752 -2320 39852
rect -2400 39688 -2392 39752
rect -2328 39688 -2320 39752
rect -2400 39592 -2320 39688
rect -2400 39528 -2392 39592
rect -2328 39528 -2320 39592
rect -2400 39432 -2320 39528
rect -2400 39368 -2392 39432
rect -2328 39368 -2320 39432
rect -2400 39272 -2320 39368
rect -2400 39208 -2392 39272
rect -2328 39208 -2320 39272
rect -2400 39112 -2320 39208
rect -2400 39048 -2392 39112
rect -2328 39048 -2320 39112
rect -2400 38952 -2320 39048
rect -2400 38888 -2392 38952
rect -2328 38888 -2320 38952
rect -2400 38792 -2320 38888
rect -2400 38728 -2392 38792
rect -2328 38728 -2320 38792
rect -2400 38632 -2320 38728
rect -2400 38568 -2392 38632
rect -2328 38568 -2320 38632
rect -2400 38472 -2320 38568
rect -2400 38408 -2392 38472
rect -2328 38408 -2320 38472
rect -2400 38312 -2320 38408
rect -2400 38248 -2392 38312
rect -2328 38248 -2320 38312
rect -2400 38152 -2320 38248
rect -2400 38088 -2392 38152
rect -2328 38088 -2320 38152
rect -2400 37992 -2320 38088
rect -2400 37928 -2392 37992
rect -2328 37928 -2320 37992
rect -2400 37832 -2320 37928
rect -2400 37768 -2392 37832
rect -2328 37768 -2320 37832
rect -2400 37668 -2320 37768
rect -2400 37612 -2388 37668
rect -2332 37612 -2320 37668
rect -2400 37512 -2320 37612
rect -2400 37448 -2392 37512
rect -2328 37448 -2320 37512
rect -2400 37352 -2320 37448
rect -2400 37288 -2392 37352
rect -2328 37288 -2320 37352
rect -2400 37192 -2320 37288
rect -2400 37128 -2392 37192
rect -2328 37128 -2320 37192
rect -2400 37032 -2320 37128
rect -2400 36968 -2392 37032
rect -2328 36968 -2320 37032
rect -2400 36872 -2320 36968
rect -2400 36808 -2392 36872
rect -2328 36808 -2320 36872
rect -2400 36712 -2320 36808
rect -2400 36648 -2392 36712
rect -2328 36648 -2320 36712
rect -2400 36552 -2320 36648
rect -2400 36488 -2392 36552
rect -2328 36488 -2320 36552
rect -2400 36392 -2320 36488
rect -2400 36328 -2392 36392
rect -2328 36328 -2320 36392
rect -2400 36068 -2320 36328
rect -2400 36012 -2388 36068
rect -2332 36012 -2320 36068
rect -2400 36000 -2320 36012
rect -2240 39908 -2160 39920
rect -2240 39852 -2228 39908
rect -2172 39852 -2160 39908
rect -2560 32412 -2548 32468
rect -2492 32412 -2480 32468
rect -2560 32400 -2480 32412
rect -2400 35752 -2320 35760
rect -2400 35688 -2392 35752
rect -2328 35688 -2320 35752
rect -2400 35592 -2320 35688
rect -2400 35528 -2392 35592
rect -2328 35528 -2320 35592
rect -2400 35432 -2320 35528
rect -2400 35368 -2392 35432
rect -2328 35368 -2320 35432
rect -2400 35272 -2320 35368
rect -2400 35208 -2392 35272
rect -2328 35208 -2320 35272
rect -2400 35112 -2320 35208
rect -2400 35048 -2392 35112
rect -2328 35048 -2320 35112
rect -2400 34952 -2320 35048
rect -2400 34888 -2392 34952
rect -2328 34888 -2320 34952
rect -2400 34792 -2320 34888
rect -2400 34728 -2392 34792
rect -2328 34728 -2320 34792
rect -2400 34632 -2320 34728
rect -2400 34568 -2392 34632
rect -2328 34568 -2320 34632
rect -2400 34472 -2320 34568
rect -2400 34408 -2392 34472
rect -2328 34408 -2320 34472
rect -2400 34312 -2320 34408
rect -2400 34248 -2392 34312
rect -2328 34248 -2320 34312
rect -2400 34152 -2320 34248
rect -2400 34088 -2392 34152
rect -2328 34088 -2320 34152
rect -2400 33992 -2320 34088
rect -2400 33928 -2392 33992
rect -2328 33928 -2320 33992
rect -2400 33832 -2320 33928
rect -2400 33768 -2392 33832
rect -2328 33768 -2320 33832
rect -2400 33672 -2320 33768
rect -2400 33608 -2392 33672
rect -2328 33608 -2320 33672
rect -2400 33512 -2320 33608
rect -2400 33448 -2392 33512
rect -2328 33448 -2320 33512
rect -2400 33272 -2320 33448
rect -2400 33208 -2392 33272
rect -2328 33208 -2320 33272
rect -2400 33112 -2320 33208
rect -2400 33048 -2392 33112
rect -2328 33048 -2320 33112
rect -2400 32948 -2320 33048
rect -2400 32892 -2388 32948
rect -2332 32892 -2320 32948
rect -2400 32628 -2320 32892
rect -2400 32572 -2388 32628
rect -2332 32572 -2320 32628
rect -2720 32252 -2708 32308
rect -2652 32252 -2640 32308
rect -2720 31988 -2640 32252
rect -2720 31932 -2708 31988
rect -2652 31932 -2640 31988
rect -2720 31920 -2640 31932
rect -2400 32308 -2320 32572
rect -2400 32252 -2388 32308
rect -2332 32252 -2320 32308
rect -2400 31988 -2320 32252
rect -2240 32148 -2160 39852
rect -2240 32092 -2228 32148
rect -2172 32092 -2160 32148
rect -2240 32080 -2160 32092
rect -2080 39752 -2000 40012
rect -2080 39688 -2072 39752
rect -2008 39688 -2000 39752
rect -2080 39592 -2000 39688
rect -2080 39528 -2072 39592
rect -2008 39528 -2000 39592
rect -2080 39432 -2000 39528
rect -2080 39368 -2072 39432
rect -2008 39368 -2000 39432
rect -2080 39272 -2000 39368
rect -2080 39208 -2072 39272
rect -2008 39208 -2000 39272
rect -2080 39112 -2000 39208
rect -2080 39048 -2072 39112
rect -2008 39048 -2000 39112
rect -2080 38952 -2000 39048
rect -2080 38888 -2072 38952
rect -2008 38888 -2000 38952
rect -2080 38792 -2000 38888
rect -2080 38728 -2072 38792
rect -2008 38728 -2000 38792
rect -2080 38632 -2000 38728
rect -2080 38568 -2072 38632
rect -2008 38568 -2000 38632
rect -2080 38472 -2000 38568
rect -2080 38408 -2072 38472
rect -2008 38408 -2000 38472
rect -2080 38312 -2000 38408
rect -2080 38248 -2072 38312
rect -2008 38248 -2000 38312
rect -2080 38152 -2000 38248
rect -2080 38088 -2072 38152
rect -2008 38088 -2000 38152
rect -2080 37992 -2000 38088
rect -2080 37928 -2072 37992
rect -2008 37928 -2000 37992
rect -2080 37832 -2000 37928
rect -2080 37768 -2072 37832
rect -2008 37768 -2000 37832
rect -2080 37668 -2000 37768
rect -2080 37612 -2068 37668
rect -2012 37612 -2000 37668
rect -2080 37512 -2000 37612
rect -2080 37448 -2072 37512
rect -2008 37448 -2000 37512
rect -2080 37352 -2000 37448
rect -2080 37288 -2072 37352
rect -2008 37288 -2000 37352
rect -2080 37192 -2000 37288
rect -2080 37128 -2072 37192
rect -2008 37128 -2000 37192
rect -2080 37032 -2000 37128
rect -2080 36968 -2072 37032
rect -2008 36968 -2000 37032
rect -2080 36872 -2000 36968
rect -2080 36808 -2072 36872
rect -2008 36808 -2000 36872
rect -2080 36712 -2000 36808
rect -2080 36648 -2072 36712
rect -2008 36648 -2000 36712
rect -2080 36552 -2000 36648
rect -2080 36488 -2072 36552
rect -2008 36488 -2000 36552
rect -2080 36392 -2000 36488
rect -2080 36328 -2072 36392
rect -2008 36328 -2000 36392
rect -2080 36068 -2000 36328
rect -1760 40068 -1680 40332
rect -1760 40012 -1748 40068
rect -1692 40012 -1680 40068
rect -1760 39752 -1680 40012
rect -1600 39908 -1520 42960
rect -1600 39852 -1588 39908
rect -1532 39852 -1520 39908
rect -1600 39840 -1520 39852
rect -1440 42868 -1360 42960
rect -1440 42812 -1428 42868
rect -1372 42812 -1360 42868
rect -1440 42548 -1360 42812
rect -1440 42492 -1428 42548
rect -1372 42492 -1360 42548
rect -1440 42228 -1360 42492
rect -1440 42172 -1428 42228
rect -1372 42172 -1360 42228
rect -1440 41908 -1360 42172
rect -1280 42068 -1200 42960
rect -1280 42012 -1268 42068
rect -1212 42012 -1200 42068
rect -1280 42000 -1200 42012
rect -1120 42868 -1040 42960
rect -1120 42812 -1108 42868
rect -1052 42812 -1040 42868
rect -1120 42548 -1040 42812
rect -1120 42492 -1108 42548
rect -1052 42492 -1040 42548
rect -1120 42228 -1040 42492
rect -1120 42172 -1108 42228
rect -1052 42172 -1040 42228
rect -1440 41852 -1428 41908
rect -1372 41852 -1360 41908
rect -1440 41748 -1360 41852
rect -1440 41692 -1428 41748
rect -1372 41692 -1360 41748
rect -1440 41588 -1360 41692
rect -1440 41532 -1428 41588
rect -1372 41532 -1360 41588
rect -1440 40868 -1360 41532
rect -1440 40812 -1428 40868
rect -1372 40812 -1360 40868
rect -1440 40708 -1360 40812
rect -1440 40652 -1428 40708
rect -1372 40652 -1360 40708
rect -1440 40388 -1360 40652
rect -1120 41908 -1040 42172
rect -1120 41852 -1108 41908
rect -1052 41852 -1040 41908
rect -1120 41748 -1040 41852
rect -1120 41692 -1108 41748
rect -1052 41692 -1040 41748
rect -1120 41588 -1040 41692
rect -1120 41532 -1108 41588
rect -1052 41532 -1040 41588
rect -1120 40868 -1040 41532
rect 41040 41348 41120 41360
rect 41040 41292 41052 41348
rect 41108 41292 41120 41348
rect 41040 41028 41120 41292
rect 41040 40972 41052 41028
rect 41108 40972 41120 41028
rect 41040 40960 41120 40972
rect 41200 41348 41280 41360
rect 41200 41292 41212 41348
rect 41268 41292 41280 41348
rect 41200 41028 41280 41292
rect 41200 40972 41212 41028
rect 41268 40972 41280 41028
rect 41200 40960 41280 40972
rect 41360 41348 41440 41360
rect 41360 41292 41372 41348
rect 41428 41292 41440 41348
rect 41360 41028 41440 41292
rect 41360 40972 41372 41028
rect 41428 40972 41440 41028
rect 41360 40960 41440 40972
rect 41520 41348 41600 41360
rect 41520 41292 41532 41348
rect 41588 41292 41600 41348
rect 41520 41028 41600 41292
rect 41520 40972 41532 41028
rect 41588 40972 41600 41028
rect 41520 40960 41600 40972
rect 41680 41348 41760 41360
rect 41680 41292 41692 41348
rect 41748 41292 41760 41348
rect 41680 41028 41760 41292
rect 41680 40972 41692 41028
rect 41748 40972 41760 41028
rect 41680 40960 41760 40972
rect 41840 41348 41920 41360
rect 41840 41292 41852 41348
rect 41908 41292 41920 41348
rect 41840 41028 41920 41292
rect 41840 40972 41852 41028
rect 41908 40972 41920 41028
rect 41840 40960 41920 40972
rect 42000 41348 42080 41360
rect 42000 41292 42012 41348
rect 42068 41292 42080 41348
rect 42000 41028 42080 41292
rect 42000 40972 42012 41028
rect 42068 40972 42080 41028
rect 42000 40960 42080 40972
rect 42160 41348 42240 41360
rect 42160 41292 42172 41348
rect 42228 41292 42240 41348
rect 42160 41028 42240 41292
rect 42160 40972 42172 41028
rect 42228 40972 42240 41028
rect 42160 40960 42240 40972
rect 42320 41348 42400 41360
rect 42320 41292 42332 41348
rect 42388 41292 42400 41348
rect 42320 41028 42400 41292
rect 42320 40972 42332 41028
rect 42388 40972 42400 41028
rect 42320 40960 42400 40972
rect 42480 41348 42560 41360
rect 42480 41292 42492 41348
rect 42548 41292 42560 41348
rect 42480 41028 42560 41292
rect 42480 40972 42492 41028
rect 42548 40972 42560 41028
rect 42480 40960 42560 40972
rect 42640 41348 42720 41360
rect 42640 41292 42652 41348
rect 42708 41292 42720 41348
rect 42640 41028 42720 41292
rect 42640 40972 42652 41028
rect 42708 40972 42720 41028
rect 42640 40960 42720 40972
rect 42800 41348 42880 41360
rect 42800 41292 42812 41348
rect 42868 41292 42880 41348
rect 42800 41028 42880 41292
rect 42800 40972 42812 41028
rect 42868 40972 42880 41028
rect 42800 40960 42880 40972
rect 42960 41348 43040 41360
rect 42960 41292 42972 41348
rect 43028 41292 43040 41348
rect 42960 41028 43040 41292
rect 42960 40972 42972 41028
rect 43028 40972 43040 41028
rect 42960 40960 43040 40972
rect 43120 41348 43200 41360
rect 43120 41292 43132 41348
rect 43188 41292 43200 41348
rect 43120 41028 43200 41292
rect 43120 40972 43132 41028
rect 43188 40972 43200 41028
rect 43120 40960 43200 40972
rect -1120 40812 -1108 40868
rect -1052 40812 -1040 40868
rect -1120 40708 -1040 40812
rect -1120 40652 -1108 40708
rect -1052 40652 -1040 40708
rect -1440 40332 -1428 40388
rect -1372 40332 -1360 40388
rect -1440 40068 -1360 40332
rect -1440 40012 -1428 40068
rect -1372 40012 -1360 40068
rect -1760 39688 -1752 39752
rect -1688 39688 -1680 39752
rect -1760 39592 -1680 39688
rect -1760 39528 -1752 39592
rect -1688 39528 -1680 39592
rect -1760 39432 -1680 39528
rect -1760 39368 -1752 39432
rect -1688 39368 -1680 39432
rect -1760 39272 -1680 39368
rect -1760 39208 -1752 39272
rect -1688 39208 -1680 39272
rect -1760 39112 -1680 39208
rect -1760 39048 -1752 39112
rect -1688 39048 -1680 39112
rect -1760 38952 -1680 39048
rect -1760 38888 -1752 38952
rect -1688 38888 -1680 38952
rect -1760 38792 -1680 38888
rect -1760 38728 -1752 38792
rect -1688 38728 -1680 38792
rect -1760 38632 -1680 38728
rect -1760 38568 -1752 38632
rect -1688 38568 -1680 38632
rect -1760 38472 -1680 38568
rect -1760 38408 -1752 38472
rect -1688 38408 -1680 38472
rect -1760 38312 -1680 38408
rect -1760 38248 -1752 38312
rect -1688 38248 -1680 38312
rect -1760 38152 -1680 38248
rect -1760 38088 -1752 38152
rect -1688 38088 -1680 38152
rect -1760 37992 -1680 38088
rect -1760 37928 -1752 37992
rect -1688 37928 -1680 37992
rect -1760 37832 -1680 37928
rect -1760 37768 -1752 37832
rect -1688 37768 -1680 37832
rect -1760 37668 -1680 37768
rect -1760 37612 -1748 37668
rect -1692 37612 -1680 37668
rect -1760 37512 -1680 37612
rect -1760 37448 -1752 37512
rect -1688 37448 -1680 37512
rect -1760 37352 -1680 37448
rect -1760 37288 -1752 37352
rect -1688 37288 -1680 37352
rect -1760 37192 -1680 37288
rect -1760 37128 -1752 37192
rect -1688 37128 -1680 37192
rect -1760 37032 -1680 37128
rect -1760 36968 -1752 37032
rect -1688 36968 -1680 37032
rect -1760 36872 -1680 36968
rect -1760 36808 -1752 36872
rect -1688 36808 -1680 36872
rect -1760 36712 -1680 36808
rect -1760 36648 -1752 36712
rect -1688 36648 -1680 36712
rect -1760 36552 -1680 36648
rect -1760 36488 -1752 36552
rect -1688 36488 -1680 36552
rect -1760 36392 -1680 36488
rect -1760 36328 -1752 36392
rect -1688 36328 -1680 36392
rect -2080 36012 -2068 36068
rect -2012 36012 -2000 36068
rect -2080 35752 -2000 36012
rect -2080 35688 -2072 35752
rect -2008 35688 -2000 35752
rect -2080 35592 -2000 35688
rect -2080 35528 -2072 35592
rect -2008 35528 -2000 35592
rect -2080 35432 -2000 35528
rect -2080 35368 -2072 35432
rect -2008 35368 -2000 35432
rect -2080 35272 -2000 35368
rect -2080 35208 -2072 35272
rect -2008 35208 -2000 35272
rect -2080 35112 -2000 35208
rect -2080 35048 -2072 35112
rect -2008 35048 -2000 35112
rect -2080 34952 -2000 35048
rect -2080 34888 -2072 34952
rect -2008 34888 -2000 34952
rect -2080 34792 -2000 34888
rect -2080 34728 -2072 34792
rect -2008 34728 -2000 34792
rect -2080 34632 -2000 34728
rect -2080 34568 -2072 34632
rect -2008 34568 -2000 34632
rect -2080 34472 -2000 34568
rect -2080 34408 -2072 34472
rect -2008 34408 -2000 34472
rect -2080 34312 -2000 34408
rect -2080 34248 -2072 34312
rect -2008 34248 -2000 34312
rect -2080 34152 -2000 34248
rect -2080 34088 -2072 34152
rect -2008 34088 -2000 34152
rect -2080 33992 -2000 34088
rect -2080 33928 -2072 33992
rect -2008 33928 -2000 33992
rect -2080 33832 -2000 33928
rect -2080 33768 -2072 33832
rect -2008 33768 -2000 33832
rect -2080 33672 -2000 33768
rect -2080 33608 -2072 33672
rect -2008 33608 -2000 33672
rect -2080 33512 -2000 33608
rect -2080 33448 -2072 33512
rect -2008 33448 -2000 33512
rect -2080 33272 -2000 33448
rect -2080 33208 -2072 33272
rect -2008 33208 -2000 33272
rect -2080 33112 -2000 33208
rect -2080 33048 -2072 33112
rect -2008 33048 -2000 33112
rect -2080 32948 -2000 33048
rect -2080 32892 -2068 32948
rect -2012 32892 -2000 32948
rect -2080 32628 -2000 32892
rect -2080 32572 -2068 32628
rect -2012 32572 -2000 32628
rect -2080 32308 -2000 32572
rect -2080 32252 -2068 32308
rect -2012 32252 -2000 32308
rect -2400 31932 -2388 31988
rect -2332 31932 -2320 31988
rect -2400 31920 -2320 31932
rect -2080 31988 -2000 32252
rect -2080 31932 -2068 31988
rect -2012 31932 -2000 31988
rect -2080 31840 -2000 31932
rect -1920 36228 -1840 36240
rect -1920 36172 -1908 36228
rect -1852 36172 -1840 36228
rect -1920 31840 -1840 36172
rect -1760 36068 -1680 36328
rect -1760 36012 -1748 36068
rect -1692 36012 -1680 36068
rect -1760 35752 -1680 36012
rect -1440 39752 -1360 40012
rect -1440 39688 -1432 39752
rect -1368 39688 -1360 39752
rect -1440 39592 -1360 39688
rect -1440 39528 -1432 39592
rect -1368 39528 -1360 39592
rect -1440 39432 -1360 39528
rect -1440 39368 -1432 39432
rect -1368 39368 -1360 39432
rect -1440 39272 -1360 39368
rect -1440 39208 -1432 39272
rect -1368 39208 -1360 39272
rect -1440 39112 -1360 39208
rect -1440 39048 -1432 39112
rect -1368 39048 -1360 39112
rect -1440 38952 -1360 39048
rect -1440 38888 -1432 38952
rect -1368 38888 -1360 38952
rect -1440 38792 -1360 38888
rect -1440 38728 -1432 38792
rect -1368 38728 -1360 38792
rect -1440 38632 -1360 38728
rect -1440 38568 -1432 38632
rect -1368 38568 -1360 38632
rect -1440 38472 -1360 38568
rect -1440 38408 -1432 38472
rect -1368 38408 -1360 38472
rect -1440 38312 -1360 38408
rect -1440 38248 -1432 38312
rect -1368 38248 -1360 38312
rect -1440 38152 -1360 38248
rect -1440 38088 -1432 38152
rect -1368 38088 -1360 38152
rect -1440 37992 -1360 38088
rect -1440 37928 -1432 37992
rect -1368 37928 -1360 37992
rect -1440 37832 -1360 37928
rect -1440 37768 -1432 37832
rect -1368 37768 -1360 37832
rect -1440 37668 -1360 37768
rect -1440 37612 -1428 37668
rect -1372 37612 -1360 37668
rect -1440 37512 -1360 37612
rect -1280 40548 -1200 40560
rect -1280 40492 -1268 40548
rect -1212 40492 -1200 40548
rect -1280 37668 -1200 40492
rect -1280 37612 -1268 37668
rect -1212 37612 -1200 37668
rect -1280 37600 -1200 37612
rect -1120 40388 -1040 40652
rect -1120 40332 -1108 40388
rect -1052 40332 -1040 40388
rect -1120 40068 -1040 40332
rect -1120 40012 -1108 40068
rect -1052 40012 -1040 40068
rect -1120 39752 -1040 40012
rect -1120 39688 -1112 39752
rect -1048 39688 -1040 39752
rect -1120 39592 -1040 39688
rect 41040 40068 41120 40080
rect 41040 40012 41052 40068
rect 41108 40012 41120 40068
rect 41040 39748 41120 40012
rect 41040 39692 41052 39748
rect 41108 39692 41120 39748
rect 41040 39680 41120 39692
rect 41200 40068 41280 40080
rect 41200 40012 41212 40068
rect 41268 40012 41280 40068
rect 41200 39748 41280 40012
rect 41200 39692 41212 39748
rect 41268 39692 41280 39748
rect 41200 39680 41280 39692
rect 41360 40068 41440 40080
rect 41360 40012 41372 40068
rect 41428 40012 41440 40068
rect 41360 39748 41440 40012
rect 41360 39692 41372 39748
rect 41428 39692 41440 39748
rect 41360 39680 41440 39692
rect 41520 40068 41600 40080
rect 41520 40012 41532 40068
rect 41588 40012 41600 40068
rect 41520 39748 41600 40012
rect 41520 39692 41532 39748
rect 41588 39692 41600 39748
rect 41520 39680 41600 39692
rect 41680 40068 41760 40080
rect 41680 40012 41692 40068
rect 41748 40012 41760 40068
rect 41680 39748 41760 40012
rect 41680 39692 41692 39748
rect 41748 39692 41760 39748
rect 41680 39680 41760 39692
rect 41840 40068 41920 40080
rect 41840 40012 41852 40068
rect 41908 40012 41920 40068
rect 41840 39748 41920 40012
rect 41840 39692 41852 39748
rect 41908 39692 41920 39748
rect 41840 39680 41920 39692
rect 42000 40068 42080 40080
rect 42000 40012 42012 40068
rect 42068 40012 42080 40068
rect 42000 39748 42080 40012
rect 42000 39692 42012 39748
rect 42068 39692 42080 39748
rect 42000 39680 42080 39692
rect 42160 40068 42240 40080
rect 42160 40012 42172 40068
rect 42228 40012 42240 40068
rect 42160 39748 42240 40012
rect 42160 39692 42172 39748
rect 42228 39692 42240 39748
rect 42160 39680 42240 39692
rect 42320 40068 42400 40080
rect 42320 40012 42332 40068
rect 42388 40012 42400 40068
rect 42320 39748 42400 40012
rect 42320 39692 42332 39748
rect 42388 39692 42400 39748
rect 42320 39680 42400 39692
rect 42480 40068 42560 40080
rect 42480 40012 42492 40068
rect 42548 40012 42560 40068
rect 42480 39748 42560 40012
rect 42480 39692 42492 39748
rect 42548 39692 42560 39748
rect 42480 39680 42560 39692
rect 42640 40068 42720 40080
rect 42640 40012 42652 40068
rect 42708 40012 42720 40068
rect 42640 39748 42720 40012
rect 42640 39692 42652 39748
rect 42708 39692 42720 39748
rect 42640 39680 42720 39692
rect 42800 40068 42880 40080
rect 42800 40012 42812 40068
rect 42868 40012 42880 40068
rect 42800 39748 42880 40012
rect 42800 39692 42812 39748
rect 42868 39692 42880 39748
rect 42800 39680 42880 39692
rect 42960 40068 43040 40080
rect 42960 40012 42972 40068
rect 43028 40012 43040 40068
rect 42960 39748 43040 40012
rect 42960 39692 42972 39748
rect 43028 39692 43040 39748
rect 42960 39680 43040 39692
rect 43120 40068 43200 40080
rect 43120 40012 43132 40068
rect 43188 40012 43200 40068
rect 43120 39748 43200 40012
rect 43120 39692 43132 39748
rect 43188 39692 43200 39748
rect 43120 39680 43200 39692
rect -1120 39528 -1112 39592
rect -1048 39528 -1040 39592
rect -1120 39432 -1040 39528
rect -1120 39368 -1112 39432
rect -1048 39368 -1040 39432
rect -1120 39272 -1040 39368
rect -1120 39208 -1112 39272
rect -1048 39208 -1040 39272
rect -1120 39112 -1040 39208
rect -1120 39048 -1112 39112
rect -1048 39048 -1040 39112
rect -1120 38952 -1040 39048
rect -1120 38888 -1112 38952
rect -1048 38888 -1040 38952
rect -1120 38792 -1040 38888
rect -1120 38728 -1112 38792
rect -1048 38728 -1040 38792
rect -1120 38632 -1040 38728
rect -1120 38568 -1112 38632
rect -1048 38568 -1040 38632
rect -1120 38472 -1040 38568
rect -1120 38408 -1112 38472
rect -1048 38408 -1040 38472
rect -1120 38312 -1040 38408
rect -1120 38248 -1112 38312
rect -1048 38248 -1040 38312
rect -1120 38152 -1040 38248
rect -1120 38088 -1112 38152
rect -1048 38088 -1040 38152
rect -1120 37992 -1040 38088
rect -1120 37928 -1112 37992
rect -1048 37928 -1040 37992
rect -1120 37832 -1040 37928
rect -1120 37768 -1112 37832
rect -1048 37768 -1040 37832
rect -1440 37448 -1432 37512
rect -1368 37448 -1360 37512
rect -1440 37352 -1360 37448
rect -1440 37288 -1432 37352
rect -1368 37288 -1360 37352
rect -1440 37192 -1360 37288
rect -1440 37128 -1432 37192
rect -1368 37128 -1360 37192
rect -1440 37032 -1360 37128
rect -1440 36968 -1432 37032
rect -1368 36968 -1360 37032
rect -1440 36872 -1360 36968
rect -1440 36808 -1432 36872
rect -1368 36808 -1360 36872
rect -1440 36712 -1360 36808
rect -1440 36648 -1432 36712
rect -1368 36648 -1360 36712
rect -1440 36552 -1360 36648
rect -1440 36488 -1432 36552
rect -1368 36488 -1360 36552
rect -1440 36392 -1360 36488
rect -1440 36328 -1432 36392
rect -1368 36328 -1360 36392
rect -1440 36068 -1360 36328
rect -1440 36012 -1428 36068
rect -1372 36012 -1360 36068
rect -1760 35688 -1752 35752
rect -1688 35688 -1680 35752
rect -1760 35592 -1680 35688
rect -1760 35528 -1752 35592
rect -1688 35528 -1680 35592
rect -1760 35432 -1680 35528
rect -1760 35368 -1752 35432
rect -1688 35368 -1680 35432
rect -1760 35272 -1680 35368
rect -1760 35208 -1752 35272
rect -1688 35208 -1680 35272
rect -1760 35112 -1680 35208
rect -1760 35048 -1752 35112
rect -1688 35048 -1680 35112
rect -1760 34952 -1680 35048
rect -1760 34888 -1752 34952
rect -1688 34888 -1680 34952
rect -1760 34792 -1680 34888
rect -1760 34728 -1752 34792
rect -1688 34728 -1680 34792
rect -1760 34632 -1680 34728
rect -1760 34568 -1752 34632
rect -1688 34568 -1680 34632
rect -1760 34472 -1680 34568
rect -1760 34408 -1752 34472
rect -1688 34408 -1680 34472
rect -1760 34312 -1680 34408
rect -1760 34248 -1752 34312
rect -1688 34248 -1680 34312
rect -1760 34152 -1680 34248
rect -1760 34088 -1752 34152
rect -1688 34088 -1680 34152
rect -1760 33992 -1680 34088
rect -1760 33928 -1752 33992
rect -1688 33928 -1680 33992
rect -1760 33832 -1680 33928
rect -1760 33768 -1752 33832
rect -1688 33768 -1680 33832
rect -1760 33672 -1680 33768
rect -1760 33608 -1752 33672
rect -1688 33608 -1680 33672
rect -1760 33512 -1680 33608
rect -1760 33448 -1752 33512
rect -1688 33448 -1680 33512
rect -1760 33272 -1680 33448
rect -1760 33208 -1752 33272
rect -1688 33208 -1680 33272
rect -1760 33112 -1680 33208
rect -1760 33048 -1752 33112
rect -1688 33048 -1680 33112
rect -1760 32948 -1680 33048
rect -1760 32892 -1748 32948
rect -1692 32892 -1680 32948
rect -1760 32628 -1680 32892
rect -1760 32572 -1748 32628
rect -1692 32572 -1680 32628
rect -1760 32308 -1680 32572
rect -1760 32252 -1748 32308
rect -1692 32252 -1680 32308
rect -1760 31988 -1680 32252
rect -1760 31932 -1748 31988
rect -1692 31932 -1680 31988
rect -1760 31840 -1680 31932
rect -1600 35908 -1520 35920
rect -1600 35852 -1588 35908
rect -1532 35852 -1520 35908
rect -1600 31840 -1520 35852
rect -1440 35752 -1360 36012
rect -1440 35688 -1432 35752
rect -1368 35688 -1360 35752
rect -1440 35592 -1360 35688
rect -1440 35528 -1432 35592
rect -1368 35528 -1360 35592
rect -1440 35432 -1360 35528
rect -1440 35368 -1432 35432
rect -1368 35368 -1360 35432
rect -1440 35272 -1360 35368
rect -1440 35208 -1432 35272
rect -1368 35208 -1360 35272
rect -1440 35112 -1360 35208
rect -1440 35048 -1432 35112
rect -1368 35048 -1360 35112
rect -1440 34952 -1360 35048
rect -1440 34888 -1432 34952
rect -1368 34888 -1360 34952
rect -1440 34792 -1360 34888
rect -1440 34728 -1432 34792
rect -1368 34728 -1360 34792
rect -1440 34632 -1360 34728
rect -1440 34568 -1432 34632
rect -1368 34568 -1360 34632
rect -1440 34472 -1360 34568
rect -1440 34408 -1432 34472
rect -1368 34408 -1360 34472
rect -1440 34312 -1360 34408
rect -1440 34248 -1432 34312
rect -1368 34248 -1360 34312
rect -1440 34152 -1360 34248
rect -1440 34088 -1432 34152
rect -1368 34088 -1360 34152
rect -1440 33992 -1360 34088
rect -1440 33928 -1432 33992
rect -1368 33928 -1360 33992
rect -1440 33832 -1360 33928
rect -1440 33768 -1432 33832
rect -1368 33768 -1360 33832
rect -1440 33672 -1360 33768
rect -1440 33608 -1432 33672
rect -1368 33608 -1360 33672
rect -1440 33512 -1360 33608
rect -1440 33448 -1432 33512
rect -1368 33448 -1360 33512
rect -1440 33272 -1360 33448
rect -1440 33208 -1432 33272
rect -1368 33208 -1360 33272
rect -1440 33112 -1360 33208
rect -1440 33048 -1432 33112
rect -1368 33048 -1360 33112
rect -1440 32948 -1360 33048
rect -1440 32892 -1428 32948
rect -1372 32892 -1360 32948
rect -1440 32628 -1360 32892
rect -1120 37512 -1040 37768
rect -1120 37448 -1112 37512
rect -1048 37448 -1040 37512
rect -1120 37352 -1040 37448
rect -1120 37288 -1112 37352
rect -1048 37288 -1040 37352
rect -1120 37192 -1040 37288
rect -1120 37128 -1112 37192
rect -1048 37128 -1040 37192
rect -1120 37032 -1040 37128
rect -1120 36968 -1112 37032
rect -1048 36968 -1040 37032
rect -1120 36872 -1040 36968
rect -1120 36808 -1112 36872
rect -1048 36808 -1040 36872
rect -1120 36712 -1040 36808
rect -1120 36648 -1112 36712
rect -1048 36648 -1040 36712
rect -1120 36552 -1040 36648
rect -1120 36488 -1112 36552
rect -1048 36488 -1040 36552
rect -1120 36392 -1040 36488
rect -1120 36328 -1112 36392
rect -1048 36328 -1040 36392
rect -1120 36068 -1040 36328
rect -1120 36012 -1108 36068
rect -1052 36012 -1040 36068
rect -1120 35752 -1040 36012
rect -1120 35688 -1112 35752
rect -1048 35688 -1040 35752
rect -1120 35592 -1040 35688
rect 41040 36068 41120 36080
rect 41040 36012 41052 36068
rect 41108 36012 41120 36068
rect 41040 35748 41120 36012
rect 41040 35692 41052 35748
rect 41108 35692 41120 35748
rect 41040 35680 41120 35692
rect 41200 36068 41280 36080
rect 41200 36012 41212 36068
rect 41268 36012 41280 36068
rect 41200 35748 41280 36012
rect 41200 35692 41212 35748
rect 41268 35692 41280 35748
rect 41200 35680 41280 35692
rect 41360 36068 41440 36080
rect 41360 36012 41372 36068
rect 41428 36012 41440 36068
rect 41360 35748 41440 36012
rect 41360 35692 41372 35748
rect 41428 35692 41440 35748
rect 41360 35680 41440 35692
rect 41520 36068 41600 36080
rect 41520 36012 41532 36068
rect 41588 36012 41600 36068
rect 41520 35748 41600 36012
rect 41520 35692 41532 35748
rect 41588 35692 41600 35748
rect 41520 35680 41600 35692
rect 41680 36068 41760 36080
rect 41680 36012 41692 36068
rect 41748 36012 41760 36068
rect 41680 35748 41760 36012
rect 41680 35692 41692 35748
rect 41748 35692 41760 35748
rect 41680 35680 41760 35692
rect 41840 36068 41920 36080
rect 41840 36012 41852 36068
rect 41908 36012 41920 36068
rect 41840 35748 41920 36012
rect 41840 35692 41852 35748
rect 41908 35692 41920 35748
rect 41840 35680 41920 35692
rect 42000 36068 42080 36080
rect 42000 36012 42012 36068
rect 42068 36012 42080 36068
rect 42000 35748 42080 36012
rect 42000 35692 42012 35748
rect 42068 35692 42080 35748
rect 42000 35680 42080 35692
rect 42160 36068 42240 36080
rect 42160 36012 42172 36068
rect 42228 36012 42240 36068
rect 42160 35748 42240 36012
rect 42160 35692 42172 35748
rect 42228 35692 42240 35748
rect 42160 35680 42240 35692
rect 42320 36068 42400 36080
rect 42320 36012 42332 36068
rect 42388 36012 42400 36068
rect 42320 35748 42400 36012
rect 42320 35692 42332 35748
rect 42388 35692 42400 35748
rect 42320 35680 42400 35692
rect 42480 36068 42560 36080
rect 42480 36012 42492 36068
rect 42548 36012 42560 36068
rect 42480 35748 42560 36012
rect 42480 35692 42492 35748
rect 42548 35692 42560 35748
rect 42480 35680 42560 35692
rect 42640 36068 42720 36080
rect 42640 36012 42652 36068
rect 42708 36012 42720 36068
rect 42640 35748 42720 36012
rect 42640 35692 42652 35748
rect 42708 35692 42720 35748
rect 42640 35680 42720 35692
rect 42800 36068 42880 36080
rect 42800 36012 42812 36068
rect 42868 36012 42880 36068
rect 42800 35748 42880 36012
rect 42800 35692 42812 35748
rect 42868 35692 42880 35748
rect 42800 35680 42880 35692
rect 42960 36068 43040 36080
rect 42960 36012 42972 36068
rect 43028 36012 43040 36068
rect 42960 35748 43040 36012
rect 42960 35692 42972 35748
rect 43028 35692 43040 35748
rect 42960 35680 43040 35692
rect 43120 36068 43200 36080
rect 43120 36012 43132 36068
rect 43188 36012 43200 36068
rect 43120 35748 43200 36012
rect 43120 35692 43132 35748
rect 43188 35692 43200 35748
rect 43120 35680 43200 35692
rect -1120 35528 -1112 35592
rect -1048 35528 -1040 35592
rect -1120 35432 -1040 35528
rect -1120 35368 -1112 35432
rect -1048 35368 -1040 35432
rect -1120 35272 -1040 35368
rect -1120 35208 -1112 35272
rect -1048 35208 -1040 35272
rect -1120 35112 -1040 35208
rect -1120 35048 -1112 35112
rect -1048 35048 -1040 35112
rect -1120 34952 -1040 35048
rect -1120 34888 -1112 34952
rect -1048 34888 -1040 34952
rect -1120 34792 -1040 34888
rect -1120 34728 -1112 34792
rect -1048 34728 -1040 34792
rect -1120 34632 -1040 34728
rect -1120 34568 -1112 34632
rect -1048 34568 -1040 34632
rect -1120 34472 -1040 34568
rect -1120 34408 -1112 34472
rect -1048 34408 -1040 34472
rect -1120 34312 -1040 34408
rect -1120 34248 -1112 34312
rect -1048 34248 -1040 34312
rect -1120 34152 -1040 34248
rect -1120 34088 -1112 34152
rect -1048 34088 -1040 34152
rect -1120 33992 -1040 34088
rect -1120 33928 -1112 33992
rect -1048 33928 -1040 33992
rect -1120 33832 -1040 33928
rect -1120 33768 -1112 33832
rect -1048 33768 -1040 33832
rect -1120 33672 -1040 33768
rect -1120 33608 -1112 33672
rect -1048 33608 -1040 33672
rect -1120 33512 -1040 33608
rect -1120 33448 -1112 33512
rect -1048 33448 -1040 33512
rect -1120 33272 -1040 33448
rect -1120 33208 -1112 33272
rect -1048 33208 -1040 33272
rect -1120 33112 -1040 33208
rect -1120 33048 -1112 33112
rect -1048 33048 -1040 33112
rect -1120 32948 -1040 33048
rect -1120 32892 -1108 32948
rect -1052 32892 -1040 32948
rect -1440 32572 -1428 32628
rect -1372 32572 -1360 32628
rect -1440 32308 -1360 32572
rect -1440 32252 -1428 32308
rect -1372 32252 -1360 32308
rect -1440 31988 -1360 32252
rect -1440 31932 -1428 31988
rect -1372 31932 -1360 31988
rect -1440 31840 -1360 31932
rect -1280 32788 -1200 32800
rect -1280 32732 -1268 32788
rect -1212 32732 -1200 32788
rect -1280 31840 -1200 32732
rect -1120 32628 -1040 32892
rect -1120 32572 -1108 32628
rect -1052 32572 -1040 32628
rect -1120 32308 -1040 32572
rect -1120 32252 -1108 32308
rect -1052 32252 -1040 32308
rect -1120 31988 -1040 32252
rect -1120 31932 -1108 31988
rect -1052 31932 -1040 31988
rect -1120 31840 -1040 31932
<< via3 >>
rect -31032 41748 -30968 41752
rect -31032 41692 -31028 41748
rect -31028 41692 -30972 41748
rect -30972 41692 -30968 41748
rect -31032 41688 -30968 41692
rect -31032 41588 -30968 41592
rect -31032 41532 -31028 41588
rect -31028 41532 -30972 41588
rect -30972 41532 -30968 41588
rect -31032 41528 -30968 41532
rect -31032 40788 -30968 40792
rect -31032 40732 -31028 40788
rect -31028 40732 -30972 40788
rect -30972 40732 -30968 40788
rect -31032 40728 -30968 40732
rect -31032 40628 -30968 40632
rect -31032 40572 -31028 40628
rect -31028 40572 -30972 40628
rect -30972 40572 -30968 40628
rect -31032 40568 -30968 40572
rect -31032 40468 -30968 40472
rect -31032 40412 -31028 40468
rect -31028 40412 -30972 40468
rect -30972 40412 -30968 40468
rect -31032 40408 -30968 40412
rect -31032 40308 -30968 40312
rect -31032 40252 -31028 40308
rect -31028 40252 -30972 40308
rect -30972 40252 -30968 40308
rect -31032 40248 -30968 40252
rect -31032 40148 -30968 40152
rect -31032 40092 -31028 40148
rect -31028 40092 -30972 40148
rect -30972 40092 -30968 40148
rect -31032 40088 -30968 40092
rect -31032 39988 -30968 39992
rect -31032 39932 -31028 39988
rect -31028 39932 -30972 39988
rect -30972 39932 -30968 39988
rect -31032 39928 -30968 39932
rect -31032 39828 -30968 39832
rect -31032 39772 -31028 39828
rect -31028 39772 -30972 39828
rect -30972 39772 -30968 39828
rect -31032 39768 -30968 39772
rect -31032 39668 -30968 39672
rect -31032 39612 -31028 39668
rect -31028 39612 -30972 39668
rect -30972 39612 -30968 39668
rect -31032 39608 -30968 39612
rect -31032 39508 -30968 39512
rect -31032 39452 -31028 39508
rect -31028 39452 -30972 39508
rect -30972 39452 -30968 39508
rect -31032 39448 -30968 39452
rect -31032 39348 -30968 39352
rect -31032 39292 -31028 39348
rect -31028 39292 -30972 39348
rect -30972 39292 -30968 39348
rect -31032 39288 -30968 39292
rect -31032 39188 -30968 39192
rect -31032 39132 -31028 39188
rect -31028 39132 -30972 39188
rect -30972 39132 -30968 39188
rect -31032 39128 -30968 39132
rect -31032 39028 -30968 39032
rect -31032 38972 -31028 39028
rect -31028 38972 -30972 39028
rect -30972 38972 -30968 39028
rect -31032 38968 -30968 38972
rect -31032 38868 -30968 38872
rect -31032 38812 -31028 38868
rect -31028 38812 -30972 38868
rect -30972 38812 -30968 38868
rect -31032 38808 -30968 38812
rect -31032 38708 -30968 38712
rect -31032 38652 -31028 38708
rect -31028 38652 -30972 38708
rect -30972 38652 -30968 38708
rect -31032 38648 -30968 38652
rect -31032 38548 -30968 38552
rect -31032 38492 -31028 38548
rect -31028 38492 -30972 38548
rect -30972 38492 -30968 38548
rect -31032 38488 -30968 38492
rect -31032 38388 -30968 38392
rect -31032 38332 -31028 38388
rect -31028 38332 -30972 38388
rect -30972 38332 -30968 38388
rect -31032 38328 -30968 38332
rect -31032 38228 -30968 38232
rect -31032 38172 -31028 38228
rect -31028 38172 -30972 38228
rect -30972 38172 -30968 38228
rect -31032 38168 -30968 38172
rect -31032 38068 -30968 38072
rect -31032 38012 -31028 38068
rect -31028 38012 -30972 38068
rect -30972 38012 -30968 38068
rect -31032 38008 -30968 38012
rect -31032 37908 -30968 37912
rect -31032 37852 -31028 37908
rect -31028 37852 -30972 37908
rect -30972 37852 -30968 37908
rect -31032 37848 -30968 37852
rect -31032 37748 -30968 37752
rect -31032 37692 -31028 37748
rect -31028 37692 -30972 37748
rect -30972 37692 -30968 37748
rect -31032 37688 -30968 37692
rect -30712 41748 -30648 41752
rect -30712 41692 -30708 41748
rect -30708 41692 -30652 41748
rect -30652 41692 -30648 41748
rect -30712 41688 -30648 41692
rect -30712 41588 -30648 41592
rect -30712 41532 -30708 41588
rect -30708 41532 -30652 41588
rect -30652 41532 -30648 41588
rect -30712 41528 -30648 41532
rect -30712 40788 -30648 40792
rect -30712 40732 -30708 40788
rect -30708 40732 -30652 40788
rect -30652 40732 -30648 40788
rect -30712 40728 -30648 40732
rect -30712 40628 -30648 40632
rect -30712 40572 -30708 40628
rect -30708 40572 -30652 40628
rect -30652 40572 -30648 40628
rect -30712 40568 -30648 40572
rect -30712 40468 -30648 40472
rect -30712 40412 -30708 40468
rect -30708 40412 -30652 40468
rect -30652 40412 -30648 40468
rect -30712 40408 -30648 40412
rect -30712 40308 -30648 40312
rect -30712 40252 -30708 40308
rect -30708 40252 -30652 40308
rect -30652 40252 -30648 40308
rect -30712 40248 -30648 40252
rect -30712 40148 -30648 40152
rect -30712 40092 -30708 40148
rect -30708 40092 -30652 40148
rect -30652 40092 -30648 40148
rect -30712 40088 -30648 40092
rect -30712 39988 -30648 39992
rect -30712 39932 -30708 39988
rect -30708 39932 -30652 39988
rect -30652 39932 -30648 39988
rect -30712 39928 -30648 39932
rect -30712 39828 -30648 39832
rect -30712 39772 -30708 39828
rect -30708 39772 -30652 39828
rect -30652 39772 -30648 39828
rect -30712 39768 -30648 39772
rect -30712 39668 -30648 39672
rect -30712 39612 -30708 39668
rect -30708 39612 -30652 39668
rect -30652 39612 -30648 39668
rect -30712 39608 -30648 39612
rect -30712 39508 -30648 39512
rect -30712 39452 -30708 39508
rect -30708 39452 -30652 39508
rect -30652 39452 -30648 39508
rect -30712 39448 -30648 39452
rect -30712 39348 -30648 39352
rect -30712 39292 -30708 39348
rect -30708 39292 -30652 39348
rect -30652 39292 -30648 39348
rect -30712 39288 -30648 39292
rect -30712 39188 -30648 39192
rect -30712 39132 -30708 39188
rect -30708 39132 -30652 39188
rect -30652 39132 -30648 39188
rect -30712 39128 -30648 39132
rect -30712 39028 -30648 39032
rect -30712 38972 -30708 39028
rect -30708 38972 -30652 39028
rect -30652 38972 -30648 39028
rect -30712 38968 -30648 38972
rect -30712 38868 -30648 38872
rect -30712 38812 -30708 38868
rect -30708 38812 -30652 38868
rect -30652 38812 -30648 38868
rect -30712 38808 -30648 38812
rect -30712 38708 -30648 38712
rect -30712 38652 -30708 38708
rect -30708 38652 -30652 38708
rect -30652 38652 -30648 38708
rect -30712 38648 -30648 38652
rect -30712 38548 -30648 38552
rect -30712 38492 -30708 38548
rect -30708 38492 -30652 38548
rect -30652 38492 -30648 38548
rect -30712 38488 -30648 38492
rect -30712 38388 -30648 38392
rect -30712 38332 -30708 38388
rect -30708 38332 -30652 38388
rect -30652 38332 -30648 38388
rect -30712 38328 -30648 38332
rect -30712 38228 -30648 38232
rect -30712 38172 -30708 38228
rect -30708 38172 -30652 38228
rect -30652 38172 -30648 38228
rect -30712 38168 -30648 38172
rect -30712 38068 -30648 38072
rect -30712 38012 -30708 38068
rect -30708 38012 -30652 38068
rect -30652 38012 -30648 38068
rect -30712 38008 -30648 38012
rect -30712 37908 -30648 37912
rect -30712 37852 -30708 37908
rect -30708 37852 -30652 37908
rect -30652 37852 -30648 37908
rect -30712 37848 -30648 37852
rect -30712 37748 -30648 37752
rect -30712 37692 -30708 37748
rect -30708 37692 -30652 37748
rect -30652 37692 -30648 37748
rect -30712 37688 -30648 37692
rect -30392 41748 -30328 41752
rect -30392 41692 -30388 41748
rect -30388 41692 -30332 41748
rect -30332 41692 -30328 41748
rect -30392 41688 -30328 41692
rect -30392 41588 -30328 41592
rect -30392 41532 -30388 41588
rect -30388 41532 -30332 41588
rect -30332 41532 -30328 41588
rect -30392 41528 -30328 41532
rect -30392 40788 -30328 40792
rect -30392 40732 -30388 40788
rect -30388 40732 -30332 40788
rect -30332 40732 -30328 40788
rect -30392 40728 -30328 40732
rect -30392 40628 -30328 40632
rect -30392 40572 -30388 40628
rect -30388 40572 -30332 40628
rect -30332 40572 -30328 40628
rect -30392 40568 -30328 40572
rect -30392 40468 -30328 40472
rect -30392 40412 -30388 40468
rect -30388 40412 -30332 40468
rect -30332 40412 -30328 40468
rect -30392 40408 -30328 40412
rect -30392 40308 -30328 40312
rect -30392 40252 -30388 40308
rect -30388 40252 -30332 40308
rect -30332 40252 -30328 40308
rect -30392 40248 -30328 40252
rect -30392 40148 -30328 40152
rect -30392 40092 -30388 40148
rect -30388 40092 -30332 40148
rect -30332 40092 -30328 40148
rect -30392 40088 -30328 40092
rect -30392 39988 -30328 39992
rect -30392 39932 -30388 39988
rect -30388 39932 -30332 39988
rect -30332 39932 -30328 39988
rect -30392 39928 -30328 39932
rect -30392 39828 -30328 39832
rect -30392 39772 -30388 39828
rect -30388 39772 -30332 39828
rect -30332 39772 -30328 39828
rect -30392 39768 -30328 39772
rect -30392 39668 -30328 39672
rect -30392 39612 -30388 39668
rect -30388 39612 -30332 39668
rect -30332 39612 -30328 39668
rect -30392 39608 -30328 39612
rect -30392 39508 -30328 39512
rect -30392 39452 -30388 39508
rect -30388 39452 -30332 39508
rect -30332 39452 -30328 39508
rect -30392 39448 -30328 39452
rect -30392 39348 -30328 39352
rect -30392 39292 -30388 39348
rect -30388 39292 -30332 39348
rect -30332 39292 -30328 39348
rect -30392 39288 -30328 39292
rect -30392 39188 -30328 39192
rect -30392 39132 -30388 39188
rect -30388 39132 -30332 39188
rect -30332 39132 -30328 39188
rect -30392 39128 -30328 39132
rect -30392 39028 -30328 39032
rect -30392 38972 -30388 39028
rect -30388 38972 -30332 39028
rect -30332 38972 -30328 39028
rect -30392 38968 -30328 38972
rect -30392 38868 -30328 38872
rect -30392 38812 -30388 38868
rect -30388 38812 -30332 38868
rect -30332 38812 -30328 38868
rect -30392 38808 -30328 38812
rect -30392 38708 -30328 38712
rect -30392 38652 -30388 38708
rect -30388 38652 -30332 38708
rect -30332 38652 -30328 38708
rect -30392 38648 -30328 38652
rect -30392 38548 -30328 38552
rect -30392 38492 -30388 38548
rect -30388 38492 -30332 38548
rect -30332 38492 -30328 38548
rect -30392 38488 -30328 38492
rect -30392 38388 -30328 38392
rect -30392 38332 -30388 38388
rect -30388 38332 -30332 38388
rect -30332 38332 -30328 38388
rect -30392 38328 -30328 38332
rect -30392 38228 -30328 38232
rect -30392 38172 -30388 38228
rect -30388 38172 -30332 38228
rect -30332 38172 -30328 38228
rect -30392 38168 -30328 38172
rect -30392 38068 -30328 38072
rect -30392 38012 -30388 38068
rect -30388 38012 -30332 38068
rect -30332 38012 -30328 38068
rect -30392 38008 -30328 38012
rect -30392 37908 -30328 37912
rect -30392 37852 -30388 37908
rect -30388 37852 -30332 37908
rect -30332 37852 -30328 37908
rect -30392 37848 -30328 37852
rect -30392 37748 -30328 37752
rect -30392 37692 -30388 37748
rect -30388 37692 -30332 37748
rect -30332 37692 -30328 37748
rect -30392 37688 -30328 37692
rect -31032 37108 -30968 37112
rect -31032 37052 -31028 37108
rect -31028 37052 -30972 37108
rect -30972 37052 -30968 37108
rect -31032 37048 -30968 37052
rect -31032 36948 -30968 36952
rect -31032 36892 -31028 36948
rect -31028 36892 -30972 36948
rect -30972 36892 -30968 36948
rect -31032 36888 -30968 36892
rect -31032 36788 -30968 36792
rect -31032 36732 -31028 36788
rect -31028 36732 -30972 36788
rect -30972 36732 -30968 36788
rect -31032 36728 -30968 36732
rect -31032 36628 -30968 36632
rect -31032 36572 -31028 36628
rect -31028 36572 -30972 36628
rect -30972 36572 -30968 36628
rect -31032 36568 -30968 36572
rect -31032 36468 -30968 36472
rect -31032 36412 -31028 36468
rect -31028 36412 -30972 36468
rect -30972 36412 -30968 36468
rect -31032 36408 -30968 36412
rect -31032 36308 -30968 36312
rect -31032 36252 -31028 36308
rect -31028 36252 -30972 36308
rect -30972 36252 -30968 36308
rect -31032 36248 -30968 36252
rect -31032 36148 -30968 36152
rect -31032 36092 -31028 36148
rect -31028 36092 -30972 36148
rect -30972 36092 -30968 36148
rect -31032 36088 -30968 36092
rect -31032 35988 -30968 35992
rect -31032 35932 -31028 35988
rect -31028 35932 -30972 35988
rect -30972 35932 -30968 35988
rect -31032 35928 -30968 35932
rect -31032 35828 -30968 35832
rect -31032 35772 -31028 35828
rect -31028 35772 -30972 35828
rect -30972 35772 -30968 35828
rect -31032 35768 -30968 35772
rect -31032 35668 -30968 35672
rect -31032 35612 -31028 35668
rect -31028 35612 -30972 35668
rect -30972 35612 -30968 35668
rect -31032 35608 -30968 35612
rect -31032 35508 -30968 35512
rect -31032 35452 -31028 35508
rect -31028 35452 -30972 35508
rect -30972 35452 -30968 35508
rect -31032 35448 -30968 35452
rect -31032 35348 -30968 35352
rect -31032 35292 -31028 35348
rect -31028 35292 -30972 35348
rect -30972 35292 -30968 35348
rect -31032 35288 -30968 35292
rect -31032 35188 -30968 35192
rect -31032 35132 -31028 35188
rect -31028 35132 -30972 35188
rect -30972 35132 -30968 35188
rect -31032 35128 -30968 35132
rect -31032 35028 -30968 35032
rect -31032 34972 -31028 35028
rect -31028 34972 -30972 35028
rect -30972 34972 -30968 35028
rect -31032 34968 -30968 34972
rect -31032 34868 -30968 34872
rect -31032 34812 -31028 34868
rect -31028 34812 -30972 34868
rect -30972 34812 -30968 34868
rect -31032 34808 -30968 34812
rect -31032 34228 -30968 34232
rect -31032 34172 -31028 34228
rect -31028 34172 -30972 34228
rect -30972 34172 -30968 34228
rect -31032 34168 -30968 34172
rect -31032 34068 -30968 34072
rect -31032 34012 -31028 34068
rect -31028 34012 -30972 34068
rect -30972 34012 -30968 34068
rect -31032 34008 -30968 34012
rect -31032 33908 -30968 33912
rect -31032 33852 -31028 33908
rect -31028 33852 -30972 33908
rect -30972 33852 -30968 33908
rect -31032 33848 -30968 33852
rect -31032 33748 -30968 33752
rect -31032 33692 -31028 33748
rect -31028 33692 -30972 33748
rect -30972 33692 -30968 33748
rect -31032 33688 -30968 33692
rect -31032 33588 -30968 33592
rect -31032 33532 -31028 33588
rect -31028 33532 -30972 33588
rect -30972 33532 -30968 33588
rect -31032 33528 -30968 33532
rect -31032 33428 -30968 33432
rect -31032 33372 -31028 33428
rect -31028 33372 -30972 33428
rect -30972 33372 -30968 33428
rect -31032 33368 -30968 33372
rect -31032 33268 -30968 33272
rect -31032 33212 -31028 33268
rect -31028 33212 -30972 33268
rect -30972 33212 -30968 33268
rect -31032 33208 -30968 33212
rect -31032 33108 -30968 33112
rect -31032 33052 -31028 33108
rect -31028 33052 -30972 33108
rect -30972 33052 -30968 33108
rect -31032 33048 -30968 33052
rect -31032 32948 -30968 32952
rect -31032 32892 -31028 32948
rect -31028 32892 -30972 32948
rect -30972 32892 -30968 32948
rect -31032 32888 -30968 32892
rect -30712 37108 -30648 37112
rect -30712 37052 -30708 37108
rect -30708 37052 -30652 37108
rect -30652 37052 -30648 37108
rect -30712 37048 -30648 37052
rect -30712 36948 -30648 36952
rect -30712 36892 -30708 36948
rect -30708 36892 -30652 36948
rect -30652 36892 -30648 36948
rect -30712 36888 -30648 36892
rect -30712 36788 -30648 36792
rect -30712 36732 -30708 36788
rect -30708 36732 -30652 36788
rect -30652 36732 -30648 36788
rect -30712 36728 -30648 36732
rect -30712 36628 -30648 36632
rect -30712 36572 -30708 36628
rect -30708 36572 -30652 36628
rect -30652 36572 -30648 36628
rect -30712 36568 -30648 36572
rect -30712 36468 -30648 36472
rect -30712 36412 -30708 36468
rect -30708 36412 -30652 36468
rect -30652 36412 -30648 36468
rect -30712 36408 -30648 36412
rect -30712 36308 -30648 36312
rect -30712 36252 -30708 36308
rect -30708 36252 -30652 36308
rect -30652 36252 -30648 36308
rect -30712 36248 -30648 36252
rect -30712 36148 -30648 36152
rect -30712 36092 -30708 36148
rect -30708 36092 -30652 36148
rect -30652 36092 -30648 36148
rect -30712 36088 -30648 36092
rect -30712 35988 -30648 35992
rect -30712 35932 -30708 35988
rect -30708 35932 -30652 35988
rect -30652 35932 -30648 35988
rect -30712 35928 -30648 35932
rect -30712 35828 -30648 35832
rect -30712 35772 -30708 35828
rect -30708 35772 -30652 35828
rect -30652 35772 -30648 35828
rect -30712 35768 -30648 35772
rect -30712 35668 -30648 35672
rect -30712 35612 -30708 35668
rect -30708 35612 -30652 35668
rect -30652 35612 -30648 35668
rect -30712 35608 -30648 35612
rect -30712 35508 -30648 35512
rect -30712 35452 -30708 35508
rect -30708 35452 -30652 35508
rect -30652 35452 -30648 35508
rect -30712 35448 -30648 35452
rect -30712 35348 -30648 35352
rect -30712 35292 -30708 35348
rect -30708 35292 -30652 35348
rect -30652 35292 -30648 35348
rect -30712 35288 -30648 35292
rect -30712 35188 -30648 35192
rect -30712 35132 -30708 35188
rect -30708 35132 -30652 35188
rect -30652 35132 -30648 35188
rect -30712 35128 -30648 35132
rect -30712 35028 -30648 35032
rect -30712 34972 -30708 35028
rect -30708 34972 -30652 35028
rect -30652 34972 -30648 35028
rect -30712 34968 -30648 34972
rect -30712 34868 -30648 34872
rect -30712 34812 -30708 34868
rect -30708 34812 -30652 34868
rect -30652 34812 -30648 34868
rect -30712 34808 -30648 34812
rect -30712 34228 -30648 34232
rect -30712 34172 -30708 34228
rect -30708 34172 -30652 34228
rect -30652 34172 -30648 34228
rect -30712 34168 -30648 34172
rect -30712 34068 -30648 34072
rect -30712 34012 -30708 34068
rect -30708 34012 -30652 34068
rect -30652 34012 -30648 34068
rect -30712 34008 -30648 34012
rect -30712 33908 -30648 33912
rect -30712 33852 -30708 33908
rect -30708 33852 -30652 33908
rect -30652 33852 -30648 33908
rect -30712 33848 -30648 33852
rect -30712 33748 -30648 33752
rect -30712 33692 -30708 33748
rect -30708 33692 -30652 33748
rect -30652 33692 -30648 33748
rect -30712 33688 -30648 33692
rect -30712 33588 -30648 33592
rect -30712 33532 -30708 33588
rect -30708 33532 -30652 33588
rect -30652 33532 -30648 33588
rect -30712 33528 -30648 33532
rect -30712 33428 -30648 33432
rect -30712 33372 -30708 33428
rect -30708 33372 -30652 33428
rect -30652 33372 -30648 33428
rect -30712 33368 -30648 33372
rect -30712 33268 -30648 33272
rect -30712 33212 -30708 33268
rect -30708 33212 -30652 33268
rect -30652 33212 -30648 33268
rect -30712 33208 -30648 33212
rect -30712 33108 -30648 33112
rect -30712 33052 -30708 33108
rect -30708 33052 -30652 33108
rect -30652 33052 -30648 33108
rect -30712 33048 -30648 33052
rect -30712 32948 -30648 32952
rect -30712 32892 -30708 32948
rect -30708 32892 -30652 32948
rect -30652 32892 -30648 32948
rect -30712 32888 -30648 32892
rect -30072 41748 -30008 41752
rect -30072 41692 -30068 41748
rect -30068 41692 -30012 41748
rect -30012 41692 -30008 41748
rect -30072 41688 -30008 41692
rect -30072 41588 -30008 41592
rect -30072 41532 -30068 41588
rect -30068 41532 -30012 41588
rect -30012 41532 -30008 41588
rect -30072 41528 -30008 41532
rect -30072 40788 -30008 40792
rect -30072 40732 -30068 40788
rect -30068 40732 -30012 40788
rect -30012 40732 -30008 40788
rect -30072 40728 -30008 40732
rect -30072 40628 -30008 40632
rect -30072 40572 -30068 40628
rect -30068 40572 -30012 40628
rect -30012 40572 -30008 40628
rect -30072 40568 -30008 40572
rect -30072 40468 -30008 40472
rect -30072 40412 -30068 40468
rect -30068 40412 -30012 40468
rect -30012 40412 -30008 40468
rect -30072 40408 -30008 40412
rect -30072 40308 -30008 40312
rect -30072 40252 -30068 40308
rect -30068 40252 -30012 40308
rect -30012 40252 -30008 40308
rect -30072 40248 -30008 40252
rect -30072 40148 -30008 40152
rect -30072 40092 -30068 40148
rect -30068 40092 -30012 40148
rect -30012 40092 -30008 40148
rect -30072 40088 -30008 40092
rect -30072 39988 -30008 39992
rect -30072 39932 -30068 39988
rect -30068 39932 -30012 39988
rect -30012 39932 -30008 39988
rect -30072 39928 -30008 39932
rect -30072 39828 -30008 39832
rect -30072 39772 -30068 39828
rect -30068 39772 -30012 39828
rect -30012 39772 -30008 39828
rect -30072 39768 -30008 39772
rect -30072 39668 -30008 39672
rect -30072 39612 -30068 39668
rect -30068 39612 -30012 39668
rect -30012 39612 -30008 39668
rect -30072 39608 -30008 39612
rect -30072 39508 -30008 39512
rect -30072 39452 -30068 39508
rect -30068 39452 -30012 39508
rect -30012 39452 -30008 39508
rect -30072 39448 -30008 39452
rect -30072 39348 -30008 39352
rect -30072 39292 -30068 39348
rect -30068 39292 -30012 39348
rect -30012 39292 -30008 39348
rect -30072 39288 -30008 39292
rect -30072 39188 -30008 39192
rect -30072 39132 -30068 39188
rect -30068 39132 -30012 39188
rect -30012 39132 -30008 39188
rect -30072 39128 -30008 39132
rect -30072 39028 -30008 39032
rect -30072 38972 -30068 39028
rect -30068 38972 -30012 39028
rect -30012 38972 -30008 39028
rect -30072 38968 -30008 38972
rect -30072 38868 -30008 38872
rect -30072 38812 -30068 38868
rect -30068 38812 -30012 38868
rect -30012 38812 -30008 38868
rect -30072 38808 -30008 38812
rect -30072 38708 -30008 38712
rect -30072 38652 -30068 38708
rect -30068 38652 -30012 38708
rect -30012 38652 -30008 38708
rect -30072 38648 -30008 38652
rect -30072 38548 -30008 38552
rect -30072 38492 -30068 38548
rect -30068 38492 -30012 38548
rect -30012 38492 -30008 38548
rect -30072 38488 -30008 38492
rect -30072 38388 -30008 38392
rect -30072 38332 -30068 38388
rect -30068 38332 -30012 38388
rect -30012 38332 -30008 38388
rect -30072 38328 -30008 38332
rect -30072 38228 -30008 38232
rect -30072 38172 -30068 38228
rect -30068 38172 -30012 38228
rect -30012 38172 -30008 38228
rect -30072 38168 -30008 38172
rect -30072 38068 -30008 38072
rect -30072 38012 -30068 38068
rect -30068 38012 -30012 38068
rect -30012 38012 -30008 38068
rect -30072 38008 -30008 38012
rect -30072 37908 -30008 37912
rect -30072 37852 -30068 37908
rect -30068 37852 -30012 37908
rect -30012 37852 -30008 37908
rect -30072 37848 -30008 37852
rect -30072 37748 -30008 37752
rect -30072 37692 -30068 37748
rect -30068 37692 -30012 37748
rect -30012 37692 -30008 37748
rect -30072 37688 -30008 37692
rect -30392 37108 -30328 37112
rect -30392 37052 -30388 37108
rect -30388 37052 -30332 37108
rect -30332 37052 -30328 37108
rect -30392 37048 -30328 37052
rect -30392 36948 -30328 36952
rect -30392 36892 -30388 36948
rect -30388 36892 -30332 36948
rect -30332 36892 -30328 36948
rect -30392 36888 -30328 36892
rect -30392 36788 -30328 36792
rect -30392 36732 -30388 36788
rect -30388 36732 -30332 36788
rect -30332 36732 -30328 36788
rect -30392 36728 -30328 36732
rect -30392 36628 -30328 36632
rect -30392 36572 -30388 36628
rect -30388 36572 -30332 36628
rect -30332 36572 -30328 36628
rect -30392 36568 -30328 36572
rect -30392 36468 -30328 36472
rect -30392 36412 -30388 36468
rect -30388 36412 -30332 36468
rect -30332 36412 -30328 36468
rect -30392 36408 -30328 36412
rect -30392 36308 -30328 36312
rect -30392 36252 -30388 36308
rect -30388 36252 -30332 36308
rect -30332 36252 -30328 36308
rect -30392 36248 -30328 36252
rect -30392 36148 -30328 36152
rect -30392 36092 -30388 36148
rect -30388 36092 -30332 36148
rect -30332 36092 -30328 36148
rect -30392 36088 -30328 36092
rect -30392 35988 -30328 35992
rect -30392 35932 -30388 35988
rect -30388 35932 -30332 35988
rect -30332 35932 -30328 35988
rect -30392 35928 -30328 35932
rect -30392 35828 -30328 35832
rect -30392 35772 -30388 35828
rect -30388 35772 -30332 35828
rect -30332 35772 -30328 35828
rect -30392 35768 -30328 35772
rect -30072 37108 -30008 37112
rect -30072 37052 -30068 37108
rect -30068 37052 -30012 37108
rect -30012 37052 -30008 37108
rect -30072 37048 -30008 37052
rect -30072 36948 -30008 36952
rect -30072 36892 -30068 36948
rect -30068 36892 -30012 36948
rect -30012 36892 -30008 36948
rect -30072 36888 -30008 36892
rect -30072 36788 -30008 36792
rect -30072 36732 -30068 36788
rect -30068 36732 -30012 36788
rect -30012 36732 -30008 36788
rect -30072 36728 -30008 36732
rect -30072 36628 -30008 36632
rect -30072 36572 -30068 36628
rect -30068 36572 -30012 36628
rect -30012 36572 -30008 36628
rect -30072 36568 -30008 36572
rect -30072 36468 -30008 36472
rect -30072 36412 -30068 36468
rect -30068 36412 -30012 36468
rect -30012 36412 -30008 36468
rect -30072 36408 -30008 36412
rect -30072 36308 -30008 36312
rect -30072 36252 -30068 36308
rect -30068 36252 -30012 36308
rect -30012 36252 -30008 36308
rect -30072 36248 -30008 36252
rect -30072 36148 -30008 36152
rect -30072 36092 -30068 36148
rect -30068 36092 -30012 36148
rect -30012 36092 -30008 36148
rect -30072 36088 -30008 36092
rect -30072 35988 -30008 35992
rect -30072 35932 -30068 35988
rect -30068 35932 -30012 35988
rect -30012 35932 -30008 35988
rect -30072 35928 -30008 35932
rect -30072 35828 -30008 35832
rect -30072 35772 -30068 35828
rect -30068 35772 -30012 35828
rect -30012 35772 -30008 35828
rect -30072 35768 -30008 35772
rect -30392 35668 -30328 35672
rect -30392 35612 -30388 35668
rect -30388 35612 -30332 35668
rect -30332 35612 -30328 35668
rect -30392 35608 -30328 35612
rect -30392 35508 -30328 35512
rect -30392 35452 -30388 35508
rect -30388 35452 -30332 35508
rect -30332 35452 -30328 35508
rect -30392 35448 -30328 35452
rect -30392 35348 -30328 35352
rect -30392 35292 -30388 35348
rect -30388 35292 -30332 35348
rect -30332 35292 -30328 35348
rect -30392 35288 -30328 35292
rect -30392 35188 -30328 35192
rect -30392 35132 -30388 35188
rect -30388 35132 -30332 35188
rect -30332 35132 -30328 35188
rect -30392 35128 -30328 35132
rect -30392 35028 -30328 35032
rect -30392 34972 -30388 35028
rect -30388 34972 -30332 35028
rect -30332 34972 -30328 35028
rect -30392 34968 -30328 34972
rect -30392 34868 -30328 34872
rect -30392 34812 -30388 34868
rect -30388 34812 -30332 34868
rect -30332 34812 -30328 34868
rect -30392 34808 -30328 34812
rect -30072 35668 -30008 35672
rect -30072 35612 -30068 35668
rect -30068 35612 -30012 35668
rect -30012 35612 -30008 35668
rect -30072 35608 -30008 35612
rect -30072 35508 -30008 35512
rect -30072 35452 -30068 35508
rect -30068 35452 -30012 35508
rect -30012 35452 -30008 35508
rect -30072 35448 -30008 35452
rect -30072 35348 -30008 35352
rect -30072 35292 -30068 35348
rect -30068 35292 -30012 35348
rect -30012 35292 -30008 35348
rect -30072 35288 -30008 35292
rect -30072 35188 -30008 35192
rect -30072 35132 -30068 35188
rect -30068 35132 -30012 35188
rect -30012 35132 -30008 35188
rect -30072 35128 -30008 35132
rect -30072 35028 -30008 35032
rect -30072 34972 -30068 35028
rect -30068 34972 -30012 35028
rect -30012 34972 -30008 35028
rect -30072 34968 -30008 34972
rect -3352 39748 -3288 39752
rect -3352 39692 -3348 39748
rect -3348 39692 -3292 39748
rect -3292 39692 -3288 39748
rect -3352 39688 -3288 39692
rect -3352 39588 -3288 39592
rect -3352 39532 -3348 39588
rect -3348 39532 -3292 39588
rect -3292 39532 -3288 39588
rect -3352 39528 -3288 39532
rect -3352 39428 -3288 39432
rect -3352 39372 -3348 39428
rect -3348 39372 -3292 39428
rect -3292 39372 -3288 39428
rect -3352 39368 -3288 39372
rect -3352 39268 -3288 39272
rect -3352 39212 -3348 39268
rect -3348 39212 -3292 39268
rect -3292 39212 -3288 39268
rect -3352 39208 -3288 39212
rect -3352 39108 -3288 39112
rect -3352 39052 -3348 39108
rect -3348 39052 -3292 39108
rect -3292 39052 -3288 39108
rect -3352 39048 -3288 39052
rect -3352 38948 -3288 38952
rect -3352 38892 -3348 38948
rect -3348 38892 -3292 38948
rect -3292 38892 -3288 38948
rect -3352 38888 -3288 38892
rect -3352 38788 -3288 38792
rect -3352 38732 -3348 38788
rect -3348 38732 -3292 38788
rect -3292 38732 -3288 38788
rect -3352 38728 -3288 38732
rect -3352 38628 -3288 38632
rect -3352 38572 -3348 38628
rect -3348 38572 -3292 38628
rect -3292 38572 -3288 38628
rect -3352 38568 -3288 38572
rect -3352 38468 -3288 38472
rect -3352 38412 -3348 38468
rect -3348 38412 -3292 38468
rect -3292 38412 -3288 38468
rect -3352 38408 -3288 38412
rect -3352 38308 -3288 38312
rect -3352 38252 -3348 38308
rect -3348 38252 -3292 38308
rect -3292 38252 -3288 38308
rect -3352 38248 -3288 38252
rect -3352 38148 -3288 38152
rect -3352 38092 -3348 38148
rect -3348 38092 -3292 38148
rect -3292 38092 -3288 38148
rect -3352 38088 -3288 38092
rect -3352 37988 -3288 37992
rect -3352 37932 -3348 37988
rect -3348 37932 -3292 37988
rect -3292 37932 -3288 37988
rect -3352 37928 -3288 37932
rect -3352 37828 -3288 37832
rect -3352 37772 -3348 37828
rect -3348 37772 -3292 37828
rect -3292 37772 -3288 37828
rect -3352 37768 -3288 37772
rect -3352 37508 -3288 37512
rect -3352 37452 -3348 37508
rect -3348 37452 -3292 37508
rect -3292 37452 -3288 37508
rect -3352 37448 -3288 37452
rect -3352 37348 -3288 37352
rect -3352 37292 -3348 37348
rect -3348 37292 -3292 37348
rect -3292 37292 -3288 37348
rect -3352 37288 -3288 37292
rect -3352 37188 -3288 37192
rect -3352 37132 -3348 37188
rect -3348 37132 -3292 37188
rect -3292 37132 -3288 37188
rect -3352 37128 -3288 37132
rect -3352 37028 -3288 37032
rect -3352 36972 -3348 37028
rect -3348 36972 -3292 37028
rect -3292 36972 -3288 37028
rect -3352 36968 -3288 36972
rect -3352 36868 -3288 36872
rect -3352 36812 -3348 36868
rect -3348 36812 -3292 36868
rect -3292 36812 -3288 36868
rect -3352 36808 -3288 36812
rect -3352 36708 -3288 36712
rect -3352 36652 -3348 36708
rect -3348 36652 -3292 36708
rect -3292 36652 -3288 36708
rect -3352 36648 -3288 36652
rect -3352 36548 -3288 36552
rect -3352 36492 -3348 36548
rect -3348 36492 -3292 36548
rect -3292 36492 -3288 36548
rect -3352 36488 -3288 36492
rect -3352 36388 -3288 36392
rect -3352 36332 -3348 36388
rect -3348 36332 -3292 36388
rect -3292 36332 -3288 36388
rect -3352 36328 -3288 36332
rect -3032 39748 -2968 39752
rect -3032 39692 -3028 39748
rect -3028 39692 -2972 39748
rect -2972 39692 -2968 39748
rect -3032 39688 -2968 39692
rect -3032 39588 -2968 39592
rect -3032 39532 -3028 39588
rect -3028 39532 -2972 39588
rect -2972 39532 -2968 39588
rect -3032 39528 -2968 39532
rect -3032 39428 -2968 39432
rect -3032 39372 -3028 39428
rect -3028 39372 -2972 39428
rect -2972 39372 -2968 39428
rect -3032 39368 -2968 39372
rect -3032 39268 -2968 39272
rect -3032 39212 -3028 39268
rect -3028 39212 -2972 39268
rect -2972 39212 -2968 39268
rect -3032 39208 -2968 39212
rect -3032 39108 -2968 39112
rect -3032 39052 -3028 39108
rect -3028 39052 -2972 39108
rect -2972 39052 -2968 39108
rect -3032 39048 -2968 39052
rect -3032 38948 -2968 38952
rect -3032 38892 -3028 38948
rect -3028 38892 -2972 38948
rect -2972 38892 -2968 38948
rect -3032 38888 -2968 38892
rect -3032 38788 -2968 38792
rect -3032 38732 -3028 38788
rect -3028 38732 -2972 38788
rect -2972 38732 -2968 38788
rect -3032 38728 -2968 38732
rect -3032 38628 -2968 38632
rect -3032 38572 -3028 38628
rect -3028 38572 -2972 38628
rect -2972 38572 -2968 38628
rect -3032 38568 -2968 38572
rect -3032 38468 -2968 38472
rect -3032 38412 -3028 38468
rect -3028 38412 -2972 38468
rect -2972 38412 -2968 38468
rect -3032 38408 -2968 38412
rect -3032 38308 -2968 38312
rect -3032 38252 -3028 38308
rect -3028 38252 -2972 38308
rect -2972 38252 -2968 38308
rect -3032 38248 -2968 38252
rect -3032 38148 -2968 38152
rect -3032 38092 -3028 38148
rect -3028 38092 -2972 38148
rect -2972 38092 -2968 38148
rect -3032 38088 -2968 38092
rect -3032 37988 -2968 37992
rect -3032 37932 -3028 37988
rect -3028 37932 -2972 37988
rect -2972 37932 -2968 37988
rect -3032 37928 -2968 37932
rect -3032 37828 -2968 37832
rect -3032 37772 -3028 37828
rect -3028 37772 -2972 37828
rect -2972 37772 -2968 37828
rect -3032 37768 -2968 37772
rect -3032 37508 -2968 37512
rect -3032 37452 -3028 37508
rect -3028 37452 -2972 37508
rect -2972 37452 -2968 37508
rect -3032 37448 -2968 37452
rect -3032 37348 -2968 37352
rect -3032 37292 -3028 37348
rect -3028 37292 -2972 37348
rect -2972 37292 -2968 37348
rect -3032 37288 -2968 37292
rect -3032 37188 -2968 37192
rect -3032 37132 -3028 37188
rect -3028 37132 -2972 37188
rect -2972 37132 -2968 37188
rect -3032 37128 -2968 37132
rect -3032 37028 -2968 37032
rect -3032 36972 -3028 37028
rect -3028 36972 -2972 37028
rect -2972 36972 -2968 37028
rect -3032 36968 -2968 36972
rect -3032 36868 -2968 36872
rect -3032 36812 -3028 36868
rect -3028 36812 -2972 36868
rect -2972 36812 -2968 36868
rect -3032 36808 -2968 36812
rect -3032 36708 -2968 36712
rect -3032 36652 -3028 36708
rect -3028 36652 -2972 36708
rect -2972 36652 -2968 36708
rect -3032 36648 -2968 36652
rect -3032 36548 -2968 36552
rect -3032 36492 -3028 36548
rect -3028 36492 -2972 36548
rect -2972 36492 -2968 36548
rect -3032 36488 -2968 36492
rect -3032 36388 -2968 36392
rect -3032 36332 -3028 36388
rect -3028 36332 -2972 36388
rect -2972 36332 -2968 36388
rect -3032 36328 -2968 36332
rect -2712 39748 -2648 39752
rect -2712 39692 -2708 39748
rect -2708 39692 -2652 39748
rect -2652 39692 -2648 39748
rect -2712 39688 -2648 39692
rect -2712 39588 -2648 39592
rect -2712 39532 -2708 39588
rect -2708 39532 -2652 39588
rect -2652 39532 -2648 39588
rect -2712 39528 -2648 39532
rect -2712 39428 -2648 39432
rect -2712 39372 -2708 39428
rect -2708 39372 -2652 39428
rect -2652 39372 -2648 39428
rect -2712 39368 -2648 39372
rect -2712 39268 -2648 39272
rect -2712 39212 -2708 39268
rect -2708 39212 -2652 39268
rect -2652 39212 -2648 39268
rect -2712 39208 -2648 39212
rect -2712 39108 -2648 39112
rect -2712 39052 -2708 39108
rect -2708 39052 -2652 39108
rect -2652 39052 -2648 39108
rect -2712 39048 -2648 39052
rect -2712 38948 -2648 38952
rect -2712 38892 -2708 38948
rect -2708 38892 -2652 38948
rect -2652 38892 -2648 38948
rect -2712 38888 -2648 38892
rect -2712 38788 -2648 38792
rect -2712 38732 -2708 38788
rect -2708 38732 -2652 38788
rect -2652 38732 -2648 38788
rect -2712 38728 -2648 38732
rect -2712 38628 -2648 38632
rect -2712 38572 -2708 38628
rect -2708 38572 -2652 38628
rect -2652 38572 -2648 38628
rect -2712 38568 -2648 38572
rect -2712 38468 -2648 38472
rect -2712 38412 -2708 38468
rect -2708 38412 -2652 38468
rect -2652 38412 -2648 38468
rect -2712 38408 -2648 38412
rect -2712 38308 -2648 38312
rect -2712 38252 -2708 38308
rect -2708 38252 -2652 38308
rect -2652 38252 -2648 38308
rect -2712 38248 -2648 38252
rect -2712 38148 -2648 38152
rect -2712 38092 -2708 38148
rect -2708 38092 -2652 38148
rect -2652 38092 -2648 38148
rect -2712 38088 -2648 38092
rect -2712 37988 -2648 37992
rect -2712 37932 -2708 37988
rect -2708 37932 -2652 37988
rect -2652 37932 -2648 37988
rect -2712 37928 -2648 37932
rect -2712 37828 -2648 37832
rect -2712 37772 -2708 37828
rect -2708 37772 -2652 37828
rect -2652 37772 -2648 37828
rect -2712 37768 -2648 37772
rect -2712 37508 -2648 37512
rect -2712 37452 -2708 37508
rect -2708 37452 -2652 37508
rect -2652 37452 -2648 37508
rect -2712 37448 -2648 37452
rect -2712 37348 -2648 37352
rect -2712 37292 -2708 37348
rect -2708 37292 -2652 37348
rect -2652 37292 -2648 37348
rect -2712 37288 -2648 37292
rect -2712 37188 -2648 37192
rect -2712 37132 -2708 37188
rect -2708 37132 -2652 37188
rect -2652 37132 -2648 37188
rect -2712 37128 -2648 37132
rect -2712 37028 -2648 37032
rect -2712 36972 -2708 37028
rect -2708 36972 -2652 37028
rect -2652 36972 -2648 37028
rect -2712 36968 -2648 36972
rect -2712 36868 -2648 36872
rect -2712 36812 -2708 36868
rect -2708 36812 -2652 36868
rect -2652 36812 -2648 36868
rect -2712 36808 -2648 36812
rect -2712 36708 -2648 36712
rect -2712 36652 -2708 36708
rect -2708 36652 -2652 36708
rect -2652 36652 -2648 36708
rect -2712 36648 -2648 36652
rect -2712 36548 -2648 36552
rect -2712 36492 -2708 36548
rect -2708 36492 -2652 36548
rect -2652 36492 -2648 36548
rect -2712 36488 -2648 36492
rect -2712 36388 -2648 36392
rect -2712 36332 -2708 36388
rect -2708 36332 -2652 36388
rect -2652 36332 -2648 36388
rect -2712 36328 -2648 36332
rect -3352 35748 -3288 35752
rect -3352 35692 -3348 35748
rect -3348 35692 -3292 35748
rect -3292 35692 -3288 35748
rect -3352 35688 -3288 35692
rect -3352 35588 -3288 35592
rect -3352 35532 -3348 35588
rect -3348 35532 -3292 35588
rect -3292 35532 -3288 35588
rect -3352 35528 -3288 35532
rect -3352 35428 -3288 35432
rect -3352 35372 -3348 35428
rect -3348 35372 -3292 35428
rect -3292 35372 -3288 35428
rect -3352 35368 -3288 35372
rect -3352 35268 -3288 35272
rect -3352 35212 -3348 35268
rect -3348 35212 -3292 35268
rect -3292 35212 -3288 35268
rect -3352 35208 -3288 35212
rect -3352 35108 -3288 35112
rect -3352 35052 -3348 35108
rect -3348 35052 -3292 35108
rect -3292 35052 -3288 35108
rect -3352 35048 -3288 35052
rect -3352 34948 -3288 34952
rect -3352 34892 -3348 34948
rect -3348 34892 -3292 34948
rect -3292 34892 -3288 34948
rect -3352 34888 -3288 34892
rect -30072 34868 -30008 34872
rect -30072 34812 -30068 34868
rect -30068 34812 -30012 34868
rect -30012 34812 -30008 34868
rect -30072 34808 -30008 34812
rect -30392 34228 -30328 34232
rect -30392 34172 -30388 34228
rect -30388 34172 -30332 34228
rect -30332 34172 -30328 34228
rect -30392 34168 -30328 34172
rect -30392 34068 -30328 34072
rect -30392 34012 -30388 34068
rect -30388 34012 -30332 34068
rect -30332 34012 -30328 34068
rect -30392 34008 -30328 34012
rect -30392 33908 -30328 33912
rect -30392 33852 -30388 33908
rect -30388 33852 -30332 33908
rect -30332 33852 -30328 33908
rect -30392 33848 -30328 33852
rect -30392 33748 -30328 33752
rect -30392 33692 -30388 33748
rect -30388 33692 -30332 33748
rect -30332 33692 -30328 33748
rect -30392 33688 -30328 33692
rect -30392 33588 -30328 33592
rect -30392 33532 -30388 33588
rect -30388 33532 -30332 33588
rect -30332 33532 -30328 33588
rect -30392 33528 -30328 33532
rect -30392 33428 -30328 33432
rect -30392 33372 -30388 33428
rect -30388 33372 -30332 33428
rect -30332 33372 -30328 33428
rect -30392 33368 -30328 33372
rect -30392 33268 -30328 33272
rect -30392 33212 -30388 33268
rect -30388 33212 -30332 33268
rect -30332 33212 -30328 33268
rect -30392 33208 -30328 33212
rect -30392 33108 -30328 33112
rect -30392 33052 -30388 33108
rect -30388 33052 -30332 33108
rect -30332 33052 -30328 33108
rect -30392 33048 -30328 33052
rect -30392 32948 -30328 32952
rect -30392 32892 -30388 32948
rect -30388 32892 -30332 32948
rect -30332 32892 -30328 32948
rect -30392 32888 -30328 32892
rect -30072 34228 -30008 34232
rect -30072 34172 -30068 34228
rect -30068 34172 -30012 34228
rect -30012 34172 -30008 34228
rect -30072 34168 -30008 34172
rect -30072 34068 -30008 34072
rect -30072 34012 -30068 34068
rect -30068 34012 -30012 34068
rect -30012 34012 -30008 34068
rect -30072 34008 -30008 34012
rect -30072 33908 -30008 33912
rect -30072 33852 -30068 33908
rect -30068 33852 -30012 33908
rect -30012 33852 -30008 33908
rect -30072 33848 -30008 33852
rect -30072 33748 -30008 33752
rect -30072 33692 -30068 33748
rect -30068 33692 -30012 33748
rect -30012 33692 -30008 33748
rect -30072 33688 -30008 33692
rect -30072 33588 -30008 33592
rect -30072 33532 -30068 33588
rect -30068 33532 -30012 33588
rect -30012 33532 -30008 33588
rect -30072 33528 -30008 33532
rect -30072 33428 -30008 33432
rect -30072 33372 -30068 33428
rect -30068 33372 -30012 33428
rect -30012 33372 -30008 33428
rect -30072 33368 -30008 33372
rect -30072 33268 -30008 33272
rect -30072 33212 -30068 33268
rect -30068 33212 -30012 33268
rect -30012 33212 -30008 33268
rect -30072 33208 -30008 33212
rect -30072 33108 -30008 33112
rect -30072 33052 -30068 33108
rect -30068 33052 -30012 33108
rect -30012 33052 -30008 33108
rect -30072 33048 -30008 33052
rect -30072 32948 -30008 32952
rect -30072 32892 -30068 32948
rect -30068 32892 -30012 32948
rect -30012 32892 -30008 32948
rect -30072 32888 -30008 32892
rect -3352 34788 -3288 34792
rect -3352 34732 -3348 34788
rect -3348 34732 -3292 34788
rect -3292 34732 -3288 34788
rect -3352 34728 -3288 34732
rect -3352 34628 -3288 34632
rect -3352 34572 -3348 34628
rect -3348 34572 -3292 34628
rect -3292 34572 -3288 34628
rect -3352 34568 -3288 34572
rect -3352 34468 -3288 34472
rect -3352 34412 -3348 34468
rect -3348 34412 -3292 34468
rect -3292 34412 -3288 34468
rect -3352 34408 -3288 34412
rect -3352 34308 -3288 34312
rect -3352 34252 -3348 34308
rect -3348 34252 -3292 34308
rect -3292 34252 -3288 34308
rect -3352 34248 -3288 34252
rect -3352 34148 -3288 34152
rect -3352 34092 -3348 34148
rect -3348 34092 -3292 34148
rect -3292 34092 -3288 34148
rect -3352 34088 -3288 34092
rect -3352 33988 -3288 33992
rect -3352 33932 -3348 33988
rect -3348 33932 -3292 33988
rect -3292 33932 -3288 33988
rect -3352 33928 -3288 33932
rect -3352 33828 -3288 33832
rect -3352 33772 -3348 33828
rect -3348 33772 -3292 33828
rect -3292 33772 -3288 33828
rect -3352 33768 -3288 33772
rect -3352 33668 -3288 33672
rect -3352 33612 -3348 33668
rect -3348 33612 -3292 33668
rect -3292 33612 -3288 33668
rect -3352 33608 -3288 33612
rect -3352 33508 -3288 33512
rect -3352 33452 -3348 33508
rect -3348 33452 -3292 33508
rect -3292 33452 -3288 33508
rect -3352 33448 -3288 33452
rect -3352 33268 -3288 33272
rect -3352 33212 -3348 33268
rect -3348 33212 -3292 33268
rect -3292 33212 -3288 33268
rect -3352 33208 -3288 33212
rect -3352 33108 -3288 33112
rect -3352 33052 -3348 33108
rect -3348 33052 -3292 33108
rect -3292 33052 -3288 33108
rect -3352 33048 -3288 33052
rect -3032 35748 -2968 35752
rect -3032 35692 -3028 35748
rect -3028 35692 -2972 35748
rect -2972 35692 -2968 35748
rect -3032 35688 -2968 35692
rect -3032 35588 -2968 35592
rect -3032 35532 -3028 35588
rect -3028 35532 -2972 35588
rect -2972 35532 -2968 35588
rect -3032 35528 -2968 35532
rect -3032 35428 -2968 35432
rect -3032 35372 -3028 35428
rect -3028 35372 -2972 35428
rect -2972 35372 -2968 35428
rect -3032 35368 -2968 35372
rect -3032 35268 -2968 35272
rect -3032 35212 -3028 35268
rect -3028 35212 -2972 35268
rect -2972 35212 -2968 35268
rect -3032 35208 -2968 35212
rect -3032 35108 -2968 35112
rect -3032 35052 -3028 35108
rect -3028 35052 -2972 35108
rect -2972 35052 -2968 35108
rect -3032 35048 -2968 35052
rect -3032 34948 -2968 34952
rect -3032 34892 -3028 34948
rect -3028 34892 -2972 34948
rect -2972 34892 -2968 34948
rect -3032 34888 -2968 34892
rect -3032 34788 -2968 34792
rect -3032 34732 -3028 34788
rect -3028 34732 -2972 34788
rect -2972 34732 -2968 34788
rect -3032 34728 -2968 34732
rect -3032 34628 -2968 34632
rect -3032 34572 -3028 34628
rect -3028 34572 -2972 34628
rect -2972 34572 -2968 34628
rect -3032 34568 -2968 34572
rect -3032 34468 -2968 34472
rect -3032 34412 -3028 34468
rect -3028 34412 -2972 34468
rect -2972 34412 -2968 34468
rect -3032 34408 -2968 34412
rect -3032 34308 -2968 34312
rect -3032 34252 -3028 34308
rect -3028 34252 -2972 34308
rect -2972 34252 -2968 34308
rect -3032 34248 -2968 34252
rect -3032 34148 -2968 34152
rect -3032 34092 -3028 34148
rect -3028 34092 -2972 34148
rect -2972 34092 -2968 34148
rect -3032 34088 -2968 34092
rect -3032 33988 -2968 33992
rect -3032 33932 -3028 33988
rect -3028 33932 -2972 33988
rect -2972 33932 -2968 33988
rect -3032 33928 -2968 33932
rect -3032 33828 -2968 33832
rect -3032 33772 -3028 33828
rect -3028 33772 -2972 33828
rect -2972 33772 -2968 33828
rect -3032 33768 -2968 33772
rect -3032 33668 -2968 33672
rect -3032 33612 -3028 33668
rect -3028 33612 -2972 33668
rect -2972 33612 -2968 33668
rect -3032 33608 -2968 33612
rect -3032 33508 -2968 33512
rect -3032 33452 -3028 33508
rect -3028 33452 -2972 33508
rect -2972 33452 -2968 33508
rect -3032 33448 -2968 33452
rect -3032 33268 -2968 33272
rect -3032 33212 -3028 33268
rect -3028 33212 -2972 33268
rect -2972 33212 -2968 33268
rect -3032 33208 -2968 33212
rect -3032 33108 -2968 33112
rect -3032 33052 -3028 33108
rect -3028 33052 -2972 33108
rect -2972 33052 -2968 33108
rect -3032 33048 -2968 33052
rect -2712 35748 -2648 35752
rect -2712 35692 -2708 35748
rect -2708 35692 -2652 35748
rect -2652 35692 -2648 35748
rect -2712 35688 -2648 35692
rect -2712 35588 -2648 35592
rect -2712 35532 -2708 35588
rect -2708 35532 -2652 35588
rect -2652 35532 -2648 35588
rect -2712 35528 -2648 35532
rect -2712 35428 -2648 35432
rect -2712 35372 -2708 35428
rect -2708 35372 -2652 35428
rect -2652 35372 -2648 35428
rect -2712 35368 -2648 35372
rect -2712 35268 -2648 35272
rect -2712 35212 -2708 35268
rect -2708 35212 -2652 35268
rect -2652 35212 -2648 35268
rect -2712 35208 -2648 35212
rect -2712 35108 -2648 35112
rect -2712 35052 -2708 35108
rect -2708 35052 -2652 35108
rect -2652 35052 -2648 35108
rect -2712 35048 -2648 35052
rect -2712 34948 -2648 34952
rect -2712 34892 -2708 34948
rect -2708 34892 -2652 34948
rect -2652 34892 -2648 34948
rect -2712 34888 -2648 34892
rect -2712 34788 -2648 34792
rect -2712 34732 -2708 34788
rect -2708 34732 -2652 34788
rect -2652 34732 -2648 34788
rect -2712 34728 -2648 34732
rect -2712 34628 -2648 34632
rect -2712 34572 -2708 34628
rect -2708 34572 -2652 34628
rect -2652 34572 -2648 34628
rect -2712 34568 -2648 34572
rect -2712 34468 -2648 34472
rect -2712 34412 -2708 34468
rect -2708 34412 -2652 34468
rect -2652 34412 -2648 34468
rect -2712 34408 -2648 34412
rect -2712 34308 -2648 34312
rect -2712 34252 -2708 34308
rect -2708 34252 -2652 34308
rect -2652 34252 -2648 34308
rect -2712 34248 -2648 34252
rect -2712 34148 -2648 34152
rect -2712 34092 -2708 34148
rect -2708 34092 -2652 34148
rect -2652 34092 -2648 34148
rect -2712 34088 -2648 34092
rect -2712 33988 -2648 33992
rect -2712 33932 -2708 33988
rect -2708 33932 -2652 33988
rect -2652 33932 -2648 33988
rect -2712 33928 -2648 33932
rect -2712 33828 -2648 33832
rect -2712 33772 -2708 33828
rect -2708 33772 -2652 33828
rect -2652 33772 -2648 33828
rect -2712 33768 -2648 33772
rect -2712 33668 -2648 33672
rect -2712 33612 -2708 33668
rect -2708 33612 -2652 33668
rect -2652 33612 -2648 33668
rect -2712 33608 -2648 33612
rect -2712 33508 -2648 33512
rect -2712 33452 -2708 33508
rect -2708 33452 -2652 33508
rect -2652 33452 -2648 33508
rect -2712 33448 -2648 33452
rect -2712 33268 -2648 33272
rect -2712 33212 -2708 33268
rect -2708 33212 -2652 33268
rect -2652 33212 -2648 33268
rect -2712 33208 -2648 33212
rect -2712 33108 -2648 33112
rect -2712 33052 -2708 33108
rect -2708 33052 -2652 33108
rect -2652 33052 -2648 33108
rect -2712 33048 -2648 33052
rect -2392 39748 -2328 39752
rect -2392 39692 -2388 39748
rect -2388 39692 -2332 39748
rect -2332 39692 -2328 39748
rect -2392 39688 -2328 39692
rect -2392 39588 -2328 39592
rect -2392 39532 -2388 39588
rect -2388 39532 -2332 39588
rect -2332 39532 -2328 39588
rect -2392 39528 -2328 39532
rect -2392 39428 -2328 39432
rect -2392 39372 -2388 39428
rect -2388 39372 -2332 39428
rect -2332 39372 -2328 39428
rect -2392 39368 -2328 39372
rect -2392 39268 -2328 39272
rect -2392 39212 -2388 39268
rect -2388 39212 -2332 39268
rect -2332 39212 -2328 39268
rect -2392 39208 -2328 39212
rect -2392 39108 -2328 39112
rect -2392 39052 -2388 39108
rect -2388 39052 -2332 39108
rect -2332 39052 -2328 39108
rect -2392 39048 -2328 39052
rect -2392 38948 -2328 38952
rect -2392 38892 -2388 38948
rect -2388 38892 -2332 38948
rect -2332 38892 -2328 38948
rect -2392 38888 -2328 38892
rect -2392 38788 -2328 38792
rect -2392 38732 -2388 38788
rect -2388 38732 -2332 38788
rect -2332 38732 -2328 38788
rect -2392 38728 -2328 38732
rect -2392 38628 -2328 38632
rect -2392 38572 -2388 38628
rect -2388 38572 -2332 38628
rect -2332 38572 -2328 38628
rect -2392 38568 -2328 38572
rect -2392 38468 -2328 38472
rect -2392 38412 -2388 38468
rect -2388 38412 -2332 38468
rect -2332 38412 -2328 38468
rect -2392 38408 -2328 38412
rect -2392 38308 -2328 38312
rect -2392 38252 -2388 38308
rect -2388 38252 -2332 38308
rect -2332 38252 -2328 38308
rect -2392 38248 -2328 38252
rect -2392 38148 -2328 38152
rect -2392 38092 -2388 38148
rect -2388 38092 -2332 38148
rect -2332 38092 -2328 38148
rect -2392 38088 -2328 38092
rect -2392 37988 -2328 37992
rect -2392 37932 -2388 37988
rect -2388 37932 -2332 37988
rect -2332 37932 -2328 37988
rect -2392 37928 -2328 37932
rect -2392 37828 -2328 37832
rect -2392 37772 -2388 37828
rect -2388 37772 -2332 37828
rect -2332 37772 -2328 37828
rect -2392 37768 -2328 37772
rect -2392 37508 -2328 37512
rect -2392 37452 -2388 37508
rect -2388 37452 -2332 37508
rect -2332 37452 -2328 37508
rect -2392 37448 -2328 37452
rect -2392 37348 -2328 37352
rect -2392 37292 -2388 37348
rect -2388 37292 -2332 37348
rect -2332 37292 -2328 37348
rect -2392 37288 -2328 37292
rect -2392 37188 -2328 37192
rect -2392 37132 -2388 37188
rect -2388 37132 -2332 37188
rect -2332 37132 -2328 37188
rect -2392 37128 -2328 37132
rect -2392 37028 -2328 37032
rect -2392 36972 -2388 37028
rect -2388 36972 -2332 37028
rect -2332 36972 -2328 37028
rect -2392 36968 -2328 36972
rect -2392 36868 -2328 36872
rect -2392 36812 -2388 36868
rect -2388 36812 -2332 36868
rect -2332 36812 -2328 36868
rect -2392 36808 -2328 36812
rect -2392 36708 -2328 36712
rect -2392 36652 -2388 36708
rect -2388 36652 -2332 36708
rect -2332 36652 -2328 36708
rect -2392 36648 -2328 36652
rect -2392 36548 -2328 36552
rect -2392 36492 -2388 36548
rect -2388 36492 -2332 36548
rect -2332 36492 -2328 36548
rect -2392 36488 -2328 36492
rect -2392 36388 -2328 36392
rect -2392 36332 -2388 36388
rect -2388 36332 -2332 36388
rect -2332 36332 -2328 36388
rect -2392 36328 -2328 36332
rect -2392 35748 -2328 35752
rect -2392 35692 -2388 35748
rect -2388 35692 -2332 35748
rect -2332 35692 -2328 35748
rect -2392 35688 -2328 35692
rect -2392 35588 -2328 35592
rect -2392 35532 -2388 35588
rect -2388 35532 -2332 35588
rect -2332 35532 -2328 35588
rect -2392 35528 -2328 35532
rect -2392 35428 -2328 35432
rect -2392 35372 -2388 35428
rect -2388 35372 -2332 35428
rect -2332 35372 -2328 35428
rect -2392 35368 -2328 35372
rect -2392 35268 -2328 35272
rect -2392 35212 -2388 35268
rect -2388 35212 -2332 35268
rect -2332 35212 -2328 35268
rect -2392 35208 -2328 35212
rect -2392 35108 -2328 35112
rect -2392 35052 -2388 35108
rect -2388 35052 -2332 35108
rect -2332 35052 -2328 35108
rect -2392 35048 -2328 35052
rect -2392 34948 -2328 34952
rect -2392 34892 -2388 34948
rect -2388 34892 -2332 34948
rect -2332 34892 -2328 34948
rect -2392 34888 -2328 34892
rect -2392 34788 -2328 34792
rect -2392 34732 -2388 34788
rect -2388 34732 -2332 34788
rect -2332 34732 -2328 34788
rect -2392 34728 -2328 34732
rect -2392 34628 -2328 34632
rect -2392 34572 -2388 34628
rect -2388 34572 -2332 34628
rect -2332 34572 -2328 34628
rect -2392 34568 -2328 34572
rect -2392 34468 -2328 34472
rect -2392 34412 -2388 34468
rect -2388 34412 -2332 34468
rect -2332 34412 -2328 34468
rect -2392 34408 -2328 34412
rect -2392 34308 -2328 34312
rect -2392 34252 -2388 34308
rect -2388 34252 -2332 34308
rect -2332 34252 -2328 34308
rect -2392 34248 -2328 34252
rect -2392 34148 -2328 34152
rect -2392 34092 -2388 34148
rect -2388 34092 -2332 34148
rect -2332 34092 -2328 34148
rect -2392 34088 -2328 34092
rect -2392 33988 -2328 33992
rect -2392 33932 -2388 33988
rect -2388 33932 -2332 33988
rect -2332 33932 -2328 33988
rect -2392 33928 -2328 33932
rect -2392 33828 -2328 33832
rect -2392 33772 -2388 33828
rect -2388 33772 -2332 33828
rect -2332 33772 -2328 33828
rect -2392 33768 -2328 33772
rect -2392 33668 -2328 33672
rect -2392 33612 -2388 33668
rect -2388 33612 -2332 33668
rect -2332 33612 -2328 33668
rect -2392 33608 -2328 33612
rect -2392 33508 -2328 33512
rect -2392 33452 -2388 33508
rect -2388 33452 -2332 33508
rect -2332 33452 -2328 33508
rect -2392 33448 -2328 33452
rect -2392 33268 -2328 33272
rect -2392 33212 -2388 33268
rect -2388 33212 -2332 33268
rect -2332 33212 -2328 33268
rect -2392 33208 -2328 33212
rect -2392 33108 -2328 33112
rect -2392 33052 -2388 33108
rect -2388 33052 -2332 33108
rect -2332 33052 -2328 33108
rect -2392 33048 -2328 33052
rect -2072 39748 -2008 39752
rect -2072 39692 -2068 39748
rect -2068 39692 -2012 39748
rect -2012 39692 -2008 39748
rect -2072 39688 -2008 39692
rect -2072 39588 -2008 39592
rect -2072 39532 -2068 39588
rect -2068 39532 -2012 39588
rect -2012 39532 -2008 39588
rect -2072 39528 -2008 39532
rect -2072 39428 -2008 39432
rect -2072 39372 -2068 39428
rect -2068 39372 -2012 39428
rect -2012 39372 -2008 39428
rect -2072 39368 -2008 39372
rect -2072 39268 -2008 39272
rect -2072 39212 -2068 39268
rect -2068 39212 -2012 39268
rect -2012 39212 -2008 39268
rect -2072 39208 -2008 39212
rect -2072 39108 -2008 39112
rect -2072 39052 -2068 39108
rect -2068 39052 -2012 39108
rect -2012 39052 -2008 39108
rect -2072 39048 -2008 39052
rect -2072 38948 -2008 38952
rect -2072 38892 -2068 38948
rect -2068 38892 -2012 38948
rect -2012 38892 -2008 38948
rect -2072 38888 -2008 38892
rect -2072 38788 -2008 38792
rect -2072 38732 -2068 38788
rect -2068 38732 -2012 38788
rect -2012 38732 -2008 38788
rect -2072 38728 -2008 38732
rect -2072 38628 -2008 38632
rect -2072 38572 -2068 38628
rect -2068 38572 -2012 38628
rect -2012 38572 -2008 38628
rect -2072 38568 -2008 38572
rect -2072 38468 -2008 38472
rect -2072 38412 -2068 38468
rect -2068 38412 -2012 38468
rect -2012 38412 -2008 38468
rect -2072 38408 -2008 38412
rect -2072 38308 -2008 38312
rect -2072 38252 -2068 38308
rect -2068 38252 -2012 38308
rect -2012 38252 -2008 38308
rect -2072 38248 -2008 38252
rect -2072 38148 -2008 38152
rect -2072 38092 -2068 38148
rect -2068 38092 -2012 38148
rect -2012 38092 -2008 38148
rect -2072 38088 -2008 38092
rect -2072 37988 -2008 37992
rect -2072 37932 -2068 37988
rect -2068 37932 -2012 37988
rect -2012 37932 -2008 37988
rect -2072 37928 -2008 37932
rect -2072 37828 -2008 37832
rect -2072 37772 -2068 37828
rect -2068 37772 -2012 37828
rect -2012 37772 -2008 37828
rect -2072 37768 -2008 37772
rect -2072 37508 -2008 37512
rect -2072 37452 -2068 37508
rect -2068 37452 -2012 37508
rect -2012 37452 -2008 37508
rect -2072 37448 -2008 37452
rect -2072 37348 -2008 37352
rect -2072 37292 -2068 37348
rect -2068 37292 -2012 37348
rect -2012 37292 -2008 37348
rect -2072 37288 -2008 37292
rect -2072 37188 -2008 37192
rect -2072 37132 -2068 37188
rect -2068 37132 -2012 37188
rect -2012 37132 -2008 37188
rect -2072 37128 -2008 37132
rect -2072 37028 -2008 37032
rect -2072 36972 -2068 37028
rect -2068 36972 -2012 37028
rect -2012 36972 -2008 37028
rect -2072 36968 -2008 36972
rect -2072 36868 -2008 36872
rect -2072 36812 -2068 36868
rect -2068 36812 -2012 36868
rect -2012 36812 -2008 36868
rect -2072 36808 -2008 36812
rect -2072 36708 -2008 36712
rect -2072 36652 -2068 36708
rect -2068 36652 -2012 36708
rect -2012 36652 -2008 36708
rect -2072 36648 -2008 36652
rect -2072 36548 -2008 36552
rect -2072 36492 -2068 36548
rect -2068 36492 -2012 36548
rect -2012 36492 -2008 36548
rect -2072 36488 -2008 36492
rect -2072 36388 -2008 36392
rect -2072 36332 -2068 36388
rect -2068 36332 -2012 36388
rect -2012 36332 -2008 36388
rect -2072 36328 -2008 36332
rect -1752 39748 -1688 39752
rect -1752 39692 -1748 39748
rect -1748 39692 -1692 39748
rect -1692 39692 -1688 39748
rect -1752 39688 -1688 39692
rect -1752 39588 -1688 39592
rect -1752 39532 -1748 39588
rect -1748 39532 -1692 39588
rect -1692 39532 -1688 39588
rect -1752 39528 -1688 39532
rect -1752 39428 -1688 39432
rect -1752 39372 -1748 39428
rect -1748 39372 -1692 39428
rect -1692 39372 -1688 39428
rect -1752 39368 -1688 39372
rect -1752 39268 -1688 39272
rect -1752 39212 -1748 39268
rect -1748 39212 -1692 39268
rect -1692 39212 -1688 39268
rect -1752 39208 -1688 39212
rect -1752 39108 -1688 39112
rect -1752 39052 -1748 39108
rect -1748 39052 -1692 39108
rect -1692 39052 -1688 39108
rect -1752 39048 -1688 39052
rect -1752 38948 -1688 38952
rect -1752 38892 -1748 38948
rect -1748 38892 -1692 38948
rect -1692 38892 -1688 38948
rect -1752 38888 -1688 38892
rect -1752 38788 -1688 38792
rect -1752 38732 -1748 38788
rect -1748 38732 -1692 38788
rect -1692 38732 -1688 38788
rect -1752 38728 -1688 38732
rect -1752 38628 -1688 38632
rect -1752 38572 -1748 38628
rect -1748 38572 -1692 38628
rect -1692 38572 -1688 38628
rect -1752 38568 -1688 38572
rect -1752 38468 -1688 38472
rect -1752 38412 -1748 38468
rect -1748 38412 -1692 38468
rect -1692 38412 -1688 38468
rect -1752 38408 -1688 38412
rect -1752 38308 -1688 38312
rect -1752 38252 -1748 38308
rect -1748 38252 -1692 38308
rect -1692 38252 -1688 38308
rect -1752 38248 -1688 38252
rect -1752 38148 -1688 38152
rect -1752 38092 -1748 38148
rect -1748 38092 -1692 38148
rect -1692 38092 -1688 38148
rect -1752 38088 -1688 38092
rect -1752 37988 -1688 37992
rect -1752 37932 -1748 37988
rect -1748 37932 -1692 37988
rect -1692 37932 -1688 37988
rect -1752 37928 -1688 37932
rect -1752 37828 -1688 37832
rect -1752 37772 -1748 37828
rect -1748 37772 -1692 37828
rect -1692 37772 -1688 37828
rect -1752 37768 -1688 37772
rect -1752 37508 -1688 37512
rect -1752 37452 -1748 37508
rect -1748 37452 -1692 37508
rect -1692 37452 -1688 37508
rect -1752 37448 -1688 37452
rect -1752 37348 -1688 37352
rect -1752 37292 -1748 37348
rect -1748 37292 -1692 37348
rect -1692 37292 -1688 37348
rect -1752 37288 -1688 37292
rect -1752 37188 -1688 37192
rect -1752 37132 -1748 37188
rect -1748 37132 -1692 37188
rect -1692 37132 -1688 37188
rect -1752 37128 -1688 37132
rect -1752 37028 -1688 37032
rect -1752 36972 -1748 37028
rect -1748 36972 -1692 37028
rect -1692 36972 -1688 37028
rect -1752 36968 -1688 36972
rect -1752 36868 -1688 36872
rect -1752 36812 -1748 36868
rect -1748 36812 -1692 36868
rect -1692 36812 -1688 36868
rect -1752 36808 -1688 36812
rect -1752 36708 -1688 36712
rect -1752 36652 -1748 36708
rect -1748 36652 -1692 36708
rect -1692 36652 -1688 36708
rect -1752 36648 -1688 36652
rect -1752 36548 -1688 36552
rect -1752 36492 -1748 36548
rect -1748 36492 -1692 36548
rect -1692 36492 -1688 36548
rect -1752 36488 -1688 36492
rect -1752 36388 -1688 36392
rect -1752 36332 -1748 36388
rect -1748 36332 -1692 36388
rect -1692 36332 -1688 36388
rect -1752 36328 -1688 36332
rect -2072 35748 -2008 35752
rect -2072 35692 -2068 35748
rect -2068 35692 -2012 35748
rect -2012 35692 -2008 35748
rect -2072 35688 -2008 35692
rect -2072 35588 -2008 35592
rect -2072 35532 -2068 35588
rect -2068 35532 -2012 35588
rect -2012 35532 -2008 35588
rect -2072 35528 -2008 35532
rect -2072 35428 -2008 35432
rect -2072 35372 -2068 35428
rect -2068 35372 -2012 35428
rect -2012 35372 -2008 35428
rect -2072 35368 -2008 35372
rect -2072 35268 -2008 35272
rect -2072 35212 -2068 35268
rect -2068 35212 -2012 35268
rect -2012 35212 -2008 35268
rect -2072 35208 -2008 35212
rect -2072 35108 -2008 35112
rect -2072 35052 -2068 35108
rect -2068 35052 -2012 35108
rect -2012 35052 -2008 35108
rect -2072 35048 -2008 35052
rect -2072 34948 -2008 34952
rect -2072 34892 -2068 34948
rect -2068 34892 -2012 34948
rect -2012 34892 -2008 34948
rect -2072 34888 -2008 34892
rect -2072 34788 -2008 34792
rect -2072 34732 -2068 34788
rect -2068 34732 -2012 34788
rect -2012 34732 -2008 34788
rect -2072 34728 -2008 34732
rect -2072 34628 -2008 34632
rect -2072 34572 -2068 34628
rect -2068 34572 -2012 34628
rect -2012 34572 -2008 34628
rect -2072 34568 -2008 34572
rect -2072 34468 -2008 34472
rect -2072 34412 -2068 34468
rect -2068 34412 -2012 34468
rect -2012 34412 -2008 34468
rect -2072 34408 -2008 34412
rect -2072 34308 -2008 34312
rect -2072 34252 -2068 34308
rect -2068 34252 -2012 34308
rect -2012 34252 -2008 34308
rect -2072 34248 -2008 34252
rect -2072 34148 -2008 34152
rect -2072 34092 -2068 34148
rect -2068 34092 -2012 34148
rect -2012 34092 -2008 34148
rect -2072 34088 -2008 34092
rect -2072 33988 -2008 33992
rect -2072 33932 -2068 33988
rect -2068 33932 -2012 33988
rect -2012 33932 -2008 33988
rect -2072 33928 -2008 33932
rect -2072 33828 -2008 33832
rect -2072 33772 -2068 33828
rect -2068 33772 -2012 33828
rect -2012 33772 -2008 33828
rect -2072 33768 -2008 33772
rect -2072 33668 -2008 33672
rect -2072 33612 -2068 33668
rect -2068 33612 -2012 33668
rect -2012 33612 -2008 33668
rect -2072 33608 -2008 33612
rect -2072 33508 -2008 33512
rect -2072 33452 -2068 33508
rect -2068 33452 -2012 33508
rect -2012 33452 -2008 33508
rect -2072 33448 -2008 33452
rect -2072 33268 -2008 33272
rect -2072 33212 -2068 33268
rect -2068 33212 -2012 33268
rect -2012 33212 -2008 33268
rect -2072 33208 -2008 33212
rect -2072 33108 -2008 33112
rect -2072 33052 -2068 33108
rect -2068 33052 -2012 33108
rect -2012 33052 -2008 33108
rect -2072 33048 -2008 33052
rect -1432 39748 -1368 39752
rect -1432 39692 -1428 39748
rect -1428 39692 -1372 39748
rect -1372 39692 -1368 39748
rect -1432 39688 -1368 39692
rect -1432 39588 -1368 39592
rect -1432 39532 -1428 39588
rect -1428 39532 -1372 39588
rect -1372 39532 -1368 39588
rect -1432 39528 -1368 39532
rect -1432 39428 -1368 39432
rect -1432 39372 -1428 39428
rect -1428 39372 -1372 39428
rect -1372 39372 -1368 39428
rect -1432 39368 -1368 39372
rect -1432 39268 -1368 39272
rect -1432 39212 -1428 39268
rect -1428 39212 -1372 39268
rect -1372 39212 -1368 39268
rect -1432 39208 -1368 39212
rect -1432 39108 -1368 39112
rect -1432 39052 -1428 39108
rect -1428 39052 -1372 39108
rect -1372 39052 -1368 39108
rect -1432 39048 -1368 39052
rect -1432 38948 -1368 38952
rect -1432 38892 -1428 38948
rect -1428 38892 -1372 38948
rect -1372 38892 -1368 38948
rect -1432 38888 -1368 38892
rect -1432 38788 -1368 38792
rect -1432 38732 -1428 38788
rect -1428 38732 -1372 38788
rect -1372 38732 -1368 38788
rect -1432 38728 -1368 38732
rect -1432 38628 -1368 38632
rect -1432 38572 -1428 38628
rect -1428 38572 -1372 38628
rect -1372 38572 -1368 38628
rect -1432 38568 -1368 38572
rect -1432 38468 -1368 38472
rect -1432 38412 -1428 38468
rect -1428 38412 -1372 38468
rect -1372 38412 -1368 38468
rect -1432 38408 -1368 38412
rect -1432 38308 -1368 38312
rect -1432 38252 -1428 38308
rect -1428 38252 -1372 38308
rect -1372 38252 -1368 38308
rect -1432 38248 -1368 38252
rect -1432 38148 -1368 38152
rect -1432 38092 -1428 38148
rect -1428 38092 -1372 38148
rect -1372 38092 -1368 38148
rect -1432 38088 -1368 38092
rect -1432 37988 -1368 37992
rect -1432 37932 -1428 37988
rect -1428 37932 -1372 37988
rect -1372 37932 -1368 37988
rect -1432 37928 -1368 37932
rect -1432 37828 -1368 37832
rect -1432 37772 -1428 37828
rect -1428 37772 -1372 37828
rect -1372 37772 -1368 37828
rect -1432 37768 -1368 37772
rect -1112 39748 -1048 39752
rect -1112 39692 -1108 39748
rect -1108 39692 -1052 39748
rect -1052 39692 -1048 39748
rect -1112 39688 -1048 39692
rect -1112 39588 -1048 39592
rect -1112 39532 -1108 39588
rect -1108 39532 -1052 39588
rect -1052 39532 -1048 39588
rect -1112 39528 -1048 39532
rect -1112 39428 -1048 39432
rect -1112 39372 -1108 39428
rect -1108 39372 -1052 39428
rect -1052 39372 -1048 39428
rect -1112 39368 -1048 39372
rect -1112 39268 -1048 39272
rect -1112 39212 -1108 39268
rect -1108 39212 -1052 39268
rect -1052 39212 -1048 39268
rect -1112 39208 -1048 39212
rect -1112 39108 -1048 39112
rect -1112 39052 -1108 39108
rect -1108 39052 -1052 39108
rect -1052 39052 -1048 39108
rect -1112 39048 -1048 39052
rect -1112 38948 -1048 38952
rect -1112 38892 -1108 38948
rect -1108 38892 -1052 38948
rect -1052 38892 -1048 38948
rect -1112 38888 -1048 38892
rect -1112 38788 -1048 38792
rect -1112 38732 -1108 38788
rect -1108 38732 -1052 38788
rect -1052 38732 -1048 38788
rect -1112 38728 -1048 38732
rect -1112 38628 -1048 38632
rect -1112 38572 -1108 38628
rect -1108 38572 -1052 38628
rect -1052 38572 -1048 38628
rect -1112 38568 -1048 38572
rect -1112 38468 -1048 38472
rect -1112 38412 -1108 38468
rect -1108 38412 -1052 38468
rect -1052 38412 -1048 38468
rect -1112 38408 -1048 38412
rect -1112 38308 -1048 38312
rect -1112 38252 -1108 38308
rect -1108 38252 -1052 38308
rect -1052 38252 -1048 38308
rect -1112 38248 -1048 38252
rect -1112 38148 -1048 38152
rect -1112 38092 -1108 38148
rect -1108 38092 -1052 38148
rect -1052 38092 -1048 38148
rect -1112 38088 -1048 38092
rect -1112 37988 -1048 37992
rect -1112 37932 -1108 37988
rect -1108 37932 -1052 37988
rect -1052 37932 -1048 37988
rect -1112 37928 -1048 37932
rect -1112 37828 -1048 37832
rect -1112 37772 -1108 37828
rect -1108 37772 -1052 37828
rect -1052 37772 -1048 37828
rect -1112 37768 -1048 37772
rect -1432 37508 -1368 37512
rect -1432 37452 -1428 37508
rect -1428 37452 -1372 37508
rect -1372 37452 -1368 37508
rect -1432 37448 -1368 37452
rect -1432 37348 -1368 37352
rect -1432 37292 -1428 37348
rect -1428 37292 -1372 37348
rect -1372 37292 -1368 37348
rect -1432 37288 -1368 37292
rect -1432 37188 -1368 37192
rect -1432 37132 -1428 37188
rect -1428 37132 -1372 37188
rect -1372 37132 -1368 37188
rect -1432 37128 -1368 37132
rect -1432 37028 -1368 37032
rect -1432 36972 -1428 37028
rect -1428 36972 -1372 37028
rect -1372 36972 -1368 37028
rect -1432 36968 -1368 36972
rect -1432 36868 -1368 36872
rect -1432 36812 -1428 36868
rect -1428 36812 -1372 36868
rect -1372 36812 -1368 36868
rect -1432 36808 -1368 36812
rect -1432 36708 -1368 36712
rect -1432 36652 -1428 36708
rect -1428 36652 -1372 36708
rect -1372 36652 -1368 36708
rect -1432 36648 -1368 36652
rect -1432 36548 -1368 36552
rect -1432 36492 -1428 36548
rect -1428 36492 -1372 36548
rect -1372 36492 -1368 36548
rect -1432 36488 -1368 36492
rect -1432 36388 -1368 36392
rect -1432 36332 -1428 36388
rect -1428 36332 -1372 36388
rect -1372 36332 -1368 36388
rect -1432 36328 -1368 36332
rect -1752 35748 -1688 35752
rect -1752 35692 -1748 35748
rect -1748 35692 -1692 35748
rect -1692 35692 -1688 35748
rect -1752 35688 -1688 35692
rect -1752 35588 -1688 35592
rect -1752 35532 -1748 35588
rect -1748 35532 -1692 35588
rect -1692 35532 -1688 35588
rect -1752 35528 -1688 35532
rect -1752 35428 -1688 35432
rect -1752 35372 -1748 35428
rect -1748 35372 -1692 35428
rect -1692 35372 -1688 35428
rect -1752 35368 -1688 35372
rect -1752 35268 -1688 35272
rect -1752 35212 -1748 35268
rect -1748 35212 -1692 35268
rect -1692 35212 -1688 35268
rect -1752 35208 -1688 35212
rect -1752 35108 -1688 35112
rect -1752 35052 -1748 35108
rect -1748 35052 -1692 35108
rect -1692 35052 -1688 35108
rect -1752 35048 -1688 35052
rect -1752 34948 -1688 34952
rect -1752 34892 -1748 34948
rect -1748 34892 -1692 34948
rect -1692 34892 -1688 34948
rect -1752 34888 -1688 34892
rect -1752 34788 -1688 34792
rect -1752 34732 -1748 34788
rect -1748 34732 -1692 34788
rect -1692 34732 -1688 34788
rect -1752 34728 -1688 34732
rect -1752 34628 -1688 34632
rect -1752 34572 -1748 34628
rect -1748 34572 -1692 34628
rect -1692 34572 -1688 34628
rect -1752 34568 -1688 34572
rect -1752 34468 -1688 34472
rect -1752 34412 -1748 34468
rect -1748 34412 -1692 34468
rect -1692 34412 -1688 34468
rect -1752 34408 -1688 34412
rect -1752 34308 -1688 34312
rect -1752 34252 -1748 34308
rect -1748 34252 -1692 34308
rect -1692 34252 -1688 34308
rect -1752 34248 -1688 34252
rect -1752 34148 -1688 34152
rect -1752 34092 -1748 34148
rect -1748 34092 -1692 34148
rect -1692 34092 -1688 34148
rect -1752 34088 -1688 34092
rect -1752 33988 -1688 33992
rect -1752 33932 -1748 33988
rect -1748 33932 -1692 33988
rect -1692 33932 -1688 33988
rect -1752 33928 -1688 33932
rect -1752 33828 -1688 33832
rect -1752 33772 -1748 33828
rect -1748 33772 -1692 33828
rect -1692 33772 -1688 33828
rect -1752 33768 -1688 33772
rect -1752 33668 -1688 33672
rect -1752 33612 -1748 33668
rect -1748 33612 -1692 33668
rect -1692 33612 -1688 33668
rect -1752 33608 -1688 33612
rect -1752 33508 -1688 33512
rect -1752 33452 -1748 33508
rect -1748 33452 -1692 33508
rect -1692 33452 -1688 33508
rect -1752 33448 -1688 33452
rect -1752 33268 -1688 33272
rect -1752 33212 -1748 33268
rect -1748 33212 -1692 33268
rect -1692 33212 -1688 33268
rect -1752 33208 -1688 33212
rect -1752 33108 -1688 33112
rect -1752 33052 -1748 33108
rect -1748 33052 -1692 33108
rect -1692 33052 -1688 33108
rect -1752 33048 -1688 33052
rect -1432 35748 -1368 35752
rect -1432 35692 -1428 35748
rect -1428 35692 -1372 35748
rect -1372 35692 -1368 35748
rect -1432 35688 -1368 35692
rect -1432 35588 -1368 35592
rect -1432 35532 -1428 35588
rect -1428 35532 -1372 35588
rect -1372 35532 -1368 35588
rect -1432 35528 -1368 35532
rect -1432 35428 -1368 35432
rect -1432 35372 -1428 35428
rect -1428 35372 -1372 35428
rect -1372 35372 -1368 35428
rect -1432 35368 -1368 35372
rect -1432 35268 -1368 35272
rect -1432 35212 -1428 35268
rect -1428 35212 -1372 35268
rect -1372 35212 -1368 35268
rect -1432 35208 -1368 35212
rect -1432 35108 -1368 35112
rect -1432 35052 -1428 35108
rect -1428 35052 -1372 35108
rect -1372 35052 -1368 35108
rect -1432 35048 -1368 35052
rect -1432 34948 -1368 34952
rect -1432 34892 -1428 34948
rect -1428 34892 -1372 34948
rect -1372 34892 -1368 34948
rect -1432 34888 -1368 34892
rect -1432 34788 -1368 34792
rect -1432 34732 -1428 34788
rect -1428 34732 -1372 34788
rect -1372 34732 -1368 34788
rect -1432 34728 -1368 34732
rect -1432 34628 -1368 34632
rect -1432 34572 -1428 34628
rect -1428 34572 -1372 34628
rect -1372 34572 -1368 34628
rect -1432 34568 -1368 34572
rect -1432 34468 -1368 34472
rect -1432 34412 -1428 34468
rect -1428 34412 -1372 34468
rect -1372 34412 -1368 34468
rect -1432 34408 -1368 34412
rect -1432 34308 -1368 34312
rect -1432 34252 -1428 34308
rect -1428 34252 -1372 34308
rect -1372 34252 -1368 34308
rect -1432 34248 -1368 34252
rect -1432 34148 -1368 34152
rect -1432 34092 -1428 34148
rect -1428 34092 -1372 34148
rect -1372 34092 -1368 34148
rect -1432 34088 -1368 34092
rect -1432 33988 -1368 33992
rect -1432 33932 -1428 33988
rect -1428 33932 -1372 33988
rect -1372 33932 -1368 33988
rect -1432 33928 -1368 33932
rect -1432 33828 -1368 33832
rect -1432 33772 -1428 33828
rect -1428 33772 -1372 33828
rect -1372 33772 -1368 33828
rect -1432 33768 -1368 33772
rect -1432 33668 -1368 33672
rect -1432 33612 -1428 33668
rect -1428 33612 -1372 33668
rect -1372 33612 -1368 33668
rect -1432 33608 -1368 33612
rect -1432 33508 -1368 33512
rect -1432 33452 -1428 33508
rect -1428 33452 -1372 33508
rect -1372 33452 -1368 33508
rect -1432 33448 -1368 33452
rect -1432 33268 -1368 33272
rect -1432 33212 -1428 33268
rect -1428 33212 -1372 33268
rect -1372 33212 -1368 33268
rect -1432 33208 -1368 33212
rect -1432 33108 -1368 33112
rect -1432 33052 -1428 33108
rect -1428 33052 -1372 33108
rect -1372 33052 -1368 33108
rect -1432 33048 -1368 33052
rect -1112 37508 -1048 37512
rect -1112 37452 -1108 37508
rect -1108 37452 -1052 37508
rect -1052 37452 -1048 37508
rect -1112 37448 -1048 37452
rect -1112 37348 -1048 37352
rect -1112 37292 -1108 37348
rect -1108 37292 -1052 37348
rect -1052 37292 -1048 37348
rect -1112 37288 -1048 37292
rect -1112 37188 -1048 37192
rect -1112 37132 -1108 37188
rect -1108 37132 -1052 37188
rect -1052 37132 -1048 37188
rect -1112 37128 -1048 37132
rect -1112 37028 -1048 37032
rect -1112 36972 -1108 37028
rect -1108 36972 -1052 37028
rect -1052 36972 -1048 37028
rect -1112 36968 -1048 36972
rect -1112 36868 -1048 36872
rect -1112 36812 -1108 36868
rect -1108 36812 -1052 36868
rect -1052 36812 -1048 36868
rect -1112 36808 -1048 36812
rect -1112 36708 -1048 36712
rect -1112 36652 -1108 36708
rect -1108 36652 -1052 36708
rect -1052 36652 -1048 36708
rect -1112 36648 -1048 36652
rect -1112 36548 -1048 36552
rect -1112 36492 -1108 36548
rect -1108 36492 -1052 36548
rect -1052 36492 -1048 36548
rect -1112 36488 -1048 36492
rect -1112 36388 -1048 36392
rect -1112 36332 -1108 36388
rect -1108 36332 -1052 36388
rect -1052 36332 -1048 36388
rect -1112 36328 -1048 36332
rect -1112 35748 -1048 35752
rect -1112 35692 -1108 35748
rect -1108 35692 -1052 35748
rect -1052 35692 -1048 35748
rect -1112 35688 -1048 35692
rect -1112 35588 -1048 35592
rect -1112 35532 -1108 35588
rect -1108 35532 -1052 35588
rect -1052 35532 -1048 35588
rect -1112 35528 -1048 35532
rect -1112 35428 -1048 35432
rect -1112 35372 -1108 35428
rect -1108 35372 -1052 35428
rect -1052 35372 -1048 35428
rect -1112 35368 -1048 35372
rect -1112 35268 -1048 35272
rect -1112 35212 -1108 35268
rect -1108 35212 -1052 35268
rect -1052 35212 -1048 35268
rect -1112 35208 -1048 35212
rect -1112 35108 -1048 35112
rect -1112 35052 -1108 35108
rect -1108 35052 -1052 35108
rect -1052 35052 -1048 35108
rect -1112 35048 -1048 35052
rect -1112 34948 -1048 34952
rect -1112 34892 -1108 34948
rect -1108 34892 -1052 34948
rect -1052 34892 -1048 34948
rect -1112 34888 -1048 34892
rect -1112 34788 -1048 34792
rect -1112 34732 -1108 34788
rect -1108 34732 -1052 34788
rect -1052 34732 -1048 34788
rect -1112 34728 -1048 34732
rect -1112 34628 -1048 34632
rect -1112 34572 -1108 34628
rect -1108 34572 -1052 34628
rect -1052 34572 -1048 34628
rect -1112 34568 -1048 34572
rect -1112 34468 -1048 34472
rect -1112 34412 -1108 34468
rect -1108 34412 -1052 34468
rect -1052 34412 -1048 34468
rect -1112 34408 -1048 34412
rect -1112 34308 -1048 34312
rect -1112 34252 -1108 34308
rect -1108 34252 -1052 34308
rect -1052 34252 -1048 34308
rect -1112 34248 -1048 34252
rect -1112 34148 -1048 34152
rect -1112 34092 -1108 34148
rect -1108 34092 -1052 34148
rect -1052 34092 -1048 34148
rect -1112 34088 -1048 34092
rect -1112 33988 -1048 33992
rect -1112 33932 -1108 33988
rect -1108 33932 -1052 33988
rect -1052 33932 -1048 33988
rect -1112 33928 -1048 33932
rect -1112 33828 -1048 33832
rect -1112 33772 -1108 33828
rect -1108 33772 -1052 33828
rect -1052 33772 -1048 33828
rect -1112 33768 -1048 33772
rect -1112 33668 -1048 33672
rect -1112 33612 -1108 33668
rect -1108 33612 -1052 33668
rect -1052 33612 -1048 33668
rect -1112 33608 -1048 33612
rect -1112 33508 -1048 33512
rect -1112 33452 -1108 33508
rect -1108 33452 -1052 33508
rect -1052 33452 -1048 33508
rect -1112 33448 -1048 33452
rect -1112 33268 -1048 33272
rect -1112 33212 -1108 33268
rect -1108 33212 -1052 33268
rect -1052 33212 -1048 33268
rect -1112 33208 -1048 33212
rect -1112 33108 -1048 33112
rect -1112 33052 -1108 33108
rect -1108 33052 -1052 33108
rect -1052 33052 -1048 33108
rect -1112 33048 -1048 33052
<< metal4 >>
rect -33120 78958 43200 79040
rect -33120 78722 -33038 78958
rect -32802 78722 42882 78958
rect 43118 78722 43200 78958
rect -33120 78640 43200 78722
rect -33120 78478 43200 78560
rect -33120 78242 -32238 78478
rect -32002 78242 42082 78478
rect 42318 78242 43200 78478
rect -33120 78160 43200 78242
rect -33120 77998 43200 78080
rect -33120 77762 -31438 77998
rect -31202 77762 41282 77998
rect 41518 77762 43200 77998
rect -33120 77680 43200 77762
rect -31520 74798 -31040 74880
rect -31520 74562 -31438 74798
rect -31202 74562 -31040 74798
rect -31520 74480 -31040 74562
rect -1040 74480 -960 74880
rect 40960 74798 41600 74880
rect 40960 74562 41282 74798
rect 41518 74562 41600 74798
rect 40960 74480 41600 74562
rect -32320 74318 -31040 74400
rect -32320 74082 -32238 74318
rect -32002 74082 -31040 74318
rect -32320 74000 -31040 74082
rect -1040 74000 -960 74400
rect 40960 74318 42400 74400
rect 40960 74082 42082 74318
rect 42318 74082 42400 74318
rect 40960 74000 42400 74082
rect 40960 73358 43200 73440
rect 40960 73122 42882 73358
rect 43118 73122 43200 73358
rect 40960 73040 43200 73122
rect -31040 41752 -30000 41760
rect -31040 41688 -31032 41752
rect -30968 41688 -30712 41752
rect -30648 41688 -30392 41752
rect -30328 41688 -30072 41752
rect -30008 41688 -30000 41752
rect -31040 41680 -30000 41688
rect -31040 41592 -30000 41600
rect -31040 41528 -31032 41592
rect -30968 41528 -30712 41592
rect -30648 41528 -30392 41592
rect -30328 41528 -30072 41592
rect -30008 41528 -30000 41592
rect -31040 41520 -30000 41528
rect -31040 40792 -30000 40800
rect -31040 40728 -31032 40792
rect -30968 40728 -30712 40792
rect -30648 40728 -30392 40792
rect -30328 40728 -30072 40792
rect -30008 40728 -30000 40792
rect -31040 40720 -30000 40728
rect -31040 40632 -30000 40640
rect -31040 40568 -31032 40632
rect -30968 40568 -30712 40632
rect -30648 40568 -30392 40632
rect -30328 40568 -30072 40632
rect -30008 40568 -30000 40632
rect -31040 40560 -30000 40568
rect -31040 40472 -30000 40480
rect -31040 40408 -31032 40472
rect -30968 40408 -30712 40472
rect -30648 40408 -30392 40472
rect -30328 40408 -30072 40472
rect -30008 40408 -30000 40472
rect -31040 40400 -30000 40408
rect -31040 40312 -30000 40320
rect -31040 40248 -31032 40312
rect -30968 40248 -30712 40312
rect -30648 40248 -30392 40312
rect -30328 40248 -30072 40312
rect -30008 40248 -30000 40312
rect -31040 40240 -30000 40248
rect -31040 40152 -30000 40160
rect -31040 40088 -31032 40152
rect -30968 40088 -30712 40152
rect -30648 40088 -30392 40152
rect -30328 40088 -30072 40152
rect -30008 40088 -30000 40152
rect -31040 40080 -30000 40088
rect -31040 39992 -30000 40000
rect -31040 39928 -31032 39992
rect -30968 39928 -30712 39992
rect -30648 39928 -30392 39992
rect -30328 39928 -30072 39992
rect -30008 39928 -30000 39992
rect -31040 39920 -30000 39928
rect -31040 39832 -30000 39840
rect -31040 39768 -31032 39832
rect -30968 39768 -30712 39832
rect -30648 39768 -30392 39832
rect -30328 39768 -30072 39832
rect -30008 39768 -30000 39832
rect -31040 39760 -30000 39768
rect -3360 39752 -1040 39760
rect -3360 39688 -3352 39752
rect -3288 39688 -3032 39752
rect -2968 39688 -2712 39752
rect -2648 39688 -2392 39752
rect -2328 39688 -2072 39752
rect -2008 39688 -1752 39752
rect -1688 39688 -1432 39752
rect -1368 39688 -1112 39752
rect -1048 39688 -1040 39752
rect -3360 39680 -1040 39688
rect -31040 39672 -30000 39680
rect -31040 39608 -31032 39672
rect -30968 39608 -30712 39672
rect -30648 39608 -30392 39672
rect -30328 39608 -30072 39672
rect -30008 39608 -30000 39672
rect -31040 39600 -30000 39608
rect -3360 39592 -1040 39600
rect -3360 39528 -3352 39592
rect -3288 39528 -3032 39592
rect -2968 39528 -2712 39592
rect -2648 39528 -2392 39592
rect -2328 39528 -2072 39592
rect -2008 39528 -1752 39592
rect -1688 39528 -1432 39592
rect -1368 39528 -1112 39592
rect -1048 39528 -1040 39592
rect -3360 39520 -1040 39528
rect -31040 39512 -30000 39520
rect -31040 39448 -31032 39512
rect -30968 39448 -30712 39512
rect -30648 39448 -30392 39512
rect -30328 39448 -30072 39512
rect -30008 39448 -30000 39512
rect -31040 39440 -30000 39448
rect -3360 39432 -1040 39440
rect -3360 39368 -3352 39432
rect -3288 39368 -3032 39432
rect -2968 39368 -2712 39432
rect -2648 39368 -2392 39432
rect -2328 39368 -2072 39432
rect -2008 39368 -1752 39432
rect -1688 39368 -1432 39432
rect -1368 39368 -1112 39432
rect -1048 39368 -1040 39432
rect -3360 39360 -1040 39368
rect -31040 39352 -30000 39360
rect -31040 39288 -31032 39352
rect -30968 39288 -30712 39352
rect -30648 39288 -30392 39352
rect -30328 39288 -30072 39352
rect -30008 39288 -30000 39352
rect -31040 39280 -30000 39288
rect -3360 39272 -1040 39280
rect -3360 39208 -3352 39272
rect -3288 39208 -3032 39272
rect -2968 39208 -2712 39272
rect -2648 39208 -2392 39272
rect -2328 39208 -2072 39272
rect -2008 39208 -1752 39272
rect -1688 39208 -1432 39272
rect -1368 39208 -1112 39272
rect -1048 39208 -1040 39272
rect -3360 39200 -1040 39208
rect -31040 39192 -30000 39200
rect -31040 39128 -31032 39192
rect -30968 39128 -30712 39192
rect -30648 39128 -30392 39192
rect -30328 39128 -30072 39192
rect -30008 39128 -30000 39192
rect -31040 39120 -30000 39128
rect -3360 39112 -1040 39120
rect -3360 39048 -3352 39112
rect -3288 39048 -3032 39112
rect -2968 39048 -2712 39112
rect -2648 39048 -2392 39112
rect -2328 39048 -2072 39112
rect -2008 39048 -1752 39112
rect -1688 39048 -1432 39112
rect -1368 39048 -1112 39112
rect -1048 39048 -1040 39112
rect -3360 39040 -1040 39048
rect -31040 39032 -30000 39040
rect -31040 38968 -31032 39032
rect -30968 38968 -30712 39032
rect -30648 38968 -30392 39032
rect -30328 38968 -30072 39032
rect -30008 38968 -30000 39032
rect -31040 38960 -30000 38968
rect -3360 38952 -1040 38960
rect -3360 38888 -3352 38952
rect -3288 38888 -3032 38952
rect -2968 38888 -2712 38952
rect -2648 38888 -2392 38952
rect -2328 38888 -2072 38952
rect -2008 38888 -1752 38952
rect -1688 38888 -1432 38952
rect -1368 38888 -1112 38952
rect -1048 38888 -1040 38952
rect -3360 38880 -1040 38888
rect -31040 38872 -30000 38880
rect -31040 38808 -31032 38872
rect -30968 38808 -30712 38872
rect -30648 38808 -30392 38872
rect -30328 38808 -30072 38872
rect -30008 38808 -30000 38872
rect -31040 38800 -30000 38808
rect -3360 38792 -1040 38800
rect -3360 38728 -3352 38792
rect -3288 38728 -3032 38792
rect -2968 38728 -2712 38792
rect -2648 38728 -2392 38792
rect -2328 38728 -2072 38792
rect -2008 38728 -1752 38792
rect -1688 38728 -1432 38792
rect -1368 38728 -1112 38792
rect -1048 38728 -1040 38792
rect -3360 38720 -1040 38728
rect -31040 38712 -30000 38720
rect -31040 38648 -31032 38712
rect -30968 38648 -30712 38712
rect -30648 38648 -30392 38712
rect -30328 38648 -30072 38712
rect -30008 38648 -30000 38712
rect -31040 38640 -30000 38648
rect -3360 38632 -1040 38640
rect -3360 38568 -3352 38632
rect -3288 38568 -3032 38632
rect -2968 38568 -2712 38632
rect -2648 38568 -2392 38632
rect -2328 38568 -2072 38632
rect -2008 38568 -1752 38632
rect -1688 38568 -1432 38632
rect -1368 38568 -1112 38632
rect -1048 38568 -1040 38632
rect -3360 38560 -1040 38568
rect -31040 38552 -30000 38560
rect -31040 38488 -31032 38552
rect -30968 38488 -30712 38552
rect -30648 38488 -30392 38552
rect -30328 38488 -30072 38552
rect -30008 38488 -30000 38552
rect -31040 38480 -30000 38488
rect -3360 38472 -1040 38480
rect -3360 38408 -3352 38472
rect -3288 38408 -3032 38472
rect -2968 38408 -2712 38472
rect -2648 38408 -2392 38472
rect -2328 38408 -2072 38472
rect -2008 38408 -1752 38472
rect -1688 38408 -1432 38472
rect -1368 38408 -1112 38472
rect -1048 38408 -1040 38472
rect -3360 38400 -1040 38408
rect -31040 38392 -30000 38400
rect -31040 38328 -31032 38392
rect -30968 38328 -30712 38392
rect -30648 38328 -30392 38392
rect -30328 38328 -30072 38392
rect -30008 38328 -30000 38392
rect -31040 38320 -30000 38328
rect -3360 38312 -1040 38320
rect -3360 38248 -3352 38312
rect -3288 38248 -3032 38312
rect -2968 38248 -2712 38312
rect -2648 38248 -2392 38312
rect -2328 38248 -2072 38312
rect -2008 38248 -1752 38312
rect -1688 38248 -1432 38312
rect -1368 38248 -1112 38312
rect -1048 38248 -1040 38312
rect -3360 38240 -1040 38248
rect -31040 38232 -30000 38240
rect -31040 38168 -31032 38232
rect -30968 38168 -30712 38232
rect -30648 38168 -30392 38232
rect -30328 38168 -30072 38232
rect -30008 38168 -30000 38232
rect -31040 38160 -30000 38168
rect -3360 38152 -1040 38160
rect -3360 38088 -3352 38152
rect -3288 38088 -3032 38152
rect -2968 38088 -2712 38152
rect -2648 38088 -2392 38152
rect -2328 38088 -2072 38152
rect -2008 38088 -1752 38152
rect -1688 38088 -1432 38152
rect -1368 38088 -1112 38152
rect -1048 38088 -1040 38152
rect -3360 38080 -1040 38088
rect -31040 38072 -30000 38080
rect -31040 38008 -31032 38072
rect -30968 38008 -30712 38072
rect -30648 38008 -30392 38072
rect -30328 38008 -30072 38072
rect -30008 38008 -30000 38072
rect -31040 38000 -30000 38008
rect -3360 37992 -1040 38000
rect -3360 37928 -3352 37992
rect -3288 37928 -3032 37992
rect -2968 37928 -2712 37992
rect -2648 37928 -2392 37992
rect -2328 37928 -2072 37992
rect -2008 37928 -1752 37992
rect -1688 37928 -1432 37992
rect -1368 37928 -1112 37992
rect -1048 37928 -1040 37992
rect -3360 37920 -1040 37928
rect -31040 37912 -30000 37920
rect -31040 37848 -31032 37912
rect -30968 37848 -30712 37912
rect -30648 37848 -30392 37912
rect -30328 37848 -30072 37912
rect -30008 37848 -30000 37912
rect -31040 37840 -30000 37848
rect -3360 37832 -1040 37840
rect -3360 37768 -3352 37832
rect -3288 37768 -3032 37832
rect -2968 37768 -2712 37832
rect -2648 37768 -2392 37832
rect -2328 37768 -2072 37832
rect -2008 37768 -1752 37832
rect -1688 37768 -1432 37832
rect -1368 37768 -1112 37832
rect -1048 37768 -1040 37832
rect -3360 37760 -1040 37768
rect -31040 37752 -30000 37760
rect -31040 37688 -31032 37752
rect -30968 37688 -30712 37752
rect -30648 37688 -30392 37752
rect -30328 37688 -30072 37752
rect -30008 37688 -30000 37752
rect -31040 37680 -30000 37688
rect -3360 37512 -1040 37520
rect -3360 37448 -3352 37512
rect -3288 37448 -3032 37512
rect -2968 37448 -2712 37512
rect -2648 37448 -2392 37512
rect -2328 37448 -2072 37512
rect -2008 37448 -1752 37512
rect -1688 37448 -1432 37512
rect -1368 37448 -1112 37512
rect -1048 37448 -1040 37512
rect -3360 37440 -1040 37448
rect -3360 37352 -1040 37360
rect -3360 37288 -3352 37352
rect -3288 37288 -3032 37352
rect -2968 37288 -2712 37352
rect -2648 37288 -2392 37352
rect -2328 37288 -2072 37352
rect -2008 37288 -1752 37352
rect -1688 37288 -1432 37352
rect -1368 37288 -1112 37352
rect -1048 37288 -1040 37352
rect -3360 37280 -1040 37288
rect -3360 37192 -1040 37200
rect -3360 37128 -3352 37192
rect -3288 37128 -3032 37192
rect -2968 37128 -2712 37192
rect -2648 37128 -2392 37192
rect -2328 37128 -2072 37192
rect -2008 37128 -1752 37192
rect -1688 37128 -1432 37192
rect -1368 37128 -1112 37192
rect -1048 37128 -1040 37192
rect -3360 37120 -1040 37128
rect -31040 37112 -30000 37120
rect -31040 37048 -31032 37112
rect -30968 37048 -30712 37112
rect -30648 37048 -30392 37112
rect -30328 37048 -30072 37112
rect -30008 37048 -30000 37112
rect -31040 37040 -30000 37048
rect -3360 37032 -1040 37040
rect -3360 36968 -3352 37032
rect -3288 36968 -3032 37032
rect -2968 36968 -2712 37032
rect -2648 36968 -2392 37032
rect -2328 36968 -2072 37032
rect -2008 36968 -1752 37032
rect -1688 36968 -1432 37032
rect -1368 36968 -1112 37032
rect -1048 36968 -1040 37032
rect -3360 36960 -1040 36968
rect -31040 36952 -30000 36960
rect -31040 36888 -31032 36952
rect -30968 36888 -30712 36952
rect -30648 36888 -30392 36952
rect -30328 36888 -30072 36952
rect -30008 36888 -30000 36952
rect -31040 36880 -30000 36888
rect -3360 36872 -1040 36880
rect -3360 36808 -3352 36872
rect -3288 36808 -3032 36872
rect -2968 36808 -2712 36872
rect -2648 36808 -2392 36872
rect -2328 36808 -2072 36872
rect -2008 36808 -1752 36872
rect -1688 36808 -1432 36872
rect -1368 36808 -1112 36872
rect -1048 36808 -1040 36872
rect -3360 36800 -1040 36808
rect -31040 36792 -30000 36800
rect -31040 36728 -31032 36792
rect -30968 36728 -30712 36792
rect -30648 36728 -30392 36792
rect -30328 36728 -30072 36792
rect -30008 36728 -30000 36792
rect -31040 36720 -30000 36728
rect -3360 36712 -1040 36720
rect -3360 36648 -3352 36712
rect -3288 36648 -3032 36712
rect -2968 36648 -2712 36712
rect -2648 36648 -2392 36712
rect -2328 36648 -2072 36712
rect -2008 36648 -1752 36712
rect -1688 36648 -1432 36712
rect -1368 36648 -1112 36712
rect -1048 36648 -1040 36712
rect -3360 36640 -1040 36648
rect -31040 36632 -30000 36640
rect -31040 36568 -31032 36632
rect -30968 36568 -30712 36632
rect -30648 36568 -30392 36632
rect -30328 36568 -30072 36632
rect -30008 36568 -30000 36632
rect -31040 36560 -30000 36568
rect -3360 36552 -1040 36560
rect -3360 36488 -3352 36552
rect -3288 36488 -3032 36552
rect -2968 36488 -2712 36552
rect -2648 36488 -2392 36552
rect -2328 36488 -2072 36552
rect -2008 36488 -1752 36552
rect -1688 36488 -1432 36552
rect -1368 36488 -1112 36552
rect -1048 36488 -1040 36552
rect -3360 36480 -1040 36488
rect -31040 36472 -30000 36480
rect -31040 36408 -31032 36472
rect -30968 36408 -30712 36472
rect -30648 36408 -30392 36472
rect -30328 36408 -30072 36472
rect -30008 36408 -30000 36472
rect -31040 36400 -30000 36408
rect -3360 36392 -1040 36400
rect -3360 36328 -3352 36392
rect -3288 36328 -3032 36392
rect -2968 36328 -2712 36392
rect -2648 36328 -2392 36392
rect -2328 36328 -2072 36392
rect -2008 36328 -1752 36392
rect -1688 36328 -1432 36392
rect -1368 36328 -1112 36392
rect -1048 36328 -1040 36392
rect -3360 36320 -1040 36328
rect -31040 36312 -30000 36320
rect -31040 36248 -31032 36312
rect -30968 36248 -30712 36312
rect -30648 36248 -30392 36312
rect -30328 36248 -30072 36312
rect -30008 36248 -30000 36312
rect -31040 36240 -30000 36248
rect -31040 36152 -30000 36160
rect -31040 36088 -31032 36152
rect -30968 36088 -30712 36152
rect -30648 36088 -30392 36152
rect -30328 36088 -30072 36152
rect -30008 36088 -30000 36152
rect -31040 36080 -30000 36088
rect -31040 35992 -30000 36000
rect -31040 35928 -31032 35992
rect -30968 35928 -30712 35992
rect -30648 35928 -30392 35992
rect -30328 35928 -30072 35992
rect -30008 35928 -30000 35992
rect -31040 35920 -30000 35928
rect -31040 35832 -30000 35840
rect -31040 35768 -31032 35832
rect -30968 35768 -30712 35832
rect -30648 35768 -30392 35832
rect -30328 35768 -30072 35832
rect -30008 35768 -30000 35832
rect -31040 35760 -30000 35768
rect -3360 35752 -1040 35760
rect -3360 35688 -3352 35752
rect -3288 35688 -3032 35752
rect -2968 35688 -2712 35752
rect -2648 35688 -2392 35752
rect -2328 35688 -2072 35752
rect -2008 35688 -1752 35752
rect -1688 35688 -1432 35752
rect -1368 35688 -1112 35752
rect -1048 35688 -1040 35752
rect -3360 35680 -1040 35688
rect -31040 35672 -30000 35680
rect -31040 35608 -31032 35672
rect -30968 35608 -30712 35672
rect -30648 35608 -30392 35672
rect -30328 35608 -30072 35672
rect -30008 35608 -30000 35672
rect -31040 35600 -30000 35608
rect -3360 35592 -1040 35600
rect -3360 35528 -3352 35592
rect -3288 35528 -3032 35592
rect -2968 35528 -2712 35592
rect -2648 35528 -2392 35592
rect -2328 35528 -2072 35592
rect -2008 35528 -1752 35592
rect -1688 35528 -1432 35592
rect -1368 35528 -1112 35592
rect -1048 35528 -1040 35592
rect -3360 35520 -1040 35528
rect -31040 35512 -30000 35520
rect -31040 35448 -31032 35512
rect -30968 35448 -30712 35512
rect -30648 35448 -30392 35512
rect -30328 35448 -30072 35512
rect -30008 35448 -30000 35512
rect -31040 35440 -30000 35448
rect -3360 35432 -1040 35440
rect -3360 35368 -3352 35432
rect -3288 35368 -3032 35432
rect -2968 35368 -2712 35432
rect -2648 35368 -2392 35432
rect -2328 35368 -2072 35432
rect -2008 35368 -1752 35432
rect -1688 35368 -1432 35432
rect -1368 35368 -1112 35432
rect -1048 35368 -1040 35432
rect -3360 35360 -1040 35368
rect -31040 35352 -30000 35360
rect -31040 35288 -31032 35352
rect -30968 35288 -30712 35352
rect -30648 35288 -30392 35352
rect -30328 35288 -30072 35352
rect -30008 35288 -30000 35352
rect -31040 35280 -30000 35288
rect -3360 35272 -1040 35280
rect -3360 35208 -3352 35272
rect -3288 35208 -3032 35272
rect -2968 35208 -2712 35272
rect -2648 35208 -2392 35272
rect -2328 35208 -2072 35272
rect -2008 35208 -1752 35272
rect -1688 35208 -1432 35272
rect -1368 35208 -1112 35272
rect -1048 35208 -1040 35272
rect -3360 35200 -1040 35208
rect -31040 35192 -30000 35200
rect -31040 35128 -31032 35192
rect -30968 35128 -30712 35192
rect -30648 35128 -30392 35192
rect -30328 35128 -30072 35192
rect -30008 35128 -30000 35192
rect -31040 35120 -30000 35128
rect -3360 35112 -1040 35120
rect -3360 35048 -3352 35112
rect -3288 35048 -3032 35112
rect -2968 35048 -2712 35112
rect -2648 35048 -2392 35112
rect -2328 35048 -2072 35112
rect -2008 35048 -1752 35112
rect -1688 35048 -1432 35112
rect -1368 35048 -1112 35112
rect -1048 35048 -1040 35112
rect -3360 35040 -1040 35048
rect -31040 35032 -30000 35040
rect -31040 34968 -31032 35032
rect -30968 34968 -30712 35032
rect -30648 34968 -30392 35032
rect -30328 34968 -30072 35032
rect -30008 34968 -30000 35032
rect -31040 34960 -30000 34968
rect -3360 34952 -1040 34960
rect -3360 34888 -3352 34952
rect -3288 34888 -3032 34952
rect -2968 34888 -2712 34952
rect -2648 34888 -2392 34952
rect -2328 34888 -2072 34952
rect -2008 34888 -1752 34952
rect -1688 34888 -1432 34952
rect -1368 34888 -1112 34952
rect -1048 34888 -1040 34952
rect -3360 34880 -1040 34888
rect -31040 34872 -30000 34880
rect -31040 34808 -31032 34872
rect -30968 34808 -30712 34872
rect -30648 34808 -30392 34872
rect -30328 34808 -30072 34872
rect -30008 34808 -30000 34872
rect -31040 34800 -30000 34808
rect -3360 34792 -1040 34800
rect -3360 34728 -3352 34792
rect -3288 34728 -3032 34792
rect -2968 34728 -2712 34792
rect -2648 34728 -2392 34792
rect -2328 34728 -2072 34792
rect -2008 34728 -1752 34792
rect -1688 34728 -1432 34792
rect -1368 34728 -1112 34792
rect -1048 34728 -1040 34792
rect -3360 34720 -1040 34728
rect -3360 34632 -1040 34640
rect -3360 34568 -3352 34632
rect -3288 34568 -3032 34632
rect -2968 34568 -2712 34632
rect -2648 34568 -2392 34632
rect -2328 34568 -2072 34632
rect -2008 34568 -1752 34632
rect -1688 34568 -1432 34632
rect -1368 34568 -1112 34632
rect -1048 34568 -1040 34632
rect -3360 34560 -1040 34568
rect -3360 34472 -1040 34480
rect -3360 34408 -3352 34472
rect -3288 34408 -3032 34472
rect -2968 34408 -2712 34472
rect -2648 34408 -2392 34472
rect -2328 34408 -2072 34472
rect -2008 34408 -1752 34472
rect -1688 34408 -1432 34472
rect -1368 34408 -1112 34472
rect -1048 34408 -1040 34472
rect -3360 34400 -1040 34408
rect -3360 34312 -1040 34320
rect -3360 34248 -3352 34312
rect -3288 34248 -3032 34312
rect -2968 34248 -2712 34312
rect -2648 34248 -2392 34312
rect -2328 34248 -2072 34312
rect -2008 34248 -1752 34312
rect -1688 34248 -1432 34312
rect -1368 34248 -1112 34312
rect -1048 34248 -1040 34312
rect -3360 34240 -1040 34248
rect -31040 34232 -30000 34240
rect -31040 34168 -31032 34232
rect -30968 34168 -30712 34232
rect -30648 34168 -30392 34232
rect -30328 34168 -30072 34232
rect -30008 34168 -30000 34232
rect -31040 34160 -30000 34168
rect -3360 34152 -1040 34160
rect -3360 34088 -3352 34152
rect -3288 34088 -3032 34152
rect -2968 34088 -2712 34152
rect -2648 34088 -2392 34152
rect -2328 34088 -2072 34152
rect -2008 34088 -1752 34152
rect -1688 34088 -1432 34152
rect -1368 34088 -1112 34152
rect -1048 34088 -1040 34152
rect -3360 34080 -1040 34088
rect -31040 34072 -30000 34080
rect -31040 34008 -31032 34072
rect -30968 34008 -30712 34072
rect -30648 34008 -30392 34072
rect -30328 34008 -30072 34072
rect -30008 34008 -30000 34072
rect -31040 34000 -30000 34008
rect -3360 33992 -1040 34000
rect -3360 33928 -3352 33992
rect -3288 33928 -3032 33992
rect -2968 33928 -2712 33992
rect -2648 33928 -2392 33992
rect -2328 33928 -2072 33992
rect -2008 33928 -1752 33992
rect -1688 33928 -1432 33992
rect -1368 33928 -1112 33992
rect -1048 33928 -1040 33992
rect -3360 33920 -1040 33928
rect -31040 33912 -30000 33920
rect -31040 33848 -31032 33912
rect -30968 33848 -30712 33912
rect -30648 33848 -30392 33912
rect -30328 33848 -30072 33912
rect -30008 33848 -30000 33912
rect -31040 33840 -30000 33848
rect -3360 33832 -1040 33840
rect -3360 33768 -3352 33832
rect -3288 33768 -3032 33832
rect -2968 33768 -2712 33832
rect -2648 33768 -2392 33832
rect -2328 33768 -2072 33832
rect -2008 33768 -1752 33832
rect -1688 33768 -1432 33832
rect -1368 33768 -1112 33832
rect -1048 33768 -1040 33832
rect -3360 33760 -1040 33768
rect -31040 33752 -30000 33760
rect -31040 33688 -31032 33752
rect -30968 33688 -30712 33752
rect -30648 33688 -30392 33752
rect -30328 33688 -30072 33752
rect -30008 33688 -30000 33752
rect -31040 33680 -30000 33688
rect -3360 33672 -1040 33680
rect -3360 33608 -3352 33672
rect -3288 33608 -3032 33672
rect -2968 33608 -2712 33672
rect -2648 33608 -2392 33672
rect -2328 33608 -2072 33672
rect -2008 33608 -1752 33672
rect -1688 33608 -1432 33672
rect -1368 33608 -1112 33672
rect -1048 33608 -1040 33672
rect -3360 33600 -1040 33608
rect -31040 33592 -30000 33600
rect -31040 33528 -31032 33592
rect -30968 33528 -30712 33592
rect -30648 33528 -30392 33592
rect -30328 33528 -30072 33592
rect -30008 33528 -30000 33592
rect -31040 33520 -30000 33528
rect -3360 33512 -1040 33520
rect -3360 33448 -3352 33512
rect -3288 33448 -3032 33512
rect -2968 33448 -2712 33512
rect -2648 33448 -2392 33512
rect -2328 33448 -2072 33512
rect -2008 33448 -1752 33512
rect -1688 33448 -1432 33512
rect -1368 33448 -1112 33512
rect -1048 33448 -1040 33512
rect -3360 33440 -1040 33448
rect -31040 33432 -30000 33440
rect -31040 33368 -31032 33432
rect -30968 33368 -30712 33432
rect -30648 33368 -30392 33432
rect -30328 33368 -30072 33432
rect -30008 33368 -30000 33432
rect -31040 33360 -30000 33368
rect -31040 33272 -30000 33280
rect -31040 33208 -31032 33272
rect -30968 33208 -30712 33272
rect -30648 33208 -30392 33272
rect -30328 33208 -30072 33272
rect -30008 33208 -30000 33272
rect -31040 33200 -30000 33208
rect -3360 33272 -1040 33280
rect -3360 33208 -3352 33272
rect -3288 33208 -3032 33272
rect -2968 33208 -2712 33272
rect -2648 33208 -2392 33272
rect -2328 33208 -2072 33272
rect -2008 33208 -1752 33272
rect -1688 33208 -1432 33272
rect -1368 33208 -1112 33272
rect -1048 33208 -1040 33272
rect -3360 33200 -1040 33208
rect -31040 33112 -30000 33120
rect -31040 33048 -31032 33112
rect -30968 33048 -30712 33112
rect -30648 33048 -30392 33112
rect -30328 33048 -30072 33112
rect -30008 33048 -30000 33112
rect -31040 33040 -30000 33048
rect -3360 33112 -1040 33120
rect -3360 33048 -3352 33112
rect -3288 33048 -3032 33112
rect -2968 33048 -2712 33112
rect -2648 33048 -2392 33112
rect -2328 33048 -2072 33112
rect -2008 33048 -1752 33112
rect -1688 33048 -1432 33112
rect -1368 33048 -1112 33112
rect -1048 33048 -1040 33112
rect -3360 33040 -1040 33048
rect -31040 32952 -30000 32960
rect -31040 32888 -31032 32952
rect -30968 32888 -30712 32952
rect -30648 32888 -30392 32952
rect -30328 32888 -30072 32952
rect -30008 32888 -30000 32952
rect -31040 32880 -30000 32888
rect -32320 718 -31040 800
rect -32320 482 -32238 718
rect -32002 482 -31040 718
rect -32320 400 -31040 482
rect -1040 400 -960 800
rect 40960 718 42400 800
rect 40960 482 42082 718
rect 42318 482 42400 718
rect 40960 400 42400 482
rect -31520 238 -31040 320
rect -31520 2 -31438 238
rect -31202 2 -31040 238
rect -31520 -80 -31040 2
rect -1040 -80 -960 320
rect 40960 238 41600 320
rect 40960 2 41282 238
rect 41518 2 41600 238
rect 40960 -80 41600 2
rect -33120 -2962 43200 -2880
rect -33120 -3198 -31438 -2962
rect -31202 -3198 41282 -2962
rect 41518 -3198 43200 -2962
rect -33120 -3280 43200 -3198
rect -33120 -3442 43200 -3360
rect -33120 -3678 -32238 -3442
rect -32002 -3678 42082 -3442
rect 42318 -3678 43200 -3442
rect -33120 -3760 43200 -3678
rect -33120 -3922 43200 -3840
rect -33120 -4158 -33038 -3922
rect -32802 -4158 42882 -3922
rect 43118 -4158 43200 -3922
rect -33120 -4240 43200 -4158
<< via4 >>
rect -33038 78722 -32802 78958
rect 42882 78722 43118 78958
rect -32238 78242 -32002 78478
rect 42082 78242 42318 78478
rect -31438 77762 -31202 77998
rect 41282 77762 41518 77998
rect -31438 74562 -31202 74798
rect 41282 74562 41518 74798
rect -32238 74082 -32002 74318
rect 42082 74082 42318 74318
rect 42882 73122 43118 73358
rect -32238 482 -32002 718
rect 42082 482 42318 718
rect -31438 2 -31202 238
rect 41282 2 41518 238
rect -31438 -3198 -31202 -2962
rect 41282 -3198 41518 -2962
rect -32238 -3678 -32002 -3442
rect 42082 -3678 42318 -3442
rect -33038 -4158 -32802 -3922
rect 42882 -4158 43118 -3922
<< metal5 >>
rect -33120 78958 -32720 79120
rect -33120 78722 -33038 78958
rect -32802 78722 -32720 78958
rect -33120 -3922 -32720 78722
rect -33120 -4158 -33038 -3922
rect -32802 -4158 -32720 -3922
rect -33120 -4240 -32720 -4158
rect -32320 78478 -31920 79120
rect -32320 78242 -32238 78478
rect -32002 78242 -31920 78478
rect -32320 74318 -31920 78242
rect -32320 74082 -32238 74318
rect -32002 74082 -31920 74318
rect -32320 718 -31920 74082
rect -32320 482 -32238 718
rect -32002 482 -31920 718
rect -32320 -3442 -31920 482
rect -32320 -3678 -32238 -3442
rect -32002 -3678 -31920 -3442
rect -32320 -4240 -31920 -3678
rect -31520 77998 -31120 79120
rect -31520 77762 -31438 77998
rect -31202 77762 -31120 77998
rect -31520 74798 -31120 77762
rect 41200 77998 41600 79040
rect 41200 77762 41282 77998
rect 41518 77762 41600 77998
rect -800 74880 -400 75360
rect 6880 74880 7280 75360
rect 11680 74880 12080 75360
rect -31520 74562 -31438 74798
rect -31202 74562 -31120 74798
rect -31520 238 -31120 74562
rect -31520 2 -31438 238
rect -31202 2 -31120 238
rect -31520 -2962 -31120 2
rect -31520 -3198 -31438 -2962
rect -31202 -3198 -31120 -2962
rect -31520 -4240 -31120 -3198
rect 41200 74798 41600 77762
rect 41200 74562 41282 74798
rect 41518 74562 41600 74798
rect 41200 238 41600 74562
rect 41200 2 41282 238
rect 41518 2 41600 238
rect 41200 -2962 41600 2
rect 41200 -3198 41282 -2962
rect 41518 -3198 41600 -2962
rect 41200 -4240 41600 -3198
rect 42000 78478 42400 79040
rect 42000 78242 42082 78478
rect 42318 78242 42400 78478
rect 42000 74318 42400 78242
rect 42000 74082 42082 74318
rect 42318 74082 42400 74318
rect 42000 718 42400 74082
rect 42000 482 42082 718
rect 42318 482 42400 718
rect 42000 -3442 42400 482
rect 42000 -3678 42082 -3442
rect 42318 -3678 42400 -3442
rect 42000 -4240 42400 -3678
rect 42800 78958 43200 79040
rect 42800 78722 42882 78958
rect 43118 78722 43200 78958
rect 42800 73358 43200 78722
rect 42800 73122 42882 73358
rect 43118 73122 43200 73358
rect 42800 -3922 43200 73122
rect 42800 -4158 42882 -3922
rect 43118 -4158 43200 -3922
rect 42800 -4240 43200 -4158
use ota  ota
timestamp 1638148091
transform 1 0 -960 0 1 4000
box -26 -6800 41946 73600
use pseudo  pseudo
timestamp 1638148091
transform 1 0 -16800 0 1 35600
box -506 -746 13066 4346
use cap1_10  cap1
timestamp 1638148091
transform -1 0 -1040 0 -1 74880
box 0 0 30000 31946
use cap1_10  cap2
timestamp 1638148091
transform 1 0 -31040 0 1 -80
box 0 0 30000 31946
<< labels >>
rlabel metal2 s -1280 40480 -1200 40560 4 q
rlabel metal2 s -1280 39840 -1200 39920 4 op
rlabel metal2 s -1280 40160 -1200 40240 4 xm
rlabel metal2 s -1280 35840 -1200 35920 4 om
rlabel metal2 s -1280 36160 -1200 36240 4 xp
rlabel metal2 s -33280 37520 -33200 37600 4 ip
port 1 nsew
rlabel metal2 s -33280 37200 -33200 37280 4 im
port 2 nsew
rlabel metal2 s 43280 39840 43360 39920 4 op
port 3 nsew
rlabel metal2 s 43280 35840 43360 35920 4 om
port 4 nsew
rlabel metal2 s -33280 34480 -33200 34560 4 fsb
port 5 nsew
rlabel metal2 s -33280 41120 -33200 41200 4 ib
port 6 nsew
rlabel metal2 s 43280 41120 43360 41200 4 ib
port 6 nsew
rlabel metal5 s -33120 79040 -32720 79120 4 vdda
port 7 nsew
rlabel metal5 s -32320 79040 -31920 79120 4 gnda
port 8 nsew
rlabel metal5 s -31520 79040 -31120 79120 4 vssa
port 9 nsew
<< end >>
