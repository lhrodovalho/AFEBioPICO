magic
tech sky130A
timestamp 1637779110
<< nwell >>
rect -180 -180 5180 780
rect -180 -900 5180 -340
<< mvnmos >>
rect 0 -1240 200 -1140
rect 320 -1240 520 -1140
rect 640 -1240 840 -1140
rect 960 -1240 1160 -1140
rect 1280 -1240 1480 -1140
rect 1600 -1240 1800 -1140
rect 1920 -1240 2120 -1140
rect 2240 -1240 2440 -1140
rect 2560 -1240 2760 -1140
rect 2880 -1240 3080 -1140
rect 3200 -1240 3400 -1140
rect 3520 -1240 3720 -1140
rect 3840 -1240 4040 -1140
rect 4160 -1240 4360 -1140
rect 4480 -1240 4680 -1140
rect 4800 -1240 5000 -1140
rect 0 -1440 200 -1340
rect 320 -1440 520 -1340
rect 640 -1440 840 -1340
rect 960 -1440 1160 -1340
rect 1280 -1440 1480 -1340
rect 1600 -1440 1800 -1340
rect 1920 -1440 2120 -1340
rect 2240 -1440 2440 -1340
rect 2560 -1440 2760 -1340
rect 2880 -1440 3080 -1340
rect 3200 -1440 3400 -1340
rect 3520 -1440 3720 -1340
rect 3840 -1440 4040 -1340
rect 4160 -1440 4360 -1340
rect 4480 -1440 4680 -1340
rect 4800 -1440 5000 -1340
<< mvpmos >>
rect 0 380 200 680
rect 320 380 520 680
rect 640 380 840 680
rect 960 380 1160 680
rect 1280 380 1480 680
rect 1600 380 1800 680
rect 1920 380 2120 680
rect 2240 380 2440 680
rect 2560 380 2760 680
rect 2880 380 3080 680
rect 3200 380 3400 680
rect 3520 380 3720 680
rect 3840 380 4040 680
rect 4160 380 4360 680
rect 4480 380 4680 680
rect 4800 380 5000 680
rect 0 -20 200 280
rect 320 -20 520 280
rect 640 -20 840 280
rect 960 -20 1160 280
rect 1280 -20 1480 280
rect 1600 -20 1800 280
rect 1920 -20 2120 280
rect 2240 -20 2440 280
rect 2560 -20 2760 280
rect 2880 -20 3080 280
rect 3200 -20 3400 280
rect 3520 -20 3720 280
rect 3840 -20 4040 280
rect 4160 -20 4360 280
rect 4480 -20 4680 280
rect 4800 -20 5000 280
rect 0 -740 200 -440
rect 320 -740 520 -440
rect 640 -740 840 -440
rect 960 -740 1160 -440
rect 1280 -740 1480 -440
rect 1600 -740 1800 -440
rect 1920 -740 2120 -440
rect 2240 -740 2440 -440
rect 2560 -740 2760 -440
rect 2880 -740 3080 -440
rect 3200 -740 3400 -440
rect 3520 -740 3720 -440
rect 3840 -740 4040 -440
rect 4160 -740 4360 -440
rect 4480 -740 4680 -440
rect 4800 -740 5000 -440
<< mvndiff >>
rect -80 -1150 0 -1140
rect -80 -1230 -75 -1150
rect -45 -1230 0 -1150
rect -80 -1240 0 -1230
rect 200 -1150 320 -1140
rect 200 -1230 245 -1150
rect 275 -1230 320 -1150
rect 200 -1240 320 -1230
rect 520 -1150 640 -1140
rect 520 -1230 565 -1150
rect 595 -1230 640 -1150
rect 520 -1240 640 -1230
rect 840 -1150 960 -1140
rect 840 -1230 885 -1150
rect 915 -1230 960 -1150
rect 840 -1240 960 -1230
rect 1160 -1150 1280 -1140
rect 1160 -1230 1205 -1150
rect 1235 -1230 1280 -1150
rect 1160 -1240 1280 -1230
rect 1480 -1150 1600 -1140
rect 1480 -1230 1525 -1150
rect 1555 -1230 1600 -1150
rect 1480 -1240 1600 -1230
rect 1800 -1150 1920 -1140
rect 1800 -1230 1845 -1150
rect 1875 -1230 1920 -1150
rect 1800 -1240 1920 -1230
rect 2120 -1150 2240 -1140
rect 2120 -1230 2165 -1150
rect 2195 -1230 2240 -1150
rect 2120 -1240 2240 -1230
rect 2440 -1150 2560 -1140
rect 2440 -1230 2485 -1150
rect 2515 -1230 2560 -1150
rect 2440 -1240 2560 -1230
rect 2760 -1150 2880 -1140
rect 2760 -1230 2805 -1150
rect 2835 -1230 2880 -1150
rect 2760 -1240 2880 -1230
rect 3080 -1150 3200 -1140
rect 3080 -1230 3125 -1150
rect 3155 -1230 3200 -1150
rect 3080 -1240 3200 -1230
rect 3400 -1150 3520 -1140
rect 3400 -1230 3445 -1150
rect 3475 -1230 3520 -1150
rect 3400 -1240 3520 -1230
rect 3720 -1150 3840 -1140
rect 3720 -1230 3765 -1150
rect 3795 -1230 3840 -1150
rect 3720 -1240 3840 -1230
rect 4040 -1150 4160 -1140
rect 4040 -1230 4085 -1150
rect 4115 -1230 4160 -1150
rect 4040 -1240 4160 -1230
rect 4360 -1150 4480 -1140
rect 4360 -1230 4405 -1150
rect 4435 -1230 4480 -1150
rect 4360 -1240 4480 -1230
rect 4680 -1150 4800 -1140
rect 4680 -1230 4725 -1150
rect 4755 -1230 4800 -1150
rect 4680 -1240 4800 -1230
rect 5000 -1150 5080 -1140
rect 5000 -1230 5045 -1150
rect 5075 -1230 5080 -1150
rect 5000 -1240 5080 -1230
rect -80 -1350 0 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 0 -1350
rect -80 -1440 0 -1430
rect 200 -1350 320 -1340
rect 200 -1430 245 -1350
rect 275 -1430 320 -1350
rect 200 -1440 320 -1430
rect 520 -1350 640 -1340
rect 520 -1430 565 -1350
rect 595 -1430 640 -1350
rect 520 -1440 640 -1430
rect 840 -1350 960 -1340
rect 840 -1430 885 -1350
rect 915 -1430 960 -1350
rect 840 -1440 960 -1430
rect 1160 -1350 1280 -1340
rect 1160 -1430 1205 -1350
rect 1235 -1430 1280 -1350
rect 1160 -1440 1280 -1430
rect 1480 -1350 1600 -1340
rect 1480 -1430 1525 -1350
rect 1555 -1430 1600 -1350
rect 1480 -1440 1600 -1430
rect 1800 -1350 1920 -1340
rect 1800 -1430 1845 -1350
rect 1875 -1430 1920 -1350
rect 1800 -1440 1920 -1430
rect 2120 -1350 2240 -1340
rect 2120 -1430 2165 -1350
rect 2195 -1430 2240 -1350
rect 2120 -1440 2240 -1430
rect 2440 -1350 2560 -1340
rect 2440 -1430 2485 -1350
rect 2515 -1430 2560 -1350
rect 2440 -1440 2560 -1430
rect 2760 -1350 2880 -1340
rect 2760 -1430 2805 -1350
rect 2835 -1430 2880 -1350
rect 2760 -1440 2880 -1430
rect 3080 -1350 3200 -1340
rect 3080 -1430 3125 -1350
rect 3155 -1430 3200 -1350
rect 3080 -1440 3200 -1430
rect 3400 -1350 3520 -1340
rect 3400 -1430 3445 -1350
rect 3475 -1430 3520 -1350
rect 3400 -1440 3520 -1430
rect 3720 -1350 3840 -1340
rect 3720 -1430 3765 -1350
rect 3795 -1430 3840 -1350
rect 3720 -1440 3840 -1430
rect 4040 -1350 4160 -1340
rect 4040 -1430 4085 -1350
rect 4115 -1430 4160 -1350
rect 4040 -1440 4160 -1430
rect 4360 -1350 4480 -1340
rect 4360 -1430 4405 -1350
rect 4435 -1430 4480 -1350
rect 4360 -1440 4480 -1430
rect 4680 -1350 4800 -1340
rect 4680 -1430 4725 -1350
rect 4755 -1430 4800 -1350
rect 4680 -1440 4800 -1430
rect 5000 -1350 5080 -1340
rect 5000 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5000 -1440 5080 -1430
<< mvpdiff >>
rect -80 670 0 680
rect -80 390 -75 670
rect -45 390 0 670
rect -80 380 0 390
rect 200 670 320 680
rect 200 390 245 670
rect 275 390 320 670
rect 200 380 320 390
rect 520 670 640 680
rect 520 390 565 670
rect 595 390 640 670
rect 520 380 640 390
rect 840 670 960 680
rect 840 390 885 670
rect 915 390 960 670
rect 840 380 960 390
rect 1160 670 1280 680
rect 1160 390 1205 670
rect 1235 390 1280 670
rect 1160 380 1280 390
rect 1480 670 1600 680
rect 1480 390 1525 670
rect 1555 390 1600 670
rect 1480 380 1600 390
rect 1800 670 1920 680
rect 1800 390 1845 670
rect 1875 390 1920 670
rect 1800 380 1920 390
rect 2120 670 2240 680
rect 2120 390 2165 670
rect 2195 390 2240 670
rect 2120 380 2240 390
rect 2440 670 2560 680
rect 2440 390 2485 670
rect 2515 390 2560 670
rect 2440 380 2560 390
rect 2760 670 2880 680
rect 2760 390 2805 670
rect 2835 390 2880 670
rect 2760 380 2880 390
rect 3080 670 3200 680
rect 3080 390 3125 670
rect 3155 390 3200 670
rect 3080 380 3200 390
rect 3400 670 3520 680
rect 3400 390 3445 670
rect 3475 390 3520 670
rect 3400 380 3520 390
rect 3720 670 3840 680
rect 3720 390 3765 670
rect 3795 390 3840 670
rect 3720 380 3840 390
rect 4040 670 4160 680
rect 4040 390 4085 670
rect 4115 390 4160 670
rect 4040 380 4160 390
rect 4360 670 4480 680
rect 4360 390 4405 670
rect 4435 390 4480 670
rect 4360 380 4480 390
rect 4680 670 4800 680
rect 4680 390 4725 670
rect 4755 390 4800 670
rect 4680 380 4800 390
rect 5000 670 5080 680
rect 5000 390 5045 670
rect 5075 390 5080 670
rect 5000 380 5080 390
rect -80 270 0 280
rect -80 -10 -75 270
rect -45 -10 0 270
rect -80 -20 0 -10
rect 200 270 320 280
rect 200 -10 245 270
rect 275 -10 320 270
rect 200 -20 320 -10
rect 520 270 640 280
rect 520 -10 565 270
rect 595 -10 640 270
rect 520 -20 640 -10
rect 840 270 960 280
rect 840 -10 885 270
rect 915 -10 960 270
rect 840 -20 960 -10
rect 1160 270 1280 280
rect 1160 -10 1205 270
rect 1235 -10 1280 270
rect 1160 -20 1280 -10
rect 1480 270 1600 280
rect 1480 -10 1525 270
rect 1555 -10 1600 270
rect 1480 -20 1600 -10
rect 1800 270 1920 280
rect 1800 -10 1845 270
rect 1875 -10 1920 270
rect 1800 -20 1920 -10
rect 2120 270 2240 280
rect 2120 -10 2165 270
rect 2195 -10 2240 270
rect 2120 -20 2240 -10
rect 2440 270 2560 280
rect 2440 -10 2485 270
rect 2515 -10 2560 270
rect 2440 -20 2560 -10
rect 2760 270 2880 280
rect 2760 -10 2805 270
rect 2835 -10 2880 270
rect 2760 -20 2880 -10
rect 3080 270 3200 280
rect 3080 -10 3125 270
rect 3155 -10 3200 270
rect 3080 -20 3200 -10
rect 3400 270 3520 280
rect 3400 -10 3445 270
rect 3475 -10 3520 270
rect 3400 -20 3520 -10
rect 3720 270 3840 280
rect 3720 -10 3765 270
rect 3795 -10 3840 270
rect 3720 -20 3840 -10
rect 4040 270 4160 280
rect 4040 -10 4085 270
rect 4115 -10 4160 270
rect 4040 -20 4160 -10
rect 4360 270 4480 280
rect 4360 -10 4405 270
rect 4435 -10 4480 270
rect 4360 -20 4480 -10
rect 4680 270 4800 280
rect 4680 -10 4725 270
rect 4755 -10 4800 270
rect 4680 -20 4800 -10
rect 5000 270 5080 280
rect 5000 -10 5045 270
rect 5075 -10 5080 270
rect 5000 -20 5080 -10
rect -80 -450 0 -440
rect -80 -730 -75 -450
rect -45 -730 0 -450
rect -80 -740 0 -730
rect 200 -450 320 -440
rect 200 -730 245 -450
rect 275 -730 320 -450
rect 200 -740 320 -730
rect 520 -450 640 -440
rect 520 -730 565 -450
rect 595 -730 640 -450
rect 520 -740 640 -730
rect 840 -450 960 -440
rect 840 -730 885 -450
rect 915 -730 960 -450
rect 840 -740 960 -730
rect 1160 -450 1280 -440
rect 1160 -730 1205 -450
rect 1235 -730 1280 -450
rect 1160 -740 1280 -730
rect 1480 -450 1600 -440
rect 1480 -730 1525 -450
rect 1555 -730 1600 -450
rect 1480 -740 1600 -730
rect 1800 -450 1920 -440
rect 1800 -730 1845 -450
rect 1875 -730 1920 -450
rect 1800 -740 1920 -730
rect 2120 -450 2240 -440
rect 2120 -730 2165 -450
rect 2195 -730 2240 -450
rect 2120 -740 2240 -730
rect 2440 -450 2560 -440
rect 2440 -730 2485 -450
rect 2515 -730 2560 -450
rect 2440 -740 2560 -730
rect 2760 -450 2880 -440
rect 2760 -730 2805 -450
rect 2835 -730 2880 -450
rect 2760 -740 2880 -730
rect 3080 -450 3200 -440
rect 3080 -730 3125 -450
rect 3155 -730 3200 -450
rect 3080 -740 3200 -730
rect 3400 -450 3520 -440
rect 3400 -730 3445 -450
rect 3475 -730 3520 -450
rect 3400 -740 3520 -730
rect 3720 -450 3840 -440
rect 3720 -730 3765 -450
rect 3795 -730 3840 -450
rect 3720 -740 3840 -730
rect 4040 -450 4160 -440
rect 4040 -730 4085 -450
rect 4115 -730 4160 -450
rect 4040 -740 4160 -730
rect 4360 -450 4480 -440
rect 4360 -730 4405 -450
rect 4435 -730 4480 -450
rect 4360 -740 4480 -730
rect 4680 -450 4800 -440
rect 4680 -730 4725 -450
rect 4755 -730 4800 -450
rect 4680 -740 4800 -730
rect 5000 -450 5080 -440
rect 5000 -730 5045 -450
rect 5075 -730 5080 -450
rect 5000 -740 5080 -730
<< mvndiffc >>
rect -75 -1230 -45 -1150
rect 245 -1230 275 -1150
rect 565 -1230 595 -1150
rect 885 -1230 915 -1150
rect 1205 -1230 1235 -1150
rect 1525 -1230 1555 -1150
rect 1845 -1230 1875 -1150
rect 2165 -1230 2195 -1150
rect 2485 -1230 2515 -1150
rect 2805 -1230 2835 -1150
rect 3125 -1230 3155 -1150
rect 3445 -1230 3475 -1150
rect 3765 -1230 3795 -1150
rect 4085 -1230 4115 -1150
rect 4405 -1230 4435 -1150
rect 4725 -1230 4755 -1150
rect 5045 -1230 5075 -1150
rect -75 -1430 -45 -1350
rect 245 -1430 275 -1350
rect 565 -1430 595 -1350
rect 885 -1430 915 -1350
rect 1205 -1430 1235 -1350
rect 1525 -1430 1555 -1350
rect 1845 -1430 1875 -1350
rect 2165 -1430 2195 -1350
rect 2485 -1430 2515 -1350
rect 2805 -1430 2835 -1350
rect 3125 -1430 3155 -1350
rect 3445 -1430 3475 -1350
rect 3765 -1430 3795 -1350
rect 4085 -1430 4115 -1350
rect 4405 -1430 4435 -1350
rect 4725 -1430 4755 -1350
rect 5045 -1430 5075 -1350
<< mvpdiffc >>
rect -75 390 -45 670
rect 245 390 275 670
rect 565 390 595 670
rect 885 390 915 670
rect 1205 390 1235 670
rect 1525 390 1555 670
rect 1845 390 1875 670
rect 2165 390 2195 670
rect 2485 390 2515 670
rect 2805 390 2835 670
rect 3125 390 3155 670
rect 3445 390 3475 670
rect 3765 390 3795 670
rect 4085 390 4115 670
rect 4405 390 4435 670
rect 4725 390 4755 670
rect 5045 390 5075 670
rect -75 -10 -45 270
rect 245 -10 275 270
rect 565 -10 595 270
rect 885 -10 915 270
rect 1205 -10 1235 270
rect 1525 -10 1555 270
rect 1845 -10 1875 270
rect 2165 -10 2195 270
rect 2485 -10 2515 270
rect 2805 -10 2835 270
rect 3125 -10 3155 270
rect 3445 -10 3475 270
rect 3765 -10 3795 270
rect 4085 -10 4115 270
rect 4405 -10 4435 270
rect 4725 -10 4755 270
rect 5045 -10 5075 270
rect -75 -730 -45 -450
rect 245 -730 275 -450
rect 565 -730 595 -450
rect 885 -730 915 -450
rect 1205 -730 1235 -450
rect 1525 -730 1555 -450
rect 1845 -730 1875 -450
rect 2165 -730 2195 -450
rect 2485 -730 2515 -450
rect 2805 -730 2835 -450
rect 3125 -730 3155 -450
rect 3445 -730 3475 -450
rect 3765 -730 3795 -450
rect 4085 -730 4115 -450
rect 4405 -730 4435 -450
rect 4725 -730 4755 -450
rect 5045 -730 5075 -450
<< psubdiff >>
rect -240 800 -180 840
rect 5180 800 5240 840
rect -240 780 -200 800
rect 5200 780 5240 800
rect -200 -240 -180 -200
rect 5180 -240 5200 -200
rect -240 -280 -200 -240
rect 5200 -280 5240 -240
rect -200 -320 -180 -280
rect 5180 -320 5200 -280
rect -200 -960 -180 -920
rect 5180 -960 5200 -920
rect -200 -1040 -180 -1000
rect 5180 -1040 5200 -1000
rect -240 -1480 -200 -1460
rect 5200 -1480 5240 -1460
rect -240 -1520 -180 -1480
rect 5180 -1520 5240 -1480
<< nsubdiff >>
rect -160 720 -100 760
rect 5100 720 5160 760
rect -160 700 -120 720
rect 5120 700 5160 720
rect -160 -120 -120 -100
rect 5120 -120 5160 -100
rect -160 -160 -100 -120
rect 5100 -160 5160 -120
rect -160 -400 -100 -360
rect 5100 -400 5160 -360
rect -160 -420 -120 -400
rect 5120 -420 5160 -400
rect -160 -840 -120 -820
rect 5120 -840 5160 -820
rect -160 -880 -100 -840
rect 5100 -880 5160 -840
<< psubdiffcont >>
rect -180 800 5180 840
rect -240 -240 -200 780
rect -180 -240 5180 -200
rect 5200 -240 5240 780
rect -240 -1460 -200 -280
rect -180 -320 5180 -280
rect -180 -960 5180 -920
rect -180 -1040 5180 -1000
rect 5200 -1460 5240 -280
rect -180 -1520 5180 -1480
<< nsubdiffcont >>
rect -100 720 5100 760
rect -160 -100 -120 700
rect 5120 -100 5160 700
rect -100 -160 5100 -120
rect -100 -400 5100 -360
rect -160 -820 -120 -420
rect 5120 -820 5160 -420
rect -100 -880 5100 -840
<< poly >>
rect 0 680 200 700
rect 320 680 520 700
rect 640 680 840 700
rect 960 680 1160 700
rect 1280 680 1480 700
rect 1600 680 1800 700
rect 1920 680 2120 700
rect 2240 680 2440 700
rect 2560 680 2760 700
rect 2880 680 3080 700
rect 3200 680 3400 700
rect 3520 680 3720 700
rect 3840 680 4040 700
rect 4160 680 4360 700
rect 4480 680 4680 700
rect 4800 680 5000 700
rect 0 280 200 380
rect 320 280 520 380
rect 640 280 840 380
rect 960 280 1160 380
rect 1280 280 1480 380
rect 1600 280 1800 380
rect 1920 280 2120 380
rect 2240 280 2440 380
rect 2560 280 2760 380
rect 2880 280 3080 380
rect 3200 280 3400 380
rect 3520 280 3720 380
rect 3840 280 4040 380
rect 4160 280 4360 380
rect 4480 280 4680 380
rect 4800 280 5000 380
rect 0 -45 200 -20
rect 0 -75 10 -45
rect 190 -75 200 -45
rect 0 -80 200 -75
rect 320 -45 520 -20
rect 320 -75 330 -45
rect 510 -75 520 -45
rect 320 -80 520 -75
rect 640 -45 840 -20
rect 640 -75 650 -45
rect 830 -75 840 -45
rect 640 -80 840 -75
rect 960 -45 1160 -20
rect 960 -75 970 -45
rect 1150 -75 1160 -45
rect 960 -80 1160 -75
rect 1280 -45 1480 -20
rect 1280 -75 1290 -45
rect 1470 -75 1480 -45
rect 1280 -80 1480 -75
rect 1600 -45 1800 -20
rect 1600 -75 1610 -45
rect 1790 -75 1800 -45
rect 1600 -80 1800 -75
rect 1920 -45 2120 -20
rect 1920 -75 1930 -45
rect 2110 -75 2120 -45
rect 1920 -80 2120 -75
rect 2240 -45 2440 -20
rect 2240 -75 2250 -45
rect 2430 -75 2440 -45
rect 2240 -80 2440 -75
rect 2560 -45 2760 -20
rect 2560 -75 2570 -45
rect 2750 -75 2760 -45
rect 2560 -80 2760 -75
rect 2880 -45 3080 -20
rect 2880 -75 2890 -45
rect 3070 -75 3080 -45
rect 2880 -80 3080 -75
rect 3200 -45 3400 -20
rect 3200 -75 3210 -45
rect 3390 -75 3400 -45
rect 3200 -80 3400 -75
rect 3520 -45 3720 -20
rect 3520 -75 3530 -45
rect 3710 -75 3720 -45
rect 3520 -80 3720 -75
rect 3840 -45 4040 -20
rect 3840 -75 3850 -45
rect 4030 -75 4040 -45
rect 3840 -80 4040 -75
rect 4160 -45 4360 -20
rect 4160 -75 4170 -45
rect 4350 -75 4360 -45
rect 4160 -80 4360 -75
rect 4480 -45 4680 -20
rect 4480 -75 4490 -45
rect 4670 -75 4680 -45
rect 4480 -80 4680 -75
rect 4800 -45 5000 -20
rect 4800 -75 4810 -45
rect 4990 -75 5000 -45
rect 4800 -80 5000 -75
rect 0 -440 200 -420
rect 320 -440 520 -420
rect 640 -440 840 -420
rect 960 -440 1160 -420
rect 1280 -440 1480 -420
rect 1600 -440 1800 -420
rect 1920 -440 2120 -420
rect 2240 -440 2440 -420
rect 2560 -440 2760 -420
rect 2880 -440 3080 -420
rect 3200 -440 3400 -420
rect 3520 -440 3720 -420
rect 3840 -440 4040 -420
rect 4160 -440 4360 -420
rect 4480 -440 4680 -420
rect 4800 -440 5000 -420
rect 0 -765 200 -740
rect 0 -795 10 -765
rect 190 -795 200 -765
rect 0 -800 200 -795
rect 320 -765 520 -740
rect 320 -795 330 -765
rect 510 -795 520 -765
rect 320 -800 520 -795
rect 640 -765 840 -740
rect 640 -795 650 -765
rect 830 -795 840 -765
rect 640 -800 840 -795
rect 960 -765 1160 -740
rect 960 -795 970 -765
rect 1150 -795 1160 -765
rect 960 -800 1160 -795
rect 1280 -765 1480 -740
rect 1280 -795 1290 -765
rect 1470 -795 1480 -765
rect 1280 -800 1480 -795
rect 1600 -765 1800 -740
rect 1600 -795 1610 -765
rect 1790 -795 1800 -765
rect 1600 -800 1800 -795
rect 1920 -765 2120 -740
rect 1920 -795 1930 -765
rect 2110 -795 2120 -765
rect 1920 -800 2120 -795
rect 2240 -765 2440 -740
rect 2240 -795 2250 -765
rect 2430 -795 2440 -765
rect 2240 -800 2440 -795
rect 2560 -765 2760 -740
rect 2560 -795 2570 -765
rect 2750 -795 2760 -765
rect 2560 -800 2760 -795
rect 2880 -765 3080 -740
rect 2880 -795 2890 -765
rect 3070 -795 3080 -765
rect 2880 -800 3080 -795
rect 3200 -765 3400 -740
rect 3200 -795 3210 -765
rect 3390 -795 3400 -765
rect 3200 -800 3400 -795
rect 3520 -765 3720 -740
rect 3520 -795 3530 -765
rect 3710 -795 3720 -765
rect 3520 -800 3720 -795
rect 3840 -765 4040 -740
rect 3840 -795 3850 -765
rect 4030 -795 4040 -765
rect 3840 -800 4040 -795
rect 4160 -765 4360 -740
rect 4160 -795 4170 -765
rect 4350 -795 4360 -765
rect 4160 -800 4360 -795
rect 4480 -765 4680 -740
rect 4480 -795 4490 -765
rect 4670 -795 4680 -765
rect 4480 -800 4680 -795
rect 4800 -765 5000 -740
rect 4800 -795 4810 -765
rect 4990 -795 5000 -765
rect 4800 -800 5000 -795
rect 0 -1085 200 -1080
rect 0 -1115 10 -1085
rect 190 -1115 200 -1085
rect 0 -1140 200 -1115
rect 320 -1085 520 -1080
rect 320 -1115 330 -1085
rect 510 -1115 520 -1085
rect 320 -1140 520 -1115
rect 640 -1085 840 -1080
rect 640 -1115 650 -1085
rect 830 -1115 840 -1085
rect 640 -1140 840 -1115
rect 960 -1085 1160 -1080
rect 960 -1115 970 -1085
rect 1150 -1115 1160 -1085
rect 960 -1140 1160 -1115
rect 1280 -1085 1480 -1080
rect 1280 -1115 1290 -1085
rect 1470 -1115 1480 -1085
rect 1280 -1140 1480 -1115
rect 1600 -1085 1800 -1080
rect 1600 -1115 1610 -1085
rect 1790 -1115 1800 -1085
rect 1600 -1140 1800 -1115
rect 1920 -1085 2120 -1080
rect 1920 -1115 1930 -1085
rect 2110 -1115 2120 -1085
rect 1920 -1140 2120 -1115
rect 2240 -1085 2440 -1080
rect 2240 -1115 2250 -1085
rect 2430 -1115 2440 -1085
rect 2240 -1140 2440 -1115
rect 2560 -1085 2760 -1080
rect 2560 -1115 2570 -1085
rect 2750 -1115 2760 -1085
rect 2560 -1140 2760 -1115
rect 2880 -1085 3080 -1080
rect 2880 -1115 2890 -1085
rect 3070 -1115 3080 -1085
rect 2880 -1140 3080 -1115
rect 3200 -1085 3400 -1080
rect 3200 -1115 3210 -1085
rect 3390 -1115 3400 -1085
rect 3200 -1140 3400 -1115
rect 3520 -1085 3720 -1080
rect 3520 -1115 3530 -1085
rect 3710 -1115 3720 -1085
rect 3520 -1140 3720 -1115
rect 3840 -1085 4040 -1080
rect 3840 -1115 3850 -1085
rect 4030 -1115 4040 -1085
rect 3840 -1140 4040 -1115
rect 4160 -1085 4360 -1080
rect 4160 -1115 4170 -1085
rect 4350 -1115 4360 -1085
rect 4160 -1140 4360 -1115
rect 4480 -1085 4680 -1080
rect 4480 -1115 4490 -1085
rect 4670 -1115 4680 -1085
rect 4480 -1140 4680 -1115
rect 4800 -1085 5000 -1080
rect 4800 -1115 4810 -1085
rect 4990 -1115 5000 -1085
rect 4800 -1140 5000 -1115
rect 0 -1340 200 -1240
rect 320 -1340 520 -1240
rect 640 -1340 840 -1240
rect 960 -1340 1160 -1240
rect 1280 -1340 1480 -1240
rect 1600 -1340 1800 -1240
rect 1920 -1340 2120 -1240
rect 2240 -1340 2440 -1240
rect 2560 -1340 2760 -1240
rect 2880 -1340 3080 -1240
rect 3200 -1340 3400 -1240
rect 3520 -1340 3720 -1240
rect 3840 -1340 4040 -1240
rect 4160 -1340 4360 -1240
rect 4480 -1340 4680 -1240
rect 4800 -1340 5000 -1240
rect 0 -1460 200 -1440
rect 320 -1460 520 -1440
rect 640 -1460 840 -1440
rect 960 -1460 1160 -1440
rect 1280 -1460 1480 -1440
rect 1600 -1460 1800 -1440
rect 1920 -1460 2120 -1440
rect 2240 -1460 2440 -1440
rect 2560 -1460 2760 -1440
rect 2880 -1460 3080 -1440
rect 3200 -1460 3400 -1440
rect 3520 -1460 3720 -1440
rect 3840 -1460 4040 -1440
rect 4160 -1460 4360 -1440
rect 4480 -1460 4680 -1440
rect 4800 -1460 5000 -1440
<< polycont >>
rect 10 -75 190 -45
rect 330 -75 510 -45
rect 650 -75 830 -45
rect 970 -75 1150 -45
rect 1290 -75 1470 -45
rect 1610 -75 1790 -45
rect 1930 -75 2110 -45
rect 2250 -75 2430 -45
rect 2570 -75 2750 -45
rect 2890 -75 3070 -45
rect 3210 -75 3390 -45
rect 3530 -75 3710 -45
rect 3850 -75 4030 -45
rect 4170 -75 4350 -45
rect 4490 -75 4670 -45
rect 4810 -75 4990 -45
rect 10 -795 190 -765
rect 330 -795 510 -765
rect 650 -795 830 -765
rect 970 -795 1150 -765
rect 1290 -795 1470 -765
rect 1610 -795 1790 -765
rect 1930 -795 2110 -765
rect 2250 -795 2430 -765
rect 2570 -795 2750 -765
rect 2890 -795 3070 -765
rect 3210 -795 3390 -765
rect 3530 -795 3710 -765
rect 3850 -795 4030 -765
rect 4170 -795 4350 -765
rect 4490 -795 4670 -765
rect 4810 -795 4990 -765
rect 10 -1115 190 -1085
rect 330 -1115 510 -1085
rect 650 -1115 830 -1085
rect 970 -1115 1150 -1085
rect 1290 -1115 1470 -1085
rect 1610 -1115 1790 -1085
rect 1930 -1115 2110 -1085
rect 2250 -1115 2430 -1085
rect 2570 -1115 2750 -1085
rect 2890 -1115 3070 -1085
rect 3210 -1115 3390 -1085
rect 3530 -1115 3710 -1085
rect 3850 -1115 4030 -1085
rect 4170 -1115 4350 -1085
rect 4490 -1115 4670 -1085
rect 4810 -1115 4990 -1085
<< locali >>
rect -240 800 -180 840
rect 5180 800 5240 840
rect -240 780 -200 800
rect 5200 780 5240 800
rect -160 720 -100 760
rect 5100 720 5160 760
rect -160 700 -120 720
rect -80 670 -40 720
rect -80 390 -75 670
rect -45 390 -40 670
rect -80 380 -40 390
rect 240 670 280 680
rect 240 390 245 670
rect 275 390 280 670
rect 240 380 280 390
rect 560 670 600 680
rect 560 390 565 670
rect 595 390 600 670
rect 560 360 600 390
rect 880 670 920 680
rect 880 390 885 670
rect 915 390 920 670
rect 880 380 920 390
rect 1200 670 1240 720
rect 1200 390 1205 670
rect 1235 390 1240 670
rect 1200 380 1240 390
rect 1520 670 1560 680
rect 1520 390 1525 670
rect 1555 390 1560 670
rect 1520 380 1560 390
rect 1840 670 1880 680
rect 1840 390 1845 670
rect 1875 390 1880 670
rect 1840 360 1880 390
rect 2160 670 2200 680
rect 2160 390 2165 670
rect 2195 390 2200 670
rect 2160 380 2200 390
rect 2480 670 2520 720
rect 2480 390 2485 670
rect 2515 390 2520 670
rect 2480 380 2520 390
rect 2800 670 2840 680
rect 2800 390 2805 670
rect 2835 390 2840 670
rect 2800 380 2840 390
rect 3120 670 3160 680
rect 3120 390 3125 670
rect 3155 390 3160 670
rect 3120 360 3160 390
rect 3440 670 3480 680
rect 3440 390 3445 670
rect 3475 390 3480 670
rect 3440 380 3480 390
rect 3760 670 3800 720
rect 3760 390 3765 670
rect 3795 390 3800 670
rect 3760 380 3800 390
rect 4080 670 4120 680
rect 4080 390 4085 670
rect 4115 390 4120 670
rect 4080 380 4120 390
rect 4400 670 4440 680
rect 4400 390 4405 670
rect 4435 390 4440 670
rect 4400 360 4440 390
rect 4720 670 4760 680
rect 4720 390 4725 670
rect 4755 390 4760 670
rect 4720 380 4760 390
rect 5040 670 5080 720
rect 5040 390 5045 670
rect 5075 390 5080 670
rect 5040 380 5080 390
rect 5120 700 5160 720
rect -80 320 5080 360
rect -80 270 -40 320
rect -80 -10 -75 270
rect -45 -10 -40 270
rect -80 -20 -40 -10
rect 240 270 280 280
rect 240 -10 245 270
rect 275 -10 280 270
rect 240 -20 280 -10
rect 560 270 600 320
rect 560 -10 565 270
rect 595 -10 600 270
rect 560 -20 600 -10
rect 880 270 920 280
rect 880 -10 885 270
rect 915 -10 920 270
rect 880 -20 920 -10
rect 1200 270 1240 320
rect 1200 -10 1205 270
rect 1235 -10 1240 270
rect 1200 -20 1240 -10
rect 1520 270 1560 280
rect 1520 -10 1525 270
rect 1555 -10 1560 270
rect 1520 -20 1560 -10
rect 1840 270 1880 320
rect 1840 -10 1845 270
rect 1875 -10 1880 270
rect 1840 -20 1880 -10
rect 2160 270 2200 280
rect 2160 -10 2165 270
rect 2195 -10 2200 270
rect 2160 -20 2200 -10
rect 2480 270 2520 320
rect 2480 -10 2485 270
rect 2515 -10 2520 270
rect 2480 -20 2520 -10
rect 2800 270 2840 280
rect 2800 -10 2805 270
rect 2835 -10 2840 270
rect 2800 -20 2840 -10
rect 3120 270 3160 320
rect 3120 -10 3125 270
rect 3155 -10 3160 270
rect 3120 -20 3160 -10
rect 3440 270 3480 280
rect 3440 -10 3445 270
rect 3475 -10 3480 270
rect 3440 -20 3480 -10
rect 3760 270 3800 320
rect 3760 -10 3765 270
rect 3795 -10 3800 270
rect 3760 -20 3800 -10
rect 4080 270 4120 280
rect 4080 -10 4085 270
rect 4115 -10 4120 270
rect 4080 -20 4120 -10
rect 4400 270 4440 320
rect 4400 -10 4405 270
rect 4435 -10 4440 270
rect 4400 -20 4440 -10
rect 4720 270 4760 280
rect 4720 -10 4725 270
rect 4755 -10 4760 270
rect 4720 -20 4760 -10
rect 5040 270 5080 320
rect 5040 -10 5045 270
rect 5075 -10 5080 270
rect 5040 -20 5080 -10
rect 0 -45 200 -40
rect 0 -75 10 -45
rect 190 -75 200 -45
rect 0 -80 200 -75
rect 320 -45 520 -40
rect 320 -75 330 -45
rect 510 -75 520 -45
rect 320 -80 520 -75
rect 640 -45 840 -40
rect 640 -75 650 -45
rect 830 -75 840 -45
rect 640 -80 840 -75
rect 960 -45 1160 -40
rect 960 -75 970 -45
rect 1150 -75 1160 -45
rect 960 -80 1160 -75
rect 1280 -45 1480 -40
rect 1280 -75 1290 -45
rect 1470 -75 1480 -45
rect 1280 -80 1480 -75
rect 1600 -45 1800 -40
rect 1600 -75 1610 -45
rect 1790 -75 1800 -45
rect 1600 -80 1800 -75
rect 1920 -45 2120 -40
rect 1920 -75 1930 -45
rect 2110 -75 2120 -45
rect 1920 -80 2120 -75
rect 2240 -45 2440 -40
rect 2240 -75 2250 -45
rect 2430 -75 2440 -45
rect 2240 -80 2440 -75
rect 2560 -45 2760 -40
rect 2560 -75 2570 -45
rect 2750 -75 2760 -45
rect 2560 -80 2760 -75
rect 2880 -45 3080 -40
rect 2880 -75 2890 -45
rect 3070 -75 3080 -45
rect 2880 -80 3080 -75
rect 3200 -45 3400 -40
rect 3200 -75 3210 -45
rect 3390 -75 3400 -45
rect 3200 -80 3400 -75
rect 3520 -45 3720 -40
rect 3520 -75 3530 -45
rect 3710 -75 3720 -45
rect 3520 -80 3720 -75
rect 3840 -45 4040 -40
rect 3840 -75 3850 -45
rect 4030 -75 4040 -45
rect 3840 -80 4040 -75
rect 4160 -45 4360 -40
rect 4160 -75 4170 -45
rect 4350 -75 4360 -45
rect 4160 -80 4360 -75
rect 4480 -45 4680 -40
rect 4480 -75 4490 -45
rect 4670 -75 4680 -45
rect 4480 -80 4680 -75
rect 4800 -45 5000 -40
rect 4800 -75 4810 -45
rect 4990 -75 5000 -45
rect 4800 -80 5000 -75
rect -160 -120 -120 -100
rect 5120 -120 5160 -100
rect -160 -160 -100 -120
rect 5100 -160 5160 -120
rect -200 -240 -180 -200
rect 5180 -240 5200 -200
rect -240 -280 -200 -240
rect 5200 -280 5240 -240
rect -200 -320 -180 -280
rect 5180 -320 5200 -280
rect -160 -400 -100 -360
rect 5100 -400 5160 -360
rect -160 -420 -120 -400
rect -80 -450 -40 -440
rect -80 -730 -75 -450
rect -45 -730 -40 -450
rect -80 -740 -40 -730
rect 240 -450 280 -400
rect 240 -730 245 -450
rect 275 -730 280 -450
rect 240 -740 280 -730
rect 560 -450 600 -440
rect 560 -730 565 -450
rect 595 -730 600 -450
rect 560 -740 600 -730
rect 880 -450 920 -400
rect 880 -730 885 -450
rect 915 -730 920 -450
rect 880 -740 920 -730
rect 1200 -450 1240 -440
rect 1200 -730 1205 -450
rect 1235 -730 1240 -450
rect 1200 -740 1240 -730
rect 1520 -450 1560 -400
rect 1520 -730 1525 -450
rect 1555 -730 1560 -450
rect 1520 -740 1560 -730
rect 1840 -450 1880 -440
rect 1840 -730 1845 -450
rect 1875 -730 1880 -450
rect 1840 -740 1880 -730
rect 2160 -450 2200 -400
rect 2160 -730 2165 -450
rect 2195 -730 2200 -450
rect 2160 -740 2200 -730
rect 2480 -450 2520 -440
rect 2480 -730 2485 -450
rect 2515 -730 2520 -450
rect 2480 -740 2520 -730
rect 2800 -450 2840 -400
rect 2800 -730 2805 -450
rect 2835 -730 2840 -450
rect 2800 -740 2840 -730
rect 3120 -450 3160 -440
rect 3120 -730 3125 -450
rect 3155 -730 3160 -450
rect 3120 -740 3160 -730
rect 3440 -450 3480 -400
rect 3440 -730 3445 -450
rect 3475 -730 3480 -450
rect 3440 -740 3480 -730
rect 3760 -450 3800 -440
rect 3760 -730 3765 -450
rect 3795 -730 3800 -450
rect 3760 -740 3800 -730
rect 4080 -450 4120 -400
rect 4080 -730 4085 -450
rect 4115 -730 4120 -450
rect 4080 -740 4120 -730
rect 4400 -450 4440 -440
rect 4400 -730 4405 -450
rect 4435 -730 4440 -450
rect 4400 -740 4440 -730
rect 4720 -450 4760 -400
rect 5120 -420 5160 -400
rect 4720 -730 4725 -450
rect 4755 -730 4760 -450
rect 4720 -740 4760 -730
rect 5040 -450 5080 -440
rect 5040 -730 5045 -450
rect 5075 -730 5080 -450
rect 5040 -740 5080 -730
rect 0 -765 200 -760
rect 0 -795 10 -765
rect 190 -795 200 -765
rect 0 -800 200 -795
rect 320 -765 520 -760
rect 320 -795 330 -765
rect 510 -795 520 -765
rect 320 -800 520 -795
rect 640 -765 840 -760
rect 640 -795 650 -765
rect 830 -795 840 -765
rect 640 -800 840 -795
rect 960 -765 1160 -760
rect 960 -795 970 -765
rect 1150 -795 1160 -765
rect 960 -800 1160 -795
rect 1280 -765 1480 -760
rect 1280 -795 1290 -765
rect 1470 -795 1480 -765
rect 1280 -800 1480 -795
rect 1600 -765 1800 -760
rect 1600 -795 1610 -765
rect 1790 -795 1800 -765
rect 1600 -800 1800 -795
rect 1920 -765 2120 -760
rect 1920 -795 1930 -765
rect 2110 -795 2120 -765
rect 1920 -800 2120 -795
rect 2240 -765 2440 -760
rect 2240 -795 2250 -765
rect 2430 -795 2440 -765
rect 2240 -800 2440 -795
rect 2560 -765 2760 -760
rect 2560 -795 2570 -765
rect 2750 -795 2760 -765
rect 2560 -800 2760 -795
rect 2880 -765 3080 -760
rect 2880 -795 2890 -765
rect 3070 -795 3080 -765
rect 2880 -800 3080 -795
rect 3200 -765 3400 -760
rect 3200 -795 3210 -765
rect 3390 -795 3400 -765
rect 3200 -800 3400 -795
rect 3520 -765 3720 -760
rect 3520 -795 3530 -765
rect 3710 -795 3720 -765
rect 3520 -800 3720 -795
rect 3840 -765 4040 -760
rect 3840 -795 3850 -765
rect 4030 -795 4040 -765
rect 3840 -800 4040 -795
rect 4160 -765 4360 -760
rect 4160 -795 4170 -765
rect 4350 -795 4360 -765
rect 4160 -800 4360 -795
rect 4480 -765 4680 -760
rect 4480 -795 4490 -765
rect 4670 -795 4680 -765
rect 4480 -800 4680 -795
rect 4800 -765 5000 -760
rect 4800 -795 4810 -765
rect 4990 -795 5000 -765
rect 4800 -800 5000 -795
rect -160 -840 -120 -820
rect 5120 -840 5160 -820
rect -160 -880 -100 -840
rect 5100 -880 5160 -840
rect -200 -960 -180 -920
rect 5180 -960 5200 -920
rect -200 -1040 -180 -1000
rect 5180 -1040 5200 -1000
rect 0 -1085 200 -1080
rect 0 -1115 10 -1085
rect 190 -1115 200 -1085
rect 0 -1120 200 -1115
rect 320 -1085 520 -1080
rect 320 -1115 330 -1085
rect 510 -1115 520 -1085
rect 320 -1120 520 -1115
rect 640 -1085 840 -1080
rect 640 -1115 650 -1085
rect 830 -1115 840 -1085
rect 640 -1120 840 -1115
rect 960 -1085 1160 -1080
rect 960 -1115 970 -1085
rect 1150 -1115 1160 -1085
rect 960 -1120 1160 -1115
rect 1280 -1085 1480 -1080
rect 1280 -1115 1290 -1085
rect 1470 -1115 1480 -1085
rect 1280 -1120 1480 -1115
rect 1600 -1085 1800 -1080
rect 1600 -1115 1610 -1085
rect 1790 -1115 1800 -1085
rect 1600 -1120 1800 -1115
rect 1920 -1085 2120 -1080
rect 1920 -1115 1930 -1085
rect 2110 -1115 2120 -1085
rect 1920 -1120 2120 -1115
rect 2240 -1085 2440 -1080
rect 2240 -1115 2250 -1085
rect 2430 -1115 2440 -1085
rect 2240 -1120 2440 -1115
rect 2560 -1085 2760 -1080
rect 2560 -1115 2570 -1085
rect 2750 -1115 2760 -1085
rect 2560 -1120 2760 -1115
rect 2880 -1085 3080 -1080
rect 2880 -1115 2890 -1085
rect 3070 -1115 3080 -1085
rect 2880 -1120 3080 -1115
rect 3200 -1085 3400 -1080
rect 3200 -1115 3210 -1085
rect 3390 -1115 3400 -1085
rect 3200 -1120 3400 -1115
rect 3520 -1085 3720 -1080
rect 3520 -1115 3530 -1085
rect 3710 -1115 3720 -1085
rect 3520 -1120 3720 -1115
rect 3840 -1085 4040 -1080
rect 3840 -1115 3850 -1085
rect 4030 -1115 4040 -1085
rect 3840 -1120 4040 -1115
rect 4160 -1085 4360 -1080
rect 4160 -1115 4170 -1085
rect 4350 -1115 4360 -1085
rect 4160 -1120 4360 -1115
rect 4480 -1085 4680 -1080
rect 4480 -1115 4490 -1085
rect 4670 -1115 4680 -1085
rect 4480 -1120 4680 -1115
rect 4800 -1085 5000 -1080
rect 4800 -1115 4810 -1085
rect 4990 -1115 5000 -1085
rect 4800 -1120 5000 -1115
rect -80 -1150 -40 -1140
rect -80 -1230 -75 -1150
rect -45 -1230 -40 -1150
rect -80 -1240 -40 -1230
rect 240 -1150 280 -1140
rect 240 -1230 245 -1150
rect 275 -1230 280 -1150
rect 240 -1280 280 -1230
rect 560 -1150 600 -1140
rect 560 -1230 565 -1150
rect 595 -1230 600 -1150
rect 560 -1240 600 -1230
rect 880 -1150 920 -1140
rect 880 -1230 885 -1150
rect 915 -1230 920 -1150
rect 880 -1280 920 -1230
rect 1200 -1150 1240 -1140
rect 1200 -1230 1205 -1150
rect 1235 -1230 1240 -1150
rect 1200 -1240 1240 -1230
rect 1520 -1150 1560 -1140
rect 1520 -1230 1525 -1150
rect 1555 -1230 1560 -1150
rect 1520 -1280 1560 -1230
rect 1840 -1150 1880 -1140
rect 1840 -1230 1845 -1150
rect 1875 -1230 1880 -1150
rect 1840 -1240 1880 -1230
rect 2160 -1150 2200 -1140
rect 2160 -1230 2165 -1150
rect 2195 -1230 2200 -1150
rect 2160 -1280 2200 -1230
rect 2480 -1150 2520 -1140
rect 2480 -1230 2485 -1150
rect 2515 -1230 2520 -1150
rect 2480 -1240 2520 -1230
rect 2800 -1150 2840 -1140
rect 2800 -1230 2805 -1150
rect 2835 -1230 2840 -1150
rect 2800 -1280 2840 -1230
rect 3120 -1150 3160 -1140
rect 3120 -1230 3125 -1150
rect 3155 -1230 3160 -1150
rect 3120 -1240 3160 -1230
rect 3440 -1150 3480 -1140
rect 3440 -1230 3445 -1150
rect 3475 -1230 3480 -1150
rect 3440 -1280 3480 -1230
rect 3760 -1150 3800 -1140
rect 3760 -1230 3765 -1150
rect 3795 -1230 3800 -1150
rect 3760 -1240 3800 -1230
rect 4080 -1150 4120 -1140
rect 4080 -1230 4085 -1150
rect 4115 -1230 4120 -1150
rect 4080 -1280 4120 -1230
rect 4400 -1150 4440 -1140
rect 4400 -1230 4405 -1150
rect 4435 -1230 4440 -1150
rect 4400 -1240 4440 -1230
rect 4720 -1150 4760 -1140
rect 4720 -1230 4725 -1150
rect 4755 -1230 4760 -1150
rect 4720 -1280 4760 -1230
rect 5040 -1150 5080 -1140
rect 5040 -1230 5045 -1150
rect 5075 -1230 5080 -1150
rect 5040 -1240 5080 -1230
rect -80 -1320 5080 -1280
rect -240 -1480 -200 -1460
rect -80 -1350 -40 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 -40 -1350
rect -80 -1480 -40 -1430
rect 240 -1350 280 -1340
rect 240 -1430 245 -1350
rect 275 -1430 280 -1350
rect 240 -1440 280 -1430
rect 560 -1350 600 -1320
rect 560 -1430 565 -1350
rect 595 -1430 600 -1350
rect 560 -1440 600 -1430
rect 880 -1350 920 -1340
rect 880 -1430 885 -1350
rect 915 -1430 920 -1350
rect 880 -1440 920 -1430
rect 1200 -1350 1240 -1340
rect 1200 -1430 1205 -1350
rect 1235 -1430 1240 -1350
rect 1200 -1480 1240 -1430
rect 1520 -1350 1560 -1340
rect 1520 -1430 1525 -1350
rect 1555 -1430 1560 -1350
rect 1520 -1440 1560 -1430
rect 1840 -1350 1880 -1320
rect 1840 -1430 1845 -1350
rect 1875 -1430 1880 -1350
rect 1840 -1440 1880 -1430
rect 2160 -1350 2200 -1340
rect 2160 -1430 2165 -1350
rect 2195 -1430 2200 -1350
rect 2160 -1440 2200 -1430
rect 2480 -1350 2520 -1340
rect 2480 -1430 2485 -1350
rect 2515 -1430 2520 -1350
rect 2480 -1480 2520 -1430
rect 2800 -1350 2840 -1340
rect 2800 -1430 2805 -1350
rect 2835 -1430 2840 -1350
rect 2800 -1440 2840 -1430
rect 3120 -1350 3160 -1320
rect 3120 -1430 3125 -1350
rect 3155 -1430 3160 -1350
rect 3120 -1440 3160 -1430
rect 3440 -1350 3480 -1340
rect 3440 -1430 3445 -1350
rect 3475 -1430 3480 -1350
rect 3440 -1440 3480 -1430
rect 3760 -1350 3800 -1340
rect 3760 -1430 3765 -1350
rect 3795 -1430 3800 -1350
rect 3760 -1480 3800 -1430
rect 4080 -1350 4120 -1340
rect 4080 -1430 4085 -1350
rect 4115 -1430 4120 -1350
rect 4080 -1440 4120 -1430
rect 4400 -1350 4440 -1320
rect 4400 -1430 4405 -1350
rect 4435 -1430 4440 -1350
rect 4400 -1440 4440 -1430
rect 4720 -1350 4760 -1340
rect 4720 -1430 4725 -1350
rect 4755 -1430 4760 -1350
rect 4720 -1440 4760 -1430
rect 5040 -1350 5080 -1340
rect 5040 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5040 -1480 5080 -1430
rect 5200 -1480 5240 -1460
rect -240 -1520 -180 -1480
rect 5180 -1520 5240 -1480
<< viali >>
rect -75 390 -45 670
rect 245 390 275 670
rect 565 390 595 670
rect 885 390 915 670
rect 1205 390 1235 670
rect 1525 390 1555 670
rect 1845 390 1875 670
rect 2165 390 2195 670
rect 2485 390 2515 670
rect 2805 390 2835 670
rect 3125 390 3155 670
rect 3445 390 3475 670
rect 3765 390 3795 670
rect 4085 390 4115 670
rect 4405 390 4435 670
rect 4725 390 4755 670
rect 5045 390 5075 670
rect -75 -10 -45 270
rect 245 -10 275 270
rect 565 -10 595 270
rect 885 -10 915 270
rect 1205 -10 1235 270
rect 1525 -10 1555 270
rect 1845 -10 1875 270
rect 2165 -10 2195 270
rect 2485 -10 2515 270
rect 2805 -10 2835 270
rect 3125 -10 3155 270
rect 3445 -10 3475 270
rect 3765 -10 3795 270
rect 4085 -10 4115 270
rect 4405 -10 4435 270
rect 4725 -10 4755 270
rect 5045 -10 5075 270
rect 10 -75 190 -45
rect 330 -75 510 -45
rect 650 -75 830 -45
rect 970 -75 1150 -45
rect 1290 -75 1470 -45
rect 1610 -75 1790 -45
rect 1930 -75 2110 -45
rect 2250 -75 2430 -45
rect 2570 -75 2750 -45
rect 2890 -75 3070 -45
rect 3210 -75 3390 -45
rect 3530 -75 3710 -45
rect 3850 -75 4030 -45
rect 4170 -75 4350 -45
rect 4490 -75 4670 -45
rect 4810 -75 4990 -45
rect -75 -730 -45 -450
rect 245 -730 275 -450
rect 565 -730 595 -450
rect 885 -730 915 -450
rect 1205 -730 1235 -450
rect 1525 -730 1555 -450
rect 1845 -730 1875 -450
rect 2165 -730 2195 -450
rect 2485 -730 2515 -450
rect 2805 -730 2835 -450
rect 3125 -730 3155 -450
rect 3445 -730 3475 -450
rect 3765 -730 3795 -450
rect 4085 -730 4115 -450
rect 4405 -730 4435 -450
rect 4725 -730 4755 -450
rect 5045 -730 5075 -450
rect 10 -795 190 -765
rect 330 -795 510 -765
rect 650 -795 830 -765
rect 970 -795 1150 -765
rect 1290 -795 1470 -765
rect 1610 -795 1790 -765
rect 1930 -795 2110 -765
rect 2250 -795 2430 -765
rect 2570 -795 2750 -765
rect 2890 -795 3070 -765
rect 3210 -795 3390 -765
rect 3530 -795 3710 -765
rect 3850 -795 4030 -765
rect 4170 -795 4350 -765
rect 4490 -795 4670 -765
rect 4810 -795 4990 -765
rect 10 -1115 190 -1085
rect 330 -1115 510 -1085
rect 650 -1115 830 -1085
rect 970 -1115 1150 -1085
rect 1290 -1115 1470 -1085
rect 1610 -1115 1790 -1085
rect 1930 -1115 2110 -1085
rect 2250 -1115 2430 -1085
rect 2570 -1115 2750 -1085
rect 2890 -1115 3070 -1085
rect 3210 -1115 3390 -1085
rect 3530 -1115 3710 -1085
rect 3850 -1115 4030 -1085
rect 4170 -1115 4350 -1085
rect 4490 -1115 4670 -1085
rect 4810 -1115 4990 -1085
rect -75 -1230 -45 -1150
rect 245 -1230 275 -1150
rect 565 -1230 595 -1150
rect 885 -1230 915 -1150
rect 1205 -1230 1235 -1150
rect 1525 -1230 1555 -1150
rect 1845 -1230 1875 -1150
rect 2165 -1230 2195 -1150
rect 2485 -1230 2515 -1150
rect 2805 -1230 2835 -1150
rect 3125 -1230 3155 -1150
rect 3445 -1230 3475 -1150
rect 3765 -1230 3795 -1150
rect 4085 -1230 4115 -1150
rect 4405 -1230 4435 -1150
rect 4725 -1230 4755 -1150
rect 5045 -1230 5075 -1150
rect -75 -1430 -45 -1350
rect 245 -1430 275 -1350
rect 565 -1430 595 -1350
rect 885 -1430 915 -1350
rect 1205 -1430 1235 -1350
rect 1525 -1430 1555 -1350
rect 1845 -1430 1875 -1350
rect 2165 -1430 2195 -1350
rect 2485 -1430 2515 -1350
rect 2805 -1430 2835 -1350
rect 3125 -1430 3155 -1350
rect 3445 -1430 3475 -1350
rect 3765 -1430 3795 -1350
rect 4085 -1430 4115 -1350
rect 4405 -1430 4435 -1350
rect 4725 -1430 4755 -1350
rect 5045 -1430 5075 -1350
<< metal1 >>
rect -80 670 -40 680
rect -80 390 -75 670
rect -45 390 -40 670
rect -80 380 -40 390
rect 240 670 280 680
rect 240 390 245 670
rect 275 390 280 670
rect 240 380 280 390
rect 560 670 600 680
rect 560 390 565 670
rect 595 390 600 670
rect 560 380 600 390
rect 880 670 920 680
rect 880 390 885 670
rect 915 390 920 670
rect 880 380 920 390
rect 1200 670 1240 680
rect 1200 390 1205 670
rect 1235 390 1240 670
rect 1200 380 1240 390
rect 1520 670 1560 680
rect 1520 390 1525 670
rect 1555 390 1560 670
rect 1520 380 1560 390
rect 1840 670 1880 680
rect 1840 390 1845 670
rect 1875 390 1880 670
rect 1840 380 1880 390
rect 2160 670 2200 680
rect 2160 390 2165 670
rect 2195 390 2200 670
rect 2160 380 2200 390
rect 2480 670 2520 680
rect 2480 390 2485 670
rect 2515 390 2520 670
rect 2480 380 2520 390
rect 2800 670 2840 680
rect 2800 390 2805 670
rect 2835 390 2840 670
rect 2800 380 2840 390
rect 3120 670 3160 680
rect 3120 390 3125 670
rect 3155 390 3160 670
rect 3120 380 3160 390
rect 3440 670 3480 680
rect 3440 390 3445 670
rect 3475 390 3480 670
rect 3440 380 3480 390
rect 3760 670 3800 680
rect 3760 390 3765 670
rect 3795 390 3800 670
rect 3760 380 3800 390
rect 4080 670 4120 680
rect 4080 390 4085 670
rect 4115 390 4120 670
rect 4080 380 4120 390
rect 4400 670 4440 680
rect 4400 390 4405 670
rect 4435 390 4440 670
rect 4400 380 4440 390
rect 4720 670 4760 680
rect 4720 390 4725 670
rect 4755 390 4760 670
rect 4720 380 4760 390
rect 5040 670 5080 680
rect 5040 390 5045 670
rect 5075 390 5080 670
rect 5040 380 5080 390
rect -80 270 -40 280
rect -80 -10 -75 270
rect -45 -10 -40 270
rect -80 -20 -40 -10
rect 240 270 280 280
rect 240 -10 245 270
rect 275 -10 280 270
rect 0 -45 200 -40
rect 0 -75 10 -45
rect 190 -75 200 -45
rect 0 -80 200 -75
rect 240 -45 280 -10
rect 560 270 600 280
rect 560 -10 565 270
rect 595 -10 600 270
rect 560 -20 600 -10
rect 880 270 920 280
rect 880 -10 885 270
rect 915 -10 920 270
rect 240 -75 245 -45
rect 275 -75 280 -45
rect -80 -450 -40 -440
rect -80 -730 -75 -450
rect -45 -730 -40 -450
rect -80 -765 -40 -730
rect 240 -450 280 -75
rect 320 -45 520 -40
rect 320 -75 330 -45
rect 510 -75 520 -45
rect 320 -80 520 -75
rect 640 -45 840 -40
rect 640 -75 650 -45
rect 830 -75 840 -45
rect 640 -80 840 -75
rect 880 -45 920 -10
rect 1200 270 1240 280
rect 1200 -10 1205 270
rect 1235 -10 1240 270
rect 1200 -20 1240 -10
rect 1520 270 1560 280
rect 1520 -10 1525 270
rect 1555 -10 1560 270
rect 880 -75 885 -45
rect 915 -75 920 -45
rect 240 -730 245 -450
rect 275 -730 280 -450
rect 240 -740 280 -730
rect 560 -450 600 -440
rect 560 -730 565 -450
rect 595 -730 600 -450
rect -80 -795 -75 -765
rect -45 -795 -40 -765
rect -80 -1150 -40 -795
rect 0 -765 200 -760
rect 0 -795 10 -765
rect 190 -795 200 -765
rect 0 -800 200 -795
rect 320 -765 520 -760
rect 320 -795 330 -765
rect 510 -795 520 -765
rect 320 -800 520 -795
rect 560 -765 600 -730
rect 880 -450 920 -75
rect 960 -45 1160 -40
rect 960 -75 970 -45
rect 1150 -75 1160 -45
rect 960 -80 1160 -75
rect 1280 -45 1480 -40
rect 1280 -75 1290 -45
rect 1470 -75 1480 -45
rect 1280 -80 1480 -75
rect 1520 -45 1560 -10
rect 1840 270 1880 280
rect 1840 -10 1845 270
rect 1875 -10 1880 270
rect 1840 -20 1880 -10
rect 2160 270 2200 280
rect 2160 -10 2165 270
rect 2195 -10 2200 270
rect 1520 -75 1525 -45
rect 1555 -75 1560 -45
rect 880 -730 885 -450
rect 915 -730 920 -450
rect 880 -740 920 -730
rect 1200 -450 1240 -440
rect 1200 -730 1205 -450
rect 1235 -730 1240 -450
rect 560 -795 565 -765
rect 595 -795 600 -765
rect 0 -1085 200 -1080
rect 0 -1115 10 -1085
rect 190 -1115 200 -1085
rect 0 -1120 200 -1115
rect 320 -1085 520 -1080
rect 320 -1115 330 -1085
rect 510 -1115 520 -1085
rect 320 -1120 520 -1115
rect -80 -1230 -75 -1150
rect -45 -1230 -40 -1150
rect -80 -1240 -40 -1230
rect 240 -1150 280 -1140
rect 240 -1230 245 -1150
rect 275 -1230 280 -1150
rect 240 -1240 280 -1230
rect 560 -1150 600 -795
rect 640 -765 840 -760
rect 640 -795 650 -765
rect 830 -795 840 -765
rect 640 -800 840 -795
rect 880 -800 920 -760
rect 960 -765 1160 -760
rect 960 -795 970 -765
rect 1150 -795 1160 -765
rect 960 -800 1160 -795
rect 1200 -765 1240 -730
rect 1520 -450 1560 -75
rect 1600 -45 1800 -40
rect 1600 -75 1610 -45
rect 1790 -75 1800 -45
rect 1600 -80 1800 -75
rect 1920 -45 2120 -40
rect 1920 -75 1930 -45
rect 2110 -75 2120 -45
rect 1920 -80 2120 -75
rect 2160 -45 2200 -10
rect 2480 270 2520 280
rect 2480 -10 2485 270
rect 2515 -10 2520 270
rect 2480 -20 2520 -10
rect 2800 270 2840 280
rect 2800 -10 2805 270
rect 2835 -10 2840 270
rect 2160 -75 2165 -45
rect 2195 -75 2200 -45
rect 1520 -730 1525 -450
rect 1555 -730 1560 -450
rect 1520 -740 1560 -730
rect 1840 -450 1880 -440
rect 1840 -730 1845 -450
rect 1875 -730 1880 -450
rect 1200 -795 1205 -765
rect 1235 -795 1240 -765
rect 640 -1085 840 -1080
rect 640 -1115 650 -1085
rect 830 -1115 840 -1085
rect 640 -1120 840 -1115
rect 960 -1085 1160 -1080
rect 960 -1115 970 -1085
rect 1150 -1115 1160 -1085
rect 960 -1120 1160 -1115
rect 560 -1230 565 -1150
rect 595 -1230 600 -1150
rect 560 -1240 600 -1230
rect 880 -1150 920 -1140
rect 880 -1230 885 -1150
rect 915 -1230 920 -1150
rect 880 -1240 920 -1230
rect 1200 -1150 1240 -795
rect 1280 -765 1480 -760
rect 1280 -795 1290 -765
rect 1470 -795 1480 -765
rect 1280 -800 1480 -795
rect 1520 -800 1560 -760
rect 1600 -765 1800 -760
rect 1600 -795 1610 -765
rect 1790 -795 1800 -765
rect 1600 -800 1800 -795
rect 1840 -765 1880 -730
rect 2160 -450 2200 -75
rect 2240 -45 2440 -40
rect 2240 -75 2250 -45
rect 2430 -75 2440 -45
rect 2240 -80 2440 -75
rect 2560 -45 2760 -40
rect 2560 -75 2570 -45
rect 2750 -75 2760 -45
rect 2560 -80 2760 -75
rect 2800 -45 2840 -10
rect 3120 270 3160 280
rect 3120 -10 3125 270
rect 3155 -10 3160 270
rect 3120 -20 3160 -10
rect 3440 270 3480 280
rect 3440 -10 3445 270
rect 3475 -10 3480 270
rect 2800 -75 2805 -45
rect 2835 -75 2840 -45
rect 2160 -730 2165 -450
rect 2195 -730 2200 -450
rect 2160 -740 2200 -730
rect 2480 -450 2520 -440
rect 2480 -730 2485 -450
rect 2515 -730 2520 -450
rect 1840 -795 1845 -765
rect 1875 -795 1880 -765
rect 1280 -1085 1480 -1080
rect 1280 -1115 1290 -1085
rect 1470 -1115 1480 -1085
rect 1280 -1120 1480 -1115
rect 1600 -1085 1800 -1080
rect 1600 -1115 1610 -1085
rect 1790 -1115 1800 -1085
rect 1600 -1120 1800 -1115
rect 1200 -1230 1205 -1150
rect 1235 -1230 1240 -1150
rect 1200 -1240 1240 -1230
rect 1520 -1150 1560 -1140
rect 1520 -1230 1525 -1150
rect 1555 -1230 1560 -1150
rect 1520 -1240 1560 -1230
rect 1840 -1150 1880 -795
rect 1920 -765 2120 -760
rect 1920 -795 1930 -765
rect 2110 -795 2120 -765
rect 1920 -800 2120 -795
rect 2160 -800 2200 -760
rect 2240 -765 2440 -760
rect 2240 -795 2250 -765
rect 2430 -795 2440 -765
rect 2240 -800 2440 -795
rect 2480 -765 2520 -730
rect 2800 -450 2840 -75
rect 2880 -45 3080 -40
rect 2880 -75 2890 -45
rect 3070 -75 3080 -45
rect 2880 -80 3080 -75
rect 3200 -45 3400 -40
rect 3200 -75 3210 -45
rect 3390 -75 3400 -45
rect 3200 -80 3400 -75
rect 3440 -45 3480 -10
rect 3760 270 3800 280
rect 3760 -10 3765 270
rect 3795 -10 3800 270
rect 3760 -20 3800 -10
rect 4080 270 4120 280
rect 4080 -10 4085 270
rect 4115 -10 4120 270
rect 3440 -75 3445 -45
rect 3475 -75 3480 -45
rect 2800 -730 2805 -450
rect 2835 -730 2840 -450
rect 2800 -740 2840 -730
rect 3120 -450 3160 -440
rect 3120 -730 3125 -450
rect 3155 -730 3160 -450
rect 2480 -795 2485 -765
rect 2515 -795 2520 -765
rect 1920 -1085 2120 -1080
rect 1920 -1115 1930 -1085
rect 2110 -1115 2120 -1085
rect 1920 -1120 2120 -1115
rect 2240 -1085 2440 -1080
rect 2240 -1115 2250 -1085
rect 2430 -1115 2440 -1085
rect 2240 -1120 2440 -1115
rect 1840 -1230 1845 -1150
rect 1875 -1230 1880 -1150
rect 1840 -1240 1880 -1230
rect 2160 -1150 2200 -1140
rect 2160 -1230 2165 -1150
rect 2195 -1230 2200 -1150
rect 2160 -1240 2200 -1230
rect 2480 -1150 2520 -795
rect 2560 -765 2760 -760
rect 2560 -795 2570 -765
rect 2750 -795 2760 -765
rect 2560 -800 2760 -795
rect 2800 -800 2840 -760
rect 2880 -765 3080 -760
rect 2880 -795 2890 -765
rect 3070 -795 3080 -765
rect 2880 -800 3080 -795
rect 3120 -765 3160 -730
rect 3440 -450 3480 -75
rect 3520 -45 3720 -40
rect 3520 -75 3530 -45
rect 3710 -75 3720 -45
rect 3520 -80 3720 -75
rect 3840 -45 4040 -40
rect 3840 -75 3850 -45
rect 4030 -75 4040 -45
rect 3840 -80 4040 -75
rect 4080 -45 4120 -10
rect 4400 270 4440 280
rect 4400 -10 4405 270
rect 4435 -10 4440 270
rect 4400 -20 4440 -10
rect 4720 270 4760 280
rect 4720 -10 4725 270
rect 4755 -10 4760 270
rect 4080 -75 4085 -45
rect 4115 -75 4120 -45
rect 3440 -730 3445 -450
rect 3475 -730 3480 -450
rect 3440 -740 3480 -730
rect 3760 -450 3800 -440
rect 3760 -730 3765 -450
rect 3795 -730 3800 -450
rect 3120 -795 3125 -765
rect 3155 -795 3160 -765
rect 2560 -1085 2760 -1080
rect 2560 -1115 2570 -1085
rect 2750 -1115 2760 -1085
rect 2560 -1120 2760 -1115
rect 2880 -1085 3080 -1080
rect 2880 -1115 2890 -1085
rect 3070 -1115 3080 -1085
rect 2880 -1120 3080 -1115
rect 2480 -1230 2485 -1150
rect 2515 -1230 2520 -1150
rect 2480 -1240 2520 -1230
rect 2800 -1150 2840 -1140
rect 2800 -1230 2805 -1150
rect 2835 -1230 2840 -1150
rect 2800 -1240 2840 -1230
rect 3120 -1150 3160 -795
rect 3200 -765 3400 -760
rect 3200 -795 3210 -765
rect 3390 -795 3400 -765
rect 3200 -800 3400 -795
rect 3440 -800 3480 -760
rect 3520 -765 3720 -760
rect 3520 -795 3530 -765
rect 3710 -795 3720 -765
rect 3520 -800 3720 -795
rect 3760 -765 3800 -730
rect 4080 -450 4120 -75
rect 4160 -45 4360 -40
rect 4160 -75 4170 -45
rect 4350 -75 4360 -45
rect 4160 -80 4360 -75
rect 4480 -45 4680 -40
rect 4480 -75 4490 -45
rect 4670 -75 4680 -45
rect 4480 -80 4680 -75
rect 4720 -45 4760 -10
rect 5040 270 5080 280
rect 5040 -10 5045 270
rect 5075 -10 5080 270
rect 5040 -20 5080 -10
rect 4720 -75 4725 -45
rect 4755 -75 4760 -45
rect 4080 -730 4085 -450
rect 4115 -730 4120 -450
rect 4080 -740 4120 -730
rect 4400 -450 4440 -440
rect 4400 -730 4405 -450
rect 4435 -730 4440 -450
rect 3760 -795 3765 -765
rect 3795 -795 3800 -765
rect 3200 -1085 3400 -1080
rect 3200 -1115 3210 -1085
rect 3390 -1115 3400 -1085
rect 3200 -1120 3400 -1115
rect 3520 -1085 3720 -1080
rect 3520 -1115 3530 -1085
rect 3710 -1115 3720 -1085
rect 3520 -1120 3720 -1115
rect 3120 -1230 3125 -1150
rect 3155 -1230 3160 -1150
rect 3120 -1240 3160 -1230
rect 3440 -1150 3480 -1140
rect 3440 -1230 3445 -1150
rect 3475 -1230 3480 -1150
rect 3440 -1240 3480 -1230
rect 3760 -1150 3800 -795
rect 3840 -765 4040 -760
rect 3840 -795 3850 -765
rect 4030 -795 4040 -765
rect 3840 -800 4040 -795
rect 4080 -800 4120 -760
rect 4160 -765 4360 -760
rect 4160 -795 4170 -765
rect 4350 -795 4360 -765
rect 4160 -800 4360 -795
rect 4400 -765 4440 -730
rect 4720 -450 4760 -75
rect 4800 -45 5000 -40
rect 4800 -75 4810 -45
rect 4990 -75 5000 -45
rect 4800 -80 5000 -75
rect 4720 -730 4725 -450
rect 4755 -730 4760 -450
rect 4720 -740 4760 -730
rect 5040 -450 5080 -440
rect 5040 -730 5045 -450
rect 5075 -730 5080 -450
rect 4400 -795 4405 -765
rect 4435 -795 4440 -765
rect 3840 -1085 4040 -1080
rect 3840 -1115 3850 -1085
rect 4030 -1115 4040 -1085
rect 3840 -1120 4040 -1115
rect 4160 -1085 4360 -1080
rect 4160 -1115 4170 -1085
rect 4350 -1115 4360 -1085
rect 4160 -1120 4360 -1115
rect 3760 -1230 3765 -1150
rect 3795 -1230 3800 -1150
rect 3760 -1240 3800 -1230
rect 4080 -1150 4120 -1140
rect 4080 -1230 4085 -1150
rect 4115 -1230 4120 -1150
rect 4080 -1240 4120 -1230
rect 4400 -1150 4440 -795
rect 4480 -765 4680 -760
rect 4480 -795 4490 -765
rect 4670 -795 4680 -765
rect 4480 -800 4680 -795
rect 4720 -800 4760 -760
rect 4800 -765 5000 -760
rect 4800 -795 4810 -765
rect 4990 -795 5000 -765
rect 4800 -800 5000 -795
rect 5040 -765 5080 -730
rect 5040 -795 5045 -765
rect 5075 -795 5080 -765
rect 4480 -1085 4680 -1080
rect 4480 -1115 4490 -1085
rect 4670 -1115 4680 -1085
rect 4480 -1120 4680 -1115
rect 4800 -1085 5000 -1080
rect 4800 -1115 4810 -1085
rect 4990 -1115 5000 -1085
rect 4800 -1120 5000 -1115
rect 4400 -1230 4405 -1150
rect 4435 -1230 4440 -1150
rect 4400 -1240 4440 -1230
rect 4720 -1150 4760 -1140
rect 4720 -1230 4725 -1150
rect 4755 -1230 4760 -1150
rect 4720 -1240 4760 -1230
rect 5040 -1150 5080 -795
rect 5040 -1230 5045 -1150
rect 5075 -1230 5080 -1150
rect 5040 -1240 5080 -1230
rect -80 -1350 -40 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 -40 -1350
rect -80 -1440 -40 -1430
rect 240 -1350 280 -1340
rect 240 -1430 245 -1350
rect 275 -1430 280 -1350
rect 240 -1440 280 -1430
rect 560 -1350 600 -1340
rect 560 -1430 565 -1350
rect 595 -1430 600 -1350
rect 560 -1440 600 -1430
rect 880 -1350 920 -1340
rect 880 -1430 885 -1350
rect 915 -1430 920 -1350
rect 880 -1440 920 -1430
rect 1200 -1350 1240 -1340
rect 1200 -1430 1205 -1350
rect 1235 -1430 1240 -1350
rect 1200 -1440 1240 -1430
rect 1520 -1350 1560 -1340
rect 1520 -1430 1525 -1350
rect 1555 -1430 1560 -1350
rect 1520 -1440 1560 -1430
rect 1840 -1350 1880 -1340
rect 1840 -1430 1845 -1350
rect 1875 -1430 1880 -1350
rect 1840 -1440 1880 -1430
rect 2160 -1350 2200 -1340
rect 2160 -1430 2165 -1350
rect 2195 -1430 2200 -1350
rect 2160 -1440 2200 -1430
rect 2480 -1350 2520 -1340
rect 2480 -1430 2485 -1350
rect 2515 -1430 2520 -1350
rect 2480 -1440 2520 -1430
rect 2800 -1350 2840 -1340
rect 2800 -1430 2805 -1350
rect 2835 -1430 2840 -1350
rect 2800 -1440 2840 -1430
rect 3120 -1350 3160 -1340
rect 3120 -1430 3125 -1350
rect 3155 -1430 3160 -1350
rect 3120 -1440 3160 -1430
rect 3440 -1350 3480 -1340
rect 3440 -1430 3445 -1350
rect 3475 -1430 3480 -1350
rect 3440 -1440 3480 -1430
rect 3760 -1350 3800 -1340
rect 3760 -1430 3765 -1350
rect 3795 -1430 3800 -1350
rect 3760 -1440 3800 -1430
rect 4080 -1350 4120 -1340
rect 4080 -1430 4085 -1350
rect 4115 -1430 4120 -1350
rect 4080 -1440 4120 -1430
rect 4400 -1350 4440 -1340
rect 4400 -1430 4405 -1350
rect 4435 -1430 4440 -1350
rect 4400 -1440 4440 -1430
rect 4720 -1350 4760 -1340
rect 4720 -1430 4725 -1350
rect 4755 -1430 4760 -1350
rect 4720 -1440 4760 -1430
rect 5040 -1350 5080 -1340
rect 5040 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5040 -1440 5080 -1430
<< via1 >>
rect -75 450 -45 630
rect 1205 450 1235 630
rect 2485 450 2515 630
rect 3765 450 3795 630
rect 5045 450 5075 630
rect 10 -75 190 -45
rect 245 -75 275 -45
rect 330 -75 510 -45
rect 650 -75 830 -45
rect 885 -75 915 -45
rect -75 -795 -45 -765
rect 10 -795 190 -765
rect 330 -795 510 -765
rect 970 -75 1150 -45
rect 1290 -75 1470 -45
rect 1525 -75 1555 -45
rect 565 -795 595 -765
rect 10 -1115 190 -1085
rect 330 -1115 510 -1085
rect 650 -795 830 -765
rect 970 -795 1150 -765
rect 1610 -75 1790 -45
rect 1930 -75 2110 -45
rect 2165 -75 2195 -45
rect 1205 -795 1235 -765
rect 650 -1115 830 -1085
rect 970 -1115 1150 -1085
rect 1290 -795 1470 -765
rect 1610 -795 1790 -765
rect 2250 -75 2430 -45
rect 2570 -75 2750 -45
rect 2805 -75 2835 -45
rect 1845 -795 1875 -765
rect 1290 -1115 1470 -1085
rect 1610 -1115 1790 -1085
rect 1930 -795 2110 -765
rect 2250 -795 2430 -765
rect 2890 -75 3070 -45
rect 3210 -75 3390 -45
rect 3445 -75 3475 -45
rect 2485 -795 2515 -765
rect 1930 -1115 2110 -1085
rect 2250 -1115 2430 -1085
rect 2570 -795 2750 -765
rect 2890 -795 3070 -765
rect 3530 -75 3710 -45
rect 3850 -75 4030 -45
rect 4085 -75 4115 -45
rect 3125 -795 3155 -765
rect 2570 -1115 2750 -1085
rect 2890 -1115 3070 -1085
rect 3210 -795 3390 -765
rect 3530 -795 3710 -765
rect 4170 -75 4350 -45
rect 4490 -75 4670 -45
rect 4725 -75 4755 -45
rect 3765 -795 3795 -765
rect 3210 -1115 3390 -1085
rect 3530 -1115 3710 -1085
rect 3850 -795 4030 -765
rect 4170 -795 4350 -765
rect 4810 -75 4990 -45
rect 4405 -795 4435 -765
rect 3850 -1115 4030 -1085
rect 4170 -1115 4350 -1085
rect 4490 -795 4670 -765
rect 4810 -795 4990 -765
rect 5045 -795 5075 -765
rect 4490 -1115 4670 -1085
rect 4810 -1115 4990 -1085
rect -75 -1430 -45 -1360
rect 1205 -1430 1235 -1360
rect 2485 -1430 2515 -1360
rect 3765 -1430 3795 -1360
rect 5045 -1430 5075 -1360
<< metal2 >>
rect -80 630 -40 640
rect -80 450 -75 630
rect -45 450 -40 630
rect -80 440 -40 450
rect 1200 630 1240 640
rect 1200 450 1205 630
rect 1235 450 1240 630
rect 1200 440 1240 450
rect 2480 630 2520 640
rect 2480 450 2485 630
rect 2515 450 2520 630
rect 2480 440 2520 450
rect 3760 630 3800 640
rect 3760 450 3765 630
rect 3795 450 3800 630
rect 3760 440 3800 450
rect 5040 630 5080 640
rect 5040 450 5045 630
rect 5075 450 5080 630
rect 5040 440 5080 450
rect -240 35 5240 40
rect -240 5 -235 35
rect -205 5 -155 35
rect -125 5 -75 35
rect -45 5 5 35
rect 35 5 85 35
rect 115 5 165 35
rect 195 5 325 35
rect 355 5 405 35
rect 435 5 485 35
rect 515 5 565 35
rect 595 5 645 35
rect 675 5 725 35
rect 755 5 805 35
rect 835 5 965 35
rect 995 5 1045 35
rect 1075 5 1125 35
rect 1155 5 1205 35
rect 1235 5 1285 35
rect 1315 5 1365 35
rect 1395 5 1445 35
rect 1475 5 1605 35
rect 1635 5 1685 35
rect 1715 5 1765 35
rect 1795 5 1845 35
rect 1875 5 1925 35
rect 1955 5 2005 35
rect 2035 5 2085 35
rect 2115 5 2245 35
rect 2275 5 2325 35
rect 2355 5 2405 35
rect 2435 5 2485 35
rect 2515 5 2565 35
rect 2595 5 2645 35
rect 2675 5 2725 35
rect 2755 5 2885 35
rect 2915 5 2965 35
rect 2995 5 3045 35
rect 3075 5 3125 35
rect 3155 5 3205 35
rect 3235 5 3285 35
rect 3315 5 3365 35
rect 3395 5 3525 35
rect 3555 5 3605 35
rect 3635 5 3685 35
rect 3715 5 3765 35
rect 3795 5 3845 35
rect 3875 5 3925 35
rect 3955 5 4005 35
rect 4035 5 4165 35
rect 4195 5 4245 35
rect 4275 5 4325 35
rect 4355 5 4405 35
rect 4435 5 4485 35
rect 4515 5 4565 35
rect 4595 5 4645 35
rect 4675 5 4805 35
rect 4835 5 4885 35
rect 4915 5 4965 35
rect 4995 5 5045 35
rect 5075 5 5125 35
rect 5155 5 5205 35
rect 5235 5 5240 35
rect -240 0 5240 5
rect -240 -45 5240 -40
rect -240 -75 10 -45
rect 190 -75 245 -45
rect 275 -75 330 -45
rect 510 -75 650 -45
rect 830 -75 885 -45
rect 915 -75 970 -45
rect 1150 -75 1290 -45
rect 1470 -75 1525 -45
rect 1555 -75 1610 -45
rect 1790 -75 1930 -45
rect 2110 -75 2165 -45
rect 2195 -75 2250 -45
rect 2430 -75 2570 -45
rect 2750 -75 2805 -45
rect 2835 -75 2890 -45
rect 3070 -75 3210 -45
rect 3390 -75 3445 -45
rect 3475 -75 3530 -45
rect 3710 -75 3850 -45
rect 4030 -75 4085 -45
rect 4115 -75 4170 -45
rect 4350 -75 4490 -45
rect 4670 -75 4725 -45
rect 4755 -75 4810 -45
rect 4990 -75 5240 -45
rect -240 -80 5240 -75
rect -240 -125 5240 -120
rect -240 -155 -235 -125
rect -205 -155 -155 -125
rect -125 -155 -75 -125
rect -45 -155 5 -125
rect 35 -155 85 -125
rect 115 -155 165 -125
rect 195 -155 325 -125
rect 355 -155 405 -125
rect 435 -155 485 -125
rect 515 -155 565 -125
rect 595 -155 645 -125
rect 675 -155 725 -125
rect 755 -155 805 -125
rect 835 -155 965 -125
rect 995 -155 1045 -125
rect 1075 -155 1125 -125
rect 1155 -155 1205 -125
rect 1235 -155 1285 -125
rect 1315 -155 1365 -125
rect 1395 -155 1445 -125
rect 1475 -155 1605 -125
rect 1635 -155 1685 -125
rect 1715 -155 1765 -125
rect 1795 -155 1845 -125
rect 1875 -155 1925 -125
rect 1955 -155 2005 -125
rect 2035 -155 2085 -125
rect 2115 -155 2245 -125
rect 2275 -155 2325 -125
rect 2355 -155 2405 -125
rect 2435 -155 2485 -125
rect 2515 -155 2565 -125
rect 2595 -155 2645 -125
rect 2675 -155 2725 -125
rect 2755 -155 2885 -125
rect 2915 -155 2965 -125
rect 2995 -155 3045 -125
rect 3075 -155 3125 -125
rect 3155 -155 3205 -125
rect 3235 -155 3285 -125
rect 3315 -155 3365 -125
rect 3395 -155 3525 -125
rect 3555 -155 3605 -125
rect 3635 -155 3685 -125
rect 3715 -155 3765 -125
rect 3795 -155 3845 -125
rect 3875 -155 3925 -125
rect 3955 -155 4005 -125
rect 4035 -155 4165 -125
rect 4195 -155 4245 -125
rect 4275 -155 4325 -125
rect 4355 -155 4405 -125
rect 4435 -155 4485 -125
rect 4515 -155 4565 -125
rect 4595 -155 4645 -125
rect 4675 -155 4805 -125
rect 4835 -155 4885 -125
rect 4915 -155 4965 -125
rect 4995 -155 5045 -125
rect 5075 -155 5125 -125
rect 5155 -155 5205 -125
rect 5235 -155 5240 -125
rect -240 -160 5240 -155
rect -240 -685 5240 -680
rect -240 -715 -235 -685
rect -205 -715 -155 -685
rect -125 -715 -75 -685
rect -45 -715 5 -685
rect 35 -715 85 -685
rect 115 -715 165 -685
rect 195 -715 245 -685
rect 275 -715 325 -685
rect 355 -715 405 -685
rect 435 -715 485 -685
rect 515 -715 565 -685
rect 595 -715 645 -685
rect 675 -715 725 -685
rect 755 -715 805 -685
rect 835 -715 885 -685
rect 915 -715 965 -685
rect 995 -715 1045 -685
rect 1075 -715 1125 -685
rect 1155 -715 1205 -685
rect 1235 -715 1285 -685
rect 1315 -715 1365 -685
rect 1395 -715 1445 -685
rect 1475 -715 1525 -685
rect 1555 -715 1605 -685
rect 1635 -715 1685 -685
rect 1715 -715 1765 -685
rect 1795 -715 1845 -685
rect 1875 -715 1925 -685
rect 1955 -715 2005 -685
rect 2035 -715 2085 -685
rect 2115 -715 2165 -685
rect 2195 -715 2245 -685
rect 2275 -715 2325 -685
rect 2355 -715 2405 -685
rect 2435 -715 2485 -685
rect 2515 -715 2565 -685
rect 2595 -715 2645 -685
rect 2675 -715 2725 -685
rect 2755 -715 2805 -685
rect 2835 -715 2885 -685
rect 2915 -715 2965 -685
rect 2995 -715 3045 -685
rect 3075 -715 3125 -685
rect 3155 -715 3205 -685
rect 3235 -715 3285 -685
rect 3315 -715 3365 -685
rect 3395 -715 3445 -685
rect 3475 -715 3525 -685
rect 3555 -715 3605 -685
rect 3635 -715 3685 -685
rect 3715 -715 3765 -685
rect 3795 -715 3845 -685
rect 3875 -715 3925 -685
rect 3955 -715 4005 -685
rect 4035 -715 4085 -685
rect 4115 -715 4165 -685
rect 4195 -715 4245 -685
rect 4275 -715 4325 -685
rect 4355 -715 4405 -685
rect 4435 -715 4485 -685
rect 4515 -715 4565 -685
rect 4595 -715 4645 -685
rect 4675 -715 4725 -685
rect 4755 -715 4805 -685
rect 4835 -715 4885 -685
rect 4915 -715 4965 -685
rect 4995 -715 5045 -685
rect 5075 -715 5125 -685
rect 5155 -715 5205 -685
rect 5235 -715 5240 -685
rect -240 -720 5240 -715
rect -240 -765 5240 -760
rect -240 -795 -75 -765
rect -45 -795 10 -765
rect 190 -795 330 -765
rect 510 -795 565 -765
rect 595 -795 650 -765
rect 830 -795 970 -765
rect 1150 -795 1205 -765
rect 1235 -795 1290 -765
rect 1470 -795 1610 -765
rect 1790 -795 1845 -765
rect 1875 -795 1930 -765
rect 2110 -795 2250 -765
rect 2430 -795 2485 -765
rect 2515 -795 2570 -765
rect 2750 -795 2890 -765
rect 3070 -795 3125 -765
rect 3155 -795 3210 -765
rect 3390 -795 3530 -765
rect 3710 -795 3765 -765
rect 3795 -795 3850 -765
rect 4030 -795 4170 -765
rect 4350 -795 4405 -765
rect 4435 -795 4490 -765
rect 4670 -795 4810 -765
rect 4990 -795 5045 -765
rect 5075 -795 5240 -765
rect -240 -800 5240 -795
rect -240 -845 5240 -840
rect -240 -875 -235 -845
rect -205 -875 -155 -845
rect -125 -875 -75 -845
rect -45 -875 5 -845
rect 35 -875 85 -845
rect 115 -875 165 -845
rect 195 -875 245 -845
rect 275 -875 325 -845
rect 355 -875 405 -845
rect 435 -875 485 -845
rect 515 -875 565 -845
rect 595 -875 645 -845
rect 675 -875 725 -845
rect 755 -875 805 -845
rect 835 -875 885 -845
rect 915 -875 965 -845
rect 995 -875 1045 -845
rect 1075 -875 1125 -845
rect 1155 -875 1205 -845
rect 1235 -875 1285 -845
rect 1315 -875 1365 -845
rect 1395 -875 1445 -845
rect 1475 -875 1525 -845
rect 1555 -875 1605 -845
rect 1635 -875 1685 -845
rect 1715 -875 1765 -845
rect 1795 -875 1845 -845
rect 1875 -875 1925 -845
rect 1955 -875 2005 -845
rect 2035 -875 2085 -845
rect 2115 -875 2165 -845
rect 2195 -875 2245 -845
rect 2275 -875 2325 -845
rect 2355 -875 2405 -845
rect 2435 -875 2485 -845
rect 2515 -875 2565 -845
rect 2595 -875 2645 -845
rect 2675 -875 2725 -845
rect 2755 -875 2805 -845
rect 2835 -875 2885 -845
rect 2915 -875 2965 -845
rect 2995 -875 3045 -845
rect 3075 -875 3125 -845
rect 3155 -875 3205 -845
rect 3235 -875 3285 -845
rect 3315 -875 3365 -845
rect 3395 -875 3445 -845
rect 3475 -875 3525 -845
rect 3555 -875 3605 -845
rect 3635 -875 3685 -845
rect 3715 -875 3765 -845
rect 3795 -875 3845 -845
rect 3875 -875 3925 -845
rect 3955 -875 4005 -845
rect 4035 -875 4085 -845
rect 4115 -875 4165 -845
rect 4195 -875 4245 -845
rect 4275 -875 4325 -845
rect 4355 -875 4405 -845
rect 4435 -875 4485 -845
rect 4515 -875 4565 -845
rect 4595 -875 4645 -845
rect 4675 -875 4725 -845
rect 4755 -875 4805 -845
rect 4835 -875 4885 -845
rect 4915 -875 4965 -845
rect 4995 -875 5045 -845
rect 5075 -875 5125 -845
rect 5155 -875 5205 -845
rect 5235 -875 5240 -845
rect -240 -880 5240 -875
rect -240 -1005 5240 -1000
rect -240 -1035 -235 -1005
rect -205 -1035 -155 -1005
rect -125 -1035 -75 -1005
rect -45 -1035 5 -1005
rect 35 -1035 85 -1005
rect 115 -1035 165 -1005
rect 195 -1035 245 -1005
rect 275 -1035 325 -1005
rect 355 -1035 405 -1005
rect 435 -1035 485 -1005
rect 515 -1035 565 -1005
rect 595 -1035 645 -1005
rect 675 -1035 725 -1005
rect 755 -1035 805 -1005
rect 835 -1035 885 -1005
rect 915 -1035 965 -1005
rect 995 -1035 1045 -1005
rect 1075 -1035 1125 -1005
rect 1155 -1035 1205 -1005
rect 1235 -1035 1285 -1005
rect 1315 -1035 1365 -1005
rect 1395 -1035 1445 -1005
rect 1475 -1035 1525 -1005
rect 1555 -1035 1605 -1005
rect 1635 -1035 1685 -1005
rect 1715 -1035 1765 -1005
rect 1795 -1035 1845 -1005
rect 1875 -1035 1925 -1005
rect 1955 -1035 2005 -1005
rect 2035 -1035 2085 -1005
rect 2115 -1035 2165 -1005
rect 2195 -1035 2245 -1005
rect 2275 -1035 2325 -1005
rect 2355 -1035 2405 -1005
rect 2435 -1035 2485 -1005
rect 2515 -1035 2565 -1005
rect 2595 -1035 2645 -1005
rect 2675 -1035 2725 -1005
rect 2755 -1035 2805 -1005
rect 2835 -1035 2885 -1005
rect 2915 -1035 2965 -1005
rect 2995 -1035 3045 -1005
rect 3075 -1035 3125 -1005
rect 3155 -1035 3205 -1005
rect 3235 -1035 3285 -1005
rect 3315 -1035 3365 -1005
rect 3395 -1035 3445 -1005
rect 3475 -1035 3525 -1005
rect 3555 -1035 3605 -1005
rect 3635 -1035 3685 -1005
rect 3715 -1035 3765 -1005
rect 3795 -1035 3845 -1005
rect 3875 -1035 3925 -1005
rect 3955 -1035 4005 -1005
rect 4035 -1035 4085 -1005
rect 4115 -1035 4165 -1005
rect 4195 -1035 4245 -1005
rect 4275 -1035 4325 -1005
rect 4355 -1035 4405 -1005
rect 4435 -1035 4485 -1005
rect 4515 -1035 4565 -1005
rect 4595 -1035 4645 -1005
rect 4675 -1035 4725 -1005
rect 4755 -1035 4805 -1005
rect 4835 -1035 4885 -1005
rect 4915 -1035 4965 -1005
rect 4995 -1035 5045 -1005
rect 5075 -1035 5125 -1005
rect 5155 -1035 5205 -1005
rect 5235 -1035 5240 -1005
rect -240 -1040 5240 -1035
rect -240 -1085 5240 -1080
rect -240 -1115 10 -1085
rect 190 -1115 330 -1085
rect 510 -1115 650 -1085
rect 830 -1115 970 -1085
rect 1150 -1115 1290 -1085
rect 1470 -1115 1610 -1085
rect 1790 -1115 1930 -1085
rect 2110 -1115 2250 -1085
rect 2430 -1115 2570 -1085
rect 2750 -1115 2890 -1085
rect 3070 -1115 3210 -1085
rect 3390 -1115 3530 -1085
rect 3710 -1115 3850 -1085
rect 4030 -1115 4170 -1085
rect 4350 -1115 4490 -1085
rect 4670 -1115 4810 -1085
rect 4990 -1115 5240 -1085
rect -240 -1120 5240 -1115
rect -240 -1165 5240 -1160
rect -240 -1195 -235 -1165
rect -205 -1195 -155 -1165
rect -125 -1195 -75 -1165
rect -45 -1195 5 -1165
rect 35 -1195 85 -1165
rect 115 -1195 165 -1165
rect 195 -1195 245 -1165
rect 275 -1195 325 -1165
rect 355 -1195 405 -1165
rect 435 -1195 485 -1165
rect 515 -1195 565 -1165
rect 595 -1195 645 -1165
rect 675 -1195 725 -1165
rect 755 -1195 805 -1165
rect 835 -1195 885 -1165
rect 915 -1195 965 -1165
rect 995 -1195 1045 -1165
rect 1075 -1195 1125 -1165
rect 1155 -1195 1205 -1165
rect 1235 -1195 1285 -1165
rect 1315 -1195 1365 -1165
rect 1395 -1195 1445 -1165
rect 1475 -1195 1525 -1165
rect 1555 -1195 1605 -1165
rect 1635 -1195 1685 -1165
rect 1715 -1195 1765 -1165
rect 1795 -1195 1845 -1165
rect 1875 -1195 1925 -1165
rect 1955 -1195 2005 -1165
rect 2035 -1195 2085 -1165
rect 2115 -1195 2165 -1165
rect 2195 -1195 2245 -1165
rect 2275 -1195 2325 -1165
rect 2355 -1195 2405 -1165
rect 2435 -1195 2485 -1165
rect 2515 -1195 2565 -1165
rect 2595 -1195 2645 -1165
rect 2675 -1195 2725 -1165
rect 2755 -1195 2805 -1165
rect 2835 -1195 2885 -1165
rect 2915 -1195 2965 -1165
rect 2995 -1195 3045 -1165
rect 3075 -1195 3125 -1165
rect 3155 -1195 3205 -1165
rect 3235 -1195 3285 -1165
rect 3315 -1195 3365 -1165
rect 3395 -1195 3445 -1165
rect 3475 -1195 3525 -1165
rect 3555 -1195 3605 -1165
rect 3635 -1195 3685 -1165
rect 3715 -1195 3765 -1165
rect 3795 -1195 3845 -1165
rect 3875 -1195 3925 -1165
rect 3955 -1195 4005 -1165
rect 4035 -1195 4085 -1165
rect 4115 -1195 4165 -1165
rect 4195 -1195 4245 -1165
rect 4275 -1195 4325 -1165
rect 4355 -1195 4405 -1165
rect 4435 -1195 4485 -1165
rect 4515 -1195 4565 -1165
rect 4595 -1195 4645 -1165
rect 4675 -1195 4725 -1165
rect 4755 -1195 4805 -1165
rect 4835 -1195 4885 -1165
rect 4915 -1195 4965 -1165
rect 4995 -1195 5045 -1165
rect 5075 -1195 5125 -1165
rect 5155 -1195 5205 -1165
rect 5235 -1195 5240 -1165
rect -240 -1200 5240 -1195
rect -80 -1430 -75 -1360
rect -45 -1430 -40 -1360
rect -80 -1440 -40 -1430
rect 1200 -1430 1205 -1360
rect 1235 -1430 1240 -1360
rect 1200 -1440 1240 -1430
rect 2480 -1430 2485 -1360
rect 2515 -1430 2520 -1360
rect 2480 -1440 2520 -1430
rect 3760 -1430 3765 -1360
rect 3795 -1430 3800 -1360
rect 3760 -1440 3800 -1430
rect 5040 -1430 5045 -1360
rect 5075 -1430 5080 -1360
rect 5040 -1440 5080 -1430
<< via2 >>
rect -75 450 -45 630
rect 1205 450 1235 630
rect 2485 450 2515 630
rect 3765 450 3795 630
rect 5045 450 5075 630
rect -235 5 -205 35
rect -155 5 -125 35
rect -75 5 -45 35
rect 5 5 35 35
rect 85 5 115 35
rect 165 5 195 35
rect 325 5 355 35
rect 405 5 435 35
rect 485 5 515 35
rect 565 5 595 35
rect 645 5 675 35
rect 725 5 755 35
rect 805 5 835 35
rect 965 5 995 35
rect 1045 5 1075 35
rect 1125 5 1155 35
rect 1205 5 1235 35
rect 1285 5 1315 35
rect 1365 5 1395 35
rect 1445 5 1475 35
rect 1605 5 1635 35
rect 1685 5 1715 35
rect 1765 5 1795 35
rect 1845 5 1875 35
rect 1925 5 1955 35
rect 2005 5 2035 35
rect 2085 5 2115 35
rect 2245 5 2275 35
rect 2325 5 2355 35
rect 2405 5 2435 35
rect 2485 5 2515 35
rect 2565 5 2595 35
rect 2645 5 2675 35
rect 2725 5 2755 35
rect 2885 5 2915 35
rect 2965 5 2995 35
rect 3045 5 3075 35
rect 3125 5 3155 35
rect 3205 5 3235 35
rect 3285 5 3315 35
rect 3365 5 3395 35
rect 3525 5 3555 35
rect 3605 5 3635 35
rect 3685 5 3715 35
rect 3765 5 3795 35
rect 3845 5 3875 35
rect 3925 5 3955 35
rect 4005 5 4035 35
rect 4165 5 4195 35
rect 4245 5 4275 35
rect 4325 5 4355 35
rect 4405 5 4435 35
rect 4485 5 4515 35
rect 4565 5 4595 35
rect 4645 5 4675 35
rect 4805 5 4835 35
rect 4885 5 4915 35
rect 4965 5 4995 35
rect 5045 5 5075 35
rect 5125 5 5155 35
rect 5205 5 5235 35
rect -235 -155 -205 -125
rect -155 -155 -125 -125
rect -75 -155 -45 -125
rect 5 -155 35 -125
rect 85 -155 115 -125
rect 165 -155 195 -125
rect 325 -155 355 -125
rect 405 -155 435 -125
rect 485 -155 515 -125
rect 565 -155 595 -125
rect 645 -155 675 -125
rect 725 -155 755 -125
rect 805 -155 835 -125
rect 965 -155 995 -125
rect 1045 -155 1075 -125
rect 1125 -155 1155 -125
rect 1205 -155 1235 -125
rect 1285 -155 1315 -125
rect 1365 -155 1395 -125
rect 1445 -155 1475 -125
rect 1605 -155 1635 -125
rect 1685 -155 1715 -125
rect 1765 -155 1795 -125
rect 1845 -155 1875 -125
rect 1925 -155 1955 -125
rect 2005 -155 2035 -125
rect 2085 -155 2115 -125
rect 2245 -155 2275 -125
rect 2325 -155 2355 -125
rect 2405 -155 2435 -125
rect 2485 -155 2515 -125
rect 2565 -155 2595 -125
rect 2645 -155 2675 -125
rect 2725 -155 2755 -125
rect 2885 -155 2915 -125
rect 2965 -155 2995 -125
rect 3045 -155 3075 -125
rect 3125 -155 3155 -125
rect 3205 -155 3235 -125
rect 3285 -155 3315 -125
rect 3365 -155 3395 -125
rect 3525 -155 3555 -125
rect 3605 -155 3635 -125
rect 3685 -155 3715 -125
rect 3765 -155 3795 -125
rect 3845 -155 3875 -125
rect 3925 -155 3955 -125
rect 4005 -155 4035 -125
rect 4165 -155 4195 -125
rect 4245 -155 4275 -125
rect 4325 -155 4355 -125
rect 4405 -155 4435 -125
rect 4485 -155 4515 -125
rect 4565 -155 4595 -125
rect 4645 -155 4675 -125
rect 4805 -155 4835 -125
rect 4885 -155 4915 -125
rect 4965 -155 4995 -125
rect 5045 -155 5075 -125
rect 5125 -155 5155 -125
rect 5205 -155 5235 -125
rect -235 -715 -205 -685
rect -155 -715 -125 -685
rect -75 -715 -45 -685
rect 5 -715 35 -685
rect 85 -715 115 -685
rect 165 -715 195 -685
rect 245 -715 275 -685
rect 325 -715 355 -685
rect 405 -715 435 -685
rect 485 -715 515 -685
rect 565 -715 595 -685
rect 645 -715 675 -685
rect 725 -715 755 -685
rect 805 -715 835 -685
rect 885 -715 915 -685
rect 965 -715 995 -685
rect 1045 -715 1075 -685
rect 1125 -715 1155 -685
rect 1205 -715 1235 -685
rect 1285 -715 1315 -685
rect 1365 -715 1395 -685
rect 1445 -715 1475 -685
rect 1525 -715 1555 -685
rect 1605 -715 1635 -685
rect 1685 -715 1715 -685
rect 1765 -715 1795 -685
rect 1845 -715 1875 -685
rect 1925 -715 1955 -685
rect 2005 -715 2035 -685
rect 2085 -715 2115 -685
rect 2165 -715 2195 -685
rect 2245 -715 2275 -685
rect 2325 -715 2355 -685
rect 2405 -715 2435 -685
rect 2485 -715 2515 -685
rect 2565 -715 2595 -685
rect 2645 -715 2675 -685
rect 2725 -715 2755 -685
rect 2805 -715 2835 -685
rect 2885 -715 2915 -685
rect 2965 -715 2995 -685
rect 3045 -715 3075 -685
rect 3125 -715 3155 -685
rect 3205 -715 3235 -685
rect 3285 -715 3315 -685
rect 3365 -715 3395 -685
rect 3445 -715 3475 -685
rect 3525 -715 3555 -685
rect 3605 -715 3635 -685
rect 3685 -715 3715 -685
rect 3765 -715 3795 -685
rect 3845 -715 3875 -685
rect 3925 -715 3955 -685
rect 4005 -715 4035 -685
rect 4085 -715 4115 -685
rect 4165 -715 4195 -685
rect 4245 -715 4275 -685
rect 4325 -715 4355 -685
rect 4405 -715 4435 -685
rect 4485 -715 4515 -685
rect 4565 -715 4595 -685
rect 4645 -715 4675 -685
rect 4725 -715 4755 -685
rect 4805 -715 4835 -685
rect 4885 -715 4915 -685
rect 4965 -715 4995 -685
rect 5045 -715 5075 -685
rect 5125 -715 5155 -685
rect 5205 -715 5235 -685
rect -235 -875 -205 -845
rect -155 -875 -125 -845
rect -75 -875 -45 -845
rect 5 -875 35 -845
rect 85 -875 115 -845
rect 165 -875 195 -845
rect 245 -875 275 -845
rect 325 -875 355 -845
rect 405 -875 435 -845
rect 485 -875 515 -845
rect 565 -875 595 -845
rect 645 -875 675 -845
rect 725 -875 755 -845
rect 805 -875 835 -845
rect 885 -875 915 -845
rect 965 -875 995 -845
rect 1045 -875 1075 -845
rect 1125 -875 1155 -845
rect 1205 -875 1235 -845
rect 1285 -875 1315 -845
rect 1365 -875 1395 -845
rect 1445 -875 1475 -845
rect 1525 -875 1555 -845
rect 1605 -875 1635 -845
rect 1685 -875 1715 -845
rect 1765 -875 1795 -845
rect 1845 -875 1875 -845
rect 1925 -875 1955 -845
rect 2005 -875 2035 -845
rect 2085 -875 2115 -845
rect 2165 -875 2195 -845
rect 2245 -875 2275 -845
rect 2325 -875 2355 -845
rect 2405 -875 2435 -845
rect 2485 -875 2515 -845
rect 2565 -875 2595 -845
rect 2645 -875 2675 -845
rect 2725 -875 2755 -845
rect 2805 -875 2835 -845
rect 2885 -875 2915 -845
rect 2965 -875 2995 -845
rect 3045 -875 3075 -845
rect 3125 -875 3155 -845
rect 3205 -875 3235 -845
rect 3285 -875 3315 -845
rect 3365 -875 3395 -845
rect 3445 -875 3475 -845
rect 3525 -875 3555 -845
rect 3605 -875 3635 -845
rect 3685 -875 3715 -845
rect 3765 -875 3795 -845
rect 3845 -875 3875 -845
rect 3925 -875 3955 -845
rect 4005 -875 4035 -845
rect 4085 -875 4115 -845
rect 4165 -875 4195 -845
rect 4245 -875 4275 -845
rect 4325 -875 4355 -845
rect 4405 -875 4435 -845
rect 4485 -875 4515 -845
rect 4565 -875 4595 -845
rect 4645 -875 4675 -845
rect 4725 -875 4755 -845
rect 4805 -875 4835 -845
rect 4885 -875 4915 -845
rect 4965 -875 4995 -845
rect 5045 -875 5075 -845
rect 5125 -875 5155 -845
rect 5205 -875 5235 -845
rect -235 -1035 -205 -1005
rect -155 -1035 -125 -1005
rect -75 -1035 -45 -1005
rect 5 -1035 35 -1005
rect 85 -1035 115 -1005
rect 165 -1035 195 -1005
rect 245 -1035 275 -1005
rect 325 -1035 355 -1005
rect 405 -1035 435 -1005
rect 485 -1035 515 -1005
rect 565 -1035 595 -1005
rect 645 -1035 675 -1005
rect 725 -1035 755 -1005
rect 805 -1035 835 -1005
rect 885 -1035 915 -1005
rect 965 -1035 995 -1005
rect 1045 -1035 1075 -1005
rect 1125 -1035 1155 -1005
rect 1205 -1035 1235 -1005
rect 1285 -1035 1315 -1005
rect 1365 -1035 1395 -1005
rect 1445 -1035 1475 -1005
rect 1525 -1035 1555 -1005
rect 1605 -1035 1635 -1005
rect 1685 -1035 1715 -1005
rect 1765 -1035 1795 -1005
rect 1845 -1035 1875 -1005
rect 1925 -1035 1955 -1005
rect 2005 -1035 2035 -1005
rect 2085 -1035 2115 -1005
rect 2165 -1035 2195 -1005
rect 2245 -1035 2275 -1005
rect 2325 -1035 2355 -1005
rect 2405 -1035 2435 -1005
rect 2485 -1035 2515 -1005
rect 2565 -1035 2595 -1005
rect 2645 -1035 2675 -1005
rect 2725 -1035 2755 -1005
rect 2805 -1035 2835 -1005
rect 2885 -1035 2915 -1005
rect 2965 -1035 2995 -1005
rect 3045 -1035 3075 -1005
rect 3125 -1035 3155 -1005
rect 3205 -1035 3235 -1005
rect 3285 -1035 3315 -1005
rect 3365 -1035 3395 -1005
rect 3445 -1035 3475 -1005
rect 3525 -1035 3555 -1005
rect 3605 -1035 3635 -1005
rect 3685 -1035 3715 -1005
rect 3765 -1035 3795 -1005
rect 3845 -1035 3875 -1005
rect 3925 -1035 3955 -1005
rect 4005 -1035 4035 -1005
rect 4085 -1035 4115 -1005
rect 4165 -1035 4195 -1005
rect 4245 -1035 4275 -1005
rect 4325 -1035 4355 -1005
rect 4405 -1035 4435 -1005
rect 4485 -1035 4515 -1005
rect 4565 -1035 4595 -1005
rect 4645 -1035 4675 -1005
rect 4725 -1035 4755 -1005
rect 4805 -1035 4835 -1005
rect 4885 -1035 4915 -1005
rect 4965 -1035 4995 -1005
rect 5045 -1035 5075 -1005
rect 5125 -1035 5155 -1005
rect 5205 -1035 5235 -1005
rect -235 -1195 -205 -1165
rect -155 -1195 -125 -1165
rect -75 -1195 -45 -1165
rect 5 -1195 35 -1165
rect 85 -1195 115 -1165
rect 165 -1195 195 -1165
rect 245 -1195 275 -1165
rect 325 -1195 355 -1165
rect 405 -1195 435 -1165
rect 485 -1195 515 -1165
rect 565 -1195 595 -1165
rect 645 -1195 675 -1165
rect 725 -1195 755 -1165
rect 805 -1195 835 -1165
rect 885 -1195 915 -1165
rect 965 -1195 995 -1165
rect 1045 -1195 1075 -1165
rect 1125 -1195 1155 -1165
rect 1205 -1195 1235 -1165
rect 1285 -1195 1315 -1165
rect 1365 -1195 1395 -1165
rect 1445 -1195 1475 -1165
rect 1525 -1195 1555 -1165
rect 1605 -1195 1635 -1165
rect 1685 -1195 1715 -1165
rect 1765 -1195 1795 -1165
rect 1845 -1195 1875 -1165
rect 1925 -1195 1955 -1165
rect 2005 -1195 2035 -1165
rect 2085 -1195 2115 -1165
rect 2165 -1195 2195 -1165
rect 2245 -1195 2275 -1165
rect 2325 -1195 2355 -1165
rect 2405 -1195 2435 -1165
rect 2485 -1195 2515 -1165
rect 2565 -1195 2595 -1165
rect 2645 -1195 2675 -1165
rect 2725 -1195 2755 -1165
rect 2805 -1195 2835 -1165
rect 2885 -1195 2915 -1165
rect 2965 -1195 2995 -1165
rect 3045 -1195 3075 -1165
rect 3125 -1195 3155 -1165
rect 3205 -1195 3235 -1165
rect 3285 -1195 3315 -1165
rect 3365 -1195 3395 -1165
rect 3445 -1195 3475 -1165
rect 3525 -1195 3555 -1165
rect 3605 -1195 3635 -1165
rect 3685 -1195 3715 -1165
rect 3765 -1195 3795 -1165
rect 3845 -1195 3875 -1165
rect 3925 -1195 3955 -1165
rect 4005 -1195 4035 -1165
rect 4085 -1195 4115 -1165
rect 4165 -1195 4195 -1165
rect 4245 -1195 4275 -1165
rect 4325 -1195 4355 -1165
rect 4405 -1195 4435 -1165
rect 4485 -1195 4515 -1165
rect 4565 -1195 4595 -1165
rect 4645 -1195 4675 -1165
rect 4725 -1195 4755 -1165
rect 4805 -1195 4835 -1165
rect 4885 -1195 4915 -1165
rect 4965 -1195 4995 -1165
rect 5045 -1195 5075 -1165
rect 5125 -1195 5155 -1165
rect 5205 -1195 5235 -1165
rect -75 -1430 -45 -1360
rect 1205 -1430 1235 -1360
rect 2485 -1430 2515 -1360
rect 3765 -1430 3795 -1360
rect 5045 -1430 5075 -1360
<< metal3 >>
rect -80 631 -40 680
rect -80 449 -76 631
rect -44 449 -40 631
rect -240 35 -200 40
rect -240 5 -235 35
rect -205 5 -200 35
rect -240 -125 -200 5
rect -240 -155 -235 -125
rect -205 -155 -200 -125
rect -240 -240 -200 -155
rect -160 35 -120 40
rect -160 5 -155 35
rect -125 5 -120 35
rect -160 -125 -120 5
rect -160 -155 -155 -125
rect -125 -155 -120 -125
rect -160 -240 -120 -155
rect -80 35 -40 449
rect 1200 631 1240 680
rect 1200 449 1204 631
rect 1236 449 1240 631
rect 1200 360 1240 449
rect 2480 631 2520 680
rect 2480 449 2484 631
rect 2516 449 2520 631
rect 2480 360 2520 449
rect 3760 631 3800 680
rect 3760 449 3764 631
rect 3796 449 3800 631
rect 3760 360 3800 449
rect 5040 631 5080 680
rect 5040 449 5044 631
rect 5076 449 5080 631
rect -80 5 -75 35
rect -45 5 -40 35
rect -80 -125 -40 5
rect -80 -155 -75 -125
rect -45 -155 -40 -125
rect -80 -240 -40 -155
rect 0 35 40 40
rect 0 5 5 35
rect 35 5 40 35
rect 0 -125 40 5
rect 0 -155 5 -125
rect 35 -155 40 -125
rect 0 -240 40 -155
rect 80 35 120 40
rect 80 5 85 35
rect 115 5 120 35
rect 80 -125 120 5
rect 80 -155 85 -125
rect 115 -155 120 -125
rect 80 -240 120 -155
rect 160 35 200 40
rect 160 5 165 35
rect 195 5 200 35
rect 160 -125 200 5
rect 160 -155 165 -125
rect 195 -155 200 -125
rect 160 -240 200 -155
rect 320 35 360 40
rect 320 5 325 35
rect 355 5 360 35
rect 320 -125 360 5
rect 320 -155 325 -125
rect 355 -155 360 -125
rect 240 -240 280 -160
rect 320 -240 360 -155
rect 400 35 440 40
rect 400 5 405 35
rect 435 5 440 35
rect 400 -125 440 5
rect 400 -155 405 -125
rect 435 -155 440 -125
rect 400 -240 440 -155
rect 480 35 520 40
rect 480 5 485 35
rect 515 5 520 35
rect 480 -125 520 5
rect 480 -155 485 -125
rect 515 -155 520 -125
rect 480 -240 520 -155
rect 560 35 600 40
rect 560 5 565 35
rect 595 5 600 35
rect 560 -125 600 5
rect 560 -155 565 -125
rect 595 -155 600 -125
rect 560 -240 600 -155
rect 640 35 680 40
rect 640 5 645 35
rect 675 5 680 35
rect 640 -125 680 5
rect 640 -155 645 -125
rect 675 -155 680 -125
rect 640 -240 680 -155
rect 720 35 760 40
rect 720 5 725 35
rect 755 5 760 35
rect 720 -125 760 5
rect 720 -155 725 -125
rect 755 -155 760 -125
rect 720 -240 760 -155
rect 800 35 840 40
rect 800 5 805 35
rect 835 5 840 35
rect 800 -125 840 5
rect 800 -155 805 -125
rect 835 -155 840 -125
rect 800 -240 840 -155
rect 960 35 1000 40
rect 960 5 965 35
rect 995 5 1000 35
rect 960 -125 1000 5
rect 960 -155 965 -125
rect 995 -155 1000 -125
rect 880 -240 920 -160
rect 960 -240 1000 -155
rect 1040 35 1080 40
rect 1040 5 1045 35
rect 1075 5 1080 35
rect 1040 -125 1080 5
rect 1040 -155 1045 -125
rect 1075 -155 1080 -125
rect 1040 -240 1080 -155
rect 1120 35 1160 40
rect 1120 5 1125 35
rect 1155 5 1160 35
rect 1120 -125 1160 5
rect 1120 -155 1125 -125
rect 1155 -155 1160 -125
rect 1120 -240 1160 -155
rect 1200 35 1240 40
rect 1200 5 1205 35
rect 1235 5 1240 35
rect 1200 -125 1240 5
rect 1200 -155 1205 -125
rect 1235 -155 1240 -125
rect 1200 -240 1240 -155
rect 1280 35 1320 40
rect 1280 5 1285 35
rect 1315 5 1320 35
rect 1280 -125 1320 5
rect 1280 -155 1285 -125
rect 1315 -155 1320 -125
rect 1280 -240 1320 -155
rect 1360 35 1400 40
rect 1360 5 1365 35
rect 1395 5 1400 35
rect 1360 -125 1400 5
rect 1360 -155 1365 -125
rect 1395 -155 1400 -125
rect 1360 -240 1400 -155
rect 1440 35 1480 40
rect 1440 5 1445 35
rect 1475 5 1480 35
rect 1440 -125 1480 5
rect 1440 -155 1445 -125
rect 1475 -155 1480 -125
rect 1440 -240 1480 -155
rect 1600 35 1640 40
rect 1600 5 1605 35
rect 1635 5 1640 35
rect 1600 -125 1640 5
rect 1600 -155 1605 -125
rect 1635 -155 1640 -125
rect 1520 -240 1560 -160
rect 1600 -240 1640 -155
rect 1680 35 1720 40
rect 1680 5 1685 35
rect 1715 5 1720 35
rect 1680 -125 1720 5
rect 1680 -155 1685 -125
rect 1715 -155 1720 -125
rect 1680 -240 1720 -155
rect 1760 35 1800 40
rect 1760 5 1765 35
rect 1795 5 1800 35
rect 1760 -125 1800 5
rect 1760 -155 1765 -125
rect 1795 -155 1800 -125
rect 1760 -240 1800 -155
rect 1840 35 1880 40
rect 1840 5 1845 35
rect 1875 5 1880 35
rect 1840 -125 1880 5
rect 1840 -155 1845 -125
rect 1875 -155 1880 -125
rect 1840 -240 1880 -155
rect 1920 35 1960 40
rect 1920 5 1925 35
rect 1955 5 1960 35
rect 1920 -125 1960 5
rect 1920 -155 1925 -125
rect 1955 -155 1960 -125
rect 1920 -240 1960 -155
rect 2000 35 2040 40
rect 2000 5 2005 35
rect 2035 5 2040 35
rect 2000 -125 2040 5
rect 2000 -155 2005 -125
rect 2035 -155 2040 -125
rect 2000 -240 2040 -155
rect 2080 35 2120 40
rect 2080 5 2085 35
rect 2115 5 2120 35
rect 2080 -125 2120 5
rect 2080 -155 2085 -125
rect 2115 -155 2120 -125
rect 2080 -240 2120 -155
rect 2240 35 2280 40
rect 2240 5 2245 35
rect 2275 5 2280 35
rect 2240 -125 2280 5
rect 2240 -155 2245 -125
rect 2275 -155 2280 -125
rect 2160 -240 2200 -160
rect 2240 -240 2280 -155
rect 2320 35 2360 40
rect 2320 5 2325 35
rect 2355 5 2360 35
rect 2320 -125 2360 5
rect 2320 -155 2325 -125
rect 2355 -155 2360 -125
rect 2320 -240 2360 -155
rect 2400 35 2440 40
rect 2400 5 2405 35
rect 2435 5 2440 35
rect 2400 -125 2440 5
rect 2400 -155 2405 -125
rect 2435 -155 2440 -125
rect 2400 -240 2440 -155
rect 2480 35 2520 40
rect 2480 5 2485 35
rect 2515 5 2520 35
rect 2480 -125 2520 5
rect 2480 -155 2485 -125
rect 2515 -155 2520 -125
rect 2480 -240 2520 -155
rect 2560 35 2600 40
rect 2560 5 2565 35
rect 2595 5 2600 35
rect 2560 -125 2600 5
rect 2560 -155 2565 -125
rect 2595 -155 2600 -125
rect 2560 -240 2600 -155
rect 2640 35 2680 40
rect 2640 5 2645 35
rect 2675 5 2680 35
rect 2640 -125 2680 5
rect 2640 -155 2645 -125
rect 2675 -155 2680 -125
rect 2640 -240 2680 -155
rect 2720 35 2760 40
rect 2720 5 2725 35
rect 2755 5 2760 35
rect 2720 -125 2760 5
rect 2720 -155 2725 -125
rect 2755 -155 2760 -125
rect 2720 -240 2760 -155
rect 2880 35 2920 40
rect 2880 5 2885 35
rect 2915 5 2920 35
rect 2880 -125 2920 5
rect 2880 -155 2885 -125
rect 2915 -155 2920 -125
rect 2800 -240 2840 -160
rect 2880 -240 2920 -155
rect 2960 35 3000 40
rect 2960 5 2965 35
rect 2995 5 3000 35
rect 2960 -125 3000 5
rect 2960 -155 2965 -125
rect 2995 -155 3000 -125
rect 2960 -240 3000 -155
rect 3040 35 3080 40
rect 3040 5 3045 35
rect 3075 5 3080 35
rect 3040 -125 3080 5
rect 3040 -155 3045 -125
rect 3075 -155 3080 -125
rect 3040 -240 3080 -155
rect 3120 35 3160 40
rect 3120 5 3125 35
rect 3155 5 3160 35
rect 3120 -125 3160 5
rect 3120 -155 3125 -125
rect 3155 -155 3160 -125
rect 3120 -240 3160 -155
rect 3200 35 3240 40
rect 3200 5 3205 35
rect 3235 5 3240 35
rect 3200 -125 3240 5
rect 3200 -155 3205 -125
rect 3235 -155 3240 -125
rect 3200 -240 3240 -155
rect 3280 35 3320 40
rect 3280 5 3285 35
rect 3315 5 3320 35
rect 3280 -125 3320 5
rect 3280 -155 3285 -125
rect 3315 -155 3320 -125
rect 3280 -240 3320 -155
rect 3360 35 3400 40
rect 3360 5 3365 35
rect 3395 5 3400 35
rect 3360 -125 3400 5
rect 3360 -155 3365 -125
rect 3395 -155 3400 -125
rect 3360 -240 3400 -155
rect 3520 35 3560 40
rect 3520 5 3525 35
rect 3555 5 3560 35
rect 3520 -125 3560 5
rect 3520 -155 3525 -125
rect 3555 -155 3560 -125
rect 3440 -240 3480 -160
rect 3520 -240 3560 -155
rect 3600 35 3640 40
rect 3600 5 3605 35
rect 3635 5 3640 35
rect 3600 -125 3640 5
rect 3600 -155 3605 -125
rect 3635 -155 3640 -125
rect 3600 -240 3640 -155
rect 3680 35 3720 40
rect 3680 5 3685 35
rect 3715 5 3720 35
rect 3680 -125 3720 5
rect 3680 -155 3685 -125
rect 3715 -155 3720 -125
rect 3680 -240 3720 -155
rect 3760 35 3800 40
rect 3760 5 3765 35
rect 3795 5 3800 35
rect 3760 -125 3800 5
rect 3760 -155 3765 -125
rect 3795 -155 3800 -125
rect 3760 -240 3800 -155
rect 3840 35 3880 40
rect 3840 5 3845 35
rect 3875 5 3880 35
rect 3840 -125 3880 5
rect 3840 -155 3845 -125
rect 3875 -155 3880 -125
rect 3840 -240 3880 -155
rect 3920 35 3960 40
rect 3920 5 3925 35
rect 3955 5 3960 35
rect 3920 -125 3960 5
rect 3920 -155 3925 -125
rect 3955 -155 3960 -125
rect 3920 -240 3960 -155
rect 4000 35 4040 40
rect 4000 5 4005 35
rect 4035 5 4040 35
rect 4000 -125 4040 5
rect 4000 -155 4005 -125
rect 4035 -155 4040 -125
rect 4000 -240 4040 -155
rect 4160 35 4200 40
rect 4160 5 4165 35
rect 4195 5 4200 35
rect 4160 -125 4200 5
rect 4160 -155 4165 -125
rect 4195 -155 4200 -125
rect 4080 -240 4120 -160
rect 4160 -240 4200 -155
rect 4240 35 4280 40
rect 4240 5 4245 35
rect 4275 5 4280 35
rect 4240 -125 4280 5
rect 4240 -155 4245 -125
rect 4275 -155 4280 -125
rect 4240 -240 4280 -155
rect 4320 35 4360 40
rect 4320 5 4325 35
rect 4355 5 4360 35
rect 4320 -125 4360 5
rect 4320 -155 4325 -125
rect 4355 -155 4360 -125
rect 4320 -240 4360 -155
rect 4400 35 4440 40
rect 4400 5 4405 35
rect 4435 5 4440 35
rect 4400 -125 4440 5
rect 4400 -155 4405 -125
rect 4435 -155 4440 -125
rect 4400 -240 4440 -155
rect 4480 35 4520 40
rect 4480 5 4485 35
rect 4515 5 4520 35
rect 4480 -125 4520 5
rect 4480 -155 4485 -125
rect 4515 -155 4520 -125
rect 4480 -240 4520 -155
rect 4560 35 4600 40
rect 4560 5 4565 35
rect 4595 5 4600 35
rect 4560 -125 4600 5
rect 4560 -155 4565 -125
rect 4595 -155 4600 -125
rect 4560 -240 4600 -155
rect 4640 35 4680 40
rect 4640 5 4645 35
rect 4675 5 4680 35
rect 4640 -125 4680 5
rect 4640 -155 4645 -125
rect 4675 -155 4680 -125
rect 4640 -240 4680 -155
rect 4800 35 4840 40
rect 4800 5 4805 35
rect 4835 5 4840 35
rect 4800 -125 4840 5
rect 4800 -155 4805 -125
rect 4835 -155 4840 -125
rect 4720 -240 4760 -160
rect 4800 -240 4840 -155
rect 4880 35 4920 40
rect 4880 5 4885 35
rect 4915 5 4920 35
rect 4880 -125 4920 5
rect 4880 -155 4885 -125
rect 4915 -155 4920 -125
rect 4880 -240 4920 -155
rect 4960 35 5000 40
rect 4960 5 4965 35
rect 4995 5 5000 35
rect 4960 -125 5000 5
rect 4960 -155 4965 -125
rect 4995 -155 5000 -125
rect 4960 -240 5000 -155
rect 5040 35 5080 449
rect 5040 5 5045 35
rect 5075 5 5080 35
rect 5040 -125 5080 5
rect 5040 -155 5045 -125
rect 5075 -155 5080 -125
rect 5040 -240 5080 -155
rect 5120 35 5160 40
rect 5120 5 5125 35
rect 5155 5 5160 35
rect 5120 -125 5160 5
rect 5120 -155 5125 -125
rect 5155 -155 5160 -125
rect 5120 -240 5160 -155
rect 5200 35 5240 40
rect 5200 5 5205 35
rect 5235 5 5240 35
rect 5200 -125 5240 5
rect 5200 -155 5205 -125
rect 5235 -155 5240 -125
rect 5200 -240 5240 -155
rect -240 -400 -200 -280
rect -160 -400 -120 -280
rect -80 -400 -40 -280
rect 0 -400 40 -280
rect 80 -400 120 -280
rect 160 -400 200 -280
rect 240 -360 280 -280
rect 320 -400 360 -280
rect 400 -400 440 -280
rect 480 -400 520 -280
rect 560 -400 600 -280
rect 640 -400 680 -280
rect 720 -400 760 -280
rect 800 -400 840 -280
rect 880 -360 920 -280
rect 960 -400 1000 -280
rect 1040 -400 1080 -280
rect 1120 -400 1160 -280
rect 1200 -400 1240 -280
rect 1280 -400 1320 -280
rect 1360 -400 1400 -280
rect 1440 -400 1480 -280
rect 1520 -360 1560 -280
rect 1600 -400 1640 -280
rect 1680 -400 1720 -280
rect 1760 -400 1800 -280
rect 1840 -400 1880 -280
rect 1920 -400 1960 -280
rect 2000 -400 2040 -280
rect 2080 -400 2120 -280
rect 2160 -360 2200 -280
rect 2240 -400 2280 -280
rect 2320 -400 2360 -280
rect 2400 -400 2440 -280
rect 2480 -400 2520 -280
rect 2560 -400 2600 -280
rect 2640 -400 2680 -280
rect 2720 -400 2760 -280
rect 2800 -360 2840 -280
rect 2880 -400 2920 -280
rect 2960 -400 3000 -280
rect 3040 -400 3080 -280
rect 3120 -400 3160 -280
rect 3200 -400 3240 -280
rect 3280 -400 3320 -280
rect 3360 -400 3400 -280
rect 3440 -360 3480 -280
rect 3520 -400 3560 -280
rect 3600 -400 3640 -280
rect 3680 -400 3720 -280
rect 3760 -400 3800 -280
rect 3840 -400 3880 -280
rect 3920 -400 3960 -280
rect 4000 -400 4040 -280
rect 4080 -360 4120 -280
rect 4160 -400 4200 -280
rect 4240 -400 4280 -280
rect 4320 -400 4360 -280
rect 4400 -400 4440 -280
rect 4480 -400 4520 -280
rect 4560 -400 4600 -280
rect 4640 -400 4680 -280
rect 4720 -360 4760 -280
rect 4800 -400 4840 -280
rect 4880 -400 4920 -280
rect 4960 -400 5000 -280
rect 5040 -400 5080 -280
rect 5120 -400 5160 -280
rect 5200 -400 5240 -280
rect -240 -685 -200 -680
rect -240 -715 -235 -685
rect -205 -715 -200 -685
rect -240 -845 -200 -715
rect -240 -875 -235 -845
rect -205 -875 -200 -845
rect -240 -1005 -200 -875
rect -240 -1035 -235 -1005
rect -205 -1035 -200 -1005
rect -240 -1165 -200 -1035
rect -240 -1195 -235 -1165
rect -205 -1195 -200 -1165
rect -240 -1360 -200 -1195
rect -160 -685 -120 -680
rect -160 -715 -155 -685
rect -125 -715 -120 -685
rect -160 -840 -120 -715
rect -80 -685 -40 -680
rect -80 -715 -75 -685
rect -45 -715 -40 -685
rect -80 -840 -40 -715
rect 0 -685 40 -680
rect 0 -715 5 -685
rect 35 -715 40 -685
rect 0 -840 40 -715
rect 80 -685 120 -680
rect 80 -715 85 -685
rect 115 -715 120 -685
rect 80 -840 120 -715
rect 160 -685 200 -680
rect 160 -715 165 -685
rect 195 -715 200 -685
rect 160 -840 200 -715
rect 240 -685 280 -680
rect 240 -715 245 -685
rect 275 -715 280 -685
rect 240 -840 280 -715
rect 320 -685 360 -680
rect 320 -715 325 -685
rect 355 -715 360 -685
rect 320 -840 360 -715
rect 400 -685 440 -680
rect 400 -715 405 -685
rect 435 -715 440 -685
rect 400 -840 440 -715
rect 480 -685 520 -680
rect 480 -715 485 -685
rect 515 -715 520 -685
rect 480 -840 520 -715
rect 560 -685 600 -680
rect 560 -715 565 -685
rect 595 -715 600 -685
rect 560 -840 600 -715
rect 640 -685 680 -680
rect 640 -715 645 -685
rect 675 -715 680 -685
rect 640 -840 680 -715
rect 720 -685 760 -680
rect 720 -715 725 -685
rect 755 -715 760 -685
rect 720 -840 760 -715
rect 800 -685 840 -680
rect 800 -715 805 -685
rect 835 -715 840 -685
rect 800 -840 840 -715
rect 880 -685 920 -680
rect 880 -715 885 -685
rect 915 -715 920 -685
rect 880 -840 920 -715
rect 960 -685 1000 -680
rect 960 -715 965 -685
rect 995 -715 1000 -685
rect 960 -840 1000 -715
rect 1040 -685 1080 -680
rect 1040 -715 1045 -685
rect 1075 -715 1080 -685
rect 1040 -840 1080 -715
rect 1120 -685 1160 -680
rect 1120 -715 1125 -685
rect 1155 -715 1160 -685
rect 1120 -840 1160 -715
rect 1200 -685 1240 -680
rect 1200 -715 1205 -685
rect 1235 -715 1240 -685
rect 1200 -840 1240 -715
rect 1280 -685 1320 -680
rect 1280 -715 1285 -685
rect 1315 -715 1320 -685
rect 1280 -840 1320 -715
rect 1360 -685 1400 -680
rect 1360 -715 1365 -685
rect 1395 -715 1400 -685
rect 1360 -840 1400 -715
rect 1440 -685 1480 -680
rect 1440 -715 1445 -685
rect 1475 -715 1480 -685
rect 1440 -840 1480 -715
rect 1520 -685 1560 -680
rect 1520 -715 1525 -685
rect 1555 -715 1560 -685
rect 1520 -840 1560 -715
rect 1600 -685 1640 -680
rect 1600 -715 1605 -685
rect 1635 -715 1640 -685
rect 1600 -840 1640 -715
rect 1680 -685 1720 -680
rect 1680 -715 1685 -685
rect 1715 -715 1720 -685
rect 1680 -840 1720 -715
rect 1760 -685 1800 -680
rect 1760 -715 1765 -685
rect 1795 -715 1800 -685
rect 1760 -840 1800 -715
rect 1840 -685 1880 -680
rect 1840 -715 1845 -685
rect 1875 -715 1880 -685
rect 1840 -840 1880 -715
rect 1920 -685 1960 -680
rect 1920 -715 1925 -685
rect 1955 -715 1960 -685
rect 1920 -840 1960 -715
rect 2000 -685 2040 -680
rect 2000 -715 2005 -685
rect 2035 -715 2040 -685
rect 2000 -840 2040 -715
rect 2080 -685 2120 -680
rect 2080 -715 2085 -685
rect 2115 -715 2120 -685
rect 2080 -840 2120 -715
rect 2160 -685 2200 -680
rect 2160 -715 2165 -685
rect 2195 -715 2200 -685
rect 2160 -840 2200 -715
rect 2240 -685 2280 -680
rect 2240 -715 2245 -685
rect 2275 -715 2280 -685
rect 2240 -840 2280 -715
rect 2320 -685 2360 -680
rect 2320 -715 2325 -685
rect 2355 -715 2360 -685
rect 2320 -840 2360 -715
rect 2400 -685 2440 -680
rect 2400 -715 2405 -685
rect 2435 -715 2440 -685
rect 2400 -840 2440 -715
rect 2480 -685 2520 -680
rect 2480 -715 2485 -685
rect 2515 -715 2520 -685
rect 2480 -840 2520 -715
rect 2560 -685 2600 -680
rect 2560 -715 2565 -685
rect 2595 -715 2600 -685
rect 2560 -840 2600 -715
rect 2640 -685 2680 -680
rect 2640 -715 2645 -685
rect 2675 -715 2680 -685
rect 2640 -840 2680 -715
rect 2720 -685 2760 -680
rect 2720 -715 2725 -685
rect 2755 -715 2760 -685
rect 2720 -840 2760 -715
rect 2800 -685 2840 -680
rect 2800 -715 2805 -685
rect 2835 -715 2840 -685
rect 2800 -840 2840 -715
rect 2880 -685 2920 -680
rect 2880 -715 2885 -685
rect 2915 -715 2920 -685
rect 2880 -840 2920 -715
rect 2960 -685 3000 -680
rect 2960 -715 2965 -685
rect 2995 -715 3000 -685
rect 2960 -840 3000 -715
rect 3040 -685 3080 -680
rect 3040 -715 3045 -685
rect 3075 -715 3080 -685
rect 3040 -840 3080 -715
rect 3120 -685 3160 -680
rect 3120 -715 3125 -685
rect 3155 -715 3160 -685
rect 3120 -840 3160 -715
rect 3200 -685 3240 -680
rect 3200 -715 3205 -685
rect 3235 -715 3240 -685
rect 3200 -840 3240 -715
rect 3280 -685 3320 -680
rect 3280 -715 3285 -685
rect 3315 -715 3320 -685
rect 3280 -840 3320 -715
rect 3360 -685 3400 -680
rect 3360 -715 3365 -685
rect 3395 -715 3400 -685
rect 3360 -840 3400 -715
rect 3440 -685 3480 -680
rect 3440 -715 3445 -685
rect 3475 -715 3480 -685
rect 3440 -840 3480 -715
rect 3520 -685 3560 -680
rect 3520 -715 3525 -685
rect 3555 -715 3560 -685
rect 3520 -840 3560 -715
rect 3600 -685 3640 -680
rect 3600 -715 3605 -685
rect 3635 -715 3640 -685
rect 3600 -840 3640 -715
rect 3680 -685 3720 -680
rect 3680 -715 3685 -685
rect 3715 -715 3720 -685
rect 3680 -840 3720 -715
rect 3760 -685 3800 -680
rect 3760 -715 3765 -685
rect 3795 -715 3800 -685
rect 3760 -840 3800 -715
rect 3840 -685 3880 -680
rect 3840 -715 3845 -685
rect 3875 -715 3880 -685
rect 3840 -840 3880 -715
rect 3920 -685 3960 -680
rect 3920 -715 3925 -685
rect 3955 -715 3960 -685
rect 3920 -840 3960 -715
rect 4000 -685 4040 -680
rect 4000 -715 4005 -685
rect 4035 -715 4040 -685
rect 4000 -840 4040 -715
rect 4080 -685 4120 -680
rect 4080 -715 4085 -685
rect 4115 -715 4120 -685
rect 4080 -840 4120 -715
rect 4160 -685 4200 -680
rect 4160 -715 4165 -685
rect 4195 -715 4200 -685
rect 4160 -840 4200 -715
rect 4240 -685 4280 -680
rect 4240 -715 4245 -685
rect 4275 -715 4280 -685
rect 4240 -840 4280 -715
rect 4320 -685 4360 -680
rect 4320 -715 4325 -685
rect 4355 -715 4360 -685
rect 4320 -840 4360 -715
rect 4400 -685 4440 -680
rect 4400 -715 4405 -685
rect 4435 -715 4440 -685
rect 4400 -840 4440 -715
rect 4480 -685 4520 -680
rect 4480 -715 4485 -685
rect 4515 -715 4520 -685
rect 4480 -840 4520 -715
rect 4560 -685 4600 -680
rect 4560 -715 4565 -685
rect 4595 -715 4600 -685
rect 4560 -840 4600 -715
rect 4640 -685 4680 -680
rect 4640 -715 4645 -685
rect 4675 -715 4680 -685
rect 4640 -840 4680 -715
rect 4720 -685 4760 -680
rect 4720 -715 4725 -685
rect 4755 -715 4760 -685
rect 4720 -840 4760 -715
rect 4800 -685 4840 -680
rect 4800 -715 4805 -685
rect 4835 -715 4840 -685
rect 4800 -840 4840 -715
rect 4880 -685 4920 -680
rect 4880 -715 4885 -685
rect 4915 -715 4920 -685
rect 4880 -840 4920 -715
rect 4960 -685 5000 -680
rect 4960 -715 4965 -685
rect 4995 -715 5000 -685
rect 4960 -840 5000 -715
rect 5040 -685 5080 -680
rect 5040 -715 5045 -685
rect 5075 -715 5080 -685
rect 5040 -840 5080 -715
rect 5120 -685 5160 -680
rect 5120 -715 5125 -685
rect 5155 -715 5160 -685
rect 5120 -840 5160 -715
rect -160 -845 5160 -840
rect -160 -875 -155 -845
rect -125 -875 -75 -845
rect -45 -875 5 -845
rect 35 -875 85 -845
rect 115 -875 165 -845
rect 195 -875 245 -845
rect 275 -875 325 -845
rect 355 -875 405 -845
rect 435 -875 485 -845
rect 515 -875 565 -845
rect 595 -875 645 -845
rect 675 -875 725 -845
rect 755 -875 805 -845
rect 835 -875 885 -845
rect 915 -875 965 -845
rect 995 -875 1045 -845
rect 1075 -875 1125 -845
rect 1155 -875 1205 -845
rect 1235 -875 1285 -845
rect 1315 -875 1365 -845
rect 1395 -875 1445 -845
rect 1475 -875 1525 -845
rect 1555 -875 1605 -845
rect 1635 -875 1685 -845
rect 1715 -875 1765 -845
rect 1795 -875 1845 -845
rect 1875 -875 1925 -845
rect 1955 -875 2005 -845
rect 2035 -875 2085 -845
rect 2115 -875 2165 -845
rect 2195 -875 2245 -845
rect 2275 -875 2325 -845
rect 2355 -875 2405 -845
rect 2435 -875 2485 -845
rect 2515 -875 2565 -845
rect 2595 -875 2645 -845
rect 2675 -875 2725 -845
rect 2755 -875 2805 -845
rect 2835 -875 2885 -845
rect 2915 -875 2965 -845
rect 2995 -875 3045 -845
rect 3075 -875 3125 -845
rect 3155 -875 3205 -845
rect 3235 -875 3285 -845
rect 3315 -875 3365 -845
rect 3395 -875 3445 -845
rect 3475 -875 3525 -845
rect 3555 -875 3605 -845
rect 3635 -875 3685 -845
rect 3715 -875 3765 -845
rect 3795 -875 3845 -845
rect 3875 -875 3925 -845
rect 3955 -875 4005 -845
rect 4035 -875 4085 -845
rect 4115 -875 4165 -845
rect 4195 -875 4245 -845
rect 4275 -875 4325 -845
rect 4355 -875 4405 -845
rect 4435 -875 4485 -845
rect 4515 -875 4565 -845
rect 4595 -875 4645 -845
rect 4675 -875 4725 -845
rect 4755 -875 4805 -845
rect 4835 -875 4885 -845
rect 4915 -875 4965 -845
rect 4995 -875 5045 -845
rect 5075 -875 5125 -845
rect 5155 -875 5160 -845
rect -160 -880 5160 -875
rect -160 -1005 -120 -880
rect -160 -1035 -155 -1005
rect -125 -1035 -120 -1005
rect -160 -1165 -120 -1035
rect -160 -1195 -155 -1165
rect -125 -1195 -120 -1165
rect -160 -1360 -120 -1195
rect -80 -1005 -40 -880
rect -80 -1035 -75 -1005
rect -45 -1035 -40 -1005
rect -80 -1165 -40 -1035
rect -80 -1195 -75 -1165
rect -45 -1195 -40 -1165
rect -80 -1349 -40 -1195
rect -80 -1431 -76 -1349
rect -44 -1431 -40 -1349
rect 0 -1005 40 -880
rect 0 -1035 5 -1005
rect 35 -1035 40 -1005
rect 0 -1165 40 -1035
rect 0 -1195 5 -1165
rect 35 -1195 40 -1165
rect 0 -1360 40 -1195
rect 80 -1005 120 -880
rect 80 -1035 85 -1005
rect 115 -1035 120 -1005
rect 80 -1165 120 -1035
rect 80 -1195 85 -1165
rect 115 -1195 120 -1165
rect 80 -1360 120 -1195
rect 160 -1005 200 -880
rect 160 -1035 165 -1005
rect 195 -1035 200 -1005
rect 160 -1165 200 -1035
rect 160 -1195 165 -1165
rect 195 -1195 200 -1165
rect 160 -1360 200 -1195
rect 240 -1005 280 -880
rect 240 -1035 245 -1005
rect 275 -1035 280 -1005
rect 240 -1165 280 -1035
rect 240 -1195 245 -1165
rect 275 -1195 280 -1165
rect 240 -1360 280 -1195
rect 320 -1005 360 -880
rect 320 -1035 325 -1005
rect 355 -1035 360 -1005
rect 320 -1165 360 -1035
rect 320 -1195 325 -1165
rect 355 -1195 360 -1165
rect 320 -1360 360 -1195
rect 400 -1005 440 -880
rect 400 -1035 405 -1005
rect 435 -1035 440 -1005
rect 400 -1165 440 -1035
rect 400 -1195 405 -1165
rect 435 -1195 440 -1165
rect 400 -1360 440 -1195
rect 480 -1005 520 -880
rect 480 -1035 485 -1005
rect 515 -1035 520 -1005
rect 480 -1165 520 -1035
rect 480 -1195 485 -1165
rect 515 -1195 520 -1165
rect 480 -1360 520 -1195
rect 560 -1005 600 -880
rect 560 -1035 565 -1005
rect 595 -1035 600 -1005
rect 560 -1165 600 -1035
rect 560 -1195 565 -1165
rect 595 -1195 600 -1165
rect 560 -1200 600 -1195
rect 640 -1005 680 -880
rect 640 -1035 645 -1005
rect 675 -1035 680 -1005
rect 640 -1165 680 -1035
rect 640 -1195 645 -1165
rect 675 -1195 680 -1165
rect 640 -1360 680 -1195
rect 720 -1005 760 -880
rect 720 -1035 725 -1005
rect 755 -1035 760 -1005
rect 720 -1165 760 -1035
rect 720 -1195 725 -1165
rect 755 -1195 760 -1165
rect 720 -1360 760 -1195
rect 800 -1005 840 -880
rect 800 -1035 805 -1005
rect 835 -1035 840 -1005
rect 800 -1165 840 -1035
rect 800 -1195 805 -1165
rect 835 -1195 840 -1165
rect 800 -1360 840 -1195
rect 880 -1005 920 -880
rect 880 -1035 885 -1005
rect 915 -1035 920 -1005
rect 880 -1165 920 -1035
rect 880 -1195 885 -1165
rect 915 -1195 920 -1165
rect 880 -1360 920 -1195
rect 960 -1005 1000 -880
rect 960 -1035 965 -1005
rect 995 -1035 1000 -1005
rect 960 -1165 1000 -1035
rect 960 -1195 965 -1165
rect 995 -1195 1000 -1165
rect 960 -1360 1000 -1195
rect 1040 -1005 1080 -880
rect 1040 -1035 1045 -1005
rect 1075 -1035 1080 -1005
rect 1040 -1165 1080 -1035
rect 1040 -1195 1045 -1165
rect 1075 -1195 1080 -1165
rect 1040 -1360 1080 -1195
rect 1120 -1005 1160 -880
rect 1120 -1035 1125 -1005
rect 1155 -1035 1160 -1005
rect 1120 -1165 1160 -1035
rect 1120 -1195 1125 -1165
rect 1155 -1195 1160 -1165
rect 1120 -1360 1160 -1195
rect 1200 -1005 1240 -880
rect 1200 -1035 1205 -1005
rect 1235 -1035 1240 -1005
rect 1200 -1165 1240 -1035
rect 1200 -1195 1205 -1165
rect 1235 -1195 1240 -1165
rect 1200 -1200 1240 -1195
rect 1280 -1005 1320 -880
rect 1280 -1035 1285 -1005
rect 1315 -1035 1320 -1005
rect 1280 -1165 1320 -1035
rect 1280 -1195 1285 -1165
rect 1315 -1195 1320 -1165
rect 1200 -1349 1240 -1280
rect -80 -1440 -40 -1431
rect 1200 -1431 1204 -1349
rect 1236 -1431 1240 -1349
rect 1280 -1360 1320 -1195
rect 1360 -1005 1400 -880
rect 1360 -1035 1365 -1005
rect 1395 -1035 1400 -1005
rect 1360 -1165 1400 -1035
rect 1360 -1195 1365 -1165
rect 1395 -1195 1400 -1165
rect 1360 -1360 1400 -1195
rect 1440 -1005 1480 -880
rect 1440 -1035 1445 -1005
rect 1475 -1035 1480 -1005
rect 1440 -1165 1480 -1035
rect 1440 -1195 1445 -1165
rect 1475 -1195 1480 -1165
rect 1440 -1360 1480 -1195
rect 1520 -1005 1560 -880
rect 1520 -1035 1525 -1005
rect 1555 -1035 1560 -1005
rect 1520 -1165 1560 -1035
rect 1520 -1195 1525 -1165
rect 1555 -1195 1560 -1165
rect 1520 -1360 1560 -1195
rect 1600 -1005 1640 -880
rect 1600 -1035 1605 -1005
rect 1635 -1035 1640 -1005
rect 1600 -1165 1640 -1035
rect 1600 -1195 1605 -1165
rect 1635 -1195 1640 -1165
rect 1600 -1360 1640 -1195
rect 1680 -1005 1720 -880
rect 1680 -1035 1685 -1005
rect 1715 -1035 1720 -1005
rect 1680 -1165 1720 -1035
rect 1680 -1195 1685 -1165
rect 1715 -1195 1720 -1165
rect 1680 -1360 1720 -1195
rect 1760 -1005 1800 -880
rect 1760 -1035 1765 -1005
rect 1795 -1035 1800 -1005
rect 1760 -1165 1800 -1035
rect 1760 -1195 1765 -1165
rect 1795 -1195 1800 -1165
rect 1760 -1360 1800 -1195
rect 1840 -1005 1880 -880
rect 1840 -1035 1845 -1005
rect 1875 -1035 1880 -1005
rect 1840 -1165 1880 -1035
rect 1840 -1195 1845 -1165
rect 1875 -1195 1880 -1165
rect 1840 -1200 1880 -1195
rect 1920 -1005 1960 -880
rect 1920 -1035 1925 -1005
rect 1955 -1035 1960 -1005
rect 1920 -1165 1960 -1035
rect 1920 -1195 1925 -1165
rect 1955 -1195 1960 -1165
rect 1920 -1360 1960 -1195
rect 2000 -1005 2040 -880
rect 2000 -1035 2005 -1005
rect 2035 -1035 2040 -1005
rect 2000 -1165 2040 -1035
rect 2000 -1195 2005 -1165
rect 2035 -1195 2040 -1165
rect 2000 -1360 2040 -1195
rect 2080 -1005 2120 -880
rect 2080 -1035 2085 -1005
rect 2115 -1035 2120 -1005
rect 2080 -1165 2120 -1035
rect 2080 -1195 2085 -1165
rect 2115 -1195 2120 -1165
rect 2080 -1360 2120 -1195
rect 2160 -1005 2200 -880
rect 2160 -1035 2165 -1005
rect 2195 -1035 2200 -1005
rect 2160 -1165 2200 -1035
rect 2160 -1195 2165 -1165
rect 2195 -1195 2200 -1165
rect 2160 -1360 2200 -1195
rect 2240 -1005 2280 -880
rect 2240 -1035 2245 -1005
rect 2275 -1035 2280 -1005
rect 2240 -1165 2280 -1035
rect 2240 -1195 2245 -1165
rect 2275 -1195 2280 -1165
rect 2240 -1360 2280 -1195
rect 2320 -1005 2360 -880
rect 2320 -1035 2325 -1005
rect 2355 -1035 2360 -1005
rect 2320 -1165 2360 -1035
rect 2320 -1195 2325 -1165
rect 2355 -1195 2360 -1165
rect 2320 -1360 2360 -1195
rect 2400 -1005 2440 -880
rect 2400 -1035 2405 -1005
rect 2435 -1035 2440 -1005
rect 2400 -1165 2440 -1035
rect 2400 -1195 2405 -1165
rect 2435 -1195 2440 -1165
rect 2400 -1360 2440 -1195
rect 2480 -1005 2520 -880
rect 2480 -1035 2485 -1005
rect 2515 -1035 2520 -1005
rect 2480 -1165 2520 -1035
rect 2480 -1195 2485 -1165
rect 2515 -1195 2520 -1165
rect 2480 -1200 2520 -1195
rect 2560 -1005 2600 -880
rect 2560 -1035 2565 -1005
rect 2595 -1035 2600 -1005
rect 2560 -1165 2600 -1035
rect 2560 -1195 2565 -1165
rect 2595 -1195 2600 -1165
rect 2480 -1349 2520 -1280
rect 1200 -1440 1240 -1431
rect 2480 -1431 2484 -1349
rect 2516 -1431 2520 -1349
rect 2560 -1360 2600 -1195
rect 2640 -1005 2680 -880
rect 2640 -1035 2645 -1005
rect 2675 -1035 2680 -1005
rect 2640 -1165 2680 -1035
rect 2640 -1195 2645 -1165
rect 2675 -1195 2680 -1165
rect 2640 -1360 2680 -1195
rect 2720 -1005 2760 -880
rect 2720 -1035 2725 -1005
rect 2755 -1035 2760 -1005
rect 2720 -1165 2760 -1035
rect 2720 -1195 2725 -1165
rect 2755 -1195 2760 -1165
rect 2720 -1360 2760 -1195
rect 2800 -1005 2840 -880
rect 2800 -1035 2805 -1005
rect 2835 -1035 2840 -1005
rect 2800 -1165 2840 -1035
rect 2800 -1195 2805 -1165
rect 2835 -1195 2840 -1165
rect 2800 -1360 2840 -1195
rect 2880 -1005 2920 -880
rect 2880 -1035 2885 -1005
rect 2915 -1035 2920 -1005
rect 2880 -1165 2920 -1035
rect 2880 -1195 2885 -1165
rect 2915 -1195 2920 -1165
rect 2880 -1360 2920 -1195
rect 2960 -1005 3000 -880
rect 2960 -1035 2965 -1005
rect 2995 -1035 3000 -1005
rect 2960 -1165 3000 -1035
rect 2960 -1195 2965 -1165
rect 2995 -1195 3000 -1165
rect 2960 -1360 3000 -1195
rect 3040 -1005 3080 -880
rect 3040 -1035 3045 -1005
rect 3075 -1035 3080 -1005
rect 3040 -1165 3080 -1035
rect 3040 -1195 3045 -1165
rect 3075 -1195 3080 -1165
rect 3040 -1360 3080 -1195
rect 3120 -1005 3160 -880
rect 3120 -1035 3125 -1005
rect 3155 -1035 3160 -1005
rect 3120 -1165 3160 -1035
rect 3120 -1195 3125 -1165
rect 3155 -1195 3160 -1165
rect 3120 -1200 3160 -1195
rect 3200 -1005 3240 -880
rect 3200 -1035 3205 -1005
rect 3235 -1035 3240 -1005
rect 3200 -1165 3240 -1035
rect 3200 -1195 3205 -1165
rect 3235 -1195 3240 -1165
rect 3200 -1360 3240 -1195
rect 3280 -1005 3320 -880
rect 3280 -1035 3285 -1005
rect 3315 -1035 3320 -1005
rect 3280 -1165 3320 -1035
rect 3280 -1195 3285 -1165
rect 3315 -1195 3320 -1165
rect 3280 -1360 3320 -1195
rect 3360 -1005 3400 -880
rect 3360 -1035 3365 -1005
rect 3395 -1035 3400 -1005
rect 3360 -1165 3400 -1035
rect 3360 -1195 3365 -1165
rect 3395 -1195 3400 -1165
rect 3360 -1360 3400 -1195
rect 3440 -1005 3480 -880
rect 3440 -1035 3445 -1005
rect 3475 -1035 3480 -1005
rect 3440 -1165 3480 -1035
rect 3440 -1195 3445 -1165
rect 3475 -1195 3480 -1165
rect 3440 -1360 3480 -1195
rect 3520 -1005 3560 -880
rect 3520 -1035 3525 -1005
rect 3555 -1035 3560 -1005
rect 3520 -1165 3560 -1035
rect 3520 -1195 3525 -1165
rect 3555 -1195 3560 -1165
rect 3520 -1360 3560 -1195
rect 3600 -1005 3640 -880
rect 3600 -1035 3605 -1005
rect 3635 -1035 3640 -1005
rect 3600 -1165 3640 -1035
rect 3600 -1195 3605 -1165
rect 3635 -1195 3640 -1165
rect 3600 -1360 3640 -1195
rect 3680 -1005 3720 -880
rect 3680 -1035 3685 -1005
rect 3715 -1035 3720 -1005
rect 3680 -1165 3720 -1035
rect 3680 -1195 3685 -1165
rect 3715 -1195 3720 -1165
rect 3680 -1360 3720 -1195
rect 3760 -1005 3800 -880
rect 3760 -1035 3765 -1005
rect 3795 -1035 3800 -1005
rect 3760 -1165 3800 -1035
rect 3760 -1195 3765 -1165
rect 3795 -1195 3800 -1165
rect 3760 -1200 3800 -1195
rect 3840 -1005 3880 -880
rect 3840 -1035 3845 -1005
rect 3875 -1035 3880 -1005
rect 3840 -1165 3880 -1035
rect 3840 -1195 3845 -1165
rect 3875 -1195 3880 -1165
rect 3760 -1349 3800 -1280
rect 2480 -1440 2520 -1431
rect 3760 -1431 3764 -1349
rect 3796 -1431 3800 -1349
rect 3840 -1360 3880 -1195
rect 3920 -1005 3960 -880
rect 3920 -1035 3925 -1005
rect 3955 -1035 3960 -1005
rect 3920 -1165 3960 -1035
rect 3920 -1195 3925 -1165
rect 3955 -1195 3960 -1165
rect 3920 -1360 3960 -1195
rect 4000 -1005 4040 -880
rect 4000 -1035 4005 -1005
rect 4035 -1035 4040 -1005
rect 4000 -1165 4040 -1035
rect 4000 -1195 4005 -1165
rect 4035 -1195 4040 -1165
rect 4000 -1360 4040 -1195
rect 4080 -1005 4120 -880
rect 4080 -1035 4085 -1005
rect 4115 -1035 4120 -1005
rect 4080 -1165 4120 -1035
rect 4080 -1195 4085 -1165
rect 4115 -1195 4120 -1165
rect 4080 -1360 4120 -1195
rect 4160 -1005 4200 -880
rect 4160 -1035 4165 -1005
rect 4195 -1035 4200 -1005
rect 4160 -1165 4200 -1035
rect 4160 -1195 4165 -1165
rect 4195 -1195 4200 -1165
rect 4160 -1360 4200 -1195
rect 4240 -1005 4280 -880
rect 4240 -1035 4245 -1005
rect 4275 -1035 4280 -1005
rect 4240 -1165 4280 -1035
rect 4240 -1195 4245 -1165
rect 4275 -1195 4280 -1165
rect 4240 -1360 4280 -1195
rect 4320 -1005 4360 -880
rect 4320 -1035 4325 -1005
rect 4355 -1035 4360 -1005
rect 4320 -1165 4360 -1035
rect 4320 -1195 4325 -1165
rect 4355 -1195 4360 -1165
rect 4320 -1360 4360 -1195
rect 4400 -1005 4440 -880
rect 4400 -1035 4405 -1005
rect 4435 -1035 4440 -1005
rect 4400 -1165 4440 -1035
rect 4400 -1195 4405 -1165
rect 4435 -1195 4440 -1165
rect 4400 -1200 4440 -1195
rect 4480 -1005 4520 -880
rect 4480 -1035 4485 -1005
rect 4515 -1035 4520 -1005
rect 4480 -1165 4520 -1035
rect 4480 -1195 4485 -1165
rect 4515 -1195 4520 -1165
rect 4480 -1360 4520 -1195
rect 4560 -1005 4600 -880
rect 4560 -1035 4565 -1005
rect 4595 -1035 4600 -1005
rect 4560 -1165 4600 -1035
rect 4560 -1195 4565 -1165
rect 4595 -1195 4600 -1165
rect 4560 -1360 4600 -1195
rect 4640 -1005 4680 -880
rect 4640 -1035 4645 -1005
rect 4675 -1035 4680 -1005
rect 4640 -1165 4680 -1035
rect 4640 -1195 4645 -1165
rect 4675 -1195 4680 -1165
rect 4640 -1360 4680 -1195
rect 4720 -1005 4760 -880
rect 4720 -1035 4725 -1005
rect 4755 -1035 4760 -1005
rect 4720 -1165 4760 -1035
rect 4720 -1195 4725 -1165
rect 4755 -1195 4760 -1165
rect 4720 -1360 4760 -1195
rect 4800 -1005 4840 -880
rect 4800 -1035 4805 -1005
rect 4835 -1035 4840 -1005
rect 4800 -1165 4840 -1035
rect 4800 -1195 4805 -1165
rect 4835 -1195 4840 -1165
rect 4800 -1360 4840 -1195
rect 4880 -1005 4920 -880
rect 4880 -1035 4885 -1005
rect 4915 -1035 4920 -1005
rect 4880 -1165 4920 -1035
rect 4880 -1195 4885 -1165
rect 4915 -1195 4920 -1165
rect 4880 -1360 4920 -1195
rect 4960 -1005 5000 -880
rect 4960 -1035 4965 -1005
rect 4995 -1035 5000 -1005
rect 4960 -1165 5000 -1035
rect 4960 -1195 4965 -1165
rect 4995 -1195 5000 -1165
rect 4960 -1360 5000 -1195
rect 5040 -1005 5080 -880
rect 5040 -1035 5045 -1005
rect 5075 -1035 5080 -1005
rect 5040 -1165 5080 -1035
rect 5040 -1195 5045 -1165
rect 5075 -1195 5080 -1165
rect 5040 -1349 5080 -1195
rect 3760 -1440 3800 -1431
rect 5040 -1431 5044 -1349
rect 5076 -1431 5080 -1349
rect 5120 -1005 5160 -880
rect 5120 -1035 5125 -1005
rect 5155 -1035 5160 -1005
rect 5120 -1165 5160 -1035
rect 5120 -1195 5125 -1165
rect 5155 -1195 5160 -1165
rect 5120 -1360 5160 -1195
rect 5200 -685 5240 -680
rect 5200 -715 5205 -685
rect 5235 -715 5240 -685
rect 5200 -845 5240 -715
rect 5200 -875 5205 -845
rect 5235 -875 5240 -845
rect 5200 -1005 5240 -875
rect 5200 -1035 5205 -1005
rect 5235 -1035 5240 -1005
rect 5200 -1165 5240 -1035
rect 5200 -1195 5205 -1165
rect 5235 -1195 5240 -1165
rect 5200 -1360 5240 -1195
rect 5040 -1440 5080 -1431
<< via3 >>
rect -76 630 -44 631
rect -76 450 -75 630
rect -75 450 -45 630
rect -45 450 -44 630
rect -76 449 -44 450
rect 1204 630 1236 631
rect 1204 450 1205 630
rect 1205 450 1235 630
rect 1235 450 1236 630
rect 1204 449 1236 450
rect 2484 630 2516 631
rect 2484 450 2485 630
rect 2485 450 2515 630
rect 2515 450 2516 630
rect 2484 449 2516 450
rect 3764 630 3796 631
rect 3764 450 3765 630
rect 3765 450 3795 630
rect 3795 450 3796 630
rect 3764 449 3796 450
rect 5044 630 5076 631
rect 5044 450 5045 630
rect 5045 450 5075 630
rect 5075 450 5076 630
rect 5044 449 5076 450
rect -76 -1360 -44 -1349
rect -76 -1430 -75 -1360
rect -75 -1430 -45 -1360
rect -45 -1430 -44 -1360
rect -76 -1431 -44 -1430
rect 1204 -1360 1236 -1349
rect 1204 -1430 1205 -1360
rect 1205 -1430 1235 -1360
rect 1235 -1430 1236 -1360
rect 1204 -1431 1236 -1430
rect 2484 -1360 2516 -1349
rect 2484 -1430 2485 -1360
rect 2485 -1430 2515 -1360
rect 2515 -1430 2516 -1360
rect 2484 -1431 2516 -1430
rect 3764 -1360 3796 -1349
rect 3764 -1430 3765 -1360
rect 3765 -1430 3795 -1360
rect 3795 -1430 3796 -1360
rect 3764 -1431 3796 -1430
rect 5044 -1360 5076 -1349
rect 5044 -1430 5045 -1360
rect 5045 -1430 5075 -1360
rect 5075 -1430 5076 -1360
rect 5044 -1431 5076 -1430
<< metal4 >>
rect -240 631 5080 640
rect -240 600 -76 631
rect -44 600 1204 631
rect 1236 600 2484 631
rect 2516 600 3764 631
rect 3796 600 5044 631
rect 5076 600 5080 631
rect -240 480 -120 600
rect 0 480 1160 600
rect 1280 480 2440 600
rect 2560 480 3720 600
rect 3840 480 5000 600
rect -240 449 -76 480
rect -44 449 1204 480
rect 1236 449 2484 480
rect 2516 449 3764 480
rect 3796 449 5044 480
rect 5076 449 5080 480
rect -240 440 5080 449
rect 5120 440 5240 640
rect -240 -1349 5240 -1320
rect -240 -1431 -76 -1349
rect -44 -1360 1204 -1349
rect -44 -1431 520 -1360
rect -240 -1480 520 -1431
rect 640 -1431 1204 -1360
rect 1236 -1360 2484 -1349
rect 1236 -1431 1800 -1360
rect 640 -1480 1800 -1431
rect 1920 -1431 2484 -1360
rect 2516 -1360 3764 -1349
rect 2516 -1431 3080 -1360
rect 1920 -1480 3080 -1431
rect 3200 -1431 3764 -1360
rect 3796 -1360 5044 -1349
rect 3796 -1431 4360 -1360
rect 3200 -1480 4360 -1431
rect 4480 -1431 5044 -1360
rect 5076 -1431 5240 -1349
rect 4480 -1480 5240 -1431
rect -240 -1520 5240 -1480
<< via4 >>
rect -120 480 -76 600
rect -76 480 -44 600
rect -44 480 0 600
rect 1160 480 1204 600
rect 1204 480 1236 600
rect 1236 480 1280 600
rect 2440 480 2484 600
rect 2484 480 2516 600
rect 2516 480 2560 600
rect 3720 480 3764 600
rect 3764 480 3796 600
rect 3796 480 3840 600
rect 5000 480 5044 600
rect 5044 480 5076 600
rect 5076 480 5120 600
rect 520 -1480 640 -1360
rect 1800 -1480 1920 -1360
rect 3080 -1480 3200 -1360
rect 4360 -1480 4480 -1360
<< metal5 >>
rect -160 600 40 840
rect -160 480 -120 600
rect 0 480 40 600
rect -160 -1520 40 480
rect 480 -1360 680 840
rect 480 -1480 520 -1360
rect 640 -1480 680 -1360
rect 480 -1520 680 -1480
rect 1120 600 1320 840
rect 1120 480 1160 600
rect 1280 480 1320 600
rect 1120 -1520 1320 480
rect 1760 -1360 1960 840
rect 1760 -1480 1800 -1360
rect 1920 -1480 1960 -1360
rect 1760 -1520 1960 -1480
rect 2400 600 2600 840
rect 2400 480 2440 600
rect 2560 480 2600 600
rect 2400 -1520 2600 480
rect 3040 -1360 3240 840
rect 3040 -1480 3080 -1360
rect 3200 -1480 3240 -1360
rect 3040 -1520 3240 -1480
rect 3680 600 3880 840
rect 3680 480 3720 600
rect 3840 480 3880 600
rect 3680 -1520 3880 480
rect 4320 -1360 4520 840
rect 4320 -1480 4360 -1360
rect 4480 -1480 4520 -1360
rect 4320 -1520 4520 -1480
rect 4960 600 5160 840
rect 4960 480 5000 600
rect 5120 480 5160 600
rect 4960 -1520 5160 480
<< labels >>
rlabel locali 2480 -1320 2520 -1280 0 xn
rlabel metal2 5200 -800 5240 -760 0 gpb
port 2 nsew
rlabel metal2 5200 -1120 5240 -1080 0 gna
port 3 nsew
rlabel metal1 240 -1440 280 -1340 0 n1
rlabel metal1 880 -1440 920 -1340 0 n2
rlabel metal1 1520 -1440 1560 -1340 0 n3
rlabel metal1 2160 -1440 2200 -1340 0 n4
rlabel metal1 2800 -1440 2840 -1340 0 n5
rlabel metal1 3440 -1440 3480 -1340 0 n6
rlabel metal1 4080 -1440 4120 -1340 0 n7
rlabel metal1 4720 -1440 4760 -1340 0 n8
rlabel locali 80 720 120 760 0 vdda
rlabel locali 2480 320 2520 360 0 xp
rlabel metal2 5200 -80 5240 -40 0 gpa
port 1 nsew
rlabel metal5 -160 800 40 840 0 vdda
port 4 nsew
rlabel metal5 480 800 680 840 0 vssa
port 5 nsew
rlabel metal1 240 380 280 680 0 p1
rlabel metal1 880 380 920 680 0 p2
rlabel metal1 1520 380 1560 680 0 p3
rlabel metal1 2160 380 2200 680 0 p4
rlabel metal1 2800 380 2840 680 0 p5
rlabel metal1 3440 380 3480 680 0 p6
rlabel metal1 4080 380 4120 680 0 p7
rlabel metal1 4720 380 4760 680 0 p8
<< end >>
