* symmetrical single-ended OTA ac testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "../mag/ota.spice"

* supply voltages
vdda vdda 0 1.8
vssa vssa 0 0.0
egnda gnda vssa vdda vssa 0.5

* input signals
vin in gnda dc 0 ac 1 SINE(0 0.4 0.5k 0 0 0)
IB ib vss 5n

* DUT
Xdut gnda in out ib vdda gnda vssa ota
CL out gnda 1p
LL out gnda 1T

.save v(in) v(out) v(ib) i(vdda)
.option gmin=1e-15
*.option rseries = 1.0e-4
.option rshunt = 1.0e9
.control

	op
	print ib i(vdda)

	ac dec 10 1m 1Meg
	plot vdb(out)
	
	noise v(out) vin dec 100 1 100
	print inoise_total onoise_total
    
.endc

.end
