magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< error_p >>
rect 8 3920 8392 3992
rect 8 3840 80 3920
rect 94 3880 8306 3906
rect 94 2760 120 3880
rect 160 3814 8240 3840
rect 160 2872 232 3814
rect 8214 2872 8240 3814
rect 160 2800 8240 2872
rect 8280 2760 8306 3880
rect 8320 2800 8392 3920
rect 94 2734 8306 2760
rect 8 2480 8392 2552
rect 8 2400 80 2480
rect 94 2440 8306 2466
rect 94 1320 120 2440
rect 160 2374 8240 2400
rect 160 1432 232 2374
rect 8214 1432 8240 2374
rect 160 1360 8240 1432
rect 8280 1320 8306 2440
rect 8320 1360 8392 2480
rect 94 1294 8306 1320
<< nwell >>
rect 120 2760 8280 3880
rect 120 1320 8280 2440
<< pwell >>
rect -26 3894 8426 4026
rect -26 2746 106 3894
rect 8294 2746 8426 3894
rect -26 2454 8426 2746
rect -26 1306 106 2454
rect 8294 1306 8426 2454
rect -26 1174 8426 1306
rect -26 534 8426 666
rect -26 106 106 534
rect 294 106 8106 534
rect 8294 106 8426 534
rect -26 -26 8426 106
<< mvnmos >>
rect 520 160 2120 360
rect 2440 160 4040 360
rect 4360 160 5960 360
rect 6280 160 7880 360
<< mvpmos >>
rect 520 3080 2120 3680
rect 2440 3080 4040 3680
rect 4360 3080 5960 3680
rect 6280 3080 7880 3680
rect 520 1640 2120 2240
rect 2440 1640 4040 2240
rect 4360 1640 5960 2240
rect 6280 1640 7880 2240
<< mvndiff >>
rect 320 311 520 360
rect 320 277 343 311
rect 377 277 520 311
rect 320 243 520 277
rect 320 209 343 243
rect 377 209 520 243
rect 320 160 520 209
rect 2120 311 2440 360
rect 2120 277 2263 311
rect 2297 277 2440 311
rect 2120 243 2440 277
rect 2120 209 2263 243
rect 2297 209 2440 243
rect 2120 160 2440 209
rect 4040 311 4360 360
rect 4040 277 4183 311
rect 4217 277 4360 311
rect 4040 243 4360 277
rect 4040 209 4183 243
rect 4217 209 4360 243
rect 4040 160 4360 209
rect 5960 311 6280 360
rect 5960 277 6103 311
rect 6137 277 6280 311
rect 5960 243 6280 277
rect 5960 209 6103 243
rect 6137 209 6280 243
rect 5960 160 6280 209
rect 7880 311 8080 360
rect 7880 277 8023 311
rect 8057 277 8080 311
rect 7880 243 8080 277
rect 7880 209 8023 243
rect 8057 209 8080 243
rect 7880 160 8080 209
<< mvpdiff >>
rect 320 3635 520 3680
rect 320 3601 343 3635
rect 377 3601 520 3635
rect 320 3567 520 3601
rect 320 3533 343 3567
rect 377 3533 520 3567
rect 320 3499 520 3533
rect 320 3465 343 3499
rect 377 3465 520 3499
rect 320 3431 520 3465
rect 320 3397 343 3431
rect 377 3397 520 3431
rect 320 3363 520 3397
rect 320 3329 343 3363
rect 377 3329 520 3363
rect 320 3295 520 3329
rect 320 3261 343 3295
rect 377 3261 520 3295
rect 320 3227 520 3261
rect 320 3193 343 3227
rect 377 3193 520 3227
rect 320 3159 520 3193
rect 320 3125 343 3159
rect 377 3125 520 3159
rect 320 3080 520 3125
rect 2120 3635 2440 3680
rect 2120 3601 2263 3635
rect 2297 3601 2440 3635
rect 2120 3567 2440 3601
rect 2120 3533 2263 3567
rect 2297 3533 2440 3567
rect 2120 3499 2440 3533
rect 2120 3465 2263 3499
rect 2297 3465 2440 3499
rect 2120 3431 2440 3465
rect 2120 3397 2263 3431
rect 2297 3397 2440 3431
rect 2120 3363 2440 3397
rect 2120 3329 2263 3363
rect 2297 3329 2440 3363
rect 2120 3295 2440 3329
rect 2120 3261 2263 3295
rect 2297 3261 2440 3295
rect 2120 3227 2440 3261
rect 2120 3193 2263 3227
rect 2297 3193 2440 3227
rect 2120 3159 2440 3193
rect 2120 3125 2263 3159
rect 2297 3125 2440 3159
rect 2120 3080 2440 3125
rect 4040 3635 4360 3680
rect 4040 3601 4183 3635
rect 4217 3601 4360 3635
rect 4040 3567 4360 3601
rect 4040 3533 4183 3567
rect 4217 3533 4360 3567
rect 4040 3499 4360 3533
rect 4040 3465 4183 3499
rect 4217 3465 4360 3499
rect 4040 3431 4360 3465
rect 4040 3397 4183 3431
rect 4217 3397 4360 3431
rect 4040 3363 4360 3397
rect 4040 3329 4183 3363
rect 4217 3329 4360 3363
rect 4040 3295 4360 3329
rect 4040 3261 4183 3295
rect 4217 3261 4360 3295
rect 4040 3227 4360 3261
rect 4040 3193 4183 3227
rect 4217 3193 4360 3227
rect 4040 3159 4360 3193
rect 4040 3125 4183 3159
rect 4217 3125 4360 3159
rect 4040 3080 4360 3125
rect 5960 3635 6280 3680
rect 5960 3601 6103 3635
rect 6137 3601 6280 3635
rect 5960 3567 6280 3601
rect 5960 3533 6103 3567
rect 6137 3533 6280 3567
rect 5960 3499 6280 3533
rect 5960 3465 6103 3499
rect 6137 3465 6280 3499
rect 5960 3431 6280 3465
rect 5960 3397 6103 3431
rect 6137 3397 6280 3431
rect 5960 3363 6280 3397
rect 5960 3329 6103 3363
rect 6137 3329 6280 3363
rect 5960 3295 6280 3329
rect 5960 3261 6103 3295
rect 6137 3261 6280 3295
rect 5960 3227 6280 3261
rect 5960 3193 6103 3227
rect 6137 3193 6280 3227
rect 5960 3159 6280 3193
rect 5960 3125 6103 3159
rect 6137 3125 6280 3159
rect 5960 3080 6280 3125
rect 7880 3635 8080 3680
rect 7880 3601 8023 3635
rect 8057 3601 8080 3635
rect 7880 3567 8080 3601
rect 7880 3533 8023 3567
rect 8057 3533 8080 3567
rect 7880 3499 8080 3533
rect 7880 3465 8023 3499
rect 8057 3465 8080 3499
rect 7880 3431 8080 3465
rect 7880 3397 8023 3431
rect 8057 3397 8080 3431
rect 7880 3363 8080 3397
rect 7880 3329 8023 3363
rect 8057 3329 8080 3363
rect 7880 3295 8080 3329
rect 7880 3261 8023 3295
rect 8057 3261 8080 3295
rect 7880 3227 8080 3261
rect 7880 3193 8023 3227
rect 8057 3193 8080 3227
rect 7880 3159 8080 3193
rect 7880 3125 8023 3159
rect 8057 3125 8080 3159
rect 7880 3080 8080 3125
rect 320 2195 520 2240
rect 320 2161 343 2195
rect 377 2161 520 2195
rect 320 2127 520 2161
rect 320 2093 343 2127
rect 377 2093 520 2127
rect 320 2059 520 2093
rect 320 2025 343 2059
rect 377 2025 520 2059
rect 320 1991 520 2025
rect 320 1957 343 1991
rect 377 1957 520 1991
rect 320 1923 520 1957
rect 320 1889 343 1923
rect 377 1889 520 1923
rect 320 1855 520 1889
rect 320 1821 343 1855
rect 377 1821 520 1855
rect 320 1787 520 1821
rect 320 1753 343 1787
rect 377 1753 520 1787
rect 320 1719 520 1753
rect 320 1685 343 1719
rect 377 1685 520 1719
rect 320 1640 520 1685
rect 2120 2195 2440 2240
rect 2120 2161 2263 2195
rect 2297 2161 2440 2195
rect 2120 2127 2440 2161
rect 2120 2093 2263 2127
rect 2297 2093 2440 2127
rect 2120 2059 2440 2093
rect 2120 2025 2263 2059
rect 2297 2025 2440 2059
rect 2120 1991 2440 2025
rect 2120 1957 2263 1991
rect 2297 1957 2440 1991
rect 2120 1923 2440 1957
rect 2120 1889 2263 1923
rect 2297 1889 2440 1923
rect 2120 1855 2440 1889
rect 2120 1821 2263 1855
rect 2297 1821 2440 1855
rect 2120 1787 2440 1821
rect 2120 1753 2263 1787
rect 2297 1753 2440 1787
rect 2120 1719 2440 1753
rect 2120 1685 2263 1719
rect 2297 1685 2440 1719
rect 2120 1640 2440 1685
rect 4040 2195 4360 2240
rect 4040 2161 4183 2195
rect 4217 2161 4360 2195
rect 4040 2127 4360 2161
rect 4040 2093 4183 2127
rect 4217 2093 4360 2127
rect 4040 2059 4360 2093
rect 4040 2025 4183 2059
rect 4217 2025 4360 2059
rect 4040 1991 4360 2025
rect 4040 1957 4183 1991
rect 4217 1957 4360 1991
rect 4040 1923 4360 1957
rect 4040 1889 4183 1923
rect 4217 1889 4360 1923
rect 4040 1855 4360 1889
rect 4040 1821 4183 1855
rect 4217 1821 4360 1855
rect 4040 1787 4360 1821
rect 4040 1753 4183 1787
rect 4217 1753 4360 1787
rect 4040 1719 4360 1753
rect 4040 1685 4183 1719
rect 4217 1685 4360 1719
rect 4040 1640 4360 1685
rect 5960 2195 6280 2240
rect 5960 2161 6103 2195
rect 6137 2161 6280 2195
rect 5960 2127 6280 2161
rect 5960 2093 6103 2127
rect 6137 2093 6280 2127
rect 5960 2059 6280 2093
rect 5960 2025 6103 2059
rect 6137 2025 6280 2059
rect 5960 1991 6280 2025
rect 5960 1957 6103 1991
rect 6137 1957 6280 1991
rect 5960 1923 6280 1957
rect 5960 1889 6103 1923
rect 6137 1889 6280 1923
rect 5960 1855 6280 1889
rect 5960 1821 6103 1855
rect 6137 1821 6280 1855
rect 5960 1787 6280 1821
rect 5960 1753 6103 1787
rect 6137 1753 6280 1787
rect 5960 1719 6280 1753
rect 5960 1685 6103 1719
rect 6137 1685 6280 1719
rect 5960 1640 6280 1685
rect 7880 2195 8080 2240
rect 7880 2161 8023 2195
rect 8057 2161 8080 2195
rect 7880 2127 8080 2161
rect 7880 2093 8023 2127
rect 8057 2093 8080 2127
rect 7880 2059 8080 2093
rect 7880 2025 8023 2059
rect 8057 2025 8080 2059
rect 7880 1991 8080 2025
rect 7880 1957 8023 1991
rect 8057 1957 8080 1991
rect 7880 1923 8080 1957
rect 7880 1889 8023 1923
rect 8057 1889 8080 1923
rect 7880 1855 8080 1889
rect 7880 1821 8023 1855
rect 8057 1821 8080 1855
rect 7880 1787 8080 1821
rect 7880 1753 8023 1787
rect 8057 1753 8080 1787
rect 7880 1719 8080 1753
rect 7880 1685 8023 1719
rect 8057 1685 8080 1719
rect 7880 1640 8080 1685
<< mvndiffc >>
rect 343 277 377 311
rect 343 209 377 243
rect 2263 277 2297 311
rect 2263 209 2297 243
rect 4183 277 4217 311
rect 4183 209 4217 243
rect 6103 277 6137 311
rect 6103 209 6137 243
rect 8023 277 8057 311
rect 8023 209 8057 243
<< mvpdiffc >>
rect 343 3601 377 3635
rect 343 3533 377 3567
rect 343 3465 377 3499
rect 343 3397 377 3431
rect 343 3329 377 3363
rect 343 3261 377 3295
rect 343 3193 377 3227
rect 343 3125 377 3159
rect 2263 3601 2297 3635
rect 2263 3533 2297 3567
rect 2263 3465 2297 3499
rect 2263 3397 2297 3431
rect 2263 3329 2297 3363
rect 2263 3261 2297 3295
rect 2263 3193 2297 3227
rect 2263 3125 2297 3159
rect 4183 3601 4217 3635
rect 4183 3533 4217 3567
rect 4183 3465 4217 3499
rect 4183 3397 4217 3431
rect 4183 3329 4217 3363
rect 4183 3261 4217 3295
rect 4183 3193 4217 3227
rect 4183 3125 4217 3159
rect 6103 3601 6137 3635
rect 6103 3533 6137 3567
rect 6103 3465 6137 3499
rect 6103 3397 6137 3431
rect 6103 3329 6137 3363
rect 6103 3261 6137 3295
rect 6103 3193 6137 3227
rect 6103 3125 6137 3159
rect 8023 3601 8057 3635
rect 8023 3533 8057 3567
rect 8023 3465 8057 3499
rect 8023 3397 8057 3431
rect 8023 3329 8057 3363
rect 8023 3261 8057 3295
rect 8023 3193 8057 3227
rect 8023 3125 8057 3159
rect 343 2161 377 2195
rect 343 2093 377 2127
rect 343 2025 377 2059
rect 343 1957 377 1991
rect 343 1889 377 1923
rect 343 1821 377 1855
rect 343 1753 377 1787
rect 343 1685 377 1719
rect 2263 2161 2297 2195
rect 2263 2093 2297 2127
rect 2263 2025 2297 2059
rect 2263 1957 2297 1991
rect 2263 1889 2297 1923
rect 2263 1821 2297 1855
rect 2263 1753 2297 1787
rect 2263 1685 2297 1719
rect 4183 2161 4217 2195
rect 4183 2093 4217 2127
rect 4183 2025 4217 2059
rect 4183 1957 4217 1991
rect 4183 1889 4217 1923
rect 4183 1821 4217 1855
rect 4183 1753 4217 1787
rect 4183 1685 4217 1719
rect 6103 2161 6137 2195
rect 6103 2093 6137 2127
rect 6103 2025 6137 2059
rect 6103 1957 6137 1991
rect 6103 1889 6137 1923
rect 6103 1821 6137 1855
rect 6103 1753 6137 1787
rect 6103 1685 6137 1719
rect 8023 2161 8057 2195
rect 8023 2093 8057 2127
rect 8023 2025 8057 2059
rect 8023 1957 8057 1991
rect 8023 1889 8057 1923
rect 8023 1821 8057 1855
rect 8023 1753 8057 1787
rect 8023 1685 8057 1719
<< psubdiff >>
rect 0 3977 8400 4000
rect 0 3943 137 3977
rect 171 3943 205 3977
rect 239 3943 273 3977
rect 307 3943 341 3977
rect 375 3943 409 3977
rect 443 3943 477 3977
rect 511 3943 545 3977
rect 579 3943 613 3977
rect 647 3943 681 3977
rect 715 3943 749 3977
rect 783 3943 817 3977
rect 851 3943 885 3977
rect 919 3943 953 3977
rect 987 3943 1021 3977
rect 1055 3943 1089 3977
rect 1123 3943 1157 3977
rect 1191 3943 1225 3977
rect 1259 3943 1293 3977
rect 1327 3943 1361 3977
rect 1395 3943 1429 3977
rect 1463 3943 1497 3977
rect 1531 3943 1565 3977
rect 1599 3943 1633 3977
rect 1667 3943 1701 3977
rect 1735 3943 1769 3977
rect 1803 3943 1837 3977
rect 1871 3943 1905 3977
rect 1939 3943 1973 3977
rect 2007 3943 2041 3977
rect 2075 3943 2109 3977
rect 2143 3943 2177 3977
rect 2211 3943 2245 3977
rect 2279 3943 2313 3977
rect 2347 3943 2381 3977
rect 2415 3943 2449 3977
rect 2483 3943 2517 3977
rect 2551 3943 2585 3977
rect 2619 3943 2653 3977
rect 2687 3943 2721 3977
rect 2755 3943 2789 3977
rect 2823 3943 2857 3977
rect 2891 3943 2925 3977
rect 2959 3943 2993 3977
rect 3027 3943 3061 3977
rect 3095 3943 3129 3977
rect 3163 3943 3197 3977
rect 3231 3943 3265 3977
rect 3299 3943 3333 3977
rect 3367 3943 3401 3977
rect 3435 3943 3469 3977
rect 3503 3943 3537 3977
rect 3571 3943 3605 3977
rect 3639 3943 3673 3977
rect 3707 3943 3741 3977
rect 3775 3943 3809 3977
rect 3843 3943 3877 3977
rect 3911 3943 3945 3977
rect 3979 3943 4013 3977
rect 4047 3943 4081 3977
rect 4115 3943 4149 3977
rect 4183 3943 4217 3977
rect 4251 3943 4285 3977
rect 4319 3943 4353 3977
rect 4387 3943 4421 3977
rect 4455 3943 4489 3977
rect 4523 3943 4557 3977
rect 4591 3943 4625 3977
rect 4659 3943 4693 3977
rect 4727 3943 4761 3977
rect 4795 3943 4829 3977
rect 4863 3943 4897 3977
rect 4931 3943 4965 3977
rect 4999 3943 5033 3977
rect 5067 3943 5101 3977
rect 5135 3943 5169 3977
rect 5203 3943 5237 3977
rect 5271 3943 5305 3977
rect 5339 3943 5373 3977
rect 5407 3943 5441 3977
rect 5475 3943 5509 3977
rect 5543 3943 5577 3977
rect 5611 3943 5645 3977
rect 5679 3943 5713 3977
rect 5747 3943 5781 3977
rect 5815 3943 5849 3977
rect 5883 3943 5917 3977
rect 5951 3943 5985 3977
rect 6019 3943 6053 3977
rect 6087 3943 6121 3977
rect 6155 3943 6189 3977
rect 6223 3943 6257 3977
rect 6291 3943 6325 3977
rect 6359 3943 6393 3977
rect 6427 3943 6461 3977
rect 6495 3943 6529 3977
rect 6563 3943 6597 3977
rect 6631 3943 6665 3977
rect 6699 3943 6733 3977
rect 6767 3943 6801 3977
rect 6835 3943 6869 3977
rect 6903 3943 6937 3977
rect 6971 3943 7005 3977
rect 7039 3943 7073 3977
rect 7107 3943 7141 3977
rect 7175 3943 7209 3977
rect 7243 3943 7277 3977
rect 7311 3943 7345 3977
rect 7379 3943 7413 3977
rect 7447 3943 7481 3977
rect 7515 3943 7549 3977
rect 7583 3943 7617 3977
rect 7651 3943 7685 3977
rect 7719 3943 7753 3977
rect 7787 3943 7821 3977
rect 7855 3943 7889 3977
rect 7923 3943 7957 3977
rect 7991 3943 8025 3977
rect 8059 3943 8093 3977
rect 8127 3943 8161 3977
rect 8195 3943 8229 3977
rect 8263 3943 8400 3977
rect 0 3920 8400 3943
rect 0 3847 80 3920
rect 0 3813 23 3847
rect 57 3813 80 3847
rect 8320 3847 8400 3920
rect 0 3779 80 3813
rect 0 3745 23 3779
rect 57 3745 80 3779
rect 0 3711 80 3745
rect 0 3677 23 3711
rect 57 3677 80 3711
rect 0 3643 80 3677
rect 0 3609 23 3643
rect 57 3609 80 3643
rect 0 3575 80 3609
rect 0 3541 23 3575
rect 57 3541 80 3575
rect 0 3507 80 3541
rect 0 3473 23 3507
rect 57 3473 80 3507
rect 0 3439 80 3473
rect 0 3405 23 3439
rect 57 3405 80 3439
rect 0 3371 80 3405
rect 0 3337 23 3371
rect 57 3337 80 3371
rect 0 3303 80 3337
rect 0 3269 23 3303
rect 57 3269 80 3303
rect 0 3235 80 3269
rect 0 3201 23 3235
rect 57 3201 80 3235
rect 0 3167 80 3201
rect 0 3133 23 3167
rect 57 3133 80 3167
rect 0 3099 80 3133
rect 0 3065 23 3099
rect 57 3065 80 3099
rect 0 3031 80 3065
rect 0 2997 23 3031
rect 57 2997 80 3031
rect 0 2963 80 2997
rect 0 2929 23 2963
rect 57 2929 80 2963
rect 0 2895 80 2929
rect 0 2861 23 2895
rect 57 2861 80 2895
rect 0 2827 80 2861
rect 0 2793 23 2827
rect 57 2793 80 2827
rect 8320 3813 8343 3847
rect 8377 3813 8400 3847
rect 8320 3779 8400 3813
rect 8320 3745 8343 3779
rect 8377 3745 8400 3779
rect 8320 3711 8400 3745
rect 8320 3677 8343 3711
rect 8377 3677 8400 3711
rect 8320 3643 8400 3677
rect 8320 3609 8343 3643
rect 8377 3609 8400 3643
rect 8320 3575 8400 3609
rect 8320 3541 8343 3575
rect 8377 3541 8400 3575
rect 8320 3507 8400 3541
rect 8320 3473 8343 3507
rect 8377 3473 8400 3507
rect 8320 3439 8400 3473
rect 8320 3405 8343 3439
rect 8377 3405 8400 3439
rect 8320 3371 8400 3405
rect 8320 3337 8343 3371
rect 8377 3337 8400 3371
rect 8320 3303 8400 3337
rect 8320 3269 8343 3303
rect 8377 3269 8400 3303
rect 8320 3235 8400 3269
rect 8320 3201 8343 3235
rect 8377 3201 8400 3235
rect 8320 3167 8400 3201
rect 8320 3133 8343 3167
rect 8377 3133 8400 3167
rect 8320 3099 8400 3133
rect 8320 3065 8343 3099
rect 8377 3065 8400 3099
rect 8320 3031 8400 3065
rect 8320 2997 8343 3031
rect 8377 2997 8400 3031
rect 8320 2963 8400 2997
rect 8320 2929 8343 2963
rect 8377 2929 8400 2963
rect 8320 2895 8400 2929
rect 8320 2861 8343 2895
rect 8377 2861 8400 2895
rect 8320 2827 8400 2861
rect 0 2720 80 2793
rect 8320 2793 8343 2827
rect 8377 2793 8400 2827
rect 8320 2720 8400 2793
rect 0 2697 8400 2720
rect 0 2663 151 2697
rect 185 2663 219 2697
rect 253 2663 287 2697
rect 321 2663 355 2697
rect 389 2663 423 2697
rect 457 2663 491 2697
rect 525 2663 559 2697
rect 593 2663 627 2697
rect 661 2663 695 2697
rect 729 2663 763 2697
rect 797 2663 831 2697
rect 865 2663 899 2697
rect 933 2663 967 2697
rect 1001 2663 1035 2697
rect 1069 2663 1103 2697
rect 1137 2663 1171 2697
rect 1205 2663 1239 2697
rect 1273 2663 1307 2697
rect 1341 2663 1375 2697
rect 1409 2663 1443 2697
rect 1477 2663 1511 2697
rect 1545 2663 1579 2697
rect 1613 2663 1647 2697
rect 1681 2663 1715 2697
rect 1749 2663 1783 2697
rect 1817 2663 1851 2697
rect 1885 2663 1919 2697
rect 1953 2663 1987 2697
rect 2021 2663 2055 2697
rect 2089 2663 2123 2697
rect 2157 2663 2191 2697
rect 2225 2663 2259 2697
rect 2293 2663 2327 2697
rect 2361 2663 2395 2697
rect 2429 2663 2463 2697
rect 2497 2663 2531 2697
rect 2565 2663 2599 2697
rect 2633 2663 2667 2697
rect 2701 2663 2735 2697
rect 2769 2663 2803 2697
rect 2837 2663 2871 2697
rect 2905 2663 2939 2697
rect 2973 2663 3007 2697
rect 3041 2663 3075 2697
rect 3109 2663 3143 2697
rect 3177 2663 3211 2697
rect 3245 2663 3279 2697
rect 3313 2663 3347 2697
rect 3381 2663 3415 2697
rect 3449 2663 3483 2697
rect 3517 2663 3551 2697
rect 3585 2663 3619 2697
rect 3653 2663 3687 2697
rect 3721 2663 3755 2697
rect 3789 2663 3823 2697
rect 3857 2663 3891 2697
rect 3925 2663 3959 2697
rect 3993 2663 4027 2697
rect 4061 2663 4095 2697
rect 4129 2663 4163 2697
rect 4197 2663 4231 2697
rect 4265 2663 4299 2697
rect 4333 2663 4367 2697
rect 4401 2663 4435 2697
rect 4469 2663 4503 2697
rect 4537 2663 4571 2697
rect 4605 2663 4639 2697
rect 4673 2663 4707 2697
rect 4741 2663 4775 2697
rect 4809 2663 4843 2697
rect 4877 2663 4911 2697
rect 4945 2663 4979 2697
rect 5013 2663 5047 2697
rect 5081 2663 5115 2697
rect 5149 2663 5183 2697
rect 5217 2663 5251 2697
rect 5285 2663 5319 2697
rect 5353 2663 5387 2697
rect 5421 2663 5455 2697
rect 5489 2663 5523 2697
rect 5557 2663 5591 2697
rect 5625 2663 5659 2697
rect 5693 2663 5727 2697
rect 5761 2663 5795 2697
rect 5829 2663 5863 2697
rect 5897 2663 5931 2697
rect 5965 2663 5999 2697
rect 6033 2663 6067 2697
rect 6101 2663 6135 2697
rect 6169 2663 6203 2697
rect 6237 2663 6271 2697
rect 6305 2663 6339 2697
rect 6373 2663 6407 2697
rect 6441 2663 6475 2697
rect 6509 2663 6543 2697
rect 6577 2663 6611 2697
rect 6645 2663 6679 2697
rect 6713 2663 6747 2697
rect 6781 2663 6815 2697
rect 6849 2663 6883 2697
rect 6917 2663 6951 2697
rect 6985 2663 7019 2697
rect 7053 2663 7087 2697
rect 7121 2663 7155 2697
rect 7189 2663 7223 2697
rect 7257 2663 7291 2697
rect 7325 2663 7359 2697
rect 7393 2663 7427 2697
rect 7461 2663 7495 2697
rect 7529 2663 7563 2697
rect 7597 2663 7631 2697
rect 7665 2663 7699 2697
rect 7733 2663 7767 2697
rect 7801 2663 7835 2697
rect 7869 2663 7903 2697
rect 7937 2663 7971 2697
rect 8005 2663 8039 2697
rect 8073 2663 8107 2697
rect 8141 2663 8175 2697
rect 8209 2663 8400 2697
rect 0 2640 8400 2663
rect 0 2537 8400 2560
rect 0 2503 151 2537
rect 185 2503 219 2537
rect 253 2503 287 2537
rect 321 2503 355 2537
rect 389 2503 423 2537
rect 457 2503 491 2537
rect 525 2503 559 2537
rect 593 2503 627 2537
rect 661 2503 695 2537
rect 729 2503 763 2537
rect 797 2503 831 2537
rect 865 2503 899 2537
rect 933 2503 967 2537
rect 1001 2503 1035 2537
rect 1069 2503 1103 2537
rect 1137 2503 1171 2537
rect 1205 2503 1239 2537
rect 1273 2503 1307 2537
rect 1341 2503 1375 2537
rect 1409 2503 1443 2537
rect 1477 2503 1511 2537
rect 1545 2503 1579 2537
rect 1613 2503 1647 2537
rect 1681 2503 1715 2537
rect 1749 2503 1783 2537
rect 1817 2503 1851 2537
rect 1885 2503 1919 2537
rect 1953 2503 1987 2537
rect 2021 2503 2055 2537
rect 2089 2503 2123 2537
rect 2157 2503 2191 2537
rect 2225 2503 2259 2537
rect 2293 2503 2327 2537
rect 2361 2503 2395 2537
rect 2429 2503 2463 2537
rect 2497 2503 2531 2537
rect 2565 2503 2599 2537
rect 2633 2503 2667 2537
rect 2701 2503 2735 2537
rect 2769 2503 2803 2537
rect 2837 2503 2871 2537
rect 2905 2503 2939 2537
rect 2973 2503 3007 2537
rect 3041 2503 3075 2537
rect 3109 2503 3143 2537
rect 3177 2503 3211 2537
rect 3245 2503 3279 2537
rect 3313 2503 3347 2537
rect 3381 2503 3415 2537
rect 3449 2503 3483 2537
rect 3517 2503 3551 2537
rect 3585 2503 3619 2537
rect 3653 2503 3687 2537
rect 3721 2503 3755 2537
rect 3789 2503 3823 2537
rect 3857 2503 3891 2537
rect 3925 2503 3959 2537
rect 3993 2503 4027 2537
rect 4061 2503 4095 2537
rect 4129 2503 4163 2537
rect 4197 2503 4231 2537
rect 4265 2503 4299 2537
rect 4333 2503 4367 2537
rect 4401 2503 4435 2537
rect 4469 2503 4503 2537
rect 4537 2503 4571 2537
rect 4605 2503 4639 2537
rect 4673 2503 4707 2537
rect 4741 2503 4775 2537
rect 4809 2503 4843 2537
rect 4877 2503 4911 2537
rect 4945 2503 4979 2537
rect 5013 2503 5047 2537
rect 5081 2503 5115 2537
rect 5149 2503 5183 2537
rect 5217 2503 5251 2537
rect 5285 2503 5319 2537
rect 5353 2503 5387 2537
rect 5421 2503 5455 2537
rect 5489 2503 5523 2537
rect 5557 2503 5591 2537
rect 5625 2503 5659 2537
rect 5693 2503 5727 2537
rect 5761 2503 5795 2537
rect 5829 2503 5863 2537
rect 5897 2503 5931 2537
rect 5965 2503 5999 2537
rect 6033 2503 6067 2537
rect 6101 2503 6135 2537
rect 6169 2503 6203 2537
rect 6237 2503 6271 2537
rect 6305 2503 6339 2537
rect 6373 2503 6407 2537
rect 6441 2503 6475 2537
rect 6509 2503 6543 2537
rect 6577 2503 6611 2537
rect 6645 2503 6679 2537
rect 6713 2503 6747 2537
rect 6781 2503 6815 2537
rect 6849 2503 6883 2537
rect 6917 2503 6951 2537
rect 6985 2503 7019 2537
rect 7053 2503 7087 2537
rect 7121 2503 7155 2537
rect 7189 2503 7223 2537
rect 7257 2503 7291 2537
rect 7325 2503 7359 2537
rect 7393 2503 7427 2537
rect 7461 2503 7495 2537
rect 7529 2503 7563 2537
rect 7597 2503 7631 2537
rect 7665 2503 7699 2537
rect 7733 2503 7767 2537
rect 7801 2503 7835 2537
rect 7869 2503 7903 2537
rect 7937 2503 7971 2537
rect 8005 2503 8039 2537
rect 8073 2503 8107 2537
rect 8141 2503 8175 2537
rect 8209 2503 8400 2537
rect 0 2480 8400 2503
rect 0 2407 80 2480
rect 0 2373 23 2407
rect 57 2373 80 2407
rect 8320 2407 8400 2480
rect 0 2339 80 2373
rect 0 2305 23 2339
rect 57 2305 80 2339
rect 0 2271 80 2305
rect 0 2237 23 2271
rect 57 2237 80 2271
rect 0 2203 80 2237
rect 0 2169 23 2203
rect 57 2169 80 2203
rect 0 2135 80 2169
rect 0 2101 23 2135
rect 57 2101 80 2135
rect 0 2067 80 2101
rect 0 2033 23 2067
rect 57 2033 80 2067
rect 0 1999 80 2033
rect 0 1965 23 1999
rect 57 1965 80 1999
rect 0 1931 80 1965
rect 0 1897 23 1931
rect 57 1897 80 1931
rect 0 1863 80 1897
rect 0 1829 23 1863
rect 57 1829 80 1863
rect 0 1795 80 1829
rect 0 1761 23 1795
rect 57 1761 80 1795
rect 0 1727 80 1761
rect 0 1693 23 1727
rect 57 1693 80 1727
rect 0 1659 80 1693
rect 0 1625 23 1659
rect 57 1625 80 1659
rect 0 1591 80 1625
rect 0 1557 23 1591
rect 57 1557 80 1591
rect 0 1523 80 1557
rect 0 1489 23 1523
rect 57 1489 80 1523
rect 0 1455 80 1489
rect 0 1421 23 1455
rect 57 1421 80 1455
rect 0 1387 80 1421
rect 0 1353 23 1387
rect 57 1353 80 1387
rect 8320 2373 8343 2407
rect 8377 2373 8400 2407
rect 8320 2339 8400 2373
rect 8320 2305 8343 2339
rect 8377 2305 8400 2339
rect 8320 2271 8400 2305
rect 8320 2237 8343 2271
rect 8377 2237 8400 2271
rect 8320 2203 8400 2237
rect 8320 2169 8343 2203
rect 8377 2169 8400 2203
rect 8320 2135 8400 2169
rect 8320 2101 8343 2135
rect 8377 2101 8400 2135
rect 8320 2067 8400 2101
rect 8320 2033 8343 2067
rect 8377 2033 8400 2067
rect 8320 1999 8400 2033
rect 8320 1965 8343 1999
rect 8377 1965 8400 1999
rect 8320 1931 8400 1965
rect 8320 1897 8343 1931
rect 8377 1897 8400 1931
rect 8320 1863 8400 1897
rect 8320 1829 8343 1863
rect 8377 1829 8400 1863
rect 8320 1795 8400 1829
rect 8320 1761 8343 1795
rect 8377 1761 8400 1795
rect 8320 1727 8400 1761
rect 8320 1693 8343 1727
rect 8377 1693 8400 1727
rect 8320 1659 8400 1693
rect 8320 1625 8343 1659
rect 8377 1625 8400 1659
rect 8320 1591 8400 1625
rect 8320 1557 8343 1591
rect 8377 1557 8400 1591
rect 8320 1523 8400 1557
rect 8320 1489 8343 1523
rect 8377 1489 8400 1523
rect 8320 1455 8400 1489
rect 8320 1421 8343 1455
rect 8377 1421 8400 1455
rect 8320 1387 8400 1421
rect 0 1280 80 1353
rect 8320 1353 8343 1387
rect 8377 1353 8400 1387
rect 8320 1280 8400 1353
rect 0 1257 8400 1280
rect 0 1223 137 1257
rect 171 1223 205 1257
rect 239 1223 273 1257
rect 307 1223 341 1257
rect 375 1223 409 1257
rect 443 1223 477 1257
rect 511 1223 545 1257
rect 579 1223 613 1257
rect 647 1223 681 1257
rect 715 1223 749 1257
rect 783 1223 817 1257
rect 851 1223 885 1257
rect 919 1223 953 1257
rect 987 1223 1021 1257
rect 1055 1223 1089 1257
rect 1123 1223 1157 1257
rect 1191 1223 1225 1257
rect 1259 1223 1293 1257
rect 1327 1223 1361 1257
rect 1395 1223 1429 1257
rect 1463 1223 1497 1257
rect 1531 1223 1565 1257
rect 1599 1223 1633 1257
rect 1667 1223 1701 1257
rect 1735 1223 1769 1257
rect 1803 1223 1837 1257
rect 1871 1223 1905 1257
rect 1939 1223 1973 1257
rect 2007 1223 2041 1257
rect 2075 1223 2109 1257
rect 2143 1223 2177 1257
rect 2211 1223 2245 1257
rect 2279 1223 2313 1257
rect 2347 1223 2381 1257
rect 2415 1223 2449 1257
rect 2483 1223 2517 1257
rect 2551 1223 2585 1257
rect 2619 1223 2653 1257
rect 2687 1223 2721 1257
rect 2755 1223 2789 1257
rect 2823 1223 2857 1257
rect 2891 1223 2925 1257
rect 2959 1223 2993 1257
rect 3027 1223 3061 1257
rect 3095 1223 3129 1257
rect 3163 1223 3197 1257
rect 3231 1223 3265 1257
rect 3299 1223 3333 1257
rect 3367 1223 3401 1257
rect 3435 1223 3469 1257
rect 3503 1223 3537 1257
rect 3571 1223 3605 1257
rect 3639 1223 3673 1257
rect 3707 1223 3741 1257
rect 3775 1223 3809 1257
rect 3843 1223 3877 1257
rect 3911 1223 3945 1257
rect 3979 1223 4013 1257
rect 4047 1223 4081 1257
rect 4115 1223 4149 1257
rect 4183 1223 4217 1257
rect 4251 1223 4285 1257
rect 4319 1223 4353 1257
rect 4387 1223 4421 1257
rect 4455 1223 4489 1257
rect 4523 1223 4557 1257
rect 4591 1223 4625 1257
rect 4659 1223 4693 1257
rect 4727 1223 4761 1257
rect 4795 1223 4829 1257
rect 4863 1223 4897 1257
rect 4931 1223 4965 1257
rect 4999 1223 5033 1257
rect 5067 1223 5101 1257
rect 5135 1223 5169 1257
rect 5203 1223 5237 1257
rect 5271 1223 5305 1257
rect 5339 1223 5373 1257
rect 5407 1223 5441 1257
rect 5475 1223 5509 1257
rect 5543 1223 5577 1257
rect 5611 1223 5645 1257
rect 5679 1223 5713 1257
rect 5747 1223 5781 1257
rect 5815 1223 5849 1257
rect 5883 1223 5917 1257
rect 5951 1223 5985 1257
rect 6019 1223 6053 1257
rect 6087 1223 6121 1257
rect 6155 1223 6189 1257
rect 6223 1223 6257 1257
rect 6291 1223 6325 1257
rect 6359 1223 6393 1257
rect 6427 1223 6461 1257
rect 6495 1223 6529 1257
rect 6563 1223 6597 1257
rect 6631 1223 6665 1257
rect 6699 1223 6733 1257
rect 6767 1223 6801 1257
rect 6835 1223 6869 1257
rect 6903 1223 6937 1257
rect 6971 1223 7005 1257
rect 7039 1223 7073 1257
rect 7107 1223 7141 1257
rect 7175 1223 7209 1257
rect 7243 1223 7277 1257
rect 7311 1223 7345 1257
rect 7379 1223 7413 1257
rect 7447 1223 7481 1257
rect 7515 1223 7549 1257
rect 7583 1223 7617 1257
rect 7651 1223 7685 1257
rect 7719 1223 7753 1257
rect 7787 1223 7821 1257
rect 7855 1223 7889 1257
rect 7923 1223 7957 1257
rect 7991 1223 8025 1257
rect 8059 1223 8093 1257
rect 8127 1223 8161 1257
rect 8195 1223 8229 1257
rect 8263 1223 8400 1257
rect 0 1200 8400 1223
rect 0 617 8400 640
rect 0 583 137 617
rect 171 583 205 617
rect 239 583 273 617
rect 307 583 341 617
rect 375 583 409 617
rect 443 583 477 617
rect 511 583 545 617
rect 579 583 613 617
rect 647 583 681 617
rect 715 583 749 617
rect 783 583 817 617
rect 851 583 885 617
rect 919 583 953 617
rect 987 583 1021 617
rect 1055 583 1089 617
rect 1123 583 1157 617
rect 1191 583 1225 617
rect 1259 583 1293 617
rect 1327 583 1361 617
rect 1395 583 1429 617
rect 1463 583 1497 617
rect 1531 583 1565 617
rect 1599 583 1633 617
rect 1667 583 1701 617
rect 1735 583 1769 617
rect 1803 583 1837 617
rect 1871 583 1905 617
rect 1939 583 1973 617
rect 2007 583 2041 617
rect 2075 583 2109 617
rect 2143 583 2177 617
rect 2211 583 2245 617
rect 2279 583 2313 617
rect 2347 583 2381 617
rect 2415 583 2449 617
rect 2483 583 2517 617
rect 2551 583 2585 617
rect 2619 583 2653 617
rect 2687 583 2721 617
rect 2755 583 2789 617
rect 2823 583 2857 617
rect 2891 583 2925 617
rect 2959 583 2993 617
rect 3027 583 3061 617
rect 3095 583 3129 617
rect 3163 583 3197 617
rect 3231 583 3265 617
rect 3299 583 3333 617
rect 3367 583 3401 617
rect 3435 583 3469 617
rect 3503 583 3537 617
rect 3571 583 3605 617
rect 3639 583 3673 617
rect 3707 583 3741 617
rect 3775 583 3809 617
rect 3843 583 3877 617
rect 3911 583 3945 617
rect 3979 583 4013 617
rect 4047 583 4081 617
rect 4115 583 4149 617
rect 4183 583 4217 617
rect 4251 583 4285 617
rect 4319 583 4353 617
rect 4387 583 4421 617
rect 4455 583 4489 617
rect 4523 583 4557 617
rect 4591 583 4625 617
rect 4659 583 4693 617
rect 4727 583 4761 617
rect 4795 583 4829 617
rect 4863 583 4897 617
rect 4931 583 4965 617
rect 4999 583 5033 617
rect 5067 583 5101 617
rect 5135 583 5169 617
rect 5203 583 5237 617
rect 5271 583 5305 617
rect 5339 583 5373 617
rect 5407 583 5441 617
rect 5475 583 5509 617
rect 5543 583 5577 617
rect 5611 583 5645 617
rect 5679 583 5713 617
rect 5747 583 5781 617
rect 5815 583 5849 617
rect 5883 583 5917 617
rect 5951 583 5985 617
rect 6019 583 6053 617
rect 6087 583 6121 617
rect 6155 583 6189 617
rect 6223 583 6257 617
rect 6291 583 6325 617
rect 6359 583 6393 617
rect 6427 583 6461 617
rect 6495 583 6529 617
rect 6563 583 6597 617
rect 6631 583 6665 617
rect 6699 583 6733 617
rect 6767 583 6801 617
rect 6835 583 6869 617
rect 6903 583 6937 617
rect 6971 583 7005 617
rect 7039 583 7073 617
rect 7107 583 7141 617
rect 7175 583 7209 617
rect 7243 583 7277 617
rect 7311 583 7345 617
rect 7379 583 7413 617
rect 7447 583 7481 617
rect 7515 583 7549 617
rect 7583 583 7617 617
rect 7651 583 7685 617
rect 7719 583 7753 617
rect 7787 583 7821 617
rect 7855 583 7889 617
rect 7923 583 7957 617
rect 7991 583 8025 617
rect 8059 583 8093 617
rect 8127 583 8161 617
rect 8195 583 8229 617
rect 8263 583 8400 617
rect 0 560 8400 583
rect 0 507 80 560
rect 0 473 23 507
rect 57 473 80 507
rect 8320 507 8400 560
rect 0 439 80 473
rect 0 405 23 439
rect 57 405 80 439
rect 0 371 80 405
rect 0 337 23 371
rect 57 337 80 371
rect 8320 473 8343 507
rect 8377 473 8400 507
rect 8320 439 8400 473
rect 8320 405 8343 439
rect 8377 405 8400 439
rect 8320 371 8400 405
rect 0 303 80 337
rect 0 269 23 303
rect 57 269 80 303
rect 0 235 80 269
rect 0 201 23 235
rect 57 201 80 235
rect 0 167 80 201
rect 0 133 23 167
rect 57 133 80 167
rect 8320 337 8343 371
rect 8377 337 8400 371
rect 8320 303 8400 337
rect 8320 269 8343 303
rect 8377 269 8400 303
rect 8320 235 8400 269
rect 8320 201 8343 235
rect 8377 201 8400 235
rect 8320 167 8400 201
rect 0 80 80 133
rect 8320 133 8343 167
rect 8377 133 8400 167
rect 8320 80 8400 133
rect 0 57 8400 80
rect 0 23 137 57
rect 171 23 205 57
rect 239 23 273 57
rect 307 23 341 57
rect 375 23 409 57
rect 443 23 477 57
rect 511 23 545 57
rect 579 23 613 57
rect 647 23 681 57
rect 715 23 749 57
rect 783 23 817 57
rect 851 23 885 57
rect 919 23 953 57
rect 987 23 1021 57
rect 1055 23 1089 57
rect 1123 23 1157 57
rect 1191 23 1225 57
rect 1259 23 1293 57
rect 1327 23 1361 57
rect 1395 23 1429 57
rect 1463 23 1497 57
rect 1531 23 1565 57
rect 1599 23 1633 57
rect 1667 23 1701 57
rect 1735 23 1769 57
rect 1803 23 1837 57
rect 1871 23 1905 57
rect 1939 23 1973 57
rect 2007 23 2041 57
rect 2075 23 2109 57
rect 2143 23 2177 57
rect 2211 23 2245 57
rect 2279 23 2313 57
rect 2347 23 2381 57
rect 2415 23 2449 57
rect 2483 23 2517 57
rect 2551 23 2585 57
rect 2619 23 2653 57
rect 2687 23 2721 57
rect 2755 23 2789 57
rect 2823 23 2857 57
rect 2891 23 2925 57
rect 2959 23 2993 57
rect 3027 23 3061 57
rect 3095 23 3129 57
rect 3163 23 3197 57
rect 3231 23 3265 57
rect 3299 23 3333 57
rect 3367 23 3401 57
rect 3435 23 3469 57
rect 3503 23 3537 57
rect 3571 23 3605 57
rect 3639 23 3673 57
rect 3707 23 3741 57
rect 3775 23 3809 57
rect 3843 23 3877 57
rect 3911 23 3945 57
rect 3979 23 4013 57
rect 4047 23 4081 57
rect 4115 23 4149 57
rect 4183 23 4217 57
rect 4251 23 4285 57
rect 4319 23 4353 57
rect 4387 23 4421 57
rect 4455 23 4489 57
rect 4523 23 4557 57
rect 4591 23 4625 57
rect 4659 23 4693 57
rect 4727 23 4761 57
rect 4795 23 4829 57
rect 4863 23 4897 57
rect 4931 23 4965 57
rect 4999 23 5033 57
rect 5067 23 5101 57
rect 5135 23 5169 57
rect 5203 23 5237 57
rect 5271 23 5305 57
rect 5339 23 5373 57
rect 5407 23 5441 57
rect 5475 23 5509 57
rect 5543 23 5577 57
rect 5611 23 5645 57
rect 5679 23 5713 57
rect 5747 23 5781 57
rect 5815 23 5849 57
rect 5883 23 5917 57
rect 5951 23 5985 57
rect 6019 23 6053 57
rect 6087 23 6121 57
rect 6155 23 6189 57
rect 6223 23 6257 57
rect 6291 23 6325 57
rect 6359 23 6393 57
rect 6427 23 6461 57
rect 6495 23 6529 57
rect 6563 23 6597 57
rect 6631 23 6665 57
rect 6699 23 6733 57
rect 6767 23 6801 57
rect 6835 23 6869 57
rect 6903 23 6937 57
rect 6971 23 7005 57
rect 7039 23 7073 57
rect 7107 23 7141 57
rect 7175 23 7209 57
rect 7243 23 7277 57
rect 7311 23 7345 57
rect 7379 23 7413 57
rect 7447 23 7481 57
rect 7515 23 7549 57
rect 7583 23 7617 57
rect 7651 23 7685 57
rect 7719 23 7753 57
rect 7787 23 7821 57
rect 7855 23 7889 57
rect 7923 23 7957 57
rect 7991 23 8025 57
rect 8059 23 8093 57
rect 8127 23 8161 57
rect 8195 23 8229 57
rect 8263 23 8400 57
rect 0 0 8400 23
<< mvnsubdiff >>
rect 160 3817 8240 3840
rect 160 3783 307 3817
rect 341 3783 375 3817
rect 409 3783 443 3817
rect 477 3783 511 3817
rect 545 3783 579 3817
rect 613 3783 647 3817
rect 681 3783 715 3817
rect 749 3783 783 3817
rect 817 3783 851 3817
rect 885 3783 919 3817
rect 953 3783 987 3817
rect 1021 3783 1055 3817
rect 1089 3783 1123 3817
rect 1157 3783 1191 3817
rect 1225 3783 1259 3817
rect 1293 3783 1327 3817
rect 1361 3783 1395 3817
rect 1429 3783 1463 3817
rect 1497 3783 1531 3817
rect 1565 3783 1599 3817
rect 1633 3783 1667 3817
rect 1701 3783 1735 3817
rect 1769 3783 1803 3817
rect 1837 3783 1871 3817
rect 1905 3783 1939 3817
rect 1973 3783 2007 3817
rect 2041 3783 2075 3817
rect 2109 3783 2143 3817
rect 2177 3783 2211 3817
rect 2245 3783 2279 3817
rect 2313 3783 2347 3817
rect 2381 3783 2415 3817
rect 2449 3783 2483 3817
rect 2517 3783 2551 3817
rect 2585 3783 2619 3817
rect 2653 3783 2687 3817
rect 2721 3783 2755 3817
rect 2789 3783 2823 3817
rect 2857 3783 2891 3817
rect 2925 3783 2959 3817
rect 2993 3783 3027 3817
rect 3061 3783 3095 3817
rect 3129 3783 3163 3817
rect 3197 3783 3231 3817
rect 3265 3783 3299 3817
rect 3333 3783 3367 3817
rect 3401 3783 3435 3817
rect 3469 3783 3503 3817
rect 3537 3783 3571 3817
rect 3605 3783 3639 3817
rect 3673 3783 3707 3817
rect 3741 3783 3775 3817
rect 3809 3783 3843 3817
rect 3877 3783 3911 3817
rect 3945 3783 3979 3817
rect 4013 3783 4047 3817
rect 4081 3783 4115 3817
rect 4149 3783 4183 3817
rect 4217 3783 4251 3817
rect 4285 3783 4319 3817
rect 4353 3783 4387 3817
rect 4421 3783 4455 3817
rect 4489 3783 4523 3817
rect 4557 3783 4591 3817
rect 4625 3783 4659 3817
rect 4693 3783 4727 3817
rect 4761 3783 4795 3817
rect 4829 3783 4863 3817
rect 4897 3783 4931 3817
rect 4965 3783 4999 3817
rect 5033 3783 5067 3817
rect 5101 3783 5135 3817
rect 5169 3783 5203 3817
rect 5237 3783 5271 3817
rect 5305 3783 5339 3817
rect 5373 3783 5407 3817
rect 5441 3783 5475 3817
rect 5509 3783 5543 3817
rect 5577 3783 5611 3817
rect 5645 3783 5679 3817
rect 5713 3783 5747 3817
rect 5781 3783 5815 3817
rect 5849 3783 5883 3817
rect 5917 3783 5951 3817
rect 5985 3783 6019 3817
rect 6053 3783 6087 3817
rect 6121 3783 6155 3817
rect 6189 3783 6223 3817
rect 6257 3783 6291 3817
rect 6325 3783 6359 3817
rect 6393 3783 6427 3817
rect 6461 3783 6495 3817
rect 6529 3783 6563 3817
rect 6597 3783 6631 3817
rect 6665 3783 6699 3817
rect 6733 3783 6767 3817
rect 6801 3783 6835 3817
rect 6869 3783 6903 3817
rect 6937 3783 6971 3817
rect 7005 3783 7039 3817
rect 7073 3783 7107 3817
rect 7141 3783 7175 3817
rect 7209 3783 7243 3817
rect 7277 3783 7311 3817
rect 7345 3783 7379 3817
rect 7413 3783 7447 3817
rect 7481 3783 7515 3817
rect 7549 3783 7583 3817
rect 7617 3783 7651 3817
rect 7685 3783 7719 3817
rect 7753 3783 7787 3817
rect 7821 3783 7855 3817
rect 7889 3783 7923 3817
rect 7957 3783 7991 3817
rect 8025 3783 8059 3817
rect 8093 3783 8240 3817
rect 160 3760 8240 3783
rect 160 3711 240 3760
rect 160 3677 183 3711
rect 217 3677 240 3711
rect 8160 3711 8240 3760
rect 160 3643 240 3677
rect 160 3609 183 3643
rect 217 3609 240 3643
rect 160 3575 240 3609
rect 160 3541 183 3575
rect 217 3541 240 3575
rect 160 3507 240 3541
rect 160 3473 183 3507
rect 217 3473 240 3507
rect 160 3439 240 3473
rect 160 3405 183 3439
rect 217 3405 240 3439
rect 160 3371 240 3405
rect 160 3337 183 3371
rect 217 3337 240 3371
rect 160 3303 240 3337
rect 160 3269 183 3303
rect 217 3269 240 3303
rect 160 3235 240 3269
rect 160 3201 183 3235
rect 217 3201 240 3235
rect 160 3167 240 3201
rect 160 3133 183 3167
rect 217 3133 240 3167
rect 160 3099 240 3133
rect 160 3065 183 3099
rect 217 3065 240 3099
rect 8160 3677 8183 3711
rect 8217 3677 8240 3711
rect 8160 3643 8240 3677
rect 8160 3609 8183 3643
rect 8217 3609 8240 3643
rect 8160 3575 8240 3609
rect 8160 3541 8183 3575
rect 8217 3541 8240 3575
rect 8160 3507 8240 3541
rect 8160 3473 8183 3507
rect 8217 3473 8240 3507
rect 8160 3439 8240 3473
rect 8160 3405 8183 3439
rect 8217 3405 8240 3439
rect 8160 3371 8240 3405
rect 8160 3337 8183 3371
rect 8217 3337 8240 3371
rect 8160 3303 8240 3337
rect 8160 3269 8183 3303
rect 8217 3269 8240 3303
rect 8160 3235 8240 3269
rect 8160 3201 8183 3235
rect 8217 3201 8240 3235
rect 8160 3167 8240 3201
rect 8160 3133 8183 3167
rect 8217 3133 8240 3167
rect 8160 3099 8240 3133
rect 160 3031 240 3065
rect 160 2997 183 3031
rect 217 2997 240 3031
rect 160 2963 240 2997
rect 160 2929 183 2963
rect 217 2929 240 2963
rect 8160 3065 8183 3099
rect 8217 3065 8240 3099
rect 8160 3031 8240 3065
rect 8160 2997 8183 3031
rect 8217 2997 8240 3031
rect 8160 2963 8240 2997
rect 160 2880 240 2929
rect 8160 2929 8183 2963
rect 8217 2929 8240 2963
rect 8160 2880 8240 2929
rect 160 2857 8240 2880
rect 160 2823 307 2857
rect 341 2823 375 2857
rect 409 2823 443 2857
rect 477 2823 511 2857
rect 545 2823 579 2857
rect 613 2823 647 2857
rect 681 2823 715 2857
rect 749 2823 783 2857
rect 817 2823 851 2857
rect 885 2823 919 2857
rect 953 2823 987 2857
rect 1021 2823 1055 2857
rect 1089 2823 1123 2857
rect 1157 2823 1191 2857
rect 1225 2823 1259 2857
rect 1293 2823 1327 2857
rect 1361 2823 1395 2857
rect 1429 2823 1463 2857
rect 1497 2823 1531 2857
rect 1565 2823 1599 2857
rect 1633 2823 1667 2857
rect 1701 2823 1735 2857
rect 1769 2823 1803 2857
rect 1837 2823 1871 2857
rect 1905 2823 1939 2857
rect 1973 2823 2007 2857
rect 2041 2823 2075 2857
rect 2109 2823 2143 2857
rect 2177 2823 2211 2857
rect 2245 2823 2279 2857
rect 2313 2823 2347 2857
rect 2381 2823 2415 2857
rect 2449 2823 2483 2857
rect 2517 2823 2551 2857
rect 2585 2823 2619 2857
rect 2653 2823 2687 2857
rect 2721 2823 2755 2857
rect 2789 2823 2823 2857
rect 2857 2823 2891 2857
rect 2925 2823 2959 2857
rect 2993 2823 3027 2857
rect 3061 2823 3095 2857
rect 3129 2823 3163 2857
rect 3197 2823 3231 2857
rect 3265 2823 3299 2857
rect 3333 2823 3367 2857
rect 3401 2823 3435 2857
rect 3469 2823 3503 2857
rect 3537 2823 3571 2857
rect 3605 2823 3639 2857
rect 3673 2823 3707 2857
rect 3741 2823 3775 2857
rect 3809 2823 3843 2857
rect 3877 2823 3911 2857
rect 3945 2823 3979 2857
rect 4013 2823 4047 2857
rect 4081 2823 4115 2857
rect 4149 2823 4183 2857
rect 4217 2823 4251 2857
rect 4285 2823 4319 2857
rect 4353 2823 4387 2857
rect 4421 2823 4455 2857
rect 4489 2823 4523 2857
rect 4557 2823 4591 2857
rect 4625 2823 4659 2857
rect 4693 2823 4727 2857
rect 4761 2823 4795 2857
rect 4829 2823 4863 2857
rect 4897 2823 4931 2857
rect 4965 2823 4999 2857
rect 5033 2823 5067 2857
rect 5101 2823 5135 2857
rect 5169 2823 5203 2857
rect 5237 2823 5271 2857
rect 5305 2823 5339 2857
rect 5373 2823 5407 2857
rect 5441 2823 5475 2857
rect 5509 2823 5543 2857
rect 5577 2823 5611 2857
rect 5645 2823 5679 2857
rect 5713 2823 5747 2857
rect 5781 2823 5815 2857
rect 5849 2823 5883 2857
rect 5917 2823 5951 2857
rect 5985 2823 6019 2857
rect 6053 2823 6087 2857
rect 6121 2823 6155 2857
rect 6189 2823 6223 2857
rect 6257 2823 6291 2857
rect 6325 2823 6359 2857
rect 6393 2823 6427 2857
rect 6461 2823 6495 2857
rect 6529 2823 6563 2857
rect 6597 2823 6631 2857
rect 6665 2823 6699 2857
rect 6733 2823 6767 2857
rect 6801 2823 6835 2857
rect 6869 2823 6903 2857
rect 6937 2823 6971 2857
rect 7005 2823 7039 2857
rect 7073 2823 7107 2857
rect 7141 2823 7175 2857
rect 7209 2823 7243 2857
rect 7277 2823 7311 2857
rect 7345 2823 7379 2857
rect 7413 2823 7447 2857
rect 7481 2823 7515 2857
rect 7549 2823 7583 2857
rect 7617 2823 7651 2857
rect 7685 2823 7719 2857
rect 7753 2823 7787 2857
rect 7821 2823 7855 2857
rect 7889 2823 7923 2857
rect 7957 2823 7991 2857
rect 8025 2823 8059 2857
rect 8093 2823 8240 2857
rect 160 2800 8240 2823
rect 160 2377 8240 2400
rect 160 2343 307 2377
rect 341 2343 375 2377
rect 409 2343 443 2377
rect 477 2343 511 2377
rect 545 2343 579 2377
rect 613 2343 647 2377
rect 681 2343 715 2377
rect 749 2343 783 2377
rect 817 2343 851 2377
rect 885 2343 919 2377
rect 953 2343 987 2377
rect 1021 2343 1055 2377
rect 1089 2343 1123 2377
rect 1157 2343 1191 2377
rect 1225 2343 1259 2377
rect 1293 2343 1327 2377
rect 1361 2343 1395 2377
rect 1429 2343 1463 2377
rect 1497 2343 1531 2377
rect 1565 2343 1599 2377
rect 1633 2343 1667 2377
rect 1701 2343 1735 2377
rect 1769 2343 1803 2377
rect 1837 2343 1871 2377
rect 1905 2343 1939 2377
rect 1973 2343 2007 2377
rect 2041 2343 2075 2377
rect 2109 2343 2143 2377
rect 2177 2343 2211 2377
rect 2245 2343 2279 2377
rect 2313 2343 2347 2377
rect 2381 2343 2415 2377
rect 2449 2343 2483 2377
rect 2517 2343 2551 2377
rect 2585 2343 2619 2377
rect 2653 2343 2687 2377
rect 2721 2343 2755 2377
rect 2789 2343 2823 2377
rect 2857 2343 2891 2377
rect 2925 2343 2959 2377
rect 2993 2343 3027 2377
rect 3061 2343 3095 2377
rect 3129 2343 3163 2377
rect 3197 2343 3231 2377
rect 3265 2343 3299 2377
rect 3333 2343 3367 2377
rect 3401 2343 3435 2377
rect 3469 2343 3503 2377
rect 3537 2343 3571 2377
rect 3605 2343 3639 2377
rect 3673 2343 3707 2377
rect 3741 2343 3775 2377
rect 3809 2343 3843 2377
rect 3877 2343 3911 2377
rect 3945 2343 3979 2377
rect 4013 2343 4047 2377
rect 4081 2343 4115 2377
rect 4149 2343 4183 2377
rect 4217 2343 4251 2377
rect 4285 2343 4319 2377
rect 4353 2343 4387 2377
rect 4421 2343 4455 2377
rect 4489 2343 4523 2377
rect 4557 2343 4591 2377
rect 4625 2343 4659 2377
rect 4693 2343 4727 2377
rect 4761 2343 4795 2377
rect 4829 2343 4863 2377
rect 4897 2343 4931 2377
rect 4965 2343 4999 2377
rect 5033 2343 5067 2377
rect 5101 2343 5135 2377
rect 5169 2343 5203 2377
rect 5237 2343 5271 2377
rect 5305 2343 5339 2377
rect 5373 2343 5407 2377
rect 5441 2343 5475 2377
rect 5509 2343 5543 2377
rect 5577 2343 5611 2377
rect 5645 2343 5679 2377
rect 5713 2343 5747 2377
rect 5781 2343 5815 2377
rect 5849 2343 5883 2377
rect 5917 2343 5951 2377
rect 5985 2343 6019 2377
rect 6053 2343 6087 2377
rect 6121 2343 6155 2377
rect 6189 2343 6223 2377
rect 6257 2343 6291 2377
rect 6325 2343 6359 2377
rect 6393 2343 6427 2377
rect 6461 2343 6495 2377
rect 6529 2343 6563 2377
rect 6597 2343 6631 2377
rect 6665 2343 6699 2377
rect 6733 2343 6767 2377
rect 6801 2343 6835 2377
rect 6869 2343 6903 2377
rect 6937 2343 6971 2377
rect 7005 2343 7039 2377
rect 7073 2343 7107 2377
rect 7141 2343 7175 2377
rect 7209 2343 7243 2377
rect 7277 2343 7311 2377
rect 7345 2343 7379 2377
rect 7413 2343 7447 2377
rect 7481 2343 7515 2377
rect 7549 2343 7583 2377
rect 7617 2343 7651 2377
rect 7685 2343 7719 2377
rect 7753 2343 7787 2377
rect 7821 2343 7855 2377
rect 7889 2343 7923 2377
rect 7957 2343 7991 2377
rect 8025 2343 8059 2377
rect 8093 2343 8240 2377
rect 160 2320 8240 2343
rect 160 2271 240 2320
rect 160 2237 183 2271
rect 217 2237 240 2271
rect 8160 2271 8240 2320
rect 160 2203 240 2237
rect 160 2169 183 2203
rect 217 2169 240 2203
rect 160 2135 240 2169
rect 160 2101 183 2135
rect 217 2101 240 2135
rect 160 2067 240 2101
rect 160 2033 183 2067
rect 217 2033 240 2067
rect 160 1999 240 2033
rect 160 1965 183 1999
rect 217 1965 240 1999
rect 160 1931 240 1965
rect 160 1897 183 1931
rect 217 1897 240 1931
rect 160 1863 240 1897
rect 160 1829 183 1863
rect 217 1829 240 1863
rect 160 1795 240 1829
rect 160 1761 183 1795
rect 217 1761 240 1795
rect 160 1727 240 1761
rect 160 1693 183 1727
rect 217 1693 240 1727
rect 160 1659 240 1693
rect 160 1625 183 1659
rect 217 1625 240 1659
rect 8160 2237 8183 2271
rect 8217 2237 8240 2271
rect 8160 2203 8240 2237
rect 8160 2169 8183 2203
rect 8217 2169 8240 2203
rect 8160 2135 8240 2169
rect 8160 2101 8183 2135
rect 8217 2101 8240 2135
rect 8160 2067 8240 2101
rect 8160 2033 8183 2067
rect 8217 2033 8240 2067
rect 8160 1999 8240 2033
rect 8160 1965 8183 1999
rect 8217 1965 8240 1999
rect 8160 1931 8240 1965
rect 8160 1897 8183 1931
rect 8217 1897 8240 1931
rect 8160 1863 8240 1897
rect 8160 1829 8183 1863
rect 8217 1829 8240 1863
rect 8160 1795 8240 1829
rect 8160 1761 8183 1795
rect 8217 1761 8240 1795
rect 8160 1727 8240 1761
rect 8160 1693 8183 1727
rect 8217 1693 8240 1727
rect 8160 1659 8240 1693
rect 160 1591 240 1625
rect 160 1557 183 1591
rect 217 1557 240 1591
rect 160 1523 240 1557
rect 160 1489 183 1523
rect 217 1489 240 1523
rect 8160 1625 8183 1659
rect 8217 1625 8240 1659
rect 8160 1591 8240 1625
rect 8160 1557 8183 1591
rect 8217 1557 8240 1591
rect 8160 1523 8240 1557
rect 160 1440 240 1489
rect 8160 1489 8183 1523
rect 8217 1489 8240 1523
rect 8160 1440 8240 1489
rect 160 1417 8240 1440
rect 160 1383 307 1417
rect 341 1383 375 1417
rect 409 1383 443 1417
rect 477 1383 511 1417
rect 545 1383 579 1417
rect 613 1383 647 1417
rect 681 1383 715 1417
rect 749 1383 783 1417
rect 817 1383 851 1417
rect 885 1383 919 1417
rect 953 1383 987 1417
rect 1021 1383 1055 1417
rect 1089 1383 1123 1417
rect 1157 1383 1191 1417
rect 1225 1383 1259 1417
rect 1293 1383 1327 1417
rect 1361 1383 1395 1417
rect 1429 1383 1463 1417
rect 1497 1383 1531 1417
rect 1565 1383 1599 1417
rect 1633 1383 1667 1417
rect 1701 1383 1735 1417
rect 1769 1383 1803 1417
rect 1837 1383 1871 1417
rect 1905 1383 1939 1417
rect 1973 1383 2007 1417
rect 2041 1383 2075 1417
rect 2109 1383 2143 1417
rect 2177 1383 2211 1417
rect 2245 1383 2279 1417
rect 2313 1383 2347 1417
rect 2381 1383 2415 1417
rect 2449 1383 2483 1417
rect 2517 1383 2551 1417
rect 2585 1383 2619 1417
rect 2653 1383 2687 1417
rect 2721 1383 2755 1417
rect 2789 1383 2823 1417
rect 2857 1383 2891 1417
rect 2925 1383 2959 1417
rect 2993 1383 3027 1417
rect 3061 1383 3095 1417
rect 3129 1383 3163 1417
rect 3197 1383 3231 1417
rect 3265 1383 3299 1417
rect 3333 1383 3367 1417
rect 3401 1383 3435 1417
rect 3469 1383 3503 1417
rect 3537 1383 3571 1417
rect 3605 1383 3639 1417
rect 3673 1383 3707 1417
rect 3741 1383 3775 1417
rect 3809 1383 3843 1417
rect 3877 1383 3911 1417
rect 3945 1383 3979 1417
rect 4013 1383 4047 1417
rect 4081 1383 4115 1417
rect 4149 1383 4183 1417
rect 4217 1383 4251 1417
rect 4285 1383 4319 1417
rect 4353 1383 4387 1417
rect 4421 1383 4455 1417
rect 4489 1383 4523 1417
rect 4557 1383 4591 1417
rect 4625 1383 4659 1417
rect 4693 1383 4727 1417
rect 4761 1383 4795 1417
rect 4829 1383 4863 1417
rect 4897 1383 4931 1417
rect 4965 1383 4999 1417
rect 5033 1383 5067 1417
rect 5101 1383 5135 1417
rect 5169 1383 5203 1417
rect 5237 1383 5271 1417
rect 5305 1383 5339 1417
rect 5373 1383 5407 1417
rect 5441 1383 5475 1417
rect 5509 1383 5543 1417
rect 5577 1383 5611 1417
rect 5645 1383 5679 1417
rect 5713 1383 5747 1417
rect 5781 1383 5815 1417
rect 5849 1383 5883 1417
rect 5917 1383 5951 1417
rect 5985 1383 6019 1417
rect 6053 1383 6087 1417
rect 6121 1383 6155 1417
rect 6189 1383 6223 1417
rect 6257 1383 6291 1417
rect 6325 1383 6359 1417
rect 6393 1383 6427 1417
rect 6461 1383 6495 1417
rect 6529 1383 6563 1417
rect 6597 1383 6631 1417
rect 6665 1383 6699 1417
rect 6733 1383 6767 1417
rect 6801 1383 6835 1417
rect 6869 1383 6903 1417
rect 6937 1383 6971 1417
rect 7005 1383 7039 1417
rect 7073 1383 7107 1417
rect 7141 1383 7175 1417
rect 7209 1383 7243 1417
rect 7277 1383 7311 1417
rect 7345 1383 7379 1417
rect 7413 1383 7447 1417
rect 7481 1383 7515 1417
rect 7549 1383 7583 1417
rect 7617 1383 7651 1417
rect 7685 1383 7719 1417
rect 7753 1383 7787 1417
rect 7821 1383 7855 1417
rect 7889 1383 7923 1417
rect 7957 1383 7991 1417
rect 8025 1383 8059 1417
rect 8093 1383 8240 1417
rect 160 1360 8240 1383
<< psubdiffcont >>
rect 137 3943 171 3977
rect 205 3943 239 3977
rect 273 3943 307 3977
rect 341 3943 375 3977
rect 409 3943 443 3977
rect 477 3943 511 3977
rect 545 3943 579 3977
rect 613 3943 647 3977
rect 681 3943 715 3977
rect 749 3943 783 3977
rect 817 3943 851 3977
rect 885 3943 919 3977
rect 953 3943 987 3977
rect 1021 3943 1055 3977
rect 1089 3943 1123 3977
rect 1157 3943 1191 3977
rect 1225 3943 1259 3977
rect 1293 3943 1327 3977
rect 1361 3943 1395 3977
rect 1429 3943 1463 3977
rect 1497 3943 1531 3977
rect 1565 3943 1599 3977
rect 1633 3943 1667 3977
rect 1701 3943 1735 3977
rect 1769 3943 1803 3977
rect 1837 3943 1871 3977
rect 1905 3943 1939 3977
rect 1973 3943 2007 3977
rect 2041 3943 2075 3977
rect 2109 3943 2143 3977
rect 2177 3943 2211 3977
rect 2245 3943 2279 3977
rect 2313 3943 2347 3977
rect 2381 3943 2415 3977
rect 2449 3943 2483 3977
rect 2517 3943 2551 3977
rect 2585 3943 2619 3977
rect 2653 3943 2687 3977
rect 2721 3943 2755 3977
rect 2789 3943 2823 3977
rect 2857 3943 2891 3977
rect 2925 3943 2959 3977
rect 2993 3943 3027 3977
rect 3061 3943 3095 3977
rect 3129 3943 3163 3977
rect 3197 3943 3231 3977
rect 3265 3943 3299 3977
rect 3333 3943 3367 3977
rect 3401 3943 3435 3977
rect 3469 3943 3503 3977
rect 3537 3943 3571 3977
rect 3605 3943 3639 3977
rect 3673 3943 3707 3977
rect 3741 3943 3775 3977
rect 3809 3943 3843 3977
rect 3877 3943 3911 3977
rect 3945 3943 3979 3977
rect 4013 3943 4047 3977
rect 4081 3943 4115 3977
rect 4149 3943 4183 3977
rect 4217 3943 4251 3977
rect 4285 3943 4319 3977
rect 4353 3943 4387 3977
rect 4421 3943 4455 3977
rect 4489 3943 4523 3977
rect 4557 3943 4591 3977
rect 4625 3943 4659 3977
rect 4693 3943 4727 3977
rect 4761 3943 4795 3977
rect 4829 3943 4863 3977
rect 4897 3943 4931 3977
rect 4965 3943 4999 3977
rect 5033 3943 5067 3977
rect 5101 3943 5135 3977
rect 5169 3943 5203 3977
rect 5237 3943 5271 3977
rect 5305 3943 5339 3977
rect 5373 3943 5407 3977
rect 5441 3943 5475 3977
rect 5509 3943 5543 3977
rect 5577 3943 5611 3977
rect 5645 3943 5679 3977
rect 5713 3943 5747 3977
rect 5781 3943 5815 3977
rect 5849 3943 5883 3977
rect 5917 3943 5951 3977
rect 5985 3943 6019 3977
rect 6053 3943 6087 3977
rect 6121 3943 6155 3977
rect 6189 3943 6223 3977
rect 6257 3943 6291 3977
rect 6325 3943 6359 3977
rect 6393 3943 6427 3977
rect 6461 3943 6495 3977
rect 6529 3943 6563 3977
rect 6597 3943 6631 3977
rect 6665 3943 6699 3977
rect 6733 3943 6767 3977
rect 6801 3943 6835 3977
rect 6869 3943 6903 3977
rect 6937 3943 6971 3977
rect 7005 3943 7039 3977
rect 7073 3943 7107 3977
rect 7141 3943 7175 3977
rect 7209 3943 7243 3977
rect 7277 3943 7311 3977
rect 7345 3943 7379 3977
rect 7413 3943 7447 3977
rect 7481 3943 7515 3977
rect 7549 3943 7583 3977
rect 7617 3943 7651 3977
rect 7685 3943 7719 3977
rect 7753 3943 7787 3977
rect 7821 3943 7855 3977
rect 7889 3943 7923 3977
rect 7957 3943 7991 3977
rect 8025 3943 8059 3977
rect 8093 3943 8127 3977
rect 8161 3943 8195 3977
rect 8229 3943 8263 3977
rect 23 3813 57 3847
rect 23 3745 57 3779
rect 23 3677 57 3711
rect 23 3609 57 3643
rect 23 3541 57 3575
rect 23 3473 57 3507
rect 23 3405 57 3439
rect 23 3337 57 3371
rect 23 3269 57 3303
rect 23 3201 57 3235
rect 23 3133 57 3167
rect 23 3065 57 3099
rect 23 2997 57 3031
rect 23 2929 57 2963
rect 23 2861 57 2895
rect 23 2793 57 2827
rect 8343 3813 8377 3847
rect 8343 3745 8377 3779
rect 8343 3677 8377 3711
rect 8343 3609 8377 3643
rect 8343 3541 8377 3575
rect 8343 3473 8377 3507
rect 8343 3405 8377 3439
rect 8343 3337 8377 3371
rect 8343 3269 8377 3303
rect 8343 3201 8377 3235
rect 8343 3133 8377 3167
rect 8343 3065 8377 3099
rect 8343 2997 8377 3031
rect 8343 2929 8377 2963
rect 8343 2861 8377 2895
rect 8343 2793 8377 2827
rect 151 2663 185 2697
rect 219 2663 253 2697
rect 287 2663 321 2697
rect 355 2663 389 2697
rect 423 2663 457 2697
rect 491 2663 525 2697
rect 559 2663 593 2697
rect 627 2663 661 2697
rect 695 2663 729 2697
rect 763 2663 797 2697
rect 831 2663 865 2697
rect 899 2663 933 2697
rect 967 2663 1001 2697
rect 1035 2663 1069 2697
rect 1103 2663 1137 2697
rect 1171 2663 1205 2697
rect 1239 2663 1273 2697
rect 1307 2663 1341 2697
rect 1375 2663 1409 2697
rect 1443 2663 1477 2697
rect 1511 2663 1545 2697
rect 1579 2663 1613 2697
rect 1647 2663 1681 2697
rect 1715 2663 1749 2697
rect 1783 2663 1817 2697
rect 1851 2663 1885 2697
rect 1919 2663 1953 2697
rect 1987 2663 2021 2697
rect 2055 2663 2089 2697
rect 2123 2663 2157 2697
rect 2191 2663 2225 2697
rect 2259 2663 2293 2697
rect 2327 2663 2361 2697
rect 2395 2663 2429 2697
rect 2463 2663 2497 2697
rect 2531 2663 2565 2697
rect 2599 2663 2633 2697
rect 2667 2663 2701 2697
rect 2735 2663 2769 2697
rect 2803 2663 2837 2697
rect 2871 2663 2905 2697
rect 2939 2663 2973 2697
rect 3007 2663 3041 2697
rect 3075 2663 3109 2697
rect 3143 2663 3177 2697
rect 3211 2663 3245 2697
rect 3279 2663 3313 2697
rect 3347 2663 3381 2697
rect 3415 2663 3449 2697
rect 3483 2663 3517 2697
rect 3551 2663 3585 2697
rect 3619 2663 3653 2697
rect 3687 2663 3721 2697
rect 3755 2663 3789 2697
rect 3823 2663 3857 2697
rect 3891 2663 3925 2697
rect 3959 2663 3993 2697
rect 4027 2663 4061 2697
rect 4095 2663 4129 2697
rect 4163 2663 4197 2697
rect 4231 2663 4265 2697
rect 4299 2663 4333 2697
rect 4367 2663 4401 2697
rect 4435 2663 4469 2697
rect 4503 2663 4537 2697
rect 4571 2663 4605 2697
rect 4639 2663 4673 2697
rect 4707 2663 4741 2697
rect 4775 2663 4809 2697
rect 4843 2663 4877 2697
rect 4911 2663 4945 2697
rect 4979 2663 5013 2697
rect 5047 2663 5081 2697
rect 5115 2663 5149 2697
rect 5183 2663 5217 2697
rect 5251 2663 5285 2697
rect 5319 2663 5353 2697
rect 5387 2663 5421 2697
rect 5455 2663 5489 2697
rect 5523 2663 5557 2697
rect 5591 2663 5625 2697
rect 5659 2663 5693 2697
rect 5727 2663 5761 2697
rect 5795 2663 5829 2697
rect 5863 2663 5897 2697
rect 5931 2663 5965 2697
rect 5999 2663 6033 2697
rect 6067 2663 6101 2697
rect 6135 2663 6169 2697
rect 6203 2663 6237 2697
rect 6271 2663 6305 2697
rect 6339 2663 6373 2697
rect 6407 2663 6441 2697
rect 6475 2663 6509 2697
rect 6543 2663 6577 2697
rect 6611 2663 6645 2697
rect 6679 2663 6713 2697
rect 6747 2663 6781 2697
rect 6815 2663 6849 2697
rect 6883 2663 6917 2697
rect 6951 2663 6985 2697
rect 7019 2663 7053 2697
rect 7087 2663 7121 2697
rect 7155 2663 7189 2697
rect 7223 2663 7257 2697
rect 7291 2663 7325 2697
rect 7359 2663 7393 2697
rect 7427 2663 7461 2697
rect 7495 2663 7529 2697
rect 7563 2663 7597 2697
rect 7631 2663 7665 2697
rect 7699 2663 7733 2697
rect 7767 2663 7801 2697
rect 7835 2663 7869 2697
rect 7903 2663 7937 2697
rect 7971 2663 8005 2697
rect 8039 2663 8073 2697
rect 8107 2663 8141 2697
rect 8175 2663 8209 2697
rect 151 2503 185 2537
rect 219 2503 253 2537
rect 287 2503 321 2537
rect 355 2503 389 2537
rect 423 2503 457 2537
rect 491 2503 525 2537
rect 559 2503 593 2537
rect 627 2503 661 2537
rect 695 2503 729 2537
rect 763 2503 797 2537
rect 831 2503 865 2537
rect 899 2503 933 2537
rect 967 2503 1001 2537
rect 1035 2503 1069 2537
rect 1103 2503 1137 2537
rect 1171 2503 1205 2537
rect 1239 2503 1273 2537
rect 1307 2503 1341 2537
rect 1375 2503 1409 2537
rect 1443 2503 1477 2537
rect 1511 2503 1545 2537
rect 1579 2503 1613 2537
rect 1647 2503 1681 2537
rect 1715 2503 1749 2537
rect 1783 2503 1817 2537
rect 1851 2503 1885 2537
rect 1919 2503 1953 2537
rect 1987 2503 2021 2537
rect 2055 2503 2089 2537
rect 2123 2503 2157 2537
rect 2191 2503 2225 2537
rect 2259 2503 2293 2537
rect 2327 2503 2361 2537
rect 2395 2503 2429 2537
rect 2463 2503 2497 2537
rect 2531 2503 2565 2537
rect 2599 2503 2633 2537
rect 2667 2503 2701 2537
rect 2735 2503 2769 2537
rect 2803 2503 2837 2537
rect 2871 2503 2905 2537
rect 2939 2503 2973 2537
rect 3007 2503 3041 2537
rect 3075 2503 3109 2537
rect 3143 2503 3177 2537
rect 3211 2503 3245 2537
rect 3279 2503 3313 2537
rect 3347 2503 3381 2537
rect 3415 2503 3449 2537
rect 3483 2503 3517 2537
rect 3551 2503 3585 2537
rect 3619 2503 3653 2537
rect 3687 2503 3721 2537
rect 3755 2503 3789 2537
rect 3823 2503 3857 2537
rect 3891 2503 3925 2537
rect 3959 2503 3993 2537
rect 4027 2503 4061 2537
rect 4095 2503 4129 2537
rect 4163 2503 4197 2537
rect 4231 2503 4265 2537
rect 4299 2503 4333 2537
rect 4367 2503 4401 2537
rect 4435 2503 4469 2537
rect 4503 2503 4537 2537
rect 4571 2503 4605 2537
rect 4639 2503 4673 2537
rect 4707 2503 4741 2537
rect 4775 2503 4809 2537
rect 4843 2503 4877 2537
rect 4911 2503 4945 2537
rect 4979 2503 5013 2537
rect 5047 2503 5081 2537
rect 5115 2503 5149 2537
rect 5183 2503 5217 2537
rect 5251 2503 5285 2537
rect 5319 2503 5353 2537
rect 5387 2503 5421 2537
rect 5455 2503 5489 2537
rect 5523 2503 5557 2537
rect 5591 2503 5625 2537
rect 5659 2503 5693 2537
rect 5727 2503 5761 2537
rect 5795 2503 5829 2537
rect 5863 2503 5897 2537
rect 5931 2503 5965 2537
rect 5999 2503 6033 2537
rect 6067 2503 6101 2537
rect 6135 2503 6169 2537
rect 6203 2503 6237 2537
rect 6271 2503 6305 2537
rect 6339 2503 6373 2537
rect 6407 2503 6441 2537
rect 6475 2503 6509 2537
rect 6543 2503 6577 2537
rect 6611 2503 6645 2537
rect 6679 2503 6713 2537
rect 6747 2503 6781 2537
rect 6815 2503 6849 2537
rect 6883 2503 6917 2537
rect 6951 2503 6985 2537
rect 7019 2503 7053 2537
rect 7087 2503 7121 2537
rect 7155 2503 7189 2537
rect 7223 2503 7257 2537
rect 7291 2503 7325 2537
rect 7359 2503 7393 2537
rect 7427 2503 7461 2537
rect 7495 2503 7529 2537
rect 7563 2503 7597 2537
rect 7631 2503 7665 2537
rect 7699 2503 7733 2537
rect 7767 2503 7801 2537
rect 7835 2503 7869 2537
rect 7903 2503 7937 2537
rect 7971 2503 8005 2537
rect 8039 2503 8073 2537
rect 8107 2503 8141 2537
rect 8175 2503 8209 2537
rect 23 2373 57 2407
rect 23 2305 57 2339
rect 23 2237 57 2271
rect 23 2169 57 2203
rect 23 2101 57 2135
rect 23 2033 57 2067
rect 23 1965 57 1999
rect 23 1897 57 1931
rect 23 1829 57 1863
rect 23 1761 57 1795
rect 23 1693 57 1727
rect 23 1625 57 1659
rect 23 1557 57 1591
rect 23 1489 57 1523
rect 23 1421 57 1455
rect 23 1353 57 1387
rect 8343 2373 8377 2407
rect 8343 2305 8377 2339
rect 8343 2237 8377 2271
rect 8343 2169 8377 2203
rect 8343 2101 8377 2135
rect 8343 2033 8377 2067
rect 8343 1965 8377 1999
rect 8343 1897 8377 1931
rect 8343 1829 8377 1863
rect 8343 1761 8377 1795
rect 8343 1693 8377 1727
rect 8343 1625 8377 1659
rect 8343 1557 8377 1591
rect 8343 1489 8377 1523
rect 8343 1421 8377 1455
rect 8343 1353 8377 1387
rect 137 1223 171 1257
rect 205 1223 239 1257
rect 273 1223 307 1257
rect 341 1223 375 1257
rect 409 1223 443 1257
rect 477 1223 511 1257
rect 545 1223 579 1257
rect 613 1223 647 1257
rect 681 1223 715 1257
rect 749 1223 783 1257
rect 817 1223 851 1257
rect 885 1223 919 1257
rect 953 1223 987 1257
rect 1021 1223 1055 1257
rect 1089 1223 1123 1257
rect 1157 1223 1191 1257
rect 1225 1223 1259 1257
rect 1293 1223 1327 1257
rect 1361 1223 1395 1257
rect 1429 1223 1463 1257
rect 1497 1223 1531 1257
rect 1565 1223 1599 1257
rect 1633 1223 1667 1257
rect 1701 1223 1735 1257
rect 1769 1223 1803 1257
rect 1837 1223 1871 1257
rect 1905 1223 1939 1257
rect 1973 1223 2007 1257
rect 2041 1223 2075 1257
rect 2109 1223 2143 1257
rect 2177 1223 2211 1257
rect 2245 1223 2279 1257
rect 2313 1223 2347 1257
rect 2381 1223 2415 1257
rect 2449 1223 2483 1257
rect 2517 1223 2551 1257
rect 2585 1223 2619 1257
rect 2653 1223 2687 1257
rect 2721 1223 2755 1257
rect 2789 1223 2823 1257
rect 2857 1223 2891 1257
rect 2925 1223 2959 1257
rect 2993 1223 3027 1257
rect 3061 1223 3095 1257
rect 3129 1223 3163 1257
rect 3197 1223 3231 1257
rect 3265 1223 3299 1257
rect 3333 1223 3367 1257
rect 3401 1223 3435 1257
rect 3469 1223 3503 1257
rect 3537 1223 3571 1257
rect 3605 1223 3639 1257
rect 3673 1223 3707 1257
rect 3741 1223 3775 1257
rect 3809 1223 3843 1257
rect 3877 1223 3911 1257
rect 3945 1223 3979 1257
rect 4013 1223 4047 1257
rect 4081 1223 4115 1257
rect 4149 1223 4183 1257
rect 4217 1223 4251 1257
rect 4285 1223 4319 1257
rect 4353 1223 4387 1257
rect 4421 1223 4455 1257
rect 4489 1223 4523 1257
rect 4557 1223 4591 1257
rect 4625 1223 4659 1257
rect 4693 1223 4727 1257
rect 4761 1223 4795 1257
rect 4829 1223 4863 1257
rect 4897 1223 4931 1257
rect 4965 1223 4999 1257
rect 5033 1223 5067 1257
rect 5101 1223 5135 1257
rect 5169 1223 5203 1257
rect 5237 1223 5271 1257
rect 5305 1223 5339 1257
rect 5373 1223 5407 1257
rect 5441 1223 5475 1257
rect 5509 1223 5543 1257
rect 5577 1223 5611 1257
rect 5645 1223 5679 1257
rect 5713 1223 5747 1257
rect 5781 1223 5815 1257
rect 5849 1223 5883 1257
rect 5917 1223 5951 1257
rect 5985 1223 6019 1257
rect 6053 1223 6087 1257
rect 6121 1223 6155 1257
rect 6189 1223 6223 1257
rect 6257 1223 6291 1257
rect 6325 1223 6359 1257
rect 6393 1223 6427 1257
rect 6461 1223 6495 1257
rect 6529 1223 6563 1257
rect 6597 1223 6631 1257
rect 6665 1223 6699 1257
rect 6733 1223 6767 1257
rect 6801 1223 6835 1257
rect 6869 1223 6903 1257
rect 6937 1223 6971 1257
rect 7005 1223 7039 1257
rect 7073 1223 7107 1257
rect 7141 1223 7175 1257
rect 7209 1223 7243 1257
rect 7277 1223 7311 1257
rect 7345 1223 7379 1257
rect 7413 1223 7447 1257
rect 7481 1223 7515 1257
rect 7549 1223 7583 1257
rect 7617 1223 7651 1257
rect 7685 1223 7719 1257
rect 7753 1223 7787 1257
rect 7821 1223 7855 1257
rect 7889 1223 7923 1257
rect 7957 1223 7991 1257
rect 8025 1223 8059 1257
rect 8093 1223 8127 1257
rect 8161 1223 8195 1257
rect 8229 1223 8263 1257
rect 137 583 171 617
rect 205 583 239 617
rect 273 583 307 617
rect 341 583 375 617
rect 409 583 443 617
rect 477 583 511 617
rect 545 583 579 617
rect 613 583 647 617
rect 681 583 715 617
rect 749 583 783 617
rect 817 583 851 617
rect 885 583 919 617
rect 953 583 987 617
rect 1021 583 1055 617
rect 1089 583 1123 617
rect 1157 583 1191 617
rect 1225 583 1259 617
rect 1293 583 1327 617
rect 1361 583 1395 617
rect 1429 583 1463 617
rect 1497 583 1531 617
rect 1565 583 1599 617
rect 1633 583 1667 617
rect 1701 583 1735 617
rect 1769 583 1803 617
rect 1837 583 1871 617
rect 1905 583 1939 617
rect 1973 583 2007 617
rect 2041 583 2075 617
rect 2109 583 2143 617
rect 2177 583 2211 617
rect 2245 583 2279 617
rect 2313 583 2347 617
rect 2381 583 2415 617
rect 2449 583 2483 617
rect 2517 583 2551 617
rect 2585 583 2619 617
rect 2653 583 2687 617
rect 2721 583 2755 617
rect 2789 583 2823 617
rect 2857 583 2891 617
rect 2925 583 2959 617
rect 2993 583 3027 617
rect 3061 583 3095 617
rect 3129 583 3163 617
rect 3197 583 3231 617
rect 3265 583 3299 617
rect 3333 583 3367 617
rect 3401 583 3435 617
rect 3469 583 3503 617
rect 3537 583 3571 617
rect 3605 583 3639 617
rect 3673 583 3707 617
rect 3741 583 3775 617
rect 3809 583 3843 617
rect 3877 583 3911 617
rect 3945 583 3979 617
rect 4013 583 4047 617
rect 4081 583 4115 617
rect 4149 583 4183 617
rect 4217 583 4251 617
rect 4285 583 4319 617
rect 4353 583 4387 617
rect 4421 583 4455 617
rect 4489 583 4523 617
rect 4557 583 4591 617
rect 4625 583 4659 617
rect 4693 583 4727 617
rect 4761 583 4795 617
rect 4829 583 4863 617
rect 4897 583 4931 617
rect 4965 583 4999 617
rect 5033 583 5067 617
rect 5101 583 5135 617
rect 5169 583 5203 617
rect 5237 583 5271 617
rect 5305 583 5339 617
rect 5373 583 5407 617
rect 5441 583 5475 617
rect 5509 583 5543 617
rect 5577 583 5611 617
rect 5645 583 5679 617
rect 5713 583 5747 617
rect 5781 583 5815 617
rect 5849 583 5883 617
rect 5917 583 5951 617
rect 5985 583 6019 617
rect 6053 583 6087 617
rect 6121 583 6155 617
rect 6189 583 6223 617
rect 6257 583 6291 617
rect 6325 583 6359 617
rect 6393 583 6427 617
rect 6461 583 6495 617
rect 6529 583 6563 617
rect 6597 583 6631 617
rect 6665 583 6699 617
rect 6733 583 6767 617
rect 6801 583 6835 617
rect 6869 583 6903 617
rect 6937 583 6971 617
rect 7005 583 7039 617
rect 7073 583 7107 617
rect 7141 583 7175 617
rect 7209 583 7243 617
rect 7277 583 7311 617
rect 7345 583 7379 617
rect 7413 583 7447 617
rect 7481 583 7515 617
rect 7549 583 7583 617
rect 7617 583 7651 617
rect 7685 583 7719 617
rect 7753 583 7787 617
rect 7821 583 7855 617
rect 7889 583 7923 617
rect 7957 583 7991 617
rect 8025 583 8059 617
rect 8093 583 8127 617
rect 8161 583 8195 617
rect 8229 583 8263 617
rect 23 473 57 507
rect 23 405 57 439
rect 23 337 57 371
rect 8343 473 8377 507
rect 8343 405 8377 439
rect 23 269 57 303
rect 23 201 57 235
rect 23 133 57 167
rect 8343 337 8377 371
rect 8343 269 8377 303
rect 8343 201 8377 235
rect 8343 133 8377 167
rect 137 23 171 57
rect 205 23 239 57
rect 273 23 307 57
rect 341 23 375 57
rect 409 23 443 57
rect 477 23 511 57
rect 545 23 579 57
rect 613 23 647 57
rect 681 23 715 57
rect 749 23 783 57
rect 817 23 851 57
rect 885 23 919 57
rect 953 23 987 57
rect 1021 23 1055 57
rect 1089 23 1123 57
rect 1157 23 1191 57
rect 1225 23 1259 57
rect 1293 23 1327 57
rect 1361 23 1395 57
rect 1429 23 1463 57
rect 1497 23 1531 57
rect 1565 23 1599 57
rect 1633 23 1667 57
rect 1701 23 1735 57
rect 1769 23 1803 57
rect 1837 23 1871 57
rect 1905 23 1939 57
rect 1973 23 2007 57
rect 2041 23 2075 57
rect 2109 23 2143 57
rect 2177 23 2211 57
rect 2245 23 2279 57
rect 2313 23 2347 57
rect 2381 23 2415 57
rect 2449 23 2483 57
rect 2517 23 2551 57
rect 2585 23 2619 57
rect 2653 23 2687 57
rect 2721 23 2755 57
rect 2789 23 2823 57
rect 2857 23 2891 57
rect 2925 23 2959 57
rect 2993 23 3027 57
rect 3061 23 3095 57
rect 3129 23 3163 57
rect 3197 23 3231 57
rect 3265 23 3299 57
rect 3333 23 3367 57
rect 3401 23 3435 57
rect 3469 23 3503 57
rect 3537 23 3571 57
rect 3605 23 3639 57
rect 3673 23 3707 57
rect 3741 23 3775 57
rect 3809 23 3843 57
rect 3877 23 3911 57
rect 3945 23 3979 57
rect 4013 23 4047 57
rect 4081 23 4115 57
rect 4149 23 4183 57
rect 4217 23 4251 57
rect 4285 23 4319 57
rect 4353 23 4387 57
rect 4421 23 4455 57
rect 4489 23 4523 57
rect 4557 23 4591 57
rect 4625 23 4659 57
rect 4693 23 4727 57
rect 4761 23 4795 57
rect 4829 23 4863 57
rect 4897 23 4931 57
rect 4965 23 4999 57
rect 5033 23 5067 57
rect 5101 23 5135 57
rect 5169 23 5203 57
rect 5237 23 5271 57
rect 5305 23 5339 57
rect 5373 23 5407 57
rect 5441 23 5475 57
rect 5509 23 5543 57
rect 5577 23 5611 57
rect 5645 23 5679 57
rect 5713 23 5747 57
rect 5781 23 5815 57
rect 5849 23 5883 57
rect 5917 23 5951 57
rect 5985 23 6019 57
rect 6053 23 6087 57
rect 6121 23 6155 57
rect 6189 23 6223 57
rect 6257 23 6291 57
rect 6325 23 6359 57
rect 6393 23 6427 57
rect 6461 23 6495 57
rect 6529 23 6563 57
rect 6597 23 6631 57
rect 6665 23 6699 57
rect 6733 23 6767 57
rect 6801 23 6835 57
rect 6869 23 6903 57
rect 6937 23 6971 57
rect 7005 23 7039 57
rect 7073 23 7107 57
rect 7141 23 7175 57
rect 7209 23 7243 57
rect 7277 23 7311 57
rect 7345 23 7379 57
rect 7413 23 7447 57
rect 7481 23 7515 57
rect 7549 23 7583 57
rect 7617 23 7651 57
rect 7685 23 7719 57
rect 7753 23 7787 57
rect 7821 23 7855 57
rect 7889 23 7923 57
rect 7957 23 7991 57
rect 8025 23 8059 57
rect 8093 23 8127 57
rect 8161 23 8195 57
rect 8229 23 8263 57
<< mvnsubdiffcont >>
rect 307 3783 341 3817
rect 375 3783 409 3817
rect 443 3783 477 3817
rect 511 3783 545 3817
rect 579 3783 613 3817
rect 647 3783 681 3817
rect 715 3783 749 3817
rect 783 3783 817 3817
rect 851 3783 885 3817
rect 919 3783 953 3817
rect 987 3783 1021 3817
rect 1055 3783 1089 3817
rect 1123 3783 1157 3817
rect 1191 3783 1225 3817
rect 1259 3783 1293 3817
rect 1327 3783 1361 3817
rect 1395 3783 1429 3817
rect 1463 3783 1497 3817
rect 1531 3783 1565 3817
rect 1599 3783 1633 3817
rect 1667 3783 1701 3817
rect 1735 3783 1769 3817
rect 1803 3783 1837 3817
rect 1871 3783 1905 3817
rect 1939 3783 1973 3817
rect 2007 3783 2041 3817
rect 2075 3783 2109 3817
rect 2143 3783 2177 3817
rect 2211 3783 2245 3817
rect 2279 3783 2313 3817
rect 2347 3783 2381 3817
rect 2415 3783 2449 3817
rect 2483 3783 2517 3817
rect 2551 3783 2585 3817
rect 2619 3783 2653 3817
rect 2687 3783 2721 3817
rect 2755 3783 2789 3817
rect 2823 3783 2857 3817
rect 2891 3783 2925 3817
rect 2959 3783 2993 3817
rect 3027 3783 3061 3817
rect 3095 3783 3129 3817
rect 3163 3783 3197 3817
rect 3231 3783 3265 3817
rect 3299 3783 3333 3817
rect 3367 3783 3401 3817
rect 3435 3783 3469 3817
rect 3503 3783 3537 3817
rect 3571 3783 3605 3817
rect 3639 3783 3673 3817
rect 3707 3783 3741 3817
rect 3775 3783 3809 3817
rect 3843 3783 3877 3817
rect 3911 3783 3945 3817
rect 3979 3783 4013 3817
rect 4047 3783 4081 3817
rect 4115 3783 4149 3817
rect 4183 3783 4217 3817
rect 4251 3783 4285 3817
rect 4319 3783 4353 3817
rect 4387 3783 4421 3817
rect 4455 3783 4489 3817
rect 4523 3783 4557 3817
rect 4591 3783 4625 3817
rect 4659 3783 4693 3817
rect 4727 3783 4761 3817
rect 4795 3783 4829 3817
rect 4863 3783 4897 3817
rect 4931 3783 4965 3817
rect 4999 3783 5033 3817
rect 5067 3783 5101 3817
rect 5135 3783 5169 3817
rect 5203 3783 5237 3817
rect 5271 3783 5305 3817
rect 5339 3783 5373 3817
rect 5407 3783 5441 3817
rect 5475 3783 5509 3817
rect 5543 3783 5577 3817
rect 5611 3783 5645 3817
rect 5679 3783 5713 3817
rect 5747 3783 5781 3817
rect 5815 3783 5849 3817
rect 5883 3783 5917 3817
rect 5951 3783 5985 3817
rect 6019 3783 6053 3817
rect 6087 3783 6121 3817
rect 6155 3783 6189 3817
rect 6223 3783 6257 3817
rect 6291 3783 6325 3817
rect 6359 3783 6393 3817
rect 6427 3783 6461 3817
rect 6495 3783 6529 3817
rect 6563 3783 6597 3817
rect 6631 3783 6665 3817
rect 6699 3783 6733 3817
rect 6767 3783 6801 3817
rect 6835 3783 6869 3817
rect 6903 3783 6937 3817
rect 6971 3783 7005 3817
rect 7039 3783 7073 3817
rect 7107 3783 7141 3817
rect 7175 3783 7209 3817
rect 7243 3783 7277 3817
rect 7311 3783 7345 3817
rect 7379 3783 7413 3817
rect 7447 3783 7481 3817
rect 7515 3783 7549 3817
rect 7583 3783 7617 3817
rect 7651 3783 7685 3817
rect 7719 3783 7753 3817
rect 7787 3783 7821 3817
rect 7855 3783 7889 3817
rect 7923 3783 7957 3817
rect 7991 3783 8025 3817
rect 8059 3783 8093 3817
rect 183 3677 217 3711
rect 183 3609 217 3643
rect 183 3541 217 3575
rect 183 3473 217 3507
rect 183 3405 217 3439
rect 183 3337 217 3371
rect 183 3269 217 3303
rect 183 3201 217 3235
rect 183 3133 217 3167
rect 183 3065 217 3099
rect 8183 3677 8217 3711
rect 8183 3609 8217 3643
rect 8183 3541 8217 3575
rect 8183 3473 8217 3507
rect 8183 3405 8217 3439
rect 8183 3337 8217 3371
rect 8183 3269 8217 3303
rect 8183 3201 8217 3235
rect 8183 3133 8217 3167
rect 183 2997 217 3031
rect 183 2929 217 2963
rect 8183 3065 8217 3099
rect 8183 2997 8217 3031
rect 8183 2929 8217 2963
rect 307 2823 341 2857
rect 375 2823 409 2857
rect 443 2823 477 2857
rect 511 2823 545 2857
rect 579 2823 613 2857
rect 647 2823 681 2857
rect 715 2823 749 2857
rect 783 2823 817 2857
rect 851 2823 885 2857
rect 919 2823 953 2857
rect 987 2823 1021 2857
rect 1055 2823 1089 2857
rect 1123 2823 1157 2857
rect 1191 2823 1225 2857
rect 1259 2823 1293 2857
rect 1327 2823 1361 2857
rect 1395 2823 1429 2857
rect 1463 2823 1497 2857
rect 1531 2823 1565 2857
rect 1599 2823 1633 2857
rect 1667 2823 1701 2857
rect 1735 2823 1769 2857
rect 1803 2823 1837 2857
rect 1871 2823 1905 2857
rect 1939 2823 1973 2857
rect 2007 2823 2041 2857
rect 2075 2823 2109 2857
rect 2143 2823 2177 2857
rect 2211 2823 2245 2857
rect 2279 2823 2313 2857
rect 2347 2823 2381 2857
rect 2415 2823 2449 2857
rect 2483 2823 2517 2857
rect 2551 2823 2585 2857
rect 2619 2823 2653 2857
rect 2687 2823 2721 2857
rect 2755 2823 2789 2857
rect 2823 2823 2857 2857
rect 2891 2823 2925 2857
rect 2959 2823 2993 2857
rect 3027 2823 3061 2857
rect 3095 2823 3129 2857
rect 3163 2823 3197 2857
rect 3231 2823 3265 2857
rect 3299 2823 3333 2857
rect 3367 2823 3401 2857
rect 3435 2823 3469 2857
rect 3503 2823 3537 2857
rect 3571 2823 3605 2857
rect 3639 2823 3673 2857
rect 3707 2823 3741 2857
rect 3775 2823 3809 2857
rect 3843 2823 3877 2857
rect 3911 2823 3945 2857
rect 3979 2823 4013 2857
rect 4047 2823 4081 2857
rect 4115 2823 4149 2857
rect 4183 2823 4217 2857
rect 4251 2823 4285 2857
rect 4319 2823 4353 2857
rect 4387 2823 4421 2857
rect 4455 2823 4489 2857
rect 4523 2823 4557 2857
rect 4591 2823 4625 2857
rect 4659 2823 4693 2857
rect 4727 2823 4761 2857
rect 4795 2823 4829 2857
rect 4863 2823 4897 2857
rect 4931 2823 4965 2857
rect 4999 2823 5033 2857
rect 5067 2823 5101 2857
rect 5135 2823 5169 2857
rect 5203 2823 5237 2857
rect 5271 2823 5305 2857
rect 5339 2823 5373 2857
rect 5407 2823 5441 2857
rect 5475 2823 5509 2857
rect 5543 2823 5577 2857
rect 5611 2823 5645 2857
rect 5679 2823 5713 2857
rect 5747 2823 5781 2857
rect 5815 2823 5849 2857
rect 5883 2823 5917 2857
rect 5951 2823 5985 2857
rect 6019 2823 6053 2857
rect 6087 2823 6121 2857
rect 6155 2823 6189 2857
rect 6223 2823 6257 2857
rect 6291 2823 6325 2857
rect 6359 2823 6393 2857
rect 6427 2823 6461 2857
rect 6495 2823 6529 2857
rect 6563 2823 6597 2857
rect 6631 2823 6665 2857
rect 6699 2823 6733 2857
rect 6767 2823 6801 2857
rect 6835 2823 6869 2857
rect 6903 2823 6937 2857
rect 6971 2823 7005 2857
rect 7039 2823 7073 2857
rect 7107 2823 7141 2857
rect 7175 2823 7209 2857
rect 7243 2823 7277 2857
rect 7311 2823 7345 2857
rect 7379 2823 7413 2857
rect 7447 2823 7481 2857
rect 7515 2823 7549 2857
rect 7583 2823 7617 2857
rect 7651 2823 7685 2857
rect 7719 2823 7753 2857
rect 7787 2823 7821 2857
rect 7855 2823 7889 2857
rect 7923 2823 7957 2857
rect 7991 2823 8025 2857
rect 8059 2823 8093 2857
rect 307 2343 341 2377
rect 375 2343 409 2377
rect 443 2343 477 2377
rect 511 2343 545 2377
rect 579 2343 613 2377
rect 647 2343 681 2377
rect 715 2343 749 2377
rect 783 2343 817 2377
rect 851 2343 885 2377
rect 919 2343 953 2377
rect 987 2343 1021 2377
rect 1055 2343 1089 2377
rect 1123 2343 1157 2377
rect 1191 2343 1225 2377
rect 1259 2343 1293 2377
rect 1327 2343 1361 2377
rect 1395 2343 1429 2377
rect 1463 2343 1497 2377
rect 1531 2343 1565 2377
rect 1599 2343 1633 2377
rect 1667 2343 1701 2377
rect 1735 2343 1769 2377
rect 1803 2343 1837 2377
rect 1871 2343 1905 2377
rect 1939 2343 1973 2377
rect 2007 2343 2041 2377
rect 2075 2343 2109 2377
rect 2143 2343 2177 2377
rect 2211 2343 2245 2377
rect 2279 2343 2313 2377
rect 2347 2343 2381 2377
rect 2415 2343 2449 2377
rect 2483 2343 2517 2377
rect 2551 2343 2585 2377
rect 2619 2343 2653 2377
rect 2687 2343 2721 2377
rect 2755 2343 2789 2377
rect 2823 2343 2857 2377
rect 2891 2343 2925 2377
rect 2959 2343 2993 2377
rect 3027 2343 3061 2377
rect 3095 2343 3129 2377
rect 3163 2343 3197 2377
rect 3231 2343 3265 2377
rect 3299 2343 3333 2377
rect 3367 2343 3401 2377
rect 3435 2343 3469 2377
rect 3503 2343 3537 2377
rect 3571 2343 3605 2377
rect 3639 2343 3673 2377
rect 3707 2343 3741 2377
rect 3775 2343 3809 2377
rect 3843 2343 3877 2377
rect 3911 2343 3945 2377
rect 3979 2343 4013 2377
rect 4047 2343 4081 2377
rect 4115 2343 4149 2377
rect 4183 2343 4217 2377
rect 4251 2343 4285 2377
rect 4319 2343 4353 2377
rect 4387 2343 4421 2377
rect 4455 2343 4489 2377
rect 4523 2343 4557 2377
rect 4591 2343 4625 2377
rect 4659 2343 4693 2377
rect 4727 2343 4761 2377
rect 4795 2343 4829 2377
rect 4863 2343 4897 2377
rect 4931 2343 4965 2377
rect 4999 2343 5033 2377
rect 5067 2343 5101 2377
rect 5135 2343 5169 2377
rect 5203 2343 5237 2377
rect 5271 2343 5305 2377
rect 5339 2343 5373 2377
rect 5407 2343 5441 2377
rect 5475 2343 5509 2377
rect 5543 2343 5577 2377
rect 5611 2343 5645 2377
rect 5679 2343 5713 2377
rect 5747 2343 5781 2377
rect 5815 2343 5849 2377
rect 5883 2343 5917 2377
rect 5951 2343 5985 2377
rect 6019 2343 6053 2377
rect 6087 2343 6121 2377
rect 6155 2343 6189 2377
rect 6223 2343 6257 2377
rect 6291 2343 6325 2377
rect 6359 2343 6393 2377
rect 6427 2343 6461 2377
rect 6495 2343 6529 2377
rect 6563 2343 6597 2377
rect 6631 2343 6665 2377
rect 6699 2343 6733 2377
rect 6767 2343 6801 2377
rect 6835 2343 6869 2377
rect 6903 2343 6937 2377
rect 6971 2343 7005 2377
rect 7039 2343 7073 2377
rect 7107 2343 7141 2377
rect 7175 2343 7209 2377
rect 7243 2343 7277 2377
rect 7311 2343 7345 2377
rect 7379 2343 7413 2377
rect 7447 2343 7481 2377
rect 7515 2343 7549 2377
rect 7583 2343 7617 2377
rect 7651 2343 7685 2377
rect 7719 2343 7753 2377
rect 7787 2343 7821 2377
rect 7855 2343 7889 2377
rect 7923 2343 7957 2377
rect 7991 2343 8025 2377
rect 8059 2343 8093 2377
rect 183 2237 217 2271
rect 183 2169 217 2203
rect 183 2101 217 2135
rect 183 2033 217 2067
rect 183 1965 217 1999
rect 183 1897 217 1931
rect 183 1829 217 1863
rect 183 1761 217 1795
rect 183 1693 217 1727
rect 183 1625 217 1659
rect 8183 2237 8217 2271
rect 8183 2169 8217 2203
rect 8183 2101 8217 2135
rect 8183 2033 8217 2067
rect 8183 1965 8217 1999
rect 8183 1897 8217 1931
rect 8183 1829 8217 1863
rect 8183 1761 8217 1795
rect 8183 1693 8217 1727
rect 183 1557 217 1591
rect 183 1489 217 1523
rect 8183 1625 8217 1659
rect 8183 1557 8217 1591
rect 8183 1489 8217 1523
rect 307 1383 341 1417
rect 375 1383 409 1417
rect 443 1383 477 1417
rect 511 1383 545 1417
rect 579 1383 613 1417
rect 647 1383 681 1417
rect 715 1383 749 1417
rect 783 1383 817 1417
rect 851 1383 885 1417
rect 919 1383 953 1417
rect 987 1383 1021 1417
rect 1055 1383 1089 1417
rect 1123 1383 1157 1417
rect 1191 1383 1225 1417
rect 1259 1383 1293 1417
rect 1327 1383 1361 1417
rect 1395 1383 1429 1417
rect 1463 1383 1497 1417
rect 1531 1383 1565 1417
rect 1599 1383 1633 1417
rect 1667 1383 1701 1417
rect 1735 1383 1769 1417
rect 1803 1383 1837 1417
rect 1871 1383 1905 1417
rect 1939 1383 1973 1417
rect 2007 1383 2041 1417
rect 2075 1383 2109 1417
rect 2143 1383 2177 1417
rect 2211 1383 2245 1417
rect 2279 1383 2313 1417
rect 2347 1383 2381 1417
rect 2415 1383 2449 1417
rect 2483 1383 2517 1417
rect 2551 1383 2585 1417
rect 2619 1383 2653 1417
rect 2687 1383 2721 1417
rect 2755 1383 2789 1417
rect 2823 1383 2857 1417
rect 2891 1383 2925 1417
rect 2959 1383 2993 1417
rect 3027 1383 3061 1417
rect 3095 1383 3129 1417
rect 3163 1383 3197 1417
rect 3231 1383 3265 1417
rect 3299 1383 3333 1417
rect 3367 1383 3401 1417
rect 3435 1383 3469 1417
rect 3503 1383 3537 1417
rect 3571 1383 3605 1417
rect 3639 1383 3673 1417
rect 3707 1383 3741 1417
rect 3775 1383 3809 1417
rect 3843 1383 3877 1417
rect 3911 1383 3945 1417
rect 3979 1383 4013 1417
rect 4047 1383 4081 1417
rect 4115 1383 4149 1417
rect 4183 1383 4217 1417
rect 4251 1383 4285 1417
rect 4319 1383 4353 1417
rect 4387 1383 4421 1417
rect 4455 1383 4489 1417
rect 4523 1383 4557 1417
rect 4591 1383 4625 1417
rect 4659 1383 4693 1417
rect 4727 1383 4761 1417
rect 4795 1383 4829 1417
rect 4863 1383 4897 1417
rect 4931 1383 4965 1417
rect 4999 1383 5033 1417
rect 5067 1383 5101 1417
rect 5135 1383 5169 1417
rect 5203 1383 5237 1417
rect 5271 1383 5305 1417
rect 5339 1383 5373 1417
rect 5407 1383 5441 1417
rect 5475 1383 5509 1417
rect 5543 1383 5577 1417
rect 5611 1383 5645 1417
rect 5679 1383 5713 1417
rect 5747 1383 5781 1417
rect 5815 1383 5849 1417
rect 5883 1383 5917 1417
rect 5951 1383 5985 1417
rect 6019 1383 6053 1417
rect 6087 1383 6121 1417
rect 6155 1383 6189 1417
rect 6223 1383 6257 1417
rect 6291 1383 6325 1417
rect 6359 1383 6393 1417
rect 6427 1383 6461 1417
rect 6495 1383 6529 1417
rect 6563 1383 6597 1417
rect 6631 1383 6665 1417
rect 6699 1383 6733 1417
rect 6767 1383 6801 1417
rect 6835 1383 6869 1417
rect 6903 1383 6937 1417
rect 6971 1383 7005 1417
rect 7039 1383 7073 1417
rect 7107 1383 7141 1417
rect 7175 1383 7209 1417
rect 7243 1383 7277 1417
rect 7311 1383 7345 1417
rect 7379 1383 7413 1417
rect 7447 1383 7481 1417
rect 7515 1383 7549 1417
rect 7583 1383 7617 1417
rect 7651 1383 7685 1417
rect 7719 1383 7753 1417
rect 7787 1383 7821 1417
rect 7855 1383 7889 1417
rect 7923 1383 7957 1417
rect 7991 1383 8025 1417
rect 8059 1383 8093 1417
<< poly >>
rect 520 3680 2120 3720
rect 2440 3680 4040 3720
rect 4360 3680 5960 3720
rect 6280 3680 7880 3720
rect 520 3017 2120 3080
rect 520 2983 555 3017
rect 589 2983 623 3017
rect 657 2983 691 3017
rect 725 2983 759 3017
rect 793 2983 827 3017
rect 861 2983 895 3017
rect 929 2983 963 3017
rect 997 2983 1031 3017
rect 1065 2983 1099 3017
rect 1133 2983 1167 3017
rect 1201 2983 1235 3017
rect 1269 2983 1303 3017
rect 1337 2983 1371 3017
rect 1405 2983 1439 3017
rect 1473 2983 1507 3017
rect 1541 2983 1575 3017
rect 1609 2983 1643 3017
rect 1677 2983 1711 3017
rect 1745 2983 1779 3017
rect 1813 2983 1847 3017
rect 1881 2983 1915 3017
rect 1949 2983 1983 3017
rect 2017 2983 2051 3017
rect 2085 2983 2120 3017
rect 520 2960 2120 2983
rect 2440 3017 4040 3080
rect 2440 2983 2475 3017
rect 2509 2983 2543 3017
rect 2577 2983 2611 3017
rect 2645 2983 2679 3017
rect 2713 2983 2747 3017
rect 2781 2983 2815 3017
rect 2849 2983 2883 3017
rect 2917 2983 2951 3017
rect 2985 2983 3019 3017
rect 3053 2983 3087 3017
rect 3121 2983 3155 3017
rect 3189 2983 3223 3017
rect 3257 2983 3291 3017
rect 3325 2983 3359 3017
rect 3393 2983 3427 3017
rect 3461 2983 3495 3017
rect 3529 2983 3563 3017
rect 3597 2983 3631 3017
rect 3665 2983 3699 3017
rect 3733 2983 3767 3017
rect 3801 2983 3835 3017
rect 3869 2983 3903 3017
rect 3937 2983 3971 3017
rect 4005 2983 4040 3017
rect 2440 2960 4040 2983
rect 4360 3017 5960 3080
rect 4360 2983 4395 3017
rect 4429 2983 4463 3017
rect 4497 2983 4531 3017
rect 4565 2983 4599 3017
rect 4633 2983 4667 3017
rect 4701 2983 4735 3017
rect 4769 2983 4803 3017
rect 4837 2983 4871 3017
rect 4905 2983 4939 3017
rect 4973 2983 5007 3017
rect 5041 2983 5075 3017
rect 5109 2983 5143 3017
rect 5177 2983 5211 3017
rect 5245 2983 5279 3017
rect 5313 2983 5347 3017
rect 5381 2983 5415 3017
rect 5449 2983 5483 3017
rect 5517 2983 5551 3017
rect 5585 2983 5619 3017
rect 5653 2983 5687 3017
rect 5721 2983 5755 3017
rect 5789 2983 5823 3017
rect 5857 2983 5891 3017
rect 5925 2983 5960 3017
rect 4360 2960 5960 2983
rect 6280 3017 7880 3080
rect 6280 2983 6315 3017
rect 6349 2983 6383 3017
rect 6417 2983 6451 3017
rect 6485 2983 6519 3017
rect 6553 2983 6587 3017
rect 6621 2983 6655 3017
rect 6689 2983 6723 3017
rect 6757 2983 6791 3017
rect 6825 2983 6859 3017
rect 6893 2983 6927 3017
rect 6961 2983 6995 3017
rect 7029 2983 7063 3017
rect 7097 2983 7131 3017
rect 7165 2983 7199 3017
rect 7233 2983 7267 3017
rect 7301 2983 7335 3017
rect 7369 2983 7403 3017
rect 7437 2983 7471 3017
rect 7505 2983 7539 3017
rect 7573 2983 7607 3017
rect 7641 2983 7675 3017
rect 7709 2983 7743 3017
rect 7777 2983 7811 3017
rect 7845 2983 7880 3017
rect 6280 2960 7880 2983
rect 520 2240 2120 2280
rect 2440 2240 4040 2280
rect 4360 2240 5960 2280
rect 6280 2240 7880 2280
rect 520 1577 2120 1640
rect 520 1543 555 1577
rect 589 1543 623 1577
rect 657 1543 691 1577
rect 725 1543 759 1577
rect 793 1543 827 1577
rect 861 1543 895 1577
rect 929 1543 963 1577
rect 997 1543 1031 1577
rect 1065 1543 1099 1577
rect 1133 1543 1167 1577
rect 1201 1543 1235 1577
rect 1269 1543 1303 1577
rect 1337 1543 1371 1577
rect 1405 1543 1439 1577
rect 1473 1543 1507 1577
rect 1541 1543 1575 1577
rect 1609 1543 1643 1577
rect 1677 1543 1711 1577
rect 1745 1543 1779 1577
rect 1813 1543 1847 1577
rect 1881 1543 1915 1577
rect 1949 1543 1983 1577
rect 2017 1543 2051 1577
rect 2085 1543 2120 1577
rect 520 1520 2120 1543
rect 2440 1577 4040 1640
rect 2440 1543 2475 1577
rect 2509 1543 2543 1577
rect 2577 1543 2611 1577
rect 2645 1543 2679 1577
rect 2713 1543 2747 1577
rect 2781 1543 2815 1577
rect 2849 1543 2883 1577
rect 2917 1543 2951 1577
rect 2985 1543 3019 1577
rect 3053 1543 3087 1577
rect 3121 1543 3155 1577
rect 3189 1543 3223 1577
rect 3257 1543 3291 1577
rect 3325 1543 3359 1577
rect 3393 1543 3427 1577
rect 3461 1543 3495 1577
rect 3529 1543 3563 1577
rect 3597 1543 3631 1577
rect 3665 1543 3699 1577
rect 3733 1543 3767 1577
rect 3801 1543 3835 1577
rect 3869 1543 3903 1577
rect 3937 1543 3971 1577
rect 4005 1543 4040 1577
rect 2440 1520 4040 1543
rect 4360 1577 5960 1640
rect 4360 1543 4395 1577
rect 4429 1543 4463 1577
rect 4497 1543 4531 1577
rect 4565 1543 4599 1577
rect 4633 1543 4667 1577
rect 4701 1543 4735 1577
rect 4769 1543 4803 1577
rect 4837 1543 4871 1577
rect 4905 1543 4939 1577
rect 4973 1543 5007 1577
rect 5041 1543 5075 1577
rect 5109 1543 5143 1577
rect 5177 1543 5211 1577
rect 5245 1543 5279 1577
rect 5313 1543 5347 1577
rect 5381 1543 5415 1577
rect 5449 1543 5483 1577
rect 5517 1543 5551 1577
rect 5585 1543 5619 1577
rect 5653 1543 5687 1577
rect 5721 1543 5755 1577
rect 5789 1543 5823 1577
rect 5857 1543 5891 1577
rect 5925 1543 5960 1577
rect 4360 1520 5960 1543
rect 6280 1577 7880 1640
rect 6280 1543 6315 1577
rect 6349 1543 6383 1577
rect 6417 1543 6451 1577
rect 6485 1543 6519 1577
rect 6553 1543 6587 1577
rect 6621 1543 6655 1577
rect 6689 1543 6723 1577
rect 6757 1543 6791 1577
rect 6825 1543 6859 1577
rect 6893 1543 6927 1577
rect 6961 1543 6995 1577
rect 7029 1543 7063 1577
rect 7097 1543 7131 1577
rect 7165 1543 7199 1577
rect 7233 1543 7267 1577
rect 7301 1543 7335 1577
rect 7369 1543 7403 1577
rect 7437 1543 7471 1577
rect 7505 1543 7539 1577
rect 7573 1543 7607 1577
rect 7641 1543 7675 1577
rect 7709 1543 7743 1577
rect 7777 1543 7811 1577
rect 7845 1543 7880 1577
rect 6280 1520 7880 1543
rect 520 457 2120 480
rect 520 423 555 457
rect 589 423 623 457
rect 657 423 691 457
rect 725 423 759 457
rect 793 423 827 457
rect 861 423 895 457
rect 929 423 963 457
rect 997 423 1031 457
rect 1065 423 1099 457
rect 1133 423 1167 457
rect 1201 423 1235 457
rect 1269 423 1303 457
rect 1337 423 1371 457
rect 1405 423 1439 457
rect 1473 423 1507 457
rect 1541 423 1575 457
rect 1609 423 1643 457
rect 1677 423 1711 457
rect 1745 423 1779 457
rect 1813 423 1847 457
rect 1881 423 1915 457
rect 1949 423 1983 457
rect 2017 423 2051 457
rect 2085 423 2120 457
rect 520 360 2120 423
rect 2440 457 4040 480
rect 2440 423 2475 457
rect 2509 423 2543 457
rect 2577 423 2611 457
rect 2645 423 2679 457
rect 2713 423 2747 457
rect 2781 423 2815 457
rect 2849 423 2883 457
rect 2917 423 2951 457
rect 2985 423 3019 457
rect 3053 423 3087 457
rect 3121 423 3155 457
rect 3189 423 3223 457
rect 3257 423 3291 457
rect 3325 423 3359 457
rect 3393 423 3427 457
rect 3461 423 3495 457
rect 3529 423 3563 457
rect 3597 423 3631 457
rect 3665 423 3699 457
rect 3733 423 3767 457
rect 3801 423 3835 457
rect 3869 423 3903 457
rect 3937 423 3971 457
rect 4005 423 4040 457
rect 2440 360 4040 423
rect 4360 457 5960 480
rect 4360 423 4395 457
rect 4429 423 4463 457
rect 4497 423 4531 457
rect 4565 423 4599 457
rect 4633 423 4667 457
rect 4701 423 4735 457
rect 4769 423 4803 457
rect 4837 423 4871 457
rect 4905 423 4939 457
rect 4973 423 5007 457
rect 5041 423 5075 457
rect 5109 423 5143 457
rect 5177 423 5211 457
rect 5245 423 5279 457
rect 5313 423 5347 457
rect 5381 423 5415 457
rect 5449 423 5483 457
rect 5517 423 5551 457
rect 5585 423 5619 457
rect 5653 423 5687 457
rect 5721 423 5755 457
rect 5789 423 5823 457
rect 5857 423 5891 457
rect 5925 423 5960 457
rect 4360 360 5960 423
rect 6280 457 7880 480
rect 6280 423 6315 457
rect 6349 423 6383 457
rect 6417 423 6451 457
rect 6485 423 6519 457
rect 6553 423 6587 457
rect 6621 423 6655 457
rect 6689 423 6723 457
rect 6757 423 6791 457
rect 6825 423 6859 457
rect 6893 423 6927 457
rect 6961 423 6995 457
rect 7029 423 7063 457
rect 7097 423 7131 457
rect 7165 423 7199 457
rect 7233 423 7267 457
rect 7301 423 7335 457
rect 7369 423 7403 457
rect 7437 423 7471 457
rect 7505 423 7539 457
rect 7573 423 7607 457
rect 7641 423 7675 457
rect 7709 423 7743 457
rect 7777 423 7811 457
rect 7845 423 7880 457
rect 6280 360 7880 423
rect 520 120 2120 160
rect 2440 120 4040 160
rect 4360 120 5960 160
rect 6280 120 7880 160
<< polycont >>
rect 555 2983 589 3017
rect 623 2983 657 3017
rect 691 2983 725 3017
rect 759 2983 793 3017
rect 827 2983 861 3017
rect 895 2983 929 3017
rect 963 2983 997 3017
rect 1031 2983 1065 3017
rect 1099 2983 1133 3017
rect 1167 2983 1201 3017
rect 1235 2983 1269 3017
rect 1303 2983 1337 3017
rect 1371 2983 1405 3017
rect 1439 2983 1473 3017
rect 1507 2983 1541 3017
rect 1575 2983 1609 3017
rect 1643 2983 1677 3017
rect 1711 2983 1745 3017
rect 1779 2983 1813 3017
rect 1847 2983 1881 3017
rect 1915 2983 1949 3017
rect 1983 2983 2017 3017
rect 2051 2983 2085 3017
rect 2475 2983 2509 3017
rect 2543 2983 2577 3017
rect 2611 2983 2645 3017
rect 2679 2983 2713 3017
rect 2747 2983 2781 3017
rect 2815 2983 2849 3017
rect 2883 2983 2917 3017
rect 2951 2983 2985 3017
rect 3019 2983 3053 3017
rect 3087 2983 3121 3017
rect 3155 2983 3189 3017
rect 3223 2983 3257 3017
rect 3291 2983 3325 3017
rect 3359 2983 3393 3017
rect 3427 2983 3461 3017
rect 3495 2983 3529 3017
rect 3563 2983 3597 3017
rect 3631 2983 3665 3017
rect 3699 2983 3733 3017
rect 3767 2983 3801 3017
rect 3835 2983 3869 3017
rect 3903 2983 3937 3017
rect 3971 2983 4005 3017
rect 4395 2983 4429 3017
rect 4463 2983 4497 3017
rect 4531 2983 4565 3017
rect 4599 2983 4633 3017
rect 4667 2983 4701 3017
rect 4735 2983 4769 3017
rect 4803 2983 4837 3017
rect 4871 2983 4905 3017
rect 4939 2983 4973 3017
rect 5007 2983 5041 3017
rect 5075 2983 5109 3017
rect 5143 2983 5177 3017
rect 5211 2983 5245 3017
rect 5279 2983 5313 3017
rect 5347 2983 5381 3017
rect 5415 2983 5449 3017
rect 5483 2983 5517 3017
rect 5551 2983 5585 3017
rect 5619 2983 5653 3017
rect 5687 2983 5721 3017
rect 5755 2983 5789 3017
rect 5823 2983 5857 3017
rect 5891 2983 5925 3017
rect 6315 2983 6349 3017
rect 6383 2983 6417 3017
rect 6451 2983 6485 3017
rect 6519 2983 6553 3017
rect 6587 2983 6621 3017
rect 6655 2983 6689 3017
rect 6723 2983 6757 3017
rect 6791 2983 6825 3017
rect 6859 2983 6893 3017
rect 6927 2983 6961 3017
rect 6995 2983 7029 3017
rect 7063 2983 7097 3017
rect 7131 2983 7165 3017
rect 7199 2983 7233 3017
rect 7267 2983 7301 3017
rect 7335 2983 7369 3017
rect 7403 2983 7437 3017
rect 7471 2983 7505 3017
rect 7539 2983 7573 3017
rect 7607 2983 7641 3017
rect 7675 2983 7709 3017
rect 7743 2983 7777 3017
rect 7811 2983 7845 3017
rect 555 1543 589 1577
rect 623 1543 657 1577
rect 691 1543 725 1577
rect 759 1543 793 1577
rect 827 1543 861 1577
rect 895 1543 929 1577
rect 963 1543 997 1577
rect 1031 1543 1065 1577
rect 1099 1543 1133 1577
rect 1167 1543 1201 1577
rect 1235 1543 1269 1577
rect 1303 1543 1337 1577
rect 1371 1543 1405 1577
rect 1439 1543 1473 1577
rect 1507 1543 1541 1577
rect 1575 1543 1609 1577
rect 1643 1543 1677 1577
rect 1711 1543 1745 1577
rect 1779 1543 1813 1577
rect 1847 1543 1881 1577
rect 1915 1543 1949 1577
rect 1983 1543 2017 1577
rect 2051 1543 2085 1577
rect 2475 1543 2509 1577
rect 2543 1543 2577 1577
rect 2611 1543 2645 1577
rect 2679 1543 2713 1577
rect 2747 1543 2781 1577
rect 2815 1543 2849 1577
rect 2883 1543 2917 1577
rect 2951 1543 2985 1577
rect 3019 1543 3053 1577
rect 3087 1543 3121 1577
rect 3155 1543 3189 1577
rect 3223 1543 3257 1577
rect 3291 1543 3325 1577
rect 3359 1543 3393 1577
rect 3427 1543 3461 1577
rect 3495 1543 3529 1577
rect 3563 1543 3597 1577
rect 3631 1543 3665 1577
rect 3699 1543 3733 1577
rect 3767 1543 3801 1577
rect 3835 1543 3869 1577
rect 3903 1543 3937 1577
rect 3971 1543 4005 1577
rect 4395 1543 4429 1577
rect 4463 1543 4497 1577
rect 4531 1543 4565 1577
rect 4599 1543 4633 1577
rect 4667 1543 4701 1577
rect 4735 1543 4769 1577
rect 4803 1543 4837 1577
rect 4871 1543 4905 1577
rect 4939 1543 4973 1577
rect 5007 1543 5041 1577
rect 5075 1543 5109 1577
rect 5143 1543 5177 1577
rect 5211 1543 5245 1577
rect 5279 1543 5313 1577
rect 5347 1543 5381 1577
rect 5415 1543 5449 1577
rect 5483 1543 5517 1577
rect 5551 1543 5585 1577
rect 5619 1543 5653 1577
rect 5687 1543 5721 1577
rect 5755 1543 5789 1577
rect 5823 1543 5857 1577
rect 5891 1543 5925 1577
rect 6315 1543 6349 1577
rect 6383 1543 6417 1577
rect 6451 1543 6485 1577
rect 6519 1543 6553 1577
rect 6587 1543 6621 1577
rect 6655 1543 6689 1577
rect 6723 1543 6757 1577
rect 6791 1543 6825 1577
rect 6859 1543 6893 1577
rect 6927 1543 6961 1577
rect 6995 1543 7029 1577
rect 7063 1543 7097 1577
rect 7131 1543 7165 1577
rect 7199 1543 7233 1577
rect 7267 1543 7301 1577
rect 7335 1543 7369 1577
rect 7403 1543 7437 1577
rect 7471 1543 7505 1577
rect 7539 1543 7573 1577
rect 7607 1543 7641 1577
rect 7675 1543 7709 1577
rect 7743 1543 7777 1577
rect 7811 1543 7845 1577
rect 555 423 589 457
rect 623 423 657 457
rect 691 423 725 457
rect 759 423 793 457
rect 827 423 861 457
rect 895 423 929 457
rect 963 423 997 457
rect 1031 423 1065 457
rect 1099 423 1133 457
rect 1167 423 1201 457
rect 1235 423 1269 457
rect 1303 423 1337 457
rect 1371 423 1405 457
rect 1439 423 1473 457
rect 1507 423 1541 457
rect 1575 423 1609 457
rect 1643 423 1677 457
rect 1711 423 1745 457
rect 1779 423 1813 457
rect 1847 423 1881 457
rect 1915 423 1949 457
rect 1983 423 2017 457
rect 2051 423 2085 457
rect 2475 423 2509 457
rect 2543 423 2577 457
rect 2611 423 2645 457
rect 2679 423 2713 457
rect 2747 423 2781 457
rect 2815 423 2849 457
rect 2883 423 2917 457
rect 2951 423 2985 457
rect 3019 423 3053 457
rect 3087 423 3121 457
rect 3155 423 3189 457
rect 3223 423 3257 457
rect 3291 423 3325 457
rect 3359 423 3393 457
rect 3427 423 3461 457
rect 3495 423 3529 457
rect 3563 423 3597 457
rect 3631 423 3665 457
rect 3699 423 3733 457
rect 3767 423 3801 457
rect 3835 423 3869 457
rect 3903 423 3937 457
rect 3971 423 4005 457
rect 4395 423 4429 457
rect 4463 423 4497 457
rect 4531 423 4565 457
rect 4599 423 4633 457
rect 4667 423 4701 457
rect 4735 423 4769 457
rect 4803 423 4837 457
rect 4871 423 4905 457
rect 4939 423 4973 457
rect 5007 423 5041 457
rect 5075 423 5109 457
rect 5143 423 5177 457
rect 5211 423 5245 457
rect 5279 423 5313 457
rect 5347 423 5381 457
rect 5415 423 5449 457
rect 5483 423 5517 457
rect 5551 423 5585 457
rect 5619 423 5653 457
rect 5687 423 5721 457
rect 5755 423 5789 457
rect 5823 423 5857 457
rect 5891 423 5925 457
rect 6315 423 6349 457
rect 6383 423 6417 457
rect 6451 423 6485 457
rect 6519 423 6553 457
rect 6587 423 6621 457
rect 6655 423 6689 457
rect 6723 423 6757 457
rect 6791 423 6825 457
rect 6859 423 6893 457
rect 6927 423 6961 457
rect 6995 423 7029 457
rect 7063 423 7097 457
rect 7131 423 7165 457
rect 7199 423 7233 457
rect 7267 423 7301 457
rect 7335 423 7369 457
rect 7403 423 7437 457
rect 7471 423 7505 457
rect 7539 423 7573 457
rect 7607 423 7641 457
rect 7675 423 7709 457
rect 7743 423 7777 457
rect 7811 423 7845 457
<< locali >>
rect 0 3977 8400 4000
rect 0 3943 137 3977
rect 171 3943 205 3977
rect 239 3943 273 3977
rect 307 3943 341 3977
rect 375 3943 409 3977
rect 443 3943 477 3977
rect 511 3943 545 3977
rect 579 3943 613 3977
rect 647 3943 681 3977
rect 715 3943 749 3977
rect 783 3943 817 3977
rect 851 3943 885 3977
rect 919 3943 953 3977
rect 987 3943 1021 3977
rect 1055 3943 1089 3977
rect 1123 3943 1157 3977
rect 1191 3943 1225 3977
rect 1259 3943 1293 3977
rect 1327 3943 1361 3977
rect 1395 3943 1429 3977
rect 1463 3943 1497 3977
rect 1531 3943 1565 3977
rect 1599 3943 1633 3977
rect 1667 3943 1701 3977
rect 1735 3943 1769 3977
rect 1803 3943 1837 3977
rect 1871 3943 1905 3977
rect 1939 3943 1973 3977
rect 2007 3943 2041 3977
rect 2075 3943 2109 3977
rect 2143 3943 2177 3977
rect 2211 3943 2245 3977
rect 2279 3943 2313 3977
rect 2347 3943 2381 3977
rect 2415 3943 2449 3977
rect 2483 3943 2517 3977
rect 2551 3943 2585 3977
rect 2619 3943 2653 3977
rect 2687 3943 2721 3977
rect 2755 3943 2789 3977
rect 2823 3943 2857 3977
rect 2891 3943 2925 3977
rect 2959 3943 2993 3977
rect 3027 3943 3061 3977
rect 3095 3943 3129 3977
rect 3163 3943 3197 3977
rect 3231 3943 3265 3977
rect 3299 3943 3333 3977
rect 3367 3943 3401 3977
rect 3435 3943 3469 3977
rect 3503 3943 3537 3977
rect 3571 3943 3605 3977
rect 3639 3943 3673 3977
rect 3707 3943 3741 3977
rect 3775 3943 3809 3977
rect 3843 3943 3877 3977
rect 3911 3943 3945 3977
rect 3979 3943 4013 3977
rect 4047 3943 4081 3977
rect 4115 3943 4149 3977
rect 4183 3943 4217 3977
rect 4251 3943 4285 3977
rect 4319 3943 4353 3977
rect 4387 3943 4421 3977
rect 4455 3943 4489 3977
rect 4523 3943 4557 3977
rect 4591 3943 4625 3977
rect 4659 3943 4693 3977
rect 4727 3943 4761 3977
rect 4795 3943 4829 3977
rect 4863 3943 4897 3977
rect 4931 3943 4965 3977
rect 4999 3943 5033 3977
rect 5067 3943 5101 3977
rect 5135 3943 5169 3977
rect 5203 3943 5237 3977
rect 5271 3943 5305 3977
rect 5339 3943 5373 3977
rect 5407 3943 5441 3977
rect 5475 3943 5509 3977
rect 5543 3943 5577 3977
rect 5611 3943 5645 3977
rect 5679 3943 5713 3977
rect 5747 3943 5781 3977
rect 5815 3943 5849 3977
rect 5883 3943 5917 3977
rect 5951 3943 5985 3977
rect 6019 3943 6053 3977
rect 6087 3943 6121 3977
rect 6155 3943 6189 3977
rect 6223 3943 6257 3977
rect 6291 3943 6325 3977
rect 6359 3943 6393 3977
rect 6427 3943 6461 3977
rect 6495 3943 6529 3977
rect 6563 3943 6597 3977
rect 6631 3943 6665 3977
rect 6699 3943 6733 3977
rect 6767 3943 6801 3977
rect 6835 3943 6869 3977
rect 6903 3943 6937 3977
rect 6971 3943 7005 3977
rect 7039 3943 7073 3977
rect 7107 3943 7141 3977
rect 7175 3943 7209 3977
rect 7243 3943 7277 3977
rect 7311 3943 7345 3977
rect 7379 3943 7413 3977
rect 7447 3943 7481 3977
rect 7515 3943 7549 3977
rect 7583 3943 7617 3977
rect 7651 3943 7685 3977
rect 7719 3943 7753 3977
rect 7787 3943 7821 3977
rect 7855 3943 7889 3977
rect 7923 3943 7957 3977
rect 7991 3943 8025 3977
rect 8059 3943 8093 3977
rect 8127 3943 8161 3977
rect 8195 3943 8229 3977
rect 8263 3943 8400 3977
rect 0 3920 8400 3943
rect 0 3847 80 3920
rect 0 3813 23 3847
rect 57 3813 80 3847
rect 8320 3847 8400 3920
rect 0 3779 80 3813
rect 0 3745 23 3779
rect 57 3745 80 3779
rect 0 3711 80 3745
rect 0 3677 23 3711
rect 57 3677 80 3711
rect 0 3643 80 3677
rect 0 3609 23 3643
rect 57 3609 80 3643
rect 0 3575 80 3609
rect 0 3541 23 3575
rect 57 3541 80 3575
rect 0 3507 80 3541
rect 0 3473 23 3507
rect 57 3473 80 3507
rect 0 3439 80 3473
rect 0 3405 23 3439
rect 57 3405 80 3439
rect 0 3371 80 3405
rect 0 3337 23 3371
rect 57 3337 80 3371
rect 0 3303 80 3337
rect 0 3269 23 3303
rect 57 3269 80 3303
rect 0 3235 80 3269
rect 0 3201 23 3235
rect 57 3201 80 3235
rect 0 3167 80 3201
rect 0 3133 23 3167
rect 57 3133 80 3167
rect 0 3099 80 3133
rect 0 3065 23 3099
rect 57 3065 80 3099
rect 0 3031 80 3065
rect 0 2997 23 3031
rect 57 2997 80 3031
rect 0 2963 80 2997
rect 0 2929 23 2963
rect 57 2929 80 2963
rect 0 2895 80 2929
rect 0 2861 23 2895
rect 57 2861 80 2895
rect 0 2827 80 2861
rect 0 2793 23 2827
rect 57 2793 80 2827
rect 160 3817 8240 3840
rect 160 3783 307 3817
rect 341 3783 375 3817
rect 409 3783 443 3817
rect 477 3783 511 3817
rect 545 3783 579 3817
rect 613 3783 647 3817
rect 681 3783 715 3817
rect 749 3783 783 3817
rect 817 3783 851 3817
rect 885 3783 919 3817
rect 953 3783 987 3817
rect 1021 3783 1055 3817
rect 1089 3783 1123 3817
rect 1157 3783 1191 3817
rect 1225 3783 1259 3817
rect 1293 3783 1327 3817
rect 1361 3783 1395 3817
rect 1429 3783 1463 3817
rect 1497 3783 1531 3817
rect 1565 3783 1599 3817
rect 1633 3783 1667 3817
rect 1701 3783 1735 3817
rect 1769 3783 1803 3817
rect 1837 3783 1871 3817
rect 1905 3783 1939 3817
rect 1973 3783 2007 3817
rect 2041 3783 2075 3817
rect 2109 3783 2143 3817
rect 2177 3783 2211 3817
rect 2245 3783 2279 3817
rect 2313 3783 2347 3817
rect 2381 3783 2415 3817
rect 2449 3783 2483 3817
rect 2517 3783 2551 3817
rect 2585 3783 2619 3817
rect 2653 3783 2687 3817
rect 2721 3783 2755 3817
rect 2789 3783 2823 3817
rect 2857 3783 2891 3817
rect 2925 3783 2959 3817
rect 2993 3783 3027 3817
rect 3061 3783 3095 3817
rect 3129 3783 3163 3817
rect 3197 3783 3231 3817
rect 3265 3783 3299 3817
rect 3333 3783 3367 3817
rect 3401 3783 3435 3817
rect 3469 3783 3503 3817
rect 3537 3783 3571 3817
rect 3605 3783 3639 3817
rect 3673 3783 3707 3817
rect 3741 3783 3775 3817
rect 3809 3783 3843 3817
rect 3877 3783 3911 3817
rect 3945 3783 3979 3817
rect 4013 3783 4047 3817
rect 4081 3783 4115 3817
rect 4149 3783 4183 3817
rect 4217 3783 4251 3817
rect 4285 3783 4319 3817
rect 4353 3783 4387 3817
rect 4421 3783 4455 3817
rect 4489 3783 4523 3817
rect 4557 3783 4591 3817
rect 4625 3783 4659 3817
rect 4693 3783 4727 3817
rect 4761 3783 4795 3817
rect 4829 3783 4863 3817
rect 4897 3783 4931 3817
rect 4965 3783 4999 3817
rect 5033 3783 5067 3817
rect 5101 3783 5135 3817
rect 5169 3783 5203 3817
rect 5237 3783 5271 3817
rect 5305 3783 5339 3817
rect 5373 3783 5407 3817
rect 5441 3783 5475 3817
rect 5509 3783 5543 3817
rect 5577 3783 5611 3817
rect 5645 3783 5679 3817
rect 5713 3783 5747 3817
rect 5781 3783 5815 3817
rect 5849 3783 5883 3817
rect 5917 3783 5951 3817
rect 5985 3783 6019 3817
rect 6053 3783 6087 3817
rect 6121 3783 6155 3817
rect 6189 3783 6223 3817
rect 6257 3783 6291 3817
rect 6325 3783 6359 3817
rect 6393 3783 6427 3817
rect 6461 3783 6495 3817
rect 6529 3783 6563 3817
rect 6597 3783 6631 3817
rect 6665 3783 6699 3817
rect 6733 3783 6767 3817
rect 6801 3783 6835 3817
rect 6869 3783 6903 3817
rect 6937 3783 6971 3817
rect 7005 3783 7039 3817
rect 7073 3783 7107 3817
rect 7141 3783 7175 3817
rect 7209 3783 7243 3817
rect 7277 3783 7311 3817
rect 7345 3783 7379 3817
rect 7413 3783 7447 3817
rect 7481 3783 7515 3817
rect 7549 3783 7583 3817
rect 7617 3783 7651 3817
rect 7685 3783 7719 3817
rect 7753 3783 7787 3817
rect 7821 3783 7855 3817
rect 7889 3783 7923 3817
rect 7957 3783 7991 3817
rect 8025 3783 8059 3817
rect 8093 3783 8240 3817
rect 160 3760 8240 3783
rect 160 3711 240 3760
rect 160 3677 183 3711
rect 217 3677 240 3711
rect 160 3643 240 3677
rect 160 3609 183 3643
rect 217 3609 240 3643
rect 160 3575 240 3609
rect 160 3541 183 3575
rect 217 3541 240 3575
rect 160 3507 240 3541
rect 160 3473 183 3507
rect 217 3473 240 3507
rect 160 3439 240 3473
rect 160 3405 183 3439
rect 217 3405 240 3439
rect 160 3371 240 3405
rect 160 3337 183 3371
rect 217 3337 240 3371
rect 160 3303 240 3337
rect 160 3269 183 3303
rect 217 3269 240 3303
rect 160 3235 240 3269
rect 160 3201 183 3235
rect 217 3201 240 3235
rect 160 3167 240 3201
rect 160 3133 183 3167
rect 217 3133 240 3167
rect 160 3099 240 3133
rect 160 3065 183 3099
rect 217 3065 240 3099
rect 320 3649 400 3680
rect 320 3601 343 3649
rect 377 3601 400 3649
rect 320 3577 400 3601
rect 320 3533 343 3577
rect 377 3533 400 3577
rect 320 3505 400 3533
rect 320 3465 343 3505
rect 377 3465 400 3505
rect 320 3433 400 3465
rect 320 3397 343 3433
rect 377 3397 400 3433
rect 320 3363 400 3397
rect 320 3327 343 3363
rect 377 3327 400 3363
rect 320 3295 400 3327
rect 320 3255 343 3295
rect 377 3255 400 3295
rect 320 3227 400 3255
rect 320 3183 343 3227
rect 377 3183 400 3227
rect 320 3159 400 3183
rect 320 3111 343 3159
rect 377 3111 400 3159
rect 320 3080 400 3111
rect 2240 3649 2320 3680
rect 2240 3601 2263 3649
rect 2297 3601 2320 3649
rect 2240 3577 2320 3601
rect 2240 3533 2263 3577
rect 2297 3533 2320 3577
rect 2240 3505 2320 3533
rect 2240 3465 2263 3505
rect 2297 3465 2320 3505
rect 2240 3433 2320 3465
rect 2240 3397 2263 3433
rect 2297 3397 2320 3433
rect 2240 3363 2320 3397
rect 2240 3327 2263 3363
rect 2297 3327 2320 3363
rect 2240 3295 2320 3327
rect 2240 3255 2263 3295
rect 2297 3255 2320 3295
rect 2240 3227 2320 3255
rect 2240 3183 2263 3227
rect 2297 3183 2320 3227
rect 2240 3159 2320 3183
rect 2240 3111 2263 3159
rect 2297 3111 2320 3159
rect 2240 3080 2320 3111
rect 4160 3649 4240 3760
rect 8160 3711 8240 3760
rect 4160 3601 4183 3649
rect 4217 3601 4240 3649
rect 4160 3577 4240 3601
rect 4160 3533 4183 3577
rect 4217 3533 4240 3577
rect 4160 3505 4240 3533
rect 4160 3465 4183 3505
rect 4217 3465 4240 3505
rect 4160 3433 4240 3465
rect 4160 3397 4183 3433
rect 4217 3397 4240 3433
rect 4160 3363 4240 3397
rect 4160 3327 4183 3363
rect 4217 3327 4240 3363
rect 4160 3295 4240 3327
rect 4160 3255 4183 3295
rect 4217 3255 4240 3295
rect 4160 3227 4240 3255
rect 4160 3183 4183 3227
rect 4217 3183 4240 3227
rect 4160 3159 4240 3183
rect 4160 3111 4183 3159
rect 4217 3111 4240 3159
rect 4160 3080 4240 3111
rect 6080 3649 6160 3680
rect 6080 3601 6103 3649
rect 6137 3601 6160 3649
rect 6080 3577 6160 3601
rect 6080 3533 6103 3577
rect 6137 3533 6160 3577
rect 6080 3505 6160 3533
rect 6080 3465 6103 3505
rect 6137 3465 6160 3505
rect 6080 3433 6160 3465
rect 6080 3397 6103 3433
rect 6137 3397 6160 3433
rect 6080 3363 6160 3397
rect 6080 3327 6103 3363
rect 6137 3327 6160 3363
rect 6080 3295 6160 3327
rect 6080 3255 6103 3295
rect 6137 3255 6160 3295
rect 6080 3227 6160 3255
rect 6080 3183 6103 3227
rect 6137 3183 6160 3227
rect 6080 3159 6160 3183
rect 6080 3111 6103 3159
rect 6137 3111 6160 3159
rect 6080 3080 6160 3111
rect 8000 3649 8080 3680
rect 8000 3601 8023 3649
rect 8057 3601 8080 3649
rect 8000 3577 8080 3601
rect 8000 3533 8023 3577
rect 8057 3533 8080 3577
rect 8000 3505 8080 3533
rect 8000 3465 8023 3505
rect 8057 3465 8080 3505
rect 8000 3433 8080 3465
rect 8000 3397 8023 3433
rect 8057 3397 8080 3433
rect 8000 3363 8080 3397
rect 8000 3327 8023 3363
rect 8057 3327 8080 3363
rect 8000 3295 8080 3327
rect 8000 3255 8023 3295
rect 8057 3255 8080 3295
rect 8000 3227 8080 3255
rect 8000 3183 8023 3227
rect 8057 3183 8080 3227
rect 8000 3159 8080 3183
rect 8000 3111 8023 3159
rect 8057 3111 8080 3159
rect 8000 3080 8080 3111
rect 8160 3677 8183 3711
rect 8217 3677 8240 3711
rect 8160 3643 8240 3677
rect 8160 3609 8183 3643
rect 8217 3609 8240 3643
rect 8160 3575 8240 3609
rect 8160 3541 8183 3575
rect 8217 3541 8240 3575
rect 8160 3507 8240 3541
rect 8160 3473 8183 3507
rect 8217 3473 8240 3507
rect 8160 3439 8240 3473
rect 8160 3405 8183 3439
rect 8217 3405 8240 3439
rect 8160 3371 8240 3405
rect 8160 3337 8183 3371
rect 8217 3337 8240 3371
rect 8160 3303 8240 3337
rect 8160 3269 8183 3303
rect 8217 3269 8240 3303
rect 8160 3235 8240 3269
rect 8160 3201 8183 3235
rect 8217 3201 8240 3235
rect 8160 3167 8240 3201
rect 8160 3133 8183 3167
rect 8217 3133 8240 3167
rect 8160 3099 8240 3133
rect 160 3031 240 3065
rect 8160 3065 8183 3099
rect 8217 3065 8240 3099
rect 160 2997 183 3031
rect 217 2997 240 3031
rect 160 2963 240 2997
rect 160 2929 183 2963
rect 217 2929 240 2963
rect 520 3017 2120 3040
rect 520 2983 547 3017
rect 589 2983 619 3017
rect 657 2983 691 3017
rect 725 2983 759 3017
rect 797 2983 827 3017
rect 869 2983 895 3017
rect 941 2983 963 3017
rect 1013 2983 1031 3017
rect 1085 2983 1099 3017
rect 1157 2983 1167 3017
rect 1229 2983 1235 3017
rect 1301 2983 1303 3017
rect 1337 2983 1339 3017
rect 1405 2983 1411 3017
rect 1473 2983 1483 3017
rect 1541 2983 1555 3017
rect 1609 2983 1627 3017
rect 1677 2983 1699 3017
rect 1745 2983 1771 3017
rect 1813 2983 1843 3017
rect 1881 2983 1915 3017
rect 1949 2983 1983 3017
rect 2021 2983 2051 3017
rect 2093 2983 2120 3017
rect 520 2960 2120 2983
rect 2440 3017 4040 3040
rect 2440 2983 2467 3017
rect 2509 2983 2539 3017
rect 2577 2983 2611 3017
rect 2645 2983 2679 3017
rect 2717 2983 2747 3017
rect 2789 2983 2815 3017
rect 2861 2983 2883 3017
rect 2933 2983 2951 3017
rect 3005 2983 3019 3017
rect 3077 2983 3087 3017
rect 3149 2983 3155 3017
rect 3221 2983 3223 3017
rect 3257 2983 3259 3017
rect 3325 2983 3331 3017
rect 3393 2983 3403 3017
rect 3461 2983 3475 3017
rect 3529 2983 3547 3017
rect 3597 2983 3619 3017
rect 3665 2983 3691 3017
rect 3733 2983 3763 3017
rect 3801 2983 3835 3017
rect 3869 2983 3903 3017
rect 3941 2983 3971 3017
rect 4013 2983 4040 3017
rect 2440 2960 4040 2983
rect 4360 3017 5960 3040
rect 4360 2983 4387 3017
rect 4429 2983 4459 3017
rect 4497 2983 4531 3017
rect 4565 2983 4599 3017
rect 4637 2983 4667 3017
rect 4709 2983 4735 3017
rect 4781 2983 4803 3017
rect 4853 2983 4871 3017
rect 4925 2983 4939 3017
rect 4997 2983 5007 3017
rect 5069 2983 5075 3017
rect 5141 2983 5143 3017
rect 5177 2983 5179 3017
rect 5245 2983 5251 3017
rect 5313 2983 5323 3017
rect 5381 2983 5395 3017
rect 5449 2983 5467 3017
rect 5517 2983 5539 3017
rect 5585 2983 5611 3017
rect 5653 2983 5683 3017
rect 5721 2983 5755 3017
rect 5789 2983 5823 3017
rect 5861 2983 5891 3017
rect 5933 2983 5960 3017
rect 4360 2960 5960 2983
rect 6280 3017 7880 3040
rect 6280 2983 6307 3017
rect 6349 2983 6379 3017
rect 6417 2983 6451 3017
rect 6485 2983 6519 3017
rect 6557 2983 6587 3017
rect 6629 2983 6655 3017
rect 6701 2983 6723 3017
rect 6773 2983 6791 3017
rect 6845 2983 6859 3017
rect 6917 2983 6927 3017
rect 6989 2983 6995 3017
rect 7061 2983 7063 3017
rect 7097 2983 7099 3017
rect 7165 2983 7171 3017
rect 7233 2983 7243 3017
rect 7301 2983 7315 3017
rect 7369 2983 7387 3017
rect 7437 2983 7459 3017
rect 7505 2983 7531 3017
rect 7573 2983 7603 3017
rect 7641 2983 7675 3017
rect 7709 2983 7743 3017
rect 7781 2983 7811 3017
rect 7853 2983 7880 3017
rect 6280 2960 7880 2983
rect 8160 3031 8240 3065
rect 8160 2997 8183 3031
rect 8217 2997 8240 3031
rect 8160 2963 8240 2997
rect 160 2880 240 2929
rect 8160 2929 8183 2963
rect 8217 2929 8240 2963
rect 8160 2880 8240 2929
rect 160 2857 8240 2880
rect 160 2823 307 2857
rect 341 2823 375 2857
rect 409 2823 443 2857
rect 477 2823 511 2857
rect 545 2823 579 2857
rect 613 2823 647 2857
rect 681 2823 715 2857
rect 749 2823 783 2857
rect 817 2823 851 2857
rect 885 2823 919 2857
rect 953 2823 987 2857
rect 1021 2823 1055 2857
rect 1089 2823 1123 2857
rect 1157 2823 1191 2857
rect 1225 2823 1259 2857
rect 1293 2823 1327 2857
rect 1361 2823 1395 2857
rect 1429 2823 1463 2857
rect 1497 2823 1531 2857
rect 1565 2823 1599 2857
rect 1633 2823 1667 2857
rect 1701 2823 1735 2857
rect 1769 2823 1803 2857
rect 1837 2823 1871 2857
rect 1905 2823 1939 2857
rect 1973 2823 2007 2857
rect 2041 2823 2075 2857
rect 2109 2823 2143 2857
rect 2177 2823 2211 2857
rect 2245 2823 2279 2857
rect 2313 2823 2347 2857
rect 2381 2823 2415 2857
rect 2449 2823 2483 2857
rect 2517 2823 2551 2857
rect 2585 2823 2619 2857
rect 2653 2823 2687 2857
rect 2721 2823 2755 2857
rect 2789 2823 2823 2857
rect 2857 2823 2891 2857
rect 2925 2823 2959 2857
rect 2993 2823 3027 2857
rect 3061 2823 3095 2857
rect 3129 2823 3163 2857
rect 3197 2823 3231 2857
rect 3265 2823 3299 2857
rect 3333 2823 3367 2857
rect 3401 2823 3435 2857
rect 3469 2823 3503 2857
rect 3537 2823 3571 2857
rect 3605 2823 3639 2857
rect 3673 2823 3707 2857
rect 3741 2823 3775 2857
rect 3809 2823 3843 2857
rect 3877 2823 3911 2857
rect 3945 2823 3979 2857
rect 4013 2823 4047 2857
rect 4081 2823 4115 2857
rect 4149 2823 4183 2857
rect 4217 2823 4251 2857
rect 4285 2823 4319 2857
rect 4353 2823 4387 2857
rect 4421 2823 4455 2857
rect 4489 2823 4523 2857
rect 4557 2823 4591 2857
rect 4625 2823 4659 2857
rect 4693 2823 4727 2857
rect 4761 2823 4795 2857
rect 4829 2823 4863 2857
rect 4897 2823 4931 2857
rect 4965 2823 4999 2857
rect 5033 2823 5067 2857
rect 5101 2823 5135 2857
rect 5169 2823 5203 2857
rect 5237 2823 5271 2857
rect 5305 2823 5339 2857
rect 5373 2823 5407 2857
rect 5441 2823 5475 2857
rect 5509 2823 5543 2857
rect 5577 2823 5611 2857
rect 5645 2823 5679 2857
rect 5713 2823 5747 2857
rect 5781 2823 5815 2857
rect 5849 2823 5883 2857
rect 5917 2823 5951 2857
rect 5985 2823 6019 2857
rect 6053 2823 6087 2857
rect 6121 2823 6155 2857
rect 6189 2823 6223 2857
rect 6257 2823 6291 2857
rect 6325 2823 6359 2857
rect 6393 2823 6427 2857
rect 6461 2823 6495 2857
rect 6529 2823 6563 2857
rect 6597 2823 6631 2857
rect 6665 2823 6699 2857
rect 6733 2823 6767 2857
rect 6801 2823 6835 2857
rect 6869 2823 6903 2857
rect 6937 2823 6971 2857
rect 7005 2823 7039 2857
rect 7073 2823 7107 2857
rect 7141 2823 7175 2857
rect 7209 2823 7243 2857
rect 7277 2823 7311 2857
rect 7345 2823 7379 2857
rect 7413 2823 7447 2857
rect 7481 2823 7515 2857
rect 7549 2823 7583 2857
rect 7617 2823 7651 2857
rect 7685 2823 7719 2857
rect 7753 2823 7787 2857
rect 7821 2823 7855 2857
rect 7889 2823 7923 2857
rect 7957 2823 7991 2857
rect 8025 2823 8059 2857
rect 8093 2823 8240 2857
rect 160 2800 8240 2823
rect 8320 3813 8343 3847
rect 8377 3813 8400 3847
rect 8320 3779 8400 3813
rect 8320 3745 8343 3779
rect 8377 3745 8400 3779
rect 8320 3711 8400 3745
rect 8320 3677 8343 3711
rect 8377 3677 8400 3711
rect 8320 3643 8400 3677
rect 8320 3609 8343 3643
rect 8377 3609 8400 3643
rect 8320 3575 8400 3609
rect 8320 3541 8343 3575
rect 8377 3541 8400 3575
rect 8320 3507 8400 3541
rect 8320 3473 8343 3507
rect 8377 3473 8400 3507
rect 8320 3439 8400 3473
rect 8320 3405 8343 3439
rect 8377 3405 8400 3439
rect 8320 3371 8400 3405
rect 8320 3337 8343 3371
rect 8377 3337 8400 3371
rect 8320 3303 8400 3337
rect 8320 3269 8343 3303
rect 8377 3269 8400 3303
rect 8320 3235 8400 3269
rect 8320 3201 8343 3235
rect 8377 3201 8400 3235
rect 8320 3167 8400 3201
rect 8320 3133 8343 3167
rect 8377 3133 8400 3167
rect 8320 3099 8400 3133
rect 8320 3065 8343 3099
rect 8377 3065 8400 3099
rect 8320 3031 8400 3065
rect 8320 2997 8343 3031
rect 8377 2997 8400 3031
rect 8320 2963 8400 2997
rect 8320 2929 8343 2963
rect 8377 2929 8400 2963
rect 8320 2895 8400 2929
rect 8320 2861 8343 2895
rect 8377 2861 8400 2895
rect 8320 2827 8400 2861
rect 0 2720 80 2793
rect 8320 2793 8343 2827
rect 8377 2793 8400 2827
rect 8320 2720 8400 2793
rect 0 2697 8400 2720
rect 0 2663 151 2697
rect 185 2663 219 2697
rect 253 2663 287 2697
rect 321 2663 355 2697
rect 389 2663 423 2697
rect 457 2663 491 2697
rect 525 2663 559 2697
rect 593 2663 627 2697
rect 661 2663 695 2697
rect 729 2663 763 2697
rect 797 2663 831 2697
rect 865 2663 899 2697
rect 933 2663 967 2697
rect 1001 2663 1035 2697
rect 1069 2663 1103 2697
rect 1137 2663 1171 2697
rect 1205 2663 1239 2697
rect 1273 2663 1307 2697
rect 1341 2663 1375 2697
rect 1409 2663 1443 2697
rect 1477 2663 1511 2697
rect 1545 2663 1579 2697
rect 1613 2663 1647 2697
rect 1681 2663 1715 2697
rect 1749 2663 1783 2697
rect 1817 2663 1851 2697
rect 1885 2663 1919 2697
rect 1953 2663 1987 2697
rect 2021 2663 2055 2697
rect 2089 2663 2123 2697
rect 2157 2663 2191 2697
rect 2225 2663 2259 2697
rect 2293 2663 2327 2697
rect 2361 2663 2395 2697
rect 2429 2663 2463 2697
rect 2497 2663 2531 2697
rect 2565 2663 2599 2697
rect 2633 2663 2667 2697
rect 2701 2663 2735 2697
rect 2769 2663 2803 2697
rect 2837 2663 2871 2697
rect 2905 2663 2939 2697
rect 2973 2663 3007 2697
rect 3041 2663 3075 2697
rect 3109 2663 3143 2697
rect 3177 2663 3211 2697
rect 3245 2663 3279 2697
rect 3313 2663 3347 2697
rect 3381 2663 3415 2697
rect 3449 2663 3483 2697
rect 3517 2663 3551 2697
rect 3585 2663 3619 2697
rect 3653 2663 3687 2697
rect 3721 2663 3755 2697
rect 3789 2663 3823 2697
rect 3857 2663 3891 2697
rect 3925 2663 3959 2697
rect 3993 2663 4027 2697
rect 4061 2663 4095 2697
rect 4129 2663 4163 2697
rect 4197 2663 4231 2697
rect 4265 2663 4299 2697
rect 4333 2663 4367 2697
rect 4401 2663 4435 2697
rect 4469 2663 4503 2697
rect 4537 2663 4571 2697
rect 4605 2663 4639 2697
rect 4673 2663 4707 2697
rect 4741 2663 4775 2697
rect 4809 2663 4843 2697
rect 4877 2663 4911 2697
rect 4945 2663 4979 2697
rect 5013 2663 5047 2697
rect 5081 2663 5115 2697
rect 5149 2663 5183 2697
rect 5217 2663 5251 2697
rect 5285 2663 5319 2697
rect 5353 2663 5387 2697
rect 5421 2663 5455 2697
rect 5489 2663 5523 2697
rect 5557 2663 5591 2697
rect 5625 2663 5659 2697
rect 5693 2663 5727 2697
rect 5761 2663 5795 2697
rect 5829 2663 5863 2697
rect 5897 2663 5931 2697
rect 5965 2663 5999 2697
rect 6033 2663 6067 2697
rect 6101 2663 6135 2697
rect 6169 2663 6203 2697
rect 6237 2663 6271 2697
rect 6305 2663 6339 2697
rect 6373 2663 6407 2697
rect 6441 2663 6475 2697
rect 6509 2663 6543 2697
rect 6577 2663 6611 2697
rect 6645 2663 6679 2697
rect 6713 2663 6747 2697
rect 6781 2663 6815 2697
rect 6849 2663 6883 2697
rect 6917 2663 6951 2697
rect 6985 2663 7019 2697
rect 7053 2663 7087 2697
rect 7121 2663 7155 2697
rect 7189 2663 7223 2697
rect 7257 2663 7291 2697
rect 7325 2663 7359 2697
rect 7393 2663 7427 2697
rect 7461 2663 7495 2697
rect 7529 2663 7563 2697
rect 7597 2663 7631 2697
rect 7665 2663 7699 2697
rect 7733 2663 7767 2697
rect 7801 2663 7835 2697
rect 7869 2663 7903 2697
rect 7937 2663 7971 2697
rect 8005 2663 8039 2697
rect 8073 2663 8107 2697
rect 8141 2663 8175 2697
rect 8209 2663 8400 2697
rect 0 2640 8400 2663
rect 0 2560 80 2640
rect 8320 2560 8400 2640
rect 0 2537 8400 2560
rect 0 2503 151 2537
rect 185 2503 219 2537
rect 253 2503 287 2537
rect 321 2503 355 2537
rect 389 2503 423 2537
rect 457 2503 491 2537
rect 525 2503 559 2537
rect 593 2503 627 2537
rect 661 2503 695 2537
rect 729 2503 763 2537
rect 797 2503 831 2537
rect 865 2503 899 2537
rect 933 2503 967 2537
rect 1001 2503 1035 2537
rect 1069 2503 1103 2537
rect 1137 2503 1171 2537
rect 1205 2503 1239 2537
rect 1273 2503 1307 2537
rect 1341 2503 1375 2537
rect 1409 2503 1443 2537
rect 1477 2503 1511 2537
rect 1545 2503 1579 2537
rect 1613 2503 1647 2537
rect 1681 2503 1715 2537
rect 1749 2503 1783 2537
rect 1817 2503 1851 2537
rect 1885 2503 1919 2537
rect 1953 2503 1987 2537
rect 2021 2503 2055 2537
rect 2089 2503 2123 2537
rect 2157 2503 2191 2537
rect 2225 2503 2259 2537
rect 2293 2503 2327 2537
rect 2361 2503 2395 2537
rect 2429 2503 2463 2537
rect 2497 2503 2531 2537
rect 2565 2503 2599 2537
rect 2633 2503 2667 2537
rect 2701 2503 2735 2537
rect 2769 2503 2803 2537
rect 2837 2503 2871 2537
rect 2905 2503 2939 2537
rect 2973 2503 3007 2537
rect 3041 2503 3075 2537
rect 3109 2503 3143 2537
rect 3177 2503 3211 2537
rect 3245 2503 3279 2537
rect 3313 2503 3347 2537
rect 3381 2503 3415 2537
rect 3449 2503 3483 2537
rect 3517 2503 3551 2537
rect 3585 2503 3619 2537
rect 3653 2503 3687 2537
rect 3721 2503 3755 2537
rect 3789 2503 3823 2537
rect 3857 2503 3891 2537
rect 3925 2503 3959 2537
rect 3993 2503 4027 2537
rect 4061 2503 4095 2537
rect 4129 2503 4163 2537
rect 4197 2503 4231 2537
rect 4265 2503 4299 2537
rect 4333 2503 4367 2537
rect 4401 2503 4435 2537
rect 4469 2503 4503 2537
rect 4537 2503 4571 2537
rect 4605 2503 4639 2537
rect 4673 2503 4707 2537
rect 4741 2503 4775 2537
rect 4809 2503 4843 2537
rect 4877 2503 4911 2537
rect 4945 2503 4979 2537
rect 5013 2503 5047 2537
rect 5081 2503 5115 2537
rect 5149 2503 5183 2537
rect 5217 2503 5251 2537
rect 5285 2503 5319 2537
rect 5353 2503 5387 2537
rect 5421 2503 5455 2537
rect 5489 2503 5523 2537
rect 5557 2503 5591 2537
rect 5625 2503 5659 2537
rect 5693 2503 5727 2537
rect 5761 2503 5795 2537
rect 5829 2503 5863 2537
rect 5897 2503 5931 2537
rect 5965 2503 5999 2537
rect 6033 2503 6067 2537
rect 6101 2503 6135 2537
rect 6169 2503 6203 2537
rect 6237 2503 6271 2537
rect 6305 2503 6339 2537
rect 6373 2503 6407 2537
rect 6441 2503 6475 2537
rect 6509 2503 6543 2537
rect 6577 2503 6611 2537
rect 6645 2503 6679 2537
rect 6713 2503 6747 2537
rect 6781 2503 6815 2537
rect 6849 2503 6883 2537
rect 6917 2503 6951 2537
rect 6985 2503 7019 2537
rect 7053 2503 7087 2537
rect 7121 2503 7155 2537
rect 7189 2503 7223 2537
rect 7257 2503 7291 2537
rect 7325 2503 7359 2537
rect 7393 2503 7427 2537
rect 7461 2503 7495 2537
rect 7529 2503 7563 2537
rect 7597 2503 7631 2537
rect 7665 2503 7699 2537
rect 7733 2503 7767 2537
rect 7801 2503 7835 2537
rect 7869 2503 7903 2537
rect 7937 2503 7971 2537
rect 8005 2503 8039 2537
rect 8073 2503 8107 2537
rect 8141 2503 8175 2537
rect 8209 2503 8400 2537
rect 0 2480 8400 2503
rect 0 2407 80 2480
rect 0 2373 23 2407
rect 57 2373 80 2407
rect 8320 2407 8400 2480
rect 0 2339 80 2373
rect 0 2305 23 2339
rect 57 2305 80 2339
rect 0 2271 80 2305
rect 0 2237 23 2271
rect 57 2237 80 2271
rect 0 2203 80 2237
rect 0 2169 23 2203
rect 57 2169 80 2203
rect 0 2135 80 2169
rect 0 2101 23 2135
rect 57 2101 80 2135
rect 0 2067 80 2101
rect 0 2033 23 2067
rect 57 2033 80 2067
rect 0 1999 80 2033
rect 0 1965 23 1999
rect 57 1965 80 1999
rect 0 1931 80 1965
rect 0 1897 23 1931
rect 57 1897 80 1931
rect 0 1863 80 1897
rect 0 1829 23 1863
rect 57 1829 80 1863
rect 0 1795 80 1829
rect 0 1761 23 1795
rect 57 1761 80 1795
rect 0 1727 80 1761
rect 0 1693 23 1727
rect 57 1693 80 1727
rect 0 1659 80 1693
rect 0 1625 23 1659
rect 57 1625 80 1659
rect 0 1591 80 1625
rect 0 1557 23 1591
rect 57 1557 80 1591
rect 0 1523 80 1557
rect 0 1489 23 1523
rect 57 1489 80 1523
rect 0 1455 80 1489
rect 0 1421 23 1455
rect 57 1421 80 1455
rect 0 1387 80 1421
rect 0 1353 23 1387
rect 57 1353 80 1387
rect 160 2377 8240 2400
rect 160 2343 307 2377
rect 341 2343 375 2377
rect 409 2343 443 2377
rect 477 2343 511 2377
rect 545 2343 579 2377
rect 613 2343 647 2377
rect 681 2343 715 2377
rect 749 2343 783 2377
rect 817 2343 851 2377
rect 885 2343 919 2377
rect 953 2343 987 2377
rect 1021 2343 1055 2377
rect 1089 2343 1123 2377
rect 1157 2343 1191 2377
rect 1225 2343 1259 2377
rect 1293 2343 1327 2377
rect 1361 2343 1395 2377
rect 1429 2343 1463 2377
rect 1497 2343 1531 2377
rect 1565 2343 1599 2377
rect 1633 2343 1667 2377
rect 1701 2343 1735 2377
rect 1769 2343 1803 2377
rect 1837 2343 1871 2377
rect 1905 2343 1939 2377
rect 1973 2343 2007 2377
rect 2041 2343 2075 2377
rect 2109 2343 2143 2377
rect 2177 2343 2211 2377
rect 2245 2343 2279 2377
rect 2313 2343 2347 2377
rect 2381 2343 2415 2377
rect 2449 2343 2483 2377
rect 2517 2343 2551 2377
rect 2585 2343 2619 2377
rect 2653 2343 2687 2377
rect 2721 2343 2755 2377
rect 2789 2343 2823 2377
rect 2857 2343 2891 2377
rect 2925 2343 2959 2377
rect 2993 2343 3027 2377
rect 3061 2343 3095 2377
rect 3129 2343 3163 2377
rect 3197 2343 3231 2377
rect 3265 2343 3299 2377
rect 3333 2343 3367 2377
rect 3401 2343 3435 2377
rect 3469 2343 3503 2377
rect 3537 2343 3571 2377
rect 3605 2343 3639 2377
rect 3673 2343 3707 2377
rect 3741 2343 3775 2377
rect 3809 2343 3843 2377
rect 3877 2343 3911 2377
rect 3945 2343 3979 2377
rect 4013 2343 4047 2377
rect 4081 2343 4115 2377
rect 4149 2343 4183 2377
rect 4217 2343 4251 2377
rect 4285 2343 4319 2377
rect 4353 2343 4387 2377
rect 4421 2343 4455 2377
rect 4489 2343 4523 2377
rect 4557 2343 4591 2377
rect 4625 2343 4659 2377
rect 4693 2343 4727 2377
rect 4761 2343 4795 2377
rect 4829 2343 4863 2377
rect 4897 2343 4931 2377
rect 4965 2343 4999 2377
rect 5033 2343 5067 2377
rect 5101 2343 5135 2377
rect 5169 2343 5203 2377
rect 5237 2343 5271 2377
rect 5305 2343 5339 2377
rect 5373 2343 5407 2377
rect 5441 2343 5475 2377
rect 5509 2343 5543 2377
rect 5577 2343 5611 2377
rect 5645 2343 5679 2377
rect 5713 2343 5747 2377
rect 5781 2343 5815 2377
rect 5849 2343 5883 2377
rect 5917 2343 5951 2377
rect 5985 2343 6019 2377
rect 6053 2343 6087 2377
rect 6121 2343 6155 2377
rect 6189 2343 6223 2377
rect 6257 2343 6291 2377
rect 6325 2343 6359 2377
rect 6393 2343 6427 2377
rect 6461 2343 6495 2377
rect 6529 2343 6563 2377
rect 6597 2343 6631 2377
rect 6665 2343 6699 2377
rect 6733 2343 6767 2377
rect 6801 2343 6835 2377
rect 6869 2343 6903 2377
rect 6937 2343 6971 2377
rect 7005 2343 7039 2377
rect 7073 2343 7107 2377
rect 7141 2343 7175 2377
rect 7209 2343 7243 2377
rect 7277 2343 7311 2377
rect 7345 2343 7379 2377
rect 7413 2343 7447 2377
rect 7481 2343 7515 2377
rect 7549 2343 7583 2377
rect 7617 2343 7651 2377
rect 7685 2343 7719 2377
rect 7753 2343 7787 2377
rect 7821 2343 7855 2377
rect 7889 2343 7923 2377
rect 7957 2343 7991 2377
rect 8025 2343 8059 2377
rect 8093 2343 8240 2377
rect 160 2320 8240 2343
rect 160 2271 240 2320
rect 160 2237 183 2271
rect 217 2237 240 2271
rect 160 2203 240 2237
rect 160 2169 183 2203
rect 217 2169 240 2203
rect 160 2135 240 2169
rect 160 2101 183 2135
rect 217 2101 240 2135
rect 160 2067 240 2101
rect 160 2033 183 2067
rect 217 2033 240 2067
rect 160 1999 240 2033
rect 160 1965 183 1999
rect 217 1965 240 1999
rect 160 1931 240 1965
rect 160 1897 183 1931
rect 217 1897 240 1931
rect 160 1863 240 1897
rect 160 1829 183 1863
rect 217 1829 240 1863
rect 160 1795 240 1829
rect 160 1761 183 1795
rect 217 1761 240 1795
rect 160 1727 240 1761
rect 160 1693 183 1727
rect 217 1693 240 1727
rect 160 1659 240 1693
rect 160 1625 183 1659
rect 217 1625 240 1659
rect 320 2209 400 2320
rect 320 2161 343 2209
rect 377 2161 400 2209
rect 320 2137 400 2161
rect 320 2093 343 2137
rect 377 2093 400 2137
rect 320 2065 400 2093
rect 320 2025 343 2065
rect 377 2025 400 2065
rect 320 1993 400 2025
rect 320 1957 343 1993
rect 377 1957 400 1993
rect 320 1923 400 1957
rect 320 1887 343 1923
rect 377 1887 400 1923
rect 320 1855 400 1887
rect 320 1815 343 1855
rect 377 1815 400 1855
rect 320 1787 400 1815
rect 320 1743 343 1787
rect 377 1743 400 1787
rect 320 1719 400 1743
rect 320 1671 343 1719
rect 377 1671 400 1719
rect 320 1640 400 1671
rect 2240 2209 2320 2240
rect 2240 2161 2263 2209
rect 2297 2161 2320 2209
rect 2240 2137 2320 2161
rect 2240 2093 2263 2137
rect 2297 2093 2320 2137
rect 2240 2065 2320 2093
rect 2240 2025 2263 2065
rect 2297 2025 2320 2065
rect 2240 1993 2320 2025
rect 2240 1957 2263 1993
rect 2297 1957 2320 1993
rect 2240 1923 2320 1957
rect 2240 1887 2263 1923
rect 2297 1887 2320 1923
rect 2240 1855 2320 1887
rect 2240 1815 2263 1855
rect 2297 1815 2320 1855
rect 2240 1787 2320 1815
rect 2240 1743 2263 1787
rect 2297 1743 2320 1787
rect 2240 1719 2320 1743
rect 2240 1671 2263 1719
rect 2297 1671 2320 1719
rect 2240 1640 2320 1671
rect 4160 2209 4240 2240
rect 4160 2161 4183 2209
rect 4217 2161 4240 2209
rect 4160 2137 4240 2161
rect 4160 2093 4183 2137
rect 4217 2093 4240 2137
rect 4160 2065 4240 2093
rect 4160 2025 4183 2065
rect 4217 2025 4240 2065
rect 4160 1993 4240 2025
rect 4160 1957 4183 1993
rect 4217 1957 4240 1993
rect 4160 1923 4240 1957
rect 4160 1887 4183 1923
rect 4217 1887 4240 1923
rect 4160 1855 4240 1887
rect 4160 1815 4183 1855
rect 4217 1815 4240 1855
rect 4160 1787 4240 1815
rect 4160 1743 4183 1787
rect 4217 1743 4240 1787
rect 4160 1719 4240 1743
rect 4160 1671 4183 1719
rect 4217 1671 4240 1719
rect 4160 1640 4240 1671
rect 6080 2209 6160 2240
rect 6080 2161 6103 2209
rect 6137 2161 6160 2209
rect 6080 2137 6160 2161
rect 6080 2093 6103 2137
rect 6137 2093 6160 2137
rect 6080 2065 6160 2093
rect 6080 2025 6103 2065
rect 6137 2025 6160 2065
rect 6080 1993 6160 2025
rect 6080 1957 6103 1993
rect 6137 1957 6160 1993
rect 6080 1923 6160 1957
rect 6080 1887 6103 1923
rect 6137 1887 6160 1923
rect 6080 1855 6160 1887
rect 6080 1815 6103 1855
rect 6137 1815 6160 1855
rect 6080 1787 6160 1815
rect 6080 1743 6103 1787
rect 6137 1743 6160 1787
rect 6080 1719 6160 1743
rect 6080 1671 6103 1719
rect 6137 1671 6160 1719
rect 6080 1640 6160 1671
rect 8000 2209 8080 2320
rect 8000 2161 8023 2209
rect 8057 2161 8080 2209
rect 8000 2137 8080 2161
rect 8000 2093 8023 2137
rect 8057 2093 8080 2137
rect 8000 2065 8080 2093
rect 8000 2025 8023 2065
rect 8057 2025 8080 2065
rect 8000 1993 8080 2025
rect 8000 1957 8023 1993
rect 8057 1957 8080 1993
rect 8000 1923 8080 1957
rect 8000 1887 8023 1923
rect 8057 1887 8080 1923
rect 8000 1855 8080 1887
rect 8000 1815 8023 1855
rect 8057 1815 8080 1855
rect 8000 1787 8080 1815
rect 8000 1743 8023 1787
rect 8057 1743 8080 1787
rect 8000 1719 8080 1743
rect 8000 1671 8023 1719
rect 8057 1671 8080 1719
rect 8000 1640 8080 1671
rect 8160 2271 8240 2320
rect 8160 2237 8183 2271
rect 8217 2237 8240 2271
rect 8160 2203 8240 2237
rect 8160 2169 8183 2203
rect 8217 2169 8240 2203
rect 8160 2135 8240 2169
rect 8160 2101 8183 2135
rect 8217 2101 8240 2135
rect 8160 2067 8240 2101
rect 8160 2033 8183 2067
rect 8217 2033 8240 2067
rect 8160 1999 8240 2033
rect 8160 1965 8183 1999
rect 8217 1965 8240 1999
rect 8160 1931 8240 1965
rect 8160 1897 8183 1931
rect 8217 1897 8240 1931
rect 8160 1863 8240 1897
rect 8160 1829 8183 1863
rect 8217 1829 8240 1863
rect 8160 1795 8240 1829
rect 8160 1761 8183 1795
rect 8217 1761 8240 1795
rect 8160 1727 8240 1761
rect 8160 1693 8183 1727
rect 8217 1693 8240 1727
rect 8160 1659 8240 1693
rect 160 1591 240 1625
rect 8160 1625 8183 1659
rect 8217 1625 8240 1659
rect 160 1557 183 1591
rect 217 1557 240 1591
rect 160 1523 240 1557
rect 160 1489 183 1523
rect 217 1489 240 1523
rect 520 1577 2120 1600
rect 520 1543 547 1577
rect 589 1543 619 1577
rect 657 1543 691 1577
rect 725 1543 759 1577
rect 797 1543 827 1577
rect 869 1543 895 1577
rect 941 1543 963 1577
rect 1013 1543 1031 1577
rect 1085 1543 1099 1577
rect 1157 1543 1167 1577
rect 1229 1543 1235 1577
rect 1301 1543 1303 1577
rect 1337 1543 1339 1577
rect 1405 1543 1411 1577
rect 1473 1543 1483 1577
rect 1541 1543 1555 1577
rect 1609 1543 1627 1577
rect 1677 1543 1699 1577
rect 1745 1543 1771 1577
rect 1813 1543 1843 1577
rect 1881 1543 1915 1577
rect 1949 1543 1983 1577
rect 2021 1543 2051 1577
rect 2093 1543 2120 1577
rect 520 1520 2120 1543
rect 2440 1577 4040 1600
rect 2440 1543 2467 1577
rect 2509 1543 2539 1577
rect 2577 1543 2611 1577
rect 2645 1543 2679 1577
rect 2717 1543 2747 1577
rect 2789 1543 2815 1577
rect 2861 1543 2883 1577
rect 2933 1543 2951 1577
rect 3005 1543 3019 1577
rect 3077 1543 3087 1577
rect 3149 1543 3155 1577
rect 3221 1543 3223 1577
rect 3257 1543 3259 1577
rect 3325 1543 3331 1577
rect 3393 1543 3403 1577
rect 3461 1543 3475 1577
rect 3529 1543 3547 1577
rect 3597 1543 3619 1577
rect 3665 1543 3691 1577
rect 3733 1543 3763 1577
rect 3801 1543 3835 1577
rect 3869 1543 3903 1577
rect 3941 1543 3971 1577
rect 4013 1543 4040 1577
rect 2440 1520 4040 1543
rect 4360 1577 5960 1600
rect 4360 1543 4387 1577
rect 4429 1543 4459 1577
rect 4497 1543 4531 1577
rect 4565 1543 4599 1577
rect 4637 1543 4667 1577
rect 4709 1543 4735 1577
rect 4781 1543 4803 1577
rect 4853 1543 4871 1577
rect 4925 1543 4939 1577
rect 4997 1543 5007 1577
rect 5069 1543 5075 1577
rect 5141 1543 5143 1577
rect 5177 1543 5179 1577
rect 5245 1543 5251 1577
rect 5313 1543 5323 1577
rect 5381 1543 5395 1577
rect 5449 1543 5467 1577
rect 5517 1543 5539 1577
rect 5585 1543 5611 1577
rect 5653 1543 5683 1577
rect 5721 1543 5755 1577
rect 5789 1543 5823 1577
rect 5861 1543 5891 1577
rect 5933 1543 5960 1577
rect 4360 1520 5960 1543
rect 6280 1577 7880 1600
rect 6280 1543 6307 1577
rect 6349 1543 6379 1577
rect 6417 1543 6451 1577
rect 6485 1543 6519 1577
rect 6557 1543 6587 1577
rect 6629 1543 6655 1577
rect 6701 1543 6723 1577
rect 6773 1543 6791 1577
rect 6845 1543 6859 1577
rect 6917 1543 6927 1577
rect 6989 1543 6995 1577
rect 7061 1543 7063 1577
rect 7097 1543 7099 1577
rect 7165 1543 7171 1577
rect 7233 1543 7243 1577
rect 7301 1543 7315 1577
rect 7369 1543 7387 1577
rect 7437 1543 7459 1577
rect 7505 1543 7531 1577
rect 7573 1543 7603 1577
rect 7641 1543 7675 1577
rect 7709 1543 7743 1577
rect 7781 1543 7811 1577
rect 7853 1543 7880 1577
rect 6280 1520 7880 1543
rect 8160 1591 8240 1625
rect 8160 1557 8183 1591
rect 8217 1557 8240 1591
rect 8160 1523 8240 1557
rect 160 1440 240 1489
rect 8160 1489 8183 1523
rect 8217 1489 8240 1523
rect 8160 1440 8240 1489
rect 160 1417 8240 1440
rect 160 1383 307 1417
rect 341 1383 375 1417
rect 409 1383 443 1417
rect 477 1383 511 1417
rect 545 1383 579 1417
rect 613 1383 647 1417
rect 681 1383 715 1417
rect 749 1383 783 1417
rect 817 1383 851 1417
rect 885 1383 919 1417
rect 953 1383 987 1417
rect 1021 1383 1055 1417
rect 1089 1383 1123 1417
rect 1157 1383 1191 1417
rect 1225 1383 1259 1417
rect 1293 1383 1327 1417
rect 1361 1383 1395 1417
rect 1429 1383 1463 1417
rect 1497 1383 1531 1417
rect 1565 1383 1599 1417
rect 1633 1383 1667 1417
rect 1701 1383 1735 1417
rect 1769 1383 1803 1417
rect 1837 1383 1871 1417
rect 1905 1383 1939 1417
rect 1973 1383 2007 1417
rect 2041 1383 2075 1417
rect 2109 1383 2143 1417
rect 2177 1383 2211 1417
rect 2245 1383 2279 1417
rect 2313 1383 2347 1417
rect 2381 1383 2415 1417
rect 2449 1383 2483 1417
rect 2517 1383 2551 1417
rect 2585 1383 2619 1417
rect 2653 1383 2687 1417
rect 2721 1383 2755 1417
rect 2789 1383 2823 1417
rect 2857 1383 2891 1417
rect 2925 1383 2959 1417
rect 2993 1383 3027 1417
rect 3061 1383 3095 1417
rect 3129 1383 3163 1417
rect 3197 1383 3231 1417
rect 3265 1383 3299 1417
rect 3333 1383 3367 1417
rect 3401 1383 3435 1417
rect 3469 1383 3503 1417
rect 3537 1383 3571 1417
rect 3605 1383 3639 1417
rect 3673 1383 3707 1417
rect 3741 1383 3775 1417
rect 3809 1383 3843 1417
rect 3877 1383 3911 1417
rect 3945 1383 3979 1417
rect 4013 1383 4047 1417
rect 4081 1383 4115 1417
rect 4149 1383 4183 1417
rect 4217 1383 4251 1417
rect 4285 1383 4319 1417
rect 4353 1383 4387 1417
rect 4421 1383 4455 1417
rect 4489 1383 4523 1417
rect 4557 1383 4591 1417
rect 4625 1383 4659 1417
rect 4693 1383 4727 1417
rect 4761 1383 4795 1417
rect 4829 1383 4863 1417
rect 4897 1383 4931 1417
rect 4965 1383 4999 1417
rect 5033 1383 5067 1417
rect 5101 1383 5135 1417
rect 5169 1383 5203 1417
rect 5237 1383 5271 1417
rect 5305 1383 5339 1417
rect 5373 1383 5407 1417
rect 5441 1383 5475 1417
rect 5509 1383 5543 1417
rect 5577 1383 5611 1417
rect 5645 1383 5679 1417
rect 5713 1383 5747 1417
rect 5781 1383 5815 1417
rect 5849 1383 5883 1417
rect 5917 1383 5951 1417
rect 5985 1383 6019 1417
rect 6053 1383 6087 1417
rect 6121 1383 6155 1417
rect 6189 1383 6223 1417
rect 6257 1383 6291 1417
rect 6325 1383 6359 1417
rect 6393 1383 6427 1417
rect 6461 1383 6495 1417
rect 6529 1383 6563 1417
rect 6597 1383 6631 1417
rect 6665 1383 6699 1417
rect 6733 1383 6767 1417
rect 6801 1383 6835 1417
rect 6869 1383 6903 1417
rect 6937 1383 6971 1417
rect 7005 1383 7039 1417
rect 7073 1383 7107 1417
rect 7141 1383 7175 1417
rect 7209 1383 7243 1417
rect 7277 1383 7311 1417
rect 7345 1383 7379 1417
rect 7413 1383 7447 1417
rect 7481 1383 7515 1417
rect 7549 1383 7583 1417
rect 7617 1383 7651 1417
rect 7685 1383 7719 1417
rect 7753 1383 7787 1417
rect 7821 1383 7855 1417
rect 7889 1383 7923 1417
rect 7957 1383 7991 1417
rect 8025 1383 8059 1417
rect 8093 1383 8240 1417
rect 160 1360 8240 1383
rect 8320 2373 8343 2407
rect 8377 2373 8400 2407
rect 8320 2339 8400 2373
rect 8320 2305 8343 2339
rect 8377 2305 8400 2339
rect 8320 2271 8400 2305
rect 8320 2237 8343 2271
rect 8377 2237 8400 2271
rect 8320 2203 8400 2237
rect 8320 2169 8343 2203
rect 8377 2169 8400 2203
rect 8320 2135 8400 2169
rect 8320 2101 8343 2135
rect 8377 2101 8400 2135
rect 8320 2067 8400 2101
rect 8320 2033 8343 2067
rect 8377 2033 8400 2067
rect 8320 1999 8400 2033
rect 8320 1965 8343 1999
rect 8377 1965 8400 1999
rect 8320 1931 8400 1965
rect 8320 1897 8343 1931
rect 8377 1897 8400 1931
rect 8320 1863 8400 1897
rect 8320 1829 8343 1863
rect 8377 1829 8400 1863
rect 8320 1795 8400 1829
rect 8320 1761 8343 1795
rect 8377 1761 8400 1795
rect 8320 1727 8400 1761
rect 8320 1693 8343 1727
rect 8377 1693 8400 1727
rect 8320 1659 8400 1693
rect 8320 1625 8343 1659
rect 8377 1625 8400 1659
rect 8320 1591 8400 1625
rect 8320 1557 8343 1591
rect 8377 1557 8400 1591
rect 8320 1523 8400 1557
rect 8320 1489 8343 1523
rect 8377 1489 8400 1523
rect 8320 1455 8400 1489
rect 8320 1421 8343 1455
rect 8377 1421 8400 1455
rect 8320 1387 8400 1421
rect 0 1280 80 1353
rect 8320 1353 8343 1387
rect 8377 1353 8400 1387
rect 8320 1280 8400 1353
rect 0 1257 8400 1280
rect 0 1223 137 1257
rect 171 1223 205 1257
rect 239 1223 273 1257
rect 307 1223 341 1257
rect 375 1223 409 1257
rect 443 1223 477 1257
rect 511 1223 545 1257
rect 579 1223 613 1257
rect 647 1223 681 1257
rect 715 1223 749 1257
rect 783 1223 817 1257
rect 851 1223 885 1257
rect 919 1223 953 1257
rect 987 1223 1021 1257
rect 1055 1223 1089 1257
rect 1123 1223 1157 1257
rect 1191 1223 1225 1257
rect 1259 1223 1293 1257
rect 1327 1223 1361 1257
rect 1395 1223 1429 1257
rect 1463 1223 1497 1257
rect 1531 1223 1565 1257
rect 1599 1223 1633 1257
rect 1667 1223 1701 1257
rect 1735 1223 1769 1257
rect 1803 1223 1837 1257
rect 1871 1223 1905 1257
rect 1939 1223 1973 1257
rect 2007 1223 2041 1257
rect 2075 1223 2109 1257
rect 2143 1223 2177 1257
rect 2211 1223 2245 1257
rect 2279 1223 2313 1257
rect 2347 1223 2381 1257
rect 2415 1223 2449 1257
rect 2483 1223 2517 1257
rect 2551 1223 2585 1257
rect 2619 1223 2653 1257
rect 2687 1223 2721 1257
rect 2755 1223 2789 1257
rect 2823 1223 2857 1257
rect 2891 1223 2925 1257
rect 2959 1223 2993 1257
rect 3027 1223 3061 1257
rect 3095 1223 3129 1257
rect 3163 1223 3197 1257
rect 3231 1223 3265 1257
rect 3299 1223 3333 1257
rect 3367 1223 3401 1257
rect 3435 1223 3469 1257
rect 3503 1223 3537 1257
rect 3571 1223 3605 1257
rect 3639 1223 3673 1257
rect 3707 1223 3741 1257
rect 3775 1223 3809 1257
rect 3843 1223 3877 1257
rect 3911 1223 3945 1257
rect 3979 1223 4013 1257
rect 4047 1223 4081 1257
rect 4115 1223 4149 1257
rect 4183 1223 4217 1257
rect 4251 1223 4285 1257
rect 4319 1223 4353 1257
rect 4387 1223 4421 1257
rect 4455 1223 4489 1257
rect 4523 1223 4557 1257
rect 4591 1223 4625 1257
rect 4659 1223 4693 1257
rect 4727 1223 4761 1257
rect 4795 1223 4829 1257
rect 4863 1223 4897 1257
rect 4931 1223 4965 1257
rect 4999 1223 5033 1257
rect 5067 1223 5101 1257
rect 5135 1223 5169 1257
rect 5203 1223 5237 1257
rect 5271 1223 5305 1257
rect 5339 1223 5373 1257
rect 5407 1223 5441 1257
rect 5475 1223 5509 1257
rect 5543 1223 5577 1257
rect 5611 1223 5645 1257
rect 5679 1223 5713 1257
rect 5747 1223 5781 1257
rect 5815 1223 5849 1257
rect 5883 1223 5917 1257
rect 5951 1223 5985 1257
rect 6019 1223 6053 1257
rect 6087 1223 6121 1257
rect 6155 1223 6189 1257
rect 6223 1223 6257 1257
rect 6291 1223 6325 1257
rect 6359 1223 6393 1257
rect 6427 1223 6461 1257
rect 6495 1223 6529 1257
rect 6563 1223 6597 1257
rect 6631 1223 6665 1257
rect 6699 1223 6733 1257
rect 6767 1223 6801 1257
rect 6835 1223 6869 1257
rect 6903 1223 6937 1257
rect 6971 1223 7005 1257
rect 7039 1223 7073 1257
rect 7107 1223 7141 1257
rect 7175 1223 7209 1257
rect 7243 1223 7277 1257
rect 7311 1223 7345 1257
rect 7379 1223 7413 1257
rect 7447 1223 7481 1257
rect 7515 1223 7549 1257
rect 7583 1223 7617 1257
rect 7651 1223 7685 1257
rect 7719 1223 7753 1257
rect 7787 1223 7821 1257
rect 7855 1223 7889 1257
rect 7923 1223 7957 1257
rect 7991 1223 8025 1257
rect 8059 1223 8093 1257
rect 8127 1223 8161 1257
rect 8195 1223 8229 1257
rect 8263 1223 8400 1257
rect 0 1200 8400 1223
rect 0 640 80 1200
rect 160 937 8240 1120
rect 160 903 183 937
rect 217 903 343 937
rect 377 903 503 937
rect 537 903 663 937
rect 697 903 823 937
rect 857 903 983 937
rect 1017 903 1143 937
rect 1177 903 1463 937
rect 1497 903 1623 937
rect 1657 903 1783 937
rect 1817 903 1943 937
rect 1977 903 2103 937
rect 2137 903 2263 937
rect 2297 903 2423 937
rect 2457 903 2583 937
rect 2617 903 2743 937
rect 2777 903 2903 937
rect 2937 903 3063 937
rect 3097 903 3383 937
rect 3417 903 3543 937
rect 3577 903 3703 937
rect 3737 903 3863 937
rect 3897 903 4023 937
rect 4057 903 4343 937
rect 4377 903 4503 937
rect 4537 903 4663 937
rect 4697 903 4823 937
rect 4857 903 4983 937
rect 5017 903 5303 937
rect 5337 903 5463 937
rect 5497 903 5623 937
rect 5657 903 5783 937
rect 5817 903 5943 937
rect 5977 903 6103 937
rect 6137 903 6263 937
rect 6297 903 6423 937
rect 6457 903 6583 937
rect 6617 903 6743 937
rect 6777 903 6903 937
rect 6937 903 7223 937
rect 7257 903 7383 937
rect 7417 903 7543 937
rect 7577 903 7703 937
rect 7737 903 7863 937
rect 7897 903 8023 937
rect 8057 903 8183 937
rect 8217 903 8240 937
rect 160 720 8240 903
rect 8320 640 8400 1200
rect 0 617 8400 640
rect 0 583 137 617
rect 171 583 205 617
rect 239 583 273 617
rect 307 583 341 617
rect 375 583 409 617
rect 443 583 477 617
rect 511 583 545 617
rect 579 583 613 617
rect 647 583 681 617
rect 715 583 749 617
rect 783 583 817 617
rect 851 583 885 617
rect 919 583 953 617
rect 987 583 1021 617
rect 1055 583 1089 617
rect 1123 583 1157 617
rect 1191 583 1225 617
rect 1259 583 1293 617
rect 1327 583 1361 617
rect 1395 583 1429 617
rect 1463 583 1497 617
rect 1531 583 1565 617
rect 1599 583 1633 617
rect 1667 583 1701 617
rect 1735 583 1769 617
rect 1803 583 1837 617
rect 1871 583 1905 617
rect 1939 583 1973 617
rect 2007 583 2041 617
rect 2075 583 2109 617
rect 2143 583 2177 617
rect 2211 583 2245 617
rect 2279 583 2313 617
rect 2347 583 2381 617
rect 2415 583 2449 617
rect 2483 583 2517 617
rect 2551 583 2585 617
rect 2619 583 2653 617
rect 2687 583 2721 617
rect 2755 583 2789 617
rect 2823 583 2857 617
rect 2891 583 2925 617
rect 2959 583 2993 617
rect 3027 583 3061 617
rect 3095 583 3129 617
rect 3163 583 3197 617
rect 3231 583 3265 617
rect 3299 583 3333 617
rect 3367 583 3401 617
rect 3435 583 3469 617
rect 3503 583 3537 617
rect 3571 583 3605 617
rect 3639 583 3673 617
rect 3707 583 3741 617
rect 3775 583 3809 617
rect 3843 583 3877 617
rect 3911 583 3945 617
rect 3979 583 4013 617
rect 4047 583 4081 617
rect 4115 583 4149 617
rect 4183 583 4217 617
rect 4251 583 4285 617
rect 4319 583 4353 617
rect 4387 583 4421 617
rect 4455 583 4489 617
rect 4523 583 4557 617
rect 4591 583 4625 617
rect 4659 583 4693 617
rect 4727 583 4761 617
rect 4795 583 4829 617
rect 4863 583 4897 617
rect 4931 583 4965 617
rect 4999 583 5033 617
rect 5067 583 5101 617
rect 5135 583 5169 617
rect 5203 583 5237 617
rect 5271 583 5305 617
rect 5339 583 5373 617
rect 5407 583 5441 617
rect 5475 583 5509 617
rect 5543 583 5577 617
rect 5611 583 5645 617
rect 5679 583 5713 617
rect 5747 583 5781 617
rect 5815 583 5849 617
rect 5883 583 5917 617
rect 5951 583 5985 617
rect 6019 583 6053 617
rect 6087 583 6121 617
rect 6155 583 6189 617
rect 6223 583 6257 617
rect 6291 583 6325 617
rect 6359 583 6393 617
rect 6427 583 6461 617
rect 6495 583 6529 617
rect 6563 583 6597 617
rect 6631 583 6665 617
rect 6699 583 6733 617
rect 6767 583 6801 617
rect 6835 583 6869 617
rect 6903 583 6937 617
rect 6971 583 7005 617
rect 7039 583 7073 617
rect 7107 583 7141 617
rect 7175 583 7209 617
rect 7243 583 7277 617
rect 7311 583 7345 617
rect 7379 583 7413 617
rect 7447 583 7481 617
rect 7515 583 7549 617
rect 7583 583 7617 617
rect 7651 583 7685 617
rect 7719 583 7753 617
rect 7787 583 7821 617
rect 7855 583 7889 617
rect 7923 583 7957 617
rect 7991 583 8025 617
rect 8059 583 8093 617
rect 8127 583 8161 617
rect 8195 583 8229 617
rect 8263 583 8400 617
rect 0 560 8400 583
rect 0 507 80 560
rect 0 473 23 507
rect 57 473 80 507
rect 8320 507 8400 560
rect 0 439 80 473
rect 0 405 23 439
rect 57 405 80 439
rect 0 371 80 405
rect 520 457 2120 480
rect 520 423 547 457
rect 589 423 619 457
rect 657 423 691 457
rect 725 423 759 457
rect 797 423 827 457
rect 869 423 895 457
rect 941 423 963 457
rect 1013 423 1031 457
rect 1085 423 1099 457
rect 1157 423 1167 457
rect 1229 423 1235 457
rect 1301 423 1303 457
rect 1337 423 1339 457
rect 1405 423 1411 457
rect 1473 423 1483 457
rect 1541 423 1555 457
rect 1609 423 1627 457
rect 1677 423 1699 457
rect 1745 423 1771 457
rect 1813 423 1843 457
rect 1881 423 1915 457
rect 1949 423 1983 457
rect 2021 423 2051 457
rect 2093 423 2120 457
rect 520 400 2120 423
rect 2440 457 4040 480
rect 2440 423 2467 457
rect 2509 423 2539 457
rect 2577 423 2611 457
rect 2645 423 2679 457
rect 2717 423 2747 457
rect 2789 423 2815 457
rect 2861 423 2883 457
rect 2933 423 2951 457
rect 3005 423 3019 457
rect 3077 423 3087 457
rect 3149 423 3155 457
rect 3221 423 3223 457
rect 3257 423 3259 457
rect 3325 423 3331 457
rect 3393 423 3403 457
rect 3461 423 3475 457
rect 3529 423 3547 457
rect 3597 423 3619 457
rect 3665 423 3691 457
rect 3733 423 3763 457
rect 3801 423 3835 457
rect 3869 423 3903 457
rect 3941 423 3971 457
rect 4013 423 4040 457
rect 2440 400 4040 423
rect 4360 457 5960 480
rect 4360 423 4387 457
rect 4429 423 4459 457
rect 4497 423 4531 457
rect 4565 423 4599 457
rect 4637 423 4667 457
rect 4709 423 4735 457
rect 4781 423 4803 457
rect 4853 423 4871 457
rect 4925 423 4939 457
rect 4997 423 5007 457
rect 5069 423 5075 457
rect 5141 423 5143 457
rect 5177 423 5179 457
rect 5245 423 5251 457
rect 5313 423 5323 457
rect 5381 423 5395 457
rect 5449 423 5467 457
rect 5517 423 5539 457
rect 5585 423 5611 457
rect 5653 423 5683 457
rect 5721 423 5755 457
rect 5789 423 5823 457
rect 5861 423 5891 457
rect 5933 423 5960 457
rect 4360 400 5960 423
rect 6280 457 7880 480
rect 6280 423 6307 457
rect 6349 423 6379 457
rect 6417 423 6451 457
rect 6485 423 6519 457
rect 6557 423 6587 457
rect 6629 423 6655 457
rect 6701 423 6723 457
rect 6773 423 6791 457
rect 6845 423 6859 457
rect 6917 423 6927 457
rect 6989 423 6995 457
rect 7061 423 7063 457
rect 7097 423 7099 457
rect 7165 423 7171 457
rect 7233 423 7243 457
rect 7301 423 7315 457
rect 7369 423 7387 457
rect 7437 423 7459 457
rect 7505 423 7531 457
rect 7573 423 7603 457
rect 7641 423 7675 457
rect 7709 423 7743 457
rect 7781 423 7811 457
rect 7853 423 7880 457
rect 6280 400 7880 423
rect 8320 473 8343 507
rect 8377 473 8400 507
rect 8320 439 8400 473
rect 8320 405 8343 439
rect 8377 405 8400 439
rect 0 337 23 371
rect 57 337 80 371
rect 8320 371 8400 405
rect 0 303 80 337
rect 0 269 23 303
rect 57 269 80 303
rect 0 235 80 269
rect 0 201 23 235
rect 57 201 80 235
rect 0 167 80 201
rect 0 133 23 167
rect 57 133 80 167
rect 0 80 80 133
rect 320 313 400 360
rect 320 277 343 313
rect 377 277 400 313
rect 320 243 400 277
rect 320 207 343 243
rect 377 207 400 243
rect 320 80 400 207
rect 2240 313 2320 360
rect 2240 277 2263 313
rect 2297 277 2320 313
rect 2240 243 2320 277
rect 2240 207 2263 243
rect 2297 207 2320 243
rect 2240 160 2320 207
rect 4160 313 4240 360
rect 4160 277 4183 313
rect 4217 277 4240 313
rect 4160 243 4240 277
rect 4160 207 4183 243
rect 4217 207 4240 243
rect 4160 160 4240 207
rect 6080 313 6160 360
rect 6080 277 6103 313
rect 6137 277 6160 313
rect 6080 243 6160 277
rect 6080 207 6103 243
rect 6137 207 6160 243
rect 6080 160 6160 207
rect 8000 313 8080 360
rect 8000 277 8023 313
rect 8057 277 8080 313
rect 8000 243 8080 277
rect 8000 207 8023 243
rect 8057 207 8080 243
rect 8000 80 8080 207
rect 8320 337 8343 371
rect 8377 337 8400 371
rect 8320 303 8400 337
rect 8320 269 8343 303
rect 8377 269 8400 303
rect 8320 235 8400 269
rect 8320 201 8343 235
rect 8377 201 8400 235
rect 8320 167 8400 201
rect 8320 133 8343 167
rect 8377 133 8400 167
rect 8320 80 8400 133
rect 0 57 8400 80
rect 0 23 137 57
rect 171 23 205 57
rect 239 23 273 57
rect 307 23 341 57
rect 375 23 409 57
rect 443 23 477 57
rect 511 23 545 57
rect 579 23 613 57
rect 647 23 681 57
rect 715 23 749 57
rect 783 23 817 57
rect 851 23 885 57
rect 919 23 953 57
rect 987 23 1021 57
rect 1055 23 1089 57
rect 1123 23 1157 57
rect 1191 23 1225 57
rect 1259 23 1293 57
rect 1327 23 1361 57
rect 1395 23 1429 57
rect 1463 23 1497 57
rect 1531 23 1565 57
rect 1599 23 1633 57
rect 1667 23 1701 57
rect 1735 23 1769 57
rect 1803 23 1837 57
rect 1871 23 1905 57
rect 1939 23 1973 57
rect 2007 23 2041 57
rect 2075 23 2109 57
rect 2143 23 2177 57
rect 2211 23 2245 57
rect 2279 23 2313 57
rect 2347 23 2381 57
rect 2415 23 2449 57
rect 2483 23 2517 57
rect 2551 23 2585 57
rect 2619 23 2653 57
rect 2687 23 2721 57
rect 2755 23 2789 57
rect 2823 23 2857 57
rect 2891 23 2925 57
rect 2959 23 2993 57
rect 3027 23 3061 57
rect 3095 23 3129 57
rect 3163 23 3197 57
rect 3231 23 3265 57
rect 3299 23 3333 57
rect 3367 23 3401 57
rect 3435 23 3469 57
rect 3503 23 3537 57
rect 3571 23 3605 57
rect 3639 23 3673 57
rect 3707 23 3741 57
rect 3775 23 3809 57
rect 3843 23 3877 57
rect 3911 23 3945 57
rect 3979 23 4013 57
rect 4047 23 4081 57
rect 4115 23 4149 57
rect 4183 23 4217 57
rect 4251 23 4285 57
rect 4319 23 4353 57
rect 4387 23 4421 57
rect 4455 23 4489 57
rect 4523 23 4557 57
rect 4591 23 4625 57
rect 4659 23 4693 57
rect 4727 23 4761 57
rect 4795 23 4829 57
rect 4863 23 4897 57
rect 4931 23 4965 57
rect 4999 23 5033 57
rect 5067 23 5101 57
rect 5135 23 5169 57
rect 5203 23 5237 57
rect 5271 23 5305 57
rect 5339 23 5373 57
rect 5407 23 5441 57
rect 5475 23 5509 57
rect 5543 23 5577 57
rect 5611 23 5645 57
rect 5679 23 5713 57
rect 5747 23 5781 57
rect 5815 23 5849 57
rect 5883 23 5917 57
rect 5951 23 5985 57
rect 6019 23 6053 57
rect 6087 23 6121 57
rect 6155 23 6189 57
rect 6223 23 6257 57
rect 6291 23 6325 57
rect 6359 23 6393 57
rect 6427 23 6461 57
rect 6495 23 6529 57
rect 6563 23 6597 57
rect 6631 23 6665 57
rect 6699 23 6733 57
rect 6767 23 6801 57
rect 6835 23 6869 57
rect 6903 23 6937 57
rect 6971 23 7005 57
rect 7039 23 7073 57
rect 7107 23 7141 57
rect 7175 23 7209 57
rect 7243 23 7277 57
rect 7311 23 7345 57
rect 7379 23 7413 57
rect 7447 23 7481 57
rect 7515 23 7549 57
rect 7583 23 7617 57
rect 7651 23 7685 57
rect 7719 23 7753 57
rect 7787 23 7821 57
rect 7855 23 7889 57
rect 7923 23 7957 57
rect 7991 23 8025 57
rect 8059 23 8093 57
rect 8127 23 8161 57
rect 8195 23 8229 57
rect 8263 23 8400 57
rect 0 0 8400 23
<< viali >>
rect 343 3635 377 3649
rect 343 3615 377 3635
rect 343 3567 377 3577
rect 343 3543 377 3567
rect 343 3499 377 3505
rect 343 3471 377 3499
rect 343 3431 377 3433
rect 343 3399 377 3431
rect 343 3329 377 3361
rect 343 3327 377 3329
rect 343 3261 377 3289
rect 343 3255 377 3261
rect 343 3193 377 3217
rect 343 3183 377 3193
rect 343 3125 377 3145
rect 343 3111 377 3125
rect 2263 3635 2297 3649
rect 2263 3615 2297 3635
rect 2263 3567 2297 3577
rect 2263 3543 2297 3567
rect 2263 3499 2297 3505
rect 2263 3471 2297 3499
rect 2263 3431 2297 3433
rect 2263 3399 2297 3431
rect 2263 3329 2297 3361
rect 2263 3327 2297 3329
rect 2263 3261 2297 3289
rect 2263 3255 2297 3261
rect 2263 3193 2297 3217
rect 2263 3183 2297 3193
rect 2263 3125 2297 3145
rect 2263 3111 2297 3125
rect 4183 3635 4217 3649
rect 4183 3615 4217 3635
rect 4183 3567 4217 3577
rect 4183 3543 4217 3567
rect 4183 3499 4217 3505
rect 4183 3471 4217 3499
rect 4183 3431 4217 3433
rect 4183 3399 4217 3431
rect 4183 3329 4217 3361
rect 4183 3327 4217 3329
rect 4183 3261 4217 3289
rect 4183 3255 4217 3261
rect 4183 3193 4217 3217
rect 4183 3183 4217 3193
rect 4183 3125 4217 3145
rect 4183 3111 4217 3125
rect 6103 3635 6137 3649
rect 6103 3615 6137 3635
rect 6103 3567 6137 3577
rect 6103 3543 6137 3567
rect 6103 3499 6137 3505
rect 6103 3471 6137 3499
rect 6103 3431 6137 3433
rect 6103 3399 6137 3431
rect 6103 3329 6137 3361
rect 6103 3327 6137 3329
rect 6103 3261 6137 3289
rect 6103 3255 6137 3261
rect 6103 3193 6137 3217
rect 6103 3183 6137 3193
rect 6103 3125 6137 3145
rect 6103 3111 6137 3125
rect 8023 3635 8057 3649
rect 8023 3615 8057 3635
rect 8023 3567 8057 3577
rect 8023 3543 8057 3567
rect 8023 3499 8057 3505
rect 8023 3471 8057 3499
rect 8023 3431 8057 3433
rect 8023 3399 8057 3431
rect 8023 3329 8057 3361
rect 8023 3327 8057 3329
rect 8023 3261 8057 3289
rect 8023 3255 8057 3261
rect 8023 3193 8057 3217
rect 8023 3183 8057 3193
rect 8023 3125 8057 3145
rect 8023 3111 8057 3125
rect 547 2983 555 3017
rect 555 2983 581 3017
rect 619 2983 623 3017
rect 623 2983 653 3017
rect 691 2983 725 3017
rect 763 2983 793 3017
rect 793 2983 797 3017
rect 835 2983 861 3017
rect 861 2983 869 3017
rect 907 2983 929 3017
rect 929 2983 941 3017
rect 979 2983 997 3017
rect 997 2983 1013 3017
rect 1051 2983 1065 3017
rect 1065 2983 1085 3017
rect 1123 2983 1133 3017
rect 1133 2983 1157 3017
rect 1195 2983 1201 3017
rect 1201 2983 1229 3017
rect 1267 2983 1269 3017
rect 1269 2983 1301 3017
rect 1339 2983 1371 3017
rect 1371 2983 1373 3017
rect 1411 2983 1439 3017
rect 1439 2983 1445 3017
rect 1483 2983 1507 3017
rect 1507 2983 1517 3017
rect 1555 2983 1575 3017
rect 1575 2983 1589 3017
rect 1627 2983 1643 3017
rect 1643 2983 1661 3017
rect 1699 2983 1711 3017
rect 1711 2983 1733 3017
rect 1771 2983 1779 3017
rect 1779 2983 1805 3017
rect 1843 2983 1847 3017
rect 1847 2983 1877 3017
rect 1915 2983 1949 3017
rect 1987 2983 2017 3017
rect 2017 2983 2021 3017
rect 2059 2983 2085 3017
rect 2085 2983 2093 3017
rect 2467 2983 2475 3017
rect 2475 2983 2501 3017
rect 2539 2983 2543 3017
rect 2543 2983 2573 3017
rect 2611 2983 2645 3017
rect 2683 2983 2713 3017
rect 2713 2983 2717 3017
rect 2755 2983 2781 3017
rect 2781 2983 2789 3017
rect 2827 2983 2849 3017
rect 2849 2983 2861 3017
rect 2899 2983 2917 3017
rect 2917 2983 2933 3017
rect 2971 2983 2985 3017
rect 2985 2983 3005 3017
rect 3043 2983 3053 3017
rect 3053 2983 3077 3017
rect 3115 2983 3121 3017
rect 3121 2983 3149 3017
rect 3187 2983 3189 3017
rect 3189 2983 3221 3017
rect 3259 2983 3291 3017
rect 3291 2983 3293 3017
rect 3331 2983 3359 3017
rect 3359 2983 3365 3017
rect 3403 2983 3427 3017
rect 3427 2983 3437 3017
rect 3475 2983 3495 3017
rect 3495 2983 3509 3017
rect 3547 2983 3563 3017
rect 3563 2983 3581 3017
rect 3619 2983 3631 3017
rect 3631 2983 3653 3017
rect 3691 2983 3699 3017
rect 3699 2983 3725 3017
rect 3763 2983 3767 3017
rect 3767 2983 3797 3017
rect 3835 2983 3869 3017
rect 3907 2983 3937 3017
rect 3937 2983 3941 3017
rect 3979 2983 4005 3017
rect 4005 2983 4013 3017
rect 4387 2983 4395 3017
rect 4395 2983 4421 3017
rect 4459 2983 4463 3017
rect 4463 2983 4493 3017
rect 4531 2983 4565 3017
rect 4603 2983 4633 3017
rect 4633 2983 4637 3017
rect 4675 2983 4701 3017
rect 4701 2983 4709 3017
rect 4747 2983 4769 3017
rect 4769 2983 4781 3017
rect 4819 2983 4837 3017
rect 4837 2983 4853 3017
rect 4891 2983 4905 3017
rect 4905 2983 4925 3017
rect 4963 2983 4973 3017
rect 4973 2983 4997 3017
rect 5035 2983 5041 3017
rect 5041 2983 5069 3017
rect 5107 2983 5109 3017
rect 5109 2983 5141 3017
rect 5179 2983 5211 3017
rect 5211 2983 5213 3017
rect 5251 2983 5279 3017
rect 5279 2983 5285 3017
rect 5323 2983 5347 3017
rect 5347 2983 5357 3017
rect 5395 2983 5415 3017
rect 5415 2983 5429 3017
rect 5467 2983 5483 3017
rect 5483 2983 5501 3017
rect 5539 2983 5551 3017
rect 5551 2983 5573 3017
rect 5611 2983 5619 3017
rect 5619 2983 5645 3017
rect 5683 2983 5687 3017
rect 5687 2983 5717 3017
rect 5755 2983 5789 3017
rect 5827 2983 5857 3017
rect 5857 2983 5861 3017
rect 5899 2983 5925 3017
rect 5925 2983 5933 3017
rect 6307 2983 6315 3017
rect 6315 2983 6341 3017
rect 6379 2983 6383 3017
rect 6383 2983 6413 3017
rect 6451 2983 6485 3017
rect 6523 2983 6553 3017
rect 6553 2983 6557 3017
rect 6595 2983 6621 3017
rect 6621 2983 6629 3017
rect 6667 2983 6689 3017
rect 6689 2983 6701 3017
rect 6739 2983 6757 3017
rect 6757 2983 6773 3017
rect 6811 2983 6825 3017
rect 6825 2983 6845 3017
rect 6883 2983 6893 3017
rect 6893 2983 6917 3017
rect 6955 2983 6961 3017
rect 6961 2983 6989 3017
rect 7027 2983 7029 3017
rect 7029 2983 7061 3017
rect 7099 2983 7131 3017
rect 7131 2983 7133 3017
rect 7171 2983 7199 3017
rect 7199 2983 7205 3017
rect 7243 2983 7267 3017
rect 7267 2983 7277 3017
rect 7315 2983 7335 3017
rect 7335 2983 7349 3017
rect 7387 2983 7403 3017
rect 7403 2983 7421 3017
rect 7459 2983 7471 3017
rect 7471 2983 7493 3017
rect 7531 2983 7539 3017
rect 7539 2983 7565 3017
rect 7603 2983 7607 3017
rect 7607 2983 7637 3017
rect 7675 2983 7709 3017
rect 7747 2983 7777 3017
rect 7777 2983 7781 3017
rect 7819 2983 7845 3017
rect 7845 2983 7853 3017
rect 343 2195 377 2209
rect 343 2175 377 2195
rect 343 2127 377 2137
rect 343 2103 377 2127
rect 343 2059 377 2065
rect 343 2031 377 2059
rect 343 1991 377 1993
rect 343 1959 377 1991
rect 343 1889 377 1921
rect 343 1887 377 1889
rect 343 1821 377 1849
rect 343 1815 377 1821
rect 343 1753 377 1777
rect 343 1743 377 1753
rect 343 1685 377 1705
rect 343 1671 377 1685
rect 2263 2195 2297 2209
rect 2263 2175 2297 2195
rect 2263 2127 2297 2137
rect 2263 2103 2297 2127
rect 2263 2059 2297 2065
rect 2263 2031 2297 2059
rect 2263 1991 2297 1993
rect 2263 1959 2297 1991
rect 2263 1889 2297 1921
rect 2263 1887 2297 1889
rect 2263 1821 2297 1849
rect 2263 1815 2297 1821
rect 2263 1753 2297 1777
rect 2263 1743 2297 1753
rect 2263 1685 2297 1705
rect 2263 1671 2297 1685
rect 4183 2195 4217 2209
rect 4183 2175 4217 2195
rect 4183 2127 4217 2137
rect 4183 2103 4217 2127
rect 4183 2059 4217 2065
rect 4183 2031 4217 2059
rect 4183 1991 4217 1993
rect 4183 1959 4217 1991
rect 4183 1889 4217 1921
rect 4183 1887 4217 1889
rect 4183 1821 4217 1849
rect 4183 1815 4217 1821
rect 4183 1753 4217 1777
rect 4183 1743 4217 1753
rect 4183 1685 4217 1705
rect 4183 1671 4217 1685
rect 6103 2195 6137 2209
rect 6103 2175 6137 2195
rect 6103 2127 6137 2137
rect 6103 2103 6137 2127
rect 6103 2059 6137 2065
rect 6103 2031 6137 2059
rect 6103 1991 6137 1993
rect 6103 1959 6137 1991
rect 6103 1889 6137 1921
rect 6103 1887 6137 1889
rect 6103 1821 6137 1849
rect 6103 1815 6137 1821
rect 6103 1753 6137 1777
rect 6103 1743 6137 1753
rect 6103 1685 6137 1705
rect 6103 1671 6137 1685
rect 8023 2195 8057 2209
rect 8023 2175 8057 2195
rect 8023 2127 8057 2137
rect 8023 2103 8057 2127
rect 8023 2059 8057 2065
rect 8023 2031 8057 2059
rect 8023 1991 8057 1993
rect 8023 1959 8057 1991
rect 8023 1889 8057 1921
rect 8023 1887 8057 1889
rect 8023 1821 8057 1849
rect 8023 1815 8057 1821
rect 8023 1753 8057 1777
rect 8023 1743 8057 1753
rect 8023 1685 8057 1705
rect 8023 1671 8057 1685
rect 547 1543 555 1577
rect 555 1543 581 1577
rect 619 1543 623 1577
rect 623 1543 653 1577
rect 691 1543 725 1577
rect 763 1543 793 1577
rect 793 1543 797 1577
rect 835 1543 861 1577
rect 861 1543 869 1577
rect 907 1543 929 1577
rect 929 1543 941 1577
rect 979 1543 997 1577
rect 997 1543 1013 1577
rect 1051 1543 1065 1577
rect 1065 1543 1085 1577
rect 1123 1543 1133 1577
rect 1133 1543 1157 1577
rect 1195 1543 1201 1577
rect 1201 1543 1229 1577
rect 1267 1543 1269 1577
rect 1269 1543 1301 1577
rect 1339 1543 1371 1577
rect 1371 1543 1373 1577
rect 1411 1543 1439 1577
rect 1439 1543 1445 1577
rect 1483 1543 1507 1577
rect 1507 1543 1517 1577
rect 1555 1543 1575 1577
rect 1575 1543 1589 1577
rect 1627 1543 1643 1577
rect 1643 1543 1661 1577
rect 1699 1543 1711 1577
rect 1711 1543 1733 1577
rect 1771 1543 1779 1577
rect 1779 1543 1805 1577
rect 1843 1543 1847 1577
rect 1847 1543 1877 1577
rect 1915 1543 1949 1577
rect 1987 1543 2017 1577
rect 2017 1543 2021 1577
rect 2059 1543 2085 1577
rect 2085 1543 2093 1577
rect 2467 1543 2475 1577
rect 2475 1543 2501 1577
rect 2539 1543 2543 1577
rect 2543 1543 2573 1577
rect 2611 1543 2645 1577
rect 2683 1543 2713 1577
rect 2713 1543 2717 1577
rect 2755 1543 2781 1577
rect 2781 1543 2789 1577
rect 2827 1543 2849 1577
rect 2849 1543 2861 1577
rect 2899 1543 2917 1577
rect 2917 1543 2933 1577
rect 2971 1543 2985 1577
rect 2985 1543 3005 1577
rect 3043 1543 3053 1577
rect 3053 1543 3077 1577
rect 3115 1543 3121 1577
rect 3121 1543 3149 1577
rect 3187 1543 3189 1577
rect 3189 1543 3221 1577
rect 3259 1543 3291 1577
rect 3291 1543 3293 1577
rect 3331 1543 3359 1577
rect 3359 1543 3365 1577
rect 3403 1543 3427 1577
rect 3427 1543 3437 1577
rect 3475 1543 3495 1577
rect 3495 1543 3509 1577
rect 3547 1543 3563 1577
rect 3563 1543 3581 1577
rect 3619 1543 3631 1577
rect 3631 1543 3653 1577
rect 3691 1543 3699 1577
rect 3699 1543 3725 1577
rect 3763 1543 3767 1577
rect 3767 1543 3797 1577
rect 3835 1543 3869 1577
rect 3907 1543 3937 1577
rect 3937 1543 3941 1577
rect 3979 1543 4005 1577
rect 4005 1543 4013 1577
rect 4387 1543 4395 1577
rect 4395 1543 4421 1577
rect 4459 1543 4463 1577
rect 4463 1543 4493 1577
rect 4531 1543 4565 1577
rect 4603 1543 4633 1577
rect 4633 1543 4637 1577
rect 4675 1543 4701 1577
rect 4701 1543 4709 1577
rect 4747 1543 4769 1577
rect 4769 1543 4781 1577
rect 4819 1543 4837 1577
rect 4837 1543 4853 1577
rect 4891 1543 4905 1577
rect 4905 1543 4925 1577
rect 4963 1543 4973 1577
rect 4973 1543 4997 1577
rect 5035 1543 5041 1577
rect 5041 1543 5069 1577
rect 5107 1543 5109 1577
rect 5109 1543 5141 1577
rect 5179 1543 5211 1577
rect 5211 1543 5213 1577
rect 5251 1543 5279 1577
rect 5279 1543 5285 1577
rect 5323 1543 5347 1577
rect 5347 1543 5357 1577
rect 5395 1543 5415 1577
rect 5415 1543 5429 1577
rect 5467 1543 5483 1577
rect 5483 1543 5501 1577
rect 5539 1543 5551 1577
rect 5551 1543 5573 1577
rect 5611 1543 5619 1577
rect 5619 1543 5645 1577
rect 5683 1543 5687 1577
rect 5687 1543 5717 1577
rect 5755 1543 5789 1577
rect 5827 1543 5857 1577
rect 5857 1543 5861 1577
rect 5899 1543 5925 1577
rect 5925 1543 5933 1577
rect 6307 1543 6315 1577
rect 6315 1543 6341 1577
rect 6379 1543 6383 1577
rect 6383 1543 6413 1577
rect 6451 1543 6485 1577
rect 6523 1543 6553 1577
rect 6553 1543 6557 1577
rect 6595 1543 6621 1577
rect 6621 1543 6629 1577
rect 6667 1543 6689 1577
rect 6689 1543 6701 1577
rect 6739 1543 6757 1577
rect 6757 1543 6773 1577
rect 6811 1543 6825 1577
rect 6825 1543 6845 1577
rect 6883 1543 6893 1577
rect 6893 1543 6917 1577
rect 6955 1543 6961 1577
rect 6961 1543 6989 1577
rect 7027 1543 7029 1577
rect 7029 1543 7061 1577
rect 7099 1543 7131 1577
rect 7131 1543 7133 1577
rect 7171 1543 7199 1577
rect 7199 1543 7205 1577
rect 7243 1543 7267 1577
rect 7267 1543 7277 1577
rect 7315 1543 7335 1577
rect 7335 1543 7349 1577
rect 7387 1543 7403 1577
rect 7403 1543 7421 1577
rect 7459 1543 7471 1577
rect 7471 1543 7493 1577
rect 7531 1543 7539 1577
rect 7539 1543 7565 1577
rect 7603 1543 7607 1577
rect 7607 1543 7637 1577
rect 7675 1543 7709 1577
rect 7747 1543 7777 1577
rect 7777 1543 7781 1577
rect 7819 1543 7845 1577
rect 7845 1543 7853 1577
rect 183 903 217 937
rect 343 903 377 937
rect 503 903 537 937
rect 663 903 697 937
rect 823 903 857 937
rect 983 903 1017 937
rect 1143 903 1177 937
rect 1463 903 1497 937
rect 1623 903 1657 937
rect 1783 903 1817 937
rect 1943 903 1977 937
rect 2103 903 2137 937
rect 2263 903 2297 937
rect 2423 903 2457 937
rect 2583 903 2617 937
rect 2743 903 2777 937
rect 2903 903 2937 937
rect 3063 903 3097 937
rect 3383 903 3417 937
rect 3543 903 3577 937
rect 3703 903 3737 937
rect 3863 903 3897 937
rect 4023 903 4057 937
rect 4343 903 4377 937
rect 4503 903 4537 937
rect 4663 903 4697 937
rect 4823 903 4857 937
rect 4983 903 5017 937
rect 5303 903 5337 937
rect 5463 903 5497 937
rect 5623 903 5657 937
rect 5783 903 5817 937
rect 5943 903 5977 937
rect 6103 903 6137 937
rect 6263 903 6297 937
rect 6423 903 6457 937
rect 6583 903 6617 937
rect 6743 903 6777 937
rect 6903 903 6937 937
rect 7223 903 7257 937
rect 7383 903 7417 937
rect 7543 903 7577 937
rect 7703 903 7737 937
rect 7863 903 7897 937
rect 8023 903 8057 937
rect 8183 903 8217 937
rect 547 423 555 457
rect 555 423 581 457
rect 619 423 623 457
rect 623 423 653 457
rect 691 423 725 457
rect 763 423 793 457
rect 793 423 797 457
rect 835 423 861 457
rect 861 423 869 457
rect 907 423 929 457
rect 929 423 941 457
rect 979 423 997 457
rect 997 423 1013 457
rect 1051 423 1065 457
rect 1065 423 1085 457
rect 1123 423 1133 457
rect 1133 423 1157 457
rect 1195 423 1201 457
rect 1201 423 1229 457
rect 1267 423 1269 457
rect 1269 423 1301 457
rect 1339 423 1371 457
rect 1371 423 1373 457
rect 1411 423 1439 457
rect 1439 423 1445 457
rect 1483 423 1507 457
rect 1507 423 1517 457
rect 1555 423 1575 457
rect 1575 423 1589 457
rect 1627 423 1643 457
rect 1643 423 1661 457
rect 1699 423 1711 457
rect 1711 423 1733 457
rect 1771 423 1779 457
rect 1779 423 1805 457
rect 1843 423 1847 457
rect 1847 423 1877 457
rect 1915 423 1949 457
rect 1987 423 2017 457
rect 2017 423 2021 457
rect 2059 423 2085 457
rect 2085 423 2093 457
rect 2467 423 2475 457
rect 2475 423 2501 457
rect 2539 423 2543 457
rect 2543 423 2573 457
rect 2611 423 2645 457
rect 2683 423 2713 457
rect 2713 423 2717 457
rect 2755 423 2781 457
rect 2781 423 2789 457
rect 2827 423 2849 457
rect 2849 423 2861 457
rect 2899 423 2917 457
rect 2917 423 2933 457
rect 2971 423 2985 457
rect 2985 423 3005 457
rect 3043 423 3053 457
rect 3053 423 3077 457
rect 3115 423 3121 457
rect 3121 423 3149 457
rect 3187 423 3189 457
rect 3189 423 3221 457
rect 3259 423 3291 457
rect 3291 423 3293 457
rect 3331 423 3359 457
rect 3359 423 3365 457
rect 3403 423 3427 457
rect 3427 423 3437 457
rect 3475 423 3495 457
rect 3495 423 3509 457
rect 3547 423 3563 457
rect 3563 423 3581 457
rect 3619 423 3631 457
rect 3631 423 3653 457
rect 3691 423 3699 457
rect 3699 423 3725 457
rect 3763 423 3767 457
rect 3767 423 3797 457
rect 3835 423 3869 457
rect 3907 423 3937 457
rect 3937 423 3941 457
rect 3979 423 4005 457
rect 4005 423 4013 457
rect 4387 423 4395 457
rect 4395 423 4421 457
rect 4459 423 4463 457
rect 4463 423 4493 457
rect 4531 423 4565 457
rect 4603 423 4633 457
rect 4633 423 4637 457
rect 4675 423 4701 457
rect 4701 423 4709 457
rect 4747 423 4769 457
rect 4769 423 4781 457
rect 4819 423 4837 457
rect 4837 423 4853 457
rect 4891 423 4905 457
rect 4905 423 4925 457
rect 4963 423 4973 457
rect 4973 423 4997 457
rect 5035 423 5041 457
rect 5041 423 5069 457
rect 5107 423 5109 457
rect 5109 423 5141 457
rect 5179 423 5211 457
rect 5211 423 5213 457
rect 5251 423 5279 457
rect 5279 423 5285 457
rect 5323 423 5347 457
rect 5347 423 5357 457
rect 5395 423 5415 457
rect 5415 423 5429 457
rect 5467 423 5483 457
rect 5483 423 5501 457
rect 5539 423 5551 457
rect 5551 423 5573 457
rect 5611 423 5619 457
rect 5619 423 5645 457
rect 5683 423 5687 457
rect 5687 423 5717 457
rect 5755 423 5789 457
rect 5827 423 5857 457
rect 5857 423 5861 457
rect 5899 423 5925 457
rect 5925 423 5933 457
rect 6307 423 6315 457
rect 6315 423 6341 457
rect 6379 423 6383 457
rect 6383 423 6413 457
rect 6451 423 6485 457
rect 6523 423 6553 457
rect 6553 423 6557 457
rect 6595 423 6621 457
rect 6621 423 6629 457
rect 6667 423 6689 457
rect 6689 423 6701 457
rect 6739 423 6757 457
rect 6757 423 6773 457
rect 6811 423 6825 457
rect 6825 423 6845 457
rect 6883 423 6893 457
rect 6893 423 6917 457
rect 6955 423 6961 457
rect 6961 423 6989 457
rect 7027 423 7029 457
rect 7029 423 7061 457
rect 7099 423 7131 457
rect 7131 423 7133 457
rect 7171 423 7199 457
rect 7199 423 7205 457
rect 7243 423 7267 457
rect 7267 423 7277 457
rect 7315 423 7335 457
rect 7335 423 7349 457
rect 7387 423 7403 457
rect 7403 423 7421 457
rect 7459 423 7471 457
rect 7471 423 7493 457
rect 7531 423 7539 457
rect 7539 423 7565 457
rect 7603 423 7607 457
rect 7607 423 7637 457
rect 7675 423 7709 457
rect 7747 423 7777 457
rect 7777 423 7781 457
rect 7819 423 7845 457
rect 7845 423 7853 457
rect 343 311 377 313
rect 343 279 377 311
rect 343 209 377 241
rect 343 207 377 209
rect 2263 311 2297 313
rect 2263 279 2297 311
rect 2263 209 2297 241
rect 2263 207 2297 209
rect 4183 311 4217 313
rect 4183 279 4217 311
rect 4183 209 4217 241
rect 4183 207 4217 209
rect 6103 311 6137 313
rect 6103 279 6137 311
rect 6103 209 6137 241
rect 6103 207 6137 209
rect 8023 311 8057 313
rect 8023 279 8057 311
rect 8023 209 8057 241
rect 8023 207 8057 209
<< metal1 >>
rect 320 3649 400 3680
rect 320 3615 343 3649
rect 377 3615 400 3649
rect 320 3577 400 3615
rect 320 3543 343 3577
rect 377 3543 400 3577
rect 320 3505 400 3543
rect 320 3471 343 3505
rect 377 3471 400 3505
rect 320 3433 400 3471
rect 320 3399 343 3433
rect 377 3399 400 3433
rect 320 3361 400 3399
rect 320 3327 343 3361
rect 377 3327 400 3361
rect 320 3289 400 3327
rect 320 3255 343 3289
rect 377 3255 400 3289
rect 320 3217 400 3255
rect 320 3183 343 3217
rect 377 3183 400 3217
rect 320 3145 400 3183
rect 320 3111 343 3145
rect 377 3111 400 3145
rect 0 2786 80 2800
rect 0 2734 14 2786
rect 66 2734 80 2786
rect 0 2466 80 2734
rect 0 2414 14 2466
rect 66 2414 80 2466
rect 0 2400 80 2414
rect 160 2786 240 2800
rect 160 2734 174 2786
rect 226 2734 240 2786
rect 160 2466 240 2734
rect 160 2414 174 2466
rect 226 2414 240 2466
rect 160 2400 240 2414
rect 320 2786 400 3111
rect 2240 3649 2320 3680
rect 2240 3615 2263 3649
rect 2297 3615 2320 3649
rect 2240 3577 2320 3615
rect 2240 3543 2263 3577
rect 2297 3543 2320 3577
rect 2240 3505 2320 3543
rect 2240 3471 2263 3505
rect 2297 3471 2320 3505
rect 2240 3433 2320 3471
rect 2240 3399 2263 3433
rect 2297 3399 2320 3433
rect 2240 3361 2320 3399
rect 2240 3327 2263 3361
rect 2297 3327 2320 3361
rect 2240 3289 2320 3327
rect 2240 3255 2263 3289
rect 2297 3255 2320 3289
rect 2240 3217 2320 3255
rect 2240 3183 2263 3217
rect 2297 3183 2320 3217
rect 2240 3145 2320 3183
rect 2240 3111 2263 3145
rect 2297 3111 2320 3145
rect 2240 3080 2320 3111
rect 4160 3649 4240 3680
rect 4160 3634 4183 3649
rect 4217 3634 4240 3649
rect 4160 3582 4174 3634
rect 4226 3582 4240 3634
rect 4160 3577 4240 3582
rect 4160 3570 4183 3577
rect 4217 3570 4240 3577
rect 4160 3518 4174 3570
rect 4226 3518 4240 3570
rect 4160 3506 4240 3518
rect 4160 3454 4174 3506
rect 4226 3454 4240 3506
rect 4160 3442 4240 3454
rect 4160 3390 4174 3442
rect 4226 3390 4240 3442
rect 4160 3378 4240 3390
rect 4160 3326 4174 3378
rect 4226 3326 4240 3378
rect 4160 3289 4240 3326
rect 4160 3255 4183 3289
rect 4217 3255 4240 3289
rect 4160 3217 4240 3255
rect 4160 3183 4183 3217
rect 4217 3183 4240 3217
rect 4160 3145 4240 3183
rect 4160 3111 4183 3145
rect 4217 3111 4240 3145
rect 4160 3080 4240 3111
rect 6080 3649 6160 3680
rect 6080 3615 6103 3649
rect 6137 3615 6160 3649
rect 6080 3577 6160 3615
rect 6080 3543 6103 3577
rect 6137 3543 6160 3577
rect 6080 3505 6160 3543
rect 6080 3471 6103 3505
rect 6137 3471 6160 3505
rect 6080 3433 6160 3471
rect 6080 3399 6103 3433
rect 6137 3399 6160 3433
rect 6080 3361 6160 3399
rect 6080 3327 6103 3361
rect 6137 3327 6160 3361
rect 6080 3289 6160 3327
rect 6080 3255 6103 3289
rect 6137 3255 6160 3289
rect 6080 3217 6160 3255
rect 6080 3183 6103 3217
rect 6137 3183 6160 3217
rect 6080 3145 6160 3183
rect 6080 3111 6103 3145
rect 6137 3111 6160 3145
rect 6080 3080 6160 3111
rect 8000 3649 8080 3680
rect 8000 3615 8023 3649
rect 8057 3615 8080 3649
rect 8000 3577 8080 3615
rect 8000 3543 8023 3577
rect 8057 3543 8080 3577
rect 8000 3505 8080 3543
rect 8000 3471 8023 3505
rect 8057 3471 8080 3505
rect 8000 3433 8080 3471
rect 8000 3399 8023 3433
rect 8057 3399 8080 3433
rect 8000 3361 8080 3399
rect 8000 3327 8023 3361
rect 8057 3327 8080 3361
rect 8000 3289 8080 3327
rect 8000 3255 8023 3289
rect 8057 3255 8080 3289
rect 8000 3217 8080 3255
rect 8000 3183 8023 3217
rect 8057 3183 8080 3217
rect 8000 3145 8080 3183
rect 8000 3111 8023 3145
rect 8057 3111 8080 3145
rect 520 3017 2120 3040
rect 520 2983 547 3017
rect 581 2983 619 3017
rect 653 2983 691 3017
rect 725 2983 763 3017
rect 797 2983 835 3017
rect 869 2983 907 3017
rect 941 2983 979 3017
rect 1013 2983 1051 3017
rect 1085 2983 1123 3017
rect 1157 2983 1195 3017
rect 1229 2983 1267 3017
rect 1301 2983 1339 3017
rect 1373 2983 1411 3017
rect 1445 2983 1483 3017
rect 1517 2983 1555 3017
rect 1589 2983 1627 3017
rect 1661 2983 1699 3017
rect 1733 2983 1771 3017
rect 1805 2983 1843 3017
rect 1877 2983 1915 3017
rect 1949 2983 1987 3017
rect 2021 2983 2059 3017
rect 2093 2983 2120 3017
rect 520 2960 2120 2983
rect 2440 3017 4040 3040
rect 2440 2983 2467 3017
rect 2501 2983 2539 3017
rect 2573 2983 2611 3017
rect 2645 2983 2683 3017
rect 2717 2983 2755 3017
rect 2789 2983 2827 3017
rect 2861 2983 2899 3017
rect 2933 2983 2971 3017
rect 3005 2983 3043 3017
rect 3077 2983 3115 3017
rect 3149 2983 3187 3017
rect 3221 2983 3259 3017
rect 3293 2983 3331 3017
rect 3365 2983 3403 3017
rect 3437 2983 3475 3017
rect 3509 2983 3547 3017
rect 3581 2983 3619 3017
rect 3653 2983 3691 3017
rect 3725 2983 3763 3017
rect 3797 2983 3835 3017
rect 3869 2983 3907 3017
rect 3941 2983 3979 3017
rect 4013 2983 4040 3017
rect 2440 2960 4040 2983
rect 4360 3017 5960 3040
rect 4360 2983 4387 3017
rect 4421 2983 4459 3017
rect 4493 2983 4531 3017
rect 4565 2983 4603 3017
rect 4637 2983 4675 3017
rect 4709 2983 4747 3017
rect 4781 2983 4819 3017
rect 4853 2983 4891 3017
rect 4925 2983 4963 3017
rect 4997 2983 5035 3017
rect 5069 2983 5107 3017
rect 5141 2983 5179 3017
rect 5213 2983 5251 3017
rect 5285 2983 5323 3017
rect 5357 2983 5395 3017
rect 5429 2983 5467 3017
rect 5501 2983 5539 3017
rect 5573 2983 5611 3017
rect 5645 2983 5683 3017
rect 5717 2983 5755 3017
rect 5789 2983 5827 3017
rect 5861 2983 5899 3017
rect 5933 2983 5960 3017
rect 4360 2960 5960 2983
rect 6280 3017 7880 3040
rect 6280 2983 6307 3017
rect 6341 2983 6379 3017
rect 6413 2983 6451 3017
rect 6485 2983 6523 3017
rect 6557 2983 6595 3017
rect 6629 2983 6667 3017
rect 6701 2983 6739 3017
rect 6773 2983 6811 3017
rect 6845 2983 6883 3017
rect 6917 2983 6955 3017
rect 6989 2983 7027 3017
rect 7061 2983 7099 3017
rect 7133 2983 7171 3017
rect 7205 2983 7243 3017
rect 7277 2983 7315 3017
rect 7349 2983 7387 3017
rect 7421 2983 7459 3017
rect 7493 2983 7531 3017
rect 7565 2983 7603 3017
rect 7637 2983 7675 3017
rect 7709 2983 7747 3017
rect 7781 2983 7819 3017
rect 7853 2983 7880 3017
rect 6280 2960 7880 2983
rect 320 2734 334 2786
rect 386 2734 400 2786
rect 320 2466 400 2734
rect 320 2414 334 2466
rect 386 2414 400 2466
rect 320 2209 400 2414
rect 480 2786 560 2800
rect 480 2734 494 2786
rect 546 2734 560 2786
rect 480 2466 560 2734
rect 480 2414 494 2466
rect 546 2414 560 2466
rect 480 2400 560 2414
rect 640 2786 720 2800
rect 640 2734 654 2786
rect 706 2734 720 2786
rect 640 2466 720 2734
rect 640 2414 654 2466
rect 706 2414 720 2466
rect 640 2400 720 2414
rect 800 2786 880 2800
rect 800 2734 814 2786
rect 866 2734 880 2786
rect 800 2466 880 2734
rect 800 2414 814 2466
rect 866 2414 880 2466
rect 800 2400 880 2414
rect 960 2786 1040 2800
rect 960 2734 974 2786
rect 1026 2734 1040 2786
rect 960 2466 1040 2734
rect 960 2414 974 2466
rect 1026 2414 1040 2466
rect 960 2400 1040 2414
rect 1120 2786 1200 2800
rect 1120 2734 1134 2786
rect 1186 2734 1200 2786
rect 1120 2466 1200 2734
rect 1280 2626 1360 2960
rect 1280 2574 1294 2626
rect 1346 2574 1360 2626
rect 1280 2560 1360 2574
rect 1440 2786 1520 2800
rect 1440 2734 1454 2786
rect 1506 2734 1520 2786
rect 1120 2414 1134 2466
rect 1186 2414 1200 2466
rect 1120 2400 1200 2414
rect 1440 2466 1520 2734
rect 1440 2414 1454 2466
rect 1506 2414 1520 2466
rect 1440 2400 1520 2414
rect 1600 2786 1680 2800
rect 1600 2734 1614 2786
rect 1666 2734 1680 2786
rect 1600 2466 1680 2734
rect 1600 2414 1614 2466
rect 1666 2414 1680 2466
rect 1600 2400 1680 2414
rect 1760 2786 1840 2800
rect 1760 2734 1774 2786
rect 1826 2734 1840 2786
rect 1760 2466 1840 2734
rect 1760 2414 1774 2466
rect 1826 2414 1840 2466
rect 1760 2400 1840 2414
rect 1920 2786 2000 2800
rect 1920 2734 1934 2786
rect 1986 2734 2000 2786
rect 1920 2466 2000 2734
rect 1920 2414 1934 2466
rect 1986 2414 2000 2466
rect 1920 2400 2000 2414
rect 2080 2786 2160 2800
rect 2080 2734 2094 2786
rect 2146 2734 2160 2786
rect 2080 2466 2160 2734
rect 2080 2414 2094 2466
rect 2146 2414 2160 2466
rect 2080 2400 2160 2414
rect 2240 2786 2320 2800
rect 2240 2734 2254 2786
rect 2306 2734 2320 2786
rect 2240 2466 2320 2734
rect 2240 2414 2254 2466
rect 2306 2414 2320 2466
rect 2240 2400 2320 2414
rect 2400 2786 2480 2800
rect 2400 2734 2414 2786
rect 2466 2734 2480 2786
rect 2400 2466 2480 2734
rect 2400 2414 2414 2466
rect 2466 2414 2480 2466
rect 2400 2400 2480 2414
rect 2560 2786 2640 2800
rect 2560 2734 2574 2786
rect 2626 2734 2640 2786
rect 2560 2466 2640 2734
rect 2560 2414 2574 2466
rect 2626 2414 2640 2466
rect 2560 2400 2640 2414
rect 2720 2786 2800 2800
rect 2720 2734 2734 2786
rect 2786 2734 2800 2786
rect 2720 2466 2800 2734
rect 2720 2414 2734 2466
rect 2786 2414 2800 2466
rect 2720 2400 2800 2414
rect 2880 2786 2960 2800
rect 2880 2734 2894 2786
rect 2946 2734 2960 2786
rect 2880 2466 2960 2734
rect 2880 2414 2894 2466
rect 2946 2414 2960 2466
rect 2880 2400 2960 2414
rect 3040 2786 3120 2800
rect 3040 2734 3054 2786
rect 3106 2734 3120 2786
rect 3040 2466 3120 2734
rect 3200 2626 3280 2960
rect 3200 2574 3214 2626
rect 3266 2574 3280 2626
rect 3200 2560 3280 2574
rect 3360 2786 3440 2800
rect 3360 2734 3374 2786
rect 3426 2734 3440 2786
rect 3040 2414 3054 2466
rect 3106 2414 3120 2466
rect 3040 2400 3120 2414
rect 3360 2466 3440 2734
rect 3360 2414 3374 2466
rect 3426 2414 3440 2466
rect 3360 2400 3440 2414
rect 3520 2786 3600 2800
rect 3520 2734 3534 2786
rect 3586 2734 3600 2786
rect 3520 2466 3600 2734
rect 3520 2414 3534 2466
rect 3586 2414 3600 2466
rect 3520 2400 3600 2414
rect 3680 2786 3760 2800
rect 3680 2734 3694 2786
rect 3746 2734 3760 2786
rect 3680 2466 3760 2734
rect 3680 2414 3694 2466
rect 3746 2414 3760 2466
rect 3680 2400 3760 2414
rect 3840 2786 3920 2800
rect 3840 2734 3854 2786
rect 3906 2734 3920 2786
rect 3840 2466 3920 2734
rect 3840 2414 3854 2466
rect 3906 2414 3920 2466
rect 3840 2400 3920 2414
rect 4000 2786 4080 2800
rect 4000 2734 4014 2786
rect 4066 2734 4080 2786
rect 4000 2466 4080 2734
rect 4000 2414 4014 2466
rect 4066 2414 4080 2466
rect 4000 2400 4080 2414
rect 4160 2786 4240 2800
rect 4160 2734 4174 2786
rect 4226 2734 4240 2786
rect 4160 2466 4240 2734
rect 4160 2414 4174 2466
rect 4226 2414 4240 2466
rect 4160 2400 4240 2414
rect 4320 2786 4400 2800
rect 4320 2734 4334 2786
rect 4386 2734 4400 2786
rect 4320 2466 4400 2734
rect 4320 2414 4334 2466
rect 4386 2414 4400 2466
rect 4320 2400 4400 2414
rect 4480 2786 4560 2800
rect 4480 2734 4494 2786
rect 4546 2734 4560 2786
rect 4480 2466 4560 2734
rect 4480 2414 4494 2466
rect 4546 2414 4560 2466
rect 4480 2400 4560 2414
rect 4640 2786 4720 2800
rect 4640 2734 4654 2786
rect 4706 2734 4720 2786
rect 4640 2466 4720 2734
rect 4640 2414 4654 2466
rect 4706 2414 4720 2466
rect 4640 2400 4720 2414
rect 4800 2786 4880 2800
rect 4800 2734 4814 2786
rect 4866 2734 4880 2786
rect 4800 2466 4880 2734
rect 4800 2414 4814 2466
rect 4866 2414 4880 2466
rect 4800 2400 4880 2414
rect 4960 2786 5040 2800
rect 4960 2734 4974 2786
rect 5026 2734 5040 2786
rect 4960 2466 5040 2734
rect 5120 2626 5200 2960
rect 5120 2574 5134 2626
rect 5186 2574 5200 2626
rect 5120 2560 5200 2574
rect 5280 2786 5360 2800
rect 5280 2734 5294 2786
rect 5346 2734 5360 2786
rect 4960 2414 4974 2466
rect 5026 2414 5040 2466
rect 4960 2400 5040 2414
rect 5280 2466 5360 2734
rect 5280 2414 5294 2466
rect 5346 2414 5360 2466
rect 5280 2400 5360 2414
rect 5440 2786 5520 2800
rect 5440 2734 5454 2786
rect 5506 2734 5520 2786
rect 5440 2466 5520 2734
rect 5440 2414 5454 2466
rect 5506 2414 5520 2466
rect 5440 2400 5520 2414
rect 5600 2786 5680 2800
rect 5600 2734 5614 2786
rect 5666 2734 5680 2786
rect 5600 2466 5680 2734
rect 5600 2414 5614 2466
rect 5666 2414 5680 2466
rect 5600 2400 5680 2414
rect 5760 2786 5840 2800
rect 5760 2734 5774 2786
rect 5826 2734 5840 2786
rect 5760 2466 5840 2734
rect 5760 2414 5774 2466
rect 5826 2414 5840 2466
rect 5760 2400 5840 2414
rect 5920 2786 6000 2800
rect 5920 2734 5934 2786
rect 5986 2734 6000 2786
rect 5920 2466 6000 2734
rect 5920 2414 5934 2466
rect 5986 2414 6000 2466
rect 5920 2400 6000 2414
rect 6080 2786 6160 2800
rect 6080 2734 6094 2786
rect 6146 2734 6160 2786
rect 6080 2466 6160 2734
rect 6080 2414 6094 2466
rect 6146 2414 6160 2466
rect 6080 2400 6160 2414
rect 6240 2786 6320 2800
rect 6240 2734 6254 2786
rect 6306 2734 6320 2786
rect 6240 2466 6320 2734
rect 6240 2414 6254 2466
rect 6306 2414 6320 2466
rect 6240 2400 6320 2414
rect 6400 2786 6480 2800
rect 6400 2734 6414 2786
rect 6466 2734 6480 2786
rect 6400 2466 6480 2734
rect 6400 2414 6414 2466
rect 6466 2414 6480 2466
rect 6400 2400 6480 2414
rect 6560 2786 6640 2800
rect 6560 2734 6574 2786
rect 6626 2734 6640 2786
rect 6560 2466 6640 2734
rect 6560 2414 6574 2466
rect 6626 2414 6640 2466
rect 6560 2400 6640 2414
rect 6720 2786 6800 2800
rect 6720 2734 6734 2786
rect 6786 2734 6800 2786
rect 6720 2466 6800 2734
rect 6720 2414 6734 2466
rect 6786 2414 6800 2466
rect 6720 2400 6800 2414
rect 6880 2786 6960 2800
rect 6880 2734 6894 2786
rect 6946 2734 6960 2786
rect 6880 2466 6960 2734
rect 7040 2626 7120 2960
rect 7040 2574 7054 2626
rect 7106 2574 7120 2626
rect 7040 2560 7120 2574
rect 7200 2786 7280 2800
rect 7200 2734 7214 2786
rect 7266 2734 7280 2786
rect 6880 2414 6894 2466
rect 6946 2414 6960 2466
rect 6880 2400 6960 2414
rect 7200 2466 7280 2734
rect 7200 2414 7214 2466
rect 7266 2414 7280 2466
rect 7200 2400 7280 2414
rect 7360 2786 7440 2800
rect 7360 2734 7374 2786
rect 7426 2734 7440 2786
rect 7360 2466 7440 2734
rect 7360 2414 7374 2466
rect 7426 2414 7440 2466
rect 7360 2400 7440 2414
rect 7520 2786 7600 2800
rect 7520 2734 7534 2786
rect 7586 2734 7600 2786
rect 7520 2466 7600 2734
rect 7520 2414 7534 2466
rect 7586 2414 7600 2466
rect 7520 2400 7600 2414
rect 7680 2786 7760 2800
rect 7680 2734 7694 2786
rect 7746 2734 7760 2786
rect 7680 2466 7760 2734
rect 7680 2414 7694 2466
rect 7746 2414 7760 2466
rect 7680 2400 7760 2414
rect 7840 2786 7920 2800
rect 7840 2734 7854 2786
rect 7906 2734 7920 2786
rect 7840 2466 7920 2734
rect 7840 2414 7854 2466
rect 7906 2414 7920 2466
rect 7840 2400 7920 2414
rect 8000 2786 8080 3111
rect 8000 2734 8014 2786
rect 8066 2734 8080 2786
rect 8000 2466 8080 2734
rect 8000 2414 8014 2466
rect 8066 2414 8080 2466
rect 320 2175 343 2209
rect 377 2175 400 2209
rect 320 2137 400 2175
rect 320 2103 343 2137
rect 377 2103 400 2137
rect 320 2065 400 2103
rect 320 2031 343 2065
rect 377 2031 400 2065
rect 320 1993 400 2031
rect 320 1959 343 1993
rect 377 1959 400 1993
rect 320 1921 400 1959
rect 320 1887 343 1921
rect 377 1887 400 1921
rect 320 1849 400 1887
rect 320 1815 343 1849
rect 377 1815 400 1849
rect 320 1777 400 1815
rect 320 1743 343 1777
rect 377 1743 400 1777
rect 320 1705 400 1743
rect 320 1671 343 1705
rect 377 1671 400 1705
rect 320 1640 400 1671
rect 2240 2209 2320 2240
rect 2240 2175 2263 2209
rect 2297 2175 2320 2209
rect 2240 2137 2320 2175
rect 2240 2103 2263 2137
rect 2297 2103 2320 2137
rect 2240 2065 2320 2103
rect 2240 2031 2263 2065
rect 2297 2031 2320 2065
rect 2240 1993 2320 2031
rect 2240 1959 2263 1993
rect 2297 1959 2320 1993
rect 2240 1921 2320 1959
rect 2240 1887 2263 1921
rect 2297 1887 2320 1921
rect 2240 1849 2320 1887
rect 2240 1815 2263 1849
rect 2297 1815 2320 1849
rect 2240 1777 2320 1815
rect 2240 1743 2263 1777
rect 2297 1743 2320 1777
rect 2240 1705 2320 1743
rect 2240 1671 2263 1705
rect 2297 1671 2320 1705
rect 2240 1640 2320 1671
rect 4160 2209 4240 2240
rect 4160 2175 4183 2209
rect 4217 2175 4240 2209
rect 4160 2137 4240 2175
rect 4160 2103 4183 2137
rect 4217 2103 4240 2137
rect 4160 2065 4240 2103
rect 4160 2031 4183 2065
rect 4217 2031 4240 2065
rect 4160 1993 4240 2031
rect 4160 1959 4183 1993
rect 4217 1959 4240 1993
rect 4160 1921 4240 1959
rect 4160 1887 4183 1921
rect 4217 1887 4240 1921
rect 4160 1849 4240 1887
rect 4160 1815 4183 1849
rect 4217 1815 4240 1849
rect 4160 1777 4240 1815
rect 4160 1743 4183 1777
rect 4217 1743 4240 1777
rect 4160 1705 4240 1743
rect 4160 1671 4183 1705
rect 4217 1671 4240 1705
rect 520 1577 2120 1600
rect 520 1543 547 1577
rect 581 1543 619 1577
rect 653 1543 691 1577
rect 725 1543 763 1577
rect 797 1543 835 1577
rect 869 1543 907 1577
rect 941 1543 979 1577
rect 1013 1543 1051 1577
rect 1085 1543 1123 1577
rect 1157 1543 1195 1577
rect 1229 1543 1267 1577
rect 1301 1543 1339 1577
rect 1373 1543 1411 1577
rect 1445 1543 1483 1577
rect 1517 1543 1555 1577
rect 1589 1543 1627 1577
rect 1661 1543 1699 1577
rect 1733 1543 1771 1577
rect 1805 1543 1843 1577
rect 1877 1543 1915 1577
rect 1949 1543 1987 1577
rect 2021 1543 2059 1577
rect 2093 1543 2120 1577
rect 520 1520 2120 1543
rect 2440 1577 4040 1600
rect 2440 1543 2467 1577
rect 2501 1543 2539 1577
rect 2573 1543 2611 1577
rect 2645 1543 2683 1577
rect 2717 1543 2755 1577
rect 2789 1543 2827 1577
rect 2861 1543 2899 1577
rect 2933 1543 2971 1577
rect 3005 1543 3043 1577
rect 3077 1543 3115 1577
rect 3149 1543 3187 1577
rect 3221 1543 3259 1577
rect 3293 1543 3331 1577
rect 3365 1543 3403 1577
rect 3437 1543 3475 1577
rect 3509 1543 3547 1577
rect 3581 1543 3619 1577
rect 3653 1543 3691 1577
rect 3725 1543 3763 1577
rect 3797 1543 3835 1577
rect 3869 1543 3907 1577
rect 3941 1543 3979 1577
rect 4013 1543 4040 1577
rect 2440 1520 4040 1543
rect 1280 1106 1360 1520
rect 1280 1054 1294 1106
rect 1346 1054 1360 1106
rect 160 946 240 960
rect 160 894 174 946
rect 226 894 240 946
rect 160 880 240 894
rect 320 937 400 960
rect 320 903 343 937
rect 377 903 400 937
rect 320 880 400 903
rect 480 937 560 960
rect 480 903 503 937
rect 537 903 560 937
rect 480 880 560 903
rect 640 937 720 960
rect 640 903 663 937
rect 697 903 720 937
rect 640 880 720 903
rect 800 937 880 960
rect 800 903 823 937
rect 857 903 880 937
rect 800 880 880 903
rect 960 937 1040 960
rect 960 903 983 937
rect 1017 903 1040 937
rect 960 880 1040 903
rect 1120 937 1200 960
rect 1120 903 1143 937
rect 1177 903 1200 937
rect 1120 880 1200 903
rect 1280 480 1360 1054
rect 3200 1106 3280 1520
rect 3200 1054 3214 1106
rect 3266 1054 3280 1106
rect 1440 937 1520 960
rect 1440 903 1463 937
rect 1497 903 1520 937
rect 1440 880 1520 903
rect 1600 937 1680 960
rect 1600 903 1623 937
rect 1657 903 1680 937
rect 1600 880 1680 903
rect 1760 937 1840 960
rect 1760 903 1783 937
rect 1817 903 1840 937
rect 1760 880 1840 903
rect 1920 937 2000 960
rect 1920 903 1943 937
rect 1977 903 2000 937
rect 1920 880 2000 903
rect 2080 937 2160 960
rect 2080 903 2103 937
rect 2137 903 2160 937
rect 2080 880 2160 903
rect 2240 937 2320 960
rect 2240 903 2263 937
rect 2297 903 2320 937
rect 2240 880 2320 903
rect 2400 937 2480 960
rect 2400 903 2423 937
rect 2457 903 2480 937
rect 2400 880 2480 903
rect 2560 937 2640 960
rect 2560 903 2583 937
rect 2617 903 2640 937
rect 2560 880 2640 903
rect 2720 937 2800 960
rect 2720 903 2743 937
rect 2777 903 2800 937
rect 2720 880 2800 903
rect 2880 937 2960 960
rect 2880 903 2903 937
rect 2937 903 2960 937
rect 2880 880 2960 903
rect 3040 937 3120 960
rect 3040 903 3063 937
rect 3097 903 3120 937
rect 3040 880 3120 903
rect 3200 480 3280 1054
rect 3360 937 3440 960
rect 3360 903 3383 937
rect 3417 903 3440 937
rect 3360 880 3440 903
rect 3520 937 3600 960
rect 3520 903 3543 937
rect 3577 903 3600 937
rect 3520 880 3600 903
rect 3680 937 3760 960
rect 3680 903 3703 937
rect 3737 903 3760 937
rect 3680 880 3760 903
rect 3840 937 3920 960
rect 3840 903 3863 937
rect 3897 903 3920 937
rect 3840 880 3920 903
rect 4000 937 4080 960
rect 4000 903 4023 937
rect 4057 903 4080 937
rect 4000 880 4080 903
rect 4160 786 4240 1671
rect 6080 2209 6160 2240
rect 6080 2175 6103 2209
rect 6137 2175 6160 2209
rect 6080 2137 6160 2175
rect 6080 2103 6103 2137
rect 6137 2103 6160 2137
rect 6080 2065 6160 2103
rect 6080 2031 6103 2065
rect 6137 2031 6160 2065
rect 6080 1993 6160 2031
rect 6080 1959 6103 1993
rect 6137 1959 6160 1993
rect 6080 1921 6160 1959
rect 6080 1887 6103 1921
rect 6137 1887 6160 1921
rect 6080 1849 6160 1887
rect 6080 1815 6103 1849
rect 6137 1815 6160 1849
rect 6080 1777 6160 1815
rect 6080 1743 6103 1777
rect 6137 1743 6160 1777
rect 6080 1705 6160 1743
rect 6080 1671 6103 1705
rect 6137 1671 6160 1705
rect 6080 1640 6160 1671
rect 8000 2209 8080 2414
rect 8160 2786 8240 2800
rect 8160 2734 8174 2786
rect 8226 2734 8240 2786
rect 8160 2466 8240 2734
rect 8160 2414 8174 2466
rect 8226 2414 8240 2466
rect 8160 2400 8240 2414
rect 8320 2786 8400 2800
rect 8320 2734 8334 2786
rect 8386 2734 8400 2786
rect 8320 2466 8400 2734
rect 8320 2414 8334 2466
rect 8386 2414 8400 2466
rect 8320 2400 8400 2414
rect 8000 2175 8023 2209
rect 8057 2175 8080 2209
rect 8000 2137 8080 2175
rect 8000 2103 8023 2137
rect 8057 2103 8080 2137
rect 8000 2065 8080 2103
rect 8000 2031 8023 2065
rect 8057 2031 8080 2065
rect 8000 1993 8080 2031
rect 8000 1959 8023 1993
rect 8057 1959 8080 1993
rect 8000 1921 8080 1959
rect 8000 1887 8023 1921
rect 8057 1887 8080 1921
rect 8000 1849 8080 1887
rect 8000 1815 8023 1849
rect 8057 1815 8080 1849
rect 8000 1777 8080 1815
rect 8000 1743 8023 1777
rect 8057 1743 8080 1777
rect 8000 1705 8080 1743
rect 8000 1671 8023 1705
rect 8057 1671 8080 1705
rect 8000 1640 8080 1671
rect 4360 1577 5960 1600
rect 4360 1543 4387 1577
rect 4421 1543 4459 1577
rect 4493 1543 4531 1577
rect 4565 1543 4603 1577
rect 4637 1543 4675 1577
rect 4709 1543 4747 1577
rect 4781 1543 4819 1577
rect 4853 1543 4891 1577
rect 4925 1543 4963 1577
rect 4997 1543 5035 1577
rect 5069 1543 5107 1577
rect 5141 1543 5179 1577
rect 5213 1543 5251 1577
rect 5285 1543 5323 1577
rect 5357 1543 5395 1577
rect 5429 1543 5467 1577
rect 5501 1543 5539 1577
rect 5573 1543 5611 1577
rect 5645 1543 5683 1577
rect 5717 1543 5755 1577
rect 5789 1543 5827 1577
rect 5861 1543 5899 1577
rect 5933 1543 5960 1577
rect 4360 1520 5960 1543
rect 6280 1577 7880 1600
rect 6280 1543 6307 1577
rect 6341 1543 6379 1577
rect 6413 1543 6451 1577
rect 6485 1543 6523 1577
rect 6557 1543 6595 1577
rect 6629 1543 6667 1577
rect 6701 1543 6739 1577
rect 6773 1543 6811 1577
rect 6845 1543 6883 1577
rect 6917 1543 6955 1577
rect 6989 1543 7027 1577
rect 7061 1543 7099 1577
rect 7133 1543 7171 1577
rect 7205 1543 7243 1577
rect 7277 1543 7315 1577
rect 7349 1543 7387 1577
rect 7421 1543 7459 1577
rect 7493 1543 7531 1577
rect 7565 1543 7603 1577
rect 7637 1543 7675 1577
rect 7709 1543 7747 1577
rect 7781 1543 7819 1577
rect 7853 1543 7880 1577
rect 6280 1520 7880 1543
rect 5120 1106 5200 1520
rect 5120 1054 5134 1106
rect 5186 1054 5200 1106
rect 4320 937 4400 960
rect 4320 903 4343 937
rect 4377 903 4400 937
rect 4320 880 4400 903
rect 4480 937 4560 960
rect 4480 903 4503 937
rect 4537 903 4560 937
rect 4480 880 4560 903
rect 4640 937 4720 960
rect 4640 903 4663 937
rect 4697 903 4720 937
rect 4640 880 4720 903
rect 4800 937 4880 960
rect 4800 903 4823 937
rect 4857 903 4880 937
rect 4800 880 4880 903
rect 4960 937 5040 960
rect 4960 903 4983 937
rect 5017 903 5040 937
rect 4960 880 5040 903
rect 4160 734 4174 786
rect 4226 734 4240 786
rect 520 457 2120 480
rect 520 423 547 457
rect 581 423 619 457
rect 653 423 691 457
rect 725 423 763 457
rect 797 423 835 457
rect 869 423 907 457
rect 941 423 979 457
rect 1013 423 1051 457
rect 1085 423 1123 457
rect 1157 423 1195 457
rect 1229 423 1267 457
rect 1301 423 1339 457
rect 1373 423 1411 457
rect 1445 423 1483 457
rect 1517 423 1555 457
rect 1589 423 1627 457
rect 1661 423 1699 457
rect 1733 423 1771 457
rect 1805 423 1843 457
rect 1877 423 1915 457
rect 1949 423 1987 457
rect 2021 423 2059 457
rect 2093 423 2120 457
rect 520 400 2120 423
rect 2440 457 4040 480
rect 2440 423 2467 457
rect 2501 423 2539 457
rect 2573 423 2611 457
rect 2645 423 2683 457
rect 2717 423 2755 457
rect 2789 423 2827 457
rect 2861 423 2899 457
rect 2933 423 2971 457
rect 3005 423 3043 457
rect 3077 423 3115 457
rect 3149 423 3187 457
rect 3221 423 3259 457
rect 3293 423 3331 457
rect 3365 423 3403 457
rect 3437 423 3475 457
rect 3509 423 3547 457
rect 3581 423 3619 457
rect 3653 423 3691 457
rect 3725 423 3763 457
rect 3797 423 3835 457
rect 3869 423 3907 457
rect 3941 423 3979 457
rect 4013 423 4040 457
rect 2440 400 4040 423
rect 320 318 400 360
rect 320 266 334 318
rect 386 266 400 318
rect 320 254 400 266
rect 320 202 334 254
rect 386 202 400 254
rect 320 160 400 202
rect 2240 313 2320 360
rect 2240 279 2263 313
rect 2297 279 2320 313
rect 2240 241 2320 279
rect 2240 207 2263 241
rect 2297 207 2320 241
rect 2240 160 2320 207
rect 4160 313 4240 734
rect 5120 480 5200 1054
rect 7040 1106 7120 1520
rect 7040 1054 7054 1106
rect 7106 1054 7120 1106
rect 5280 937 5360 960
rect 5280 903 5303 937
rect 5337 903 5360 937
rect 5280 880 5360 903
rect 5440 937 5520 960
rect 5440 903 5463 937
rect 5497 903 5520 937
rect 5440 880 5520 903
rect 5600 937 5680 960
rect 5600 903 5623 937
rect 5657 903 5680 937
rect 5600 880 5680 903
rect 5760 937 5840 960
rect 5760 903 5783 937
rect 5817 903 5840 937
rect 5760 880 5840 903
rect 5920 937 6000 960
rect 5920 903 5943 937
rect 5977 903 6000 937
rect 5920 880 6000 903
rect 6080 937 6160 960
rect 6080 903 6103 937
rect 6137 903 6160 937
rect 6080 880 6160 903
rect 6240 937 6320 960
rect 6240 903 6263 937
rect 6297 903 6320 937
rect 6240 880 6320 903
rect 6400 937 6480 960
rect 6400 903 6423 937
rect 6457 903 6480 937
rect 6400 880 6480 903
rect 6560 937 6640 960
rect 6560 903 6583 937
rect 6617 903 6640 937
rect 6560 880 6640 903
rect 6720 937 6800 960
rect 6720 903 6743 937
rect 6777 903 6800 937
rect 6720 880 6800 903
rect 6880 937 6960 960
rect 6880 903 6903 937
rect 6937 903 6960 937
rect 6880 880 6960 903
rect 7040 480 7120 1054
rect 7200 937 7280 960
rect 7200 903 7223 937
rect 7257 903 7280 937
rect 7200 880 7280 903
rect 7360 937 7440 960
rect 7360 903 7383 937
rect 7417 903 7440 937
rect 7360 880 7440 903
rect 7520 937 7600 960
rect 7520 903 7543 937
rect 7577 903 7600 937
rect 7520 880 7600 903
rect 7680 937 7760 960
rect 7680 903 7703 937
rect 7737 903 7760 937
rect 7680 880 7760 903
rect 7840 937 7920 960
rect 7840 903 7863 937
rect 7897 903 7920 937
rect 7840 880 7920 903
rect 8000 937 8080 960
rect 8000 903 8023 937
rect 8057 903 8080 937
rect 8000 880 8080 903
rect 8160 937 8240 960
rect 8160 903 8183 937
rect 8217 903 8240 937
rect 8160 880 8240 903
rect 4360 457 5960 480
rect 4360 423 4387 457
rect 4421 423 4459 457
rect 4493 423 4531 457
rect 4565 423 4603 457
rect 4637 423 4675 457
rect 4709 423 4747 457
rect 4781 423 4819 457
rect 4853 423 4891 457
rect 4925 423 4963 457
rect 4997 423 5035 457
rect 5069 423 5107 457
rect 5141 423 5179 457
rect 5213 423 5251 457
rect 5285 423 5323 457
rect 5357 423 5395 457
rect 5429 423 5467 457
rect 5501 423 5539 457
rect 5573 423 5611 457
rect 5645 423 5683 457
rect 5717 423 5755 457
rect 5789 423 5827 457
rect 5861 423 5899 457
rect 5933 423 5960 457
rect 4360 400 5960 423
rect 6280 457 7880 480
rect 6280 423 6307 457
rect 6341 423 6379 457
rect 6413 423 6451 457
rect 6485 423 6523 457
rect 6557 423 6595 457
rect 6629 423 6667 457
rect 6701 423 6739 457
rect 6773 423 6811 457
rect 6845 423 6883 457
rect 6917 423 6955 457
rect 6989 423 7027 457
rect 7061 423 7099 457
rect 7133 423 7171 457
rect 7205 423 7243 457
rect 7277 423 7315 457
rect 7349 423 7387 457
rect 7421 423 7459 457
rect 7493 423 7531 457
rect 7565 423 7603 457
rect 7637 423 7675 457
rect 7709 423 7747 457
rect 7781 423 7819 457
rect 7853 423 7880 457
rect 6280 400 7880 423
rect 4160 279 4183 313
rect 4217 279 4240 313
rect 4160 241 4240 279
rect 4160 207 4183 241
rect 4217 207 4240 241
rect 4160 160 4240 207
rect 6080 313 6160 360
rect 6080 279 6103 313
rect 6137 279 6160 313
rect 6080 241 6160 279
rect 6080 207 6103 241
rect 6137 207 6160 241
rect 6080 160 6160 207
rect 8000 318 8080 360
rect 8000 266 8014 318
rect 8066 266 8080 318
rect 8000 254 8080 266
rect 8000 202 8014 254
rect 8066 202 8080 254
rect 8000 160 8080 202
<< via1 >>
rect 14 2734 66 2786
rect 14 2414 66 2466
rect 174 2734 226 2786
rect 174 2414 226 2466
rect 4174 3615 4183 3634
rect 4183 3615 4217 3634
rect 4217 3615 4226 3634
rect 4174 3582 4226 3615
rect 4174 3543 4183 3570
rect 4183 3543 4217 3570
rect 4217 3543 4226 3570
rect 4174 3518 4226 3543
rect 4174 3505 4226 3506
rect 4174 3471 4183 3505
rect 4183 3471 4217 3505
rect 4217 3471 4226 3505
rect 4174 3454 4226 3471
rect 4174 3433 4226 3442
rect 4174 3399 4183 3433
rect 4183 3399 4217 3433
rect 4217 3399 4226 3433
rect 4174 3390 4226 3399
rect 4174 3361 4226 3378
rect 4174 3327 4183 3361
rect 4183 3327 4217 3361
rect 4217 3327 4226 3361
rect 4174 3326 4226 3327
rect 334 2734 386 2786
rect 334 2414 386 2466
rect 494 2734 546 2786
rect 494 2414 546 2466
rect 654 2734 706 2786
rect 654 2414 706 2466
rect 814 2734 866 2786
rect 814 2414 866 2466
rect 974 2734 1026 2786
rect 974 2414 1026 2466
rect 1134 2734 1186 2786
rect 1294 2574 1346 2626
rect 1454 2734 1506 2786
rect 1134 2414 1186 2466
rect 1454 2414 1506 2466
rect 1614 2734 1666 2786
rect 1614 2414 1666 2466
rect 1774 2734 1826 2786
rect 1774 2414 1826 2466
rect 1934 2734 1986 2786
rect 1934 2414 1986 2466
rect 2094 2734 2146 2786
rect 2094 2414 2146 2466
rect 2254 2734 2306 2786
rect 2254 2414 2306 2466
rect 2414 2734 2466 2786
rect 2414 2414 2466 2466
rect 2574 2734 2626 2786
rect 2574 2414 2626 2466
rect 2734 2734 2786 2786
rect 2734 2414 2786 2466
rect 2894 2734 2946 2786
rect 2894 2414 2946 2466
rect 3054 2734 3106 2786
rect 3214 2574 3266 2626
rect 3374 2734 3426 2786
rect 3054 2414 3106 2466
rect 3374 2414 3426 2466
rect 3534 2734 3586 2786
rect 3534 2414 3586 2466
rect 3694 2734 3746 2786
rect 3694 2414 3746 2466
rect 3854 2734 3906 2786
rect 3854 2414 3906 2466
rect 4014 2734 4066 2786
rect 4014 2414 4066 2466
rect 4174 2734 4226 2786
rect 4174 2414 4226 2466
rect 4334 2734 4386 2786
rect 4334 2414 4386 2466
rect 4494 2734 4546 2786
rect 4494 2414 4546 2466
rect 4654 2734 4706 2786
rect 4654 2414 4706 2466
rect 4814 2734 4866 2786
rect 4814 2414 4866 2466
rect 4974 2734 5026 2786
rect 5134 2574 5186 2626
rect 5294 2734 5346 2786
rect 4974 2414 5026 2466
rect 5294 2414 5346 2466
rect 5454 2734 5506 2786
rect 5454 2414 5506 2466
rect 5614 2734 5666 2786
rect 5614 2414 5666 2466
rect 5774 2734 5826 2786
rect 5774 2414 5826 2466
rect 5934 2734 5986 2786
rect 5934 2414 5986 2466
rect 6094 2734 6146 2786
rect 6094 2414 6146 2466
rect 6254 2734 6306 2786
rect 6254 2414 6306 2466
rect 6414 2734 6466 2786
rect 6414 2414 6466 2466
rect 6574 2734 6626 2786
rect 6574 2414 6626 2466
rect 6734 2734 6786 2786
rect 6734 2414 6786 2466
rect 6894 2734 6946 2786
rect 7054 2574 7106 2626
rect 7214 2734 7266 2786
rect 6894 2414 6946 2466
rect 7214 2414 7266 2466
rect 7374 2734 7426 2786
rect 7374 2414 7426 2466
rect 7534 2734 7586 2786
rect 7534 2414 7586 2466
rect 7694 2734 7746 2786
rect 7694 2414 7746 2466
rect 7854 2734 7906 2786
rect 7854 2414 7906 2466
rect 8014 2734 8066 2786
rect 8014 2414 8066 2466
rect 1294 1054 1346 1106
rect 174 937 226 946
rect 174 903 183 937
rect 183 903 217 937
rect 217 903 226 937
rect 174 894 226 903
rect 3214 1054 3266 1106
rect 8174 2734 8226 2786
rect 8174 2414 8226 2466
rect 8334 2734 8386 2786
rect 8334 2414 8386 2466
rect 5134 1054 5186 1106
rect 4174 734 4226 786
rect 334 313 386 318
rect 334 279 343 313
rect 343 279 377 313
rect 377 279 386 313
rect 334 266 386 279
rect 334 241 386 254
rect 334 207 343 241
rect 343 207 377 241
rect 377 207 386 241
rect 334 202 386 207
rect 7054 1054 7106 1106
rect 8014 313 8066 318
rect 8014 279 8023 313
rect 8023 279 8057 313
rect 8057 279 8066 313
rect 8014 266 8066 279
rect 8014 241 8066 254
rect 8014 207 8023 241
rect 8023 207 8057 241
rect 8057 207 8066 241
rect 8014 202 8066 207
<< metal2 >>
rect 4160 3634 4240 3680
rect 4160 3628 4174 3634
rect 4226 3628 4240 3634
rect 4160 3572 4172 3628
rect 4228 3572 4240 3628
rect 4160 3570 4240 3572
rect 4160 3548 4174 3570
rect 4226 3548 4240 3570
rect 4160 3492 4172 3548
rect 4228 3492 4240 3548
rect 4160 3468 4174 3492
rect 4226 3468 4240 3492
rect 4160 3412 4172 3468
rect 4228 3412 4240 3468
rect 4160 3390 4174 3412
rect 4226 3390 4240 3412
rect 4160 3388 4240 3390
rect 4160 3332 4172 3388
rect 4228 3332 4240 3388
rect 4160 3326 4174 3332
rect 4226 3326 4240 3332
rect 4160 3280 4240 3326
rect 0 2788 8400 2800
rect 0 2732 12 2788
rect 68 2732 172 2788
rect 228 2732 332 2788
rect 388 2732 492 2788
rect 548 2732 652 2788
rect 708 2732 812 2788
rect 868 2732 972 2788
rect 1028 2732 1132 2788
rect 1188 2732 1452 2788
rect 1508 2732 1612 2788
rect 1668 2732 1772 2788
rect 1828 2732 1932 2788
rect 1988 2732 2092 2788
rect 2148 2732 2252 2788
rect 2308 2732 2412 2788
rect 2468 2732 2572 2788
rect 2628 2732 2732 2788
rect 2788 2732 2892 2788
rect 2948 2732 3052 2788
rect 3108 2732 3372 2788
rect 3428 2732 3532 2788
rect 3588 2732 3692 2788
rect 3748 2732 3852 2788
rect 3908 2732 4012 2788
rect 4068 2732 4172 2788
rect 4228 2732 4332 2788
rect 4388 2732 4492 2788
rect 4548 2732 4652 2788
rect 4708 2732 4812 2788
rect 4868 2732 4972 2788
rect 5028 2732 5292 2788
rect 5348 2732 5452 2788
rect 5508 2732 5612 2788
rect 5668 2732 5772 2788
rect 5828 2732 5932 2788
rect 5988 2732 6092 2788
rect 6148 2732 6252 2788
rect 6308 2732 6412 2788
rect 6468 2732 6572 2788
rect 6628 2732 6732 2788
rect 6788 2732 6892 2788
rect 6948 2732 7212 2788
rect 7268 2732 7372 2788
rect 7428 2732 7532 2788
rect 7588 2732 7692 2788
rect 7748 2732 7852 2788
rect 7908 2732 8012 2788
rect 8068 2732 8172 2788
rect 8228 2732 8332 2788
rect 8388 2732 8400 2788
rect 0 2720 8400 2732
rect 0 2626 8400 2640
rect 0 2574 1294 2626
rect 1346 2574 3214 2626
rect 3266 2574 5134 2626
rect 5186 2574 7054 2626
rect 7106 2574 8400 2626
rect 0 2560 8400 2574
rect 0 2468 8400 2480
rect 0 2412 12 2468
rect 68 2412 172 2468
rect 228 2412 332 2468
rect 388 2412 492 2468
rect 548 2412 652 2468
rect 708 2412 812 2468
rect 868 2412 972 2468
rect 1028 2412 1132 2468
rect 1188 2412 1452 2468
rect 1508 2412 1612 2468
rect 1668 2412 1772 2468
rect 1828 2412 1932 2468
rect 1988 2412 2092 2468
rect 2148 2412 2252 2468
rect 2308 2412 2412 2468
rect 2468 2412 2572 2468
rect 2628 2412 2732 2468
rect 2788 2412 2892 2468
rect 2948 2412 3052 2468
rect 3108 2412 3372 2468
rect 3428 2412 3532 2468
rect 3588 2412 3692 2468
rect 3748 2412 3852 2468
rect 3908 2412 4012 2468
rect 4068 2412 4172 2468
rect 4228 2412 4332 2468
rect 4388 2412 4492 2468
rect 4548 2412 4652 2468
rect 4708 2412 4812 2468
rect 4868 2412 4972 2468
rect 5028 2412 5292 2468
rect 5348 2412 5452 2468
rect 5508 2412 5612 2468
rect 5668 2412 5772 2468
rect 5828 2412 5932 2468
rect 5988 2412 6092 2468
rect 6148 2412 6252 2468
rect 6308 2412 6412 2468
rect 6468 2412 6572 2468
rect 6628 2412 6732 2468
rect 6788 2412 6892 2468
rect 6948 2412 7212 2468
rect 7268 2412 7372 2468
rect 7428 2412 7532 2468
rect 7588 2412 7692 2468
rect 7748 2412 7852 2468
rect 7908 2412 8012 2468
rect 8068 2412 8172 2468
rect 8228 2412 8332 2468
rect 8388 2412 8400 2468
rect 0 2400 8400 2412
rect 0 1268 8400 1280
rect 0 1212 172 1268
rect 228 1212 332 1268
rect 388 1212 492 1268
rect 548 1212 652 1268
rect 708 1212 812 1268
rect 868 1212 972 1268
rect 1028 1212 1132 1268
rect 1188 1212 1452 1268
rect 1508 1212 1612 1268
rect 1668 1212 1772 1268
rect 1828 1212 1932 1268
rect 1988 1212 2092 1268
rect 2148 1212 2252 1268
rect 2308 1212 2412 1268
rect 2468 1212 2572 1268
rect 2628 1212 2732 1268
rect 2788 1212 2892 1268
rect 2948 1212 3052 1268
rect 3108 1212 3372 1268
rect 3428 1212 3532 1268
rect 3588 1212 3692 1268
rect 3748 1212 3852 1268
rect 3908 1212 4012 1268
rect 4068 1212 4332 1268
rect 4388 1212 4492 1268
rect 4548 1212 4652 1268
rect 4708 1212 4812 1268
rect 4868 1212 4972 1268
rect 5028 1212 5292 1268
rect 5348 1212 5452 1268
rect 5508 1212 5612 1268
rect 5668 1212 5772 1268
rect 5828 1212 5932 1268
rect 5988 1212 6092 1268
rect 6148 1212 6252 1268
rect 6308 1212 6412 1268
rect 6468 1212 6572 1268
rect 6628 1212 6732 1268
rect 6788 1212 6892 1268
rect 6948 1212 7212 1268
rect 7268 1212 7372 1268
rect 7428 1212 7532 1268
rect 7588 1212 7692 1268
rect 7748 1212 7852 1268
rect 7908 1212 8012 1268
rect 8068 1212 8172 1268
rect 8228 1212 8400 1268
rect 0 1200 8400 1212
rect 0 1106 8400 1120
rect 0 1054 1294 1106
rect 1346 1054 3214 1106
rect 3266 1054 5134 1106
rect 5186 1054 7054 1106
rect 7106 1054 8400 1106
rect 0 1040 8400 1054
rect 0 948 8400 960
rect 0 892 172 948
rect 228 892 332 948
rect 388 892 492 948
rect 548 892 652 948
rect 708 892 812 948
rect 868 892 972 948
rect 1028 892 1132 948
rect 1188 892 1452 948
rect 1508 892 1612 948
rect 1668 892 1772 948
rect 1828 892 1932 948
rect 1988 892 2092 948
rect 2148 892 2252 948
rect 2308 892 2412 948
rect 2468 892 2572 948
rect 2628 892 2732 948
rect 2788 892 2892 948
rect 2948 892 3052 948
rect 3108 892 3372 948
rect 3428 892 3532 948
rect 3588 892 3692 948
rect 3748 892 3852 948
rect 3908 892 4012 948
rect 4068 892 4332 948
rect 4388 892 4492 948
rect 4548 892 4652 948
rect 4708 892 4812 948
rect 4868 892 4972 948
rect 5028 892 5292 948
rect 5348 892 5452 948
rect 5508 892 5612 948
rect 5668 892 5772 948
rect 5828 892 5932 948
rect 5988 892 6092 948
rect 6148 892 6252 948
rect 6308 892 6412 948
rect 6468 892 6572 948
rect 6628 892 6732 948
rect 6788 892 6892 948
rect 6948 892 7212 948
rect 7268 892 7372 948
rect 7428 892 7532 948
rect 7588 892 7692 948
rect 7748 892 7852 948
rect 7908 892 8012 948
rect 8068 892 8172 948
rect 8228 892 8400 948
rect 0 880 8400 892
rect 0 786 8400 800
rect 0 734 4174 786
rect 4226 734 8400 786
rect 0 720 8400 734
rect 0 628 8400 640
rect 0 572 172 628
rect 228 572 332 628
rect 388 572 492 628
rect 548 572 652 628
rect 708 572 812 628
rect 868 572 972 628
rect 1028 572 1132 628
rect 1188 572 1452 628
rect 1508 572 1612 628
rect 1668 572 1772 628
rect 1828 572 1932 628
rect 1988 572 2092 628
rect 2148 572 2252 628
rect 2308 572 2412 628
rect 2468 572 2572 628
rect 2628 572 2732 628
rect 2788 572 2892 628
rect 2948 572 3052 628
rect 3108 572 3372 628
rect 3428 572 3532 628
rect 3588 572 3692 628
rect 3748 572 3852 628
rect 3908 572 4012 628
rect 4068 572 4332 628
rect 4388 572 4492 628
rect 4548 572 4652 628
rect 4708 572 4812 628
rect 4868 572 4972 628
rect 5028 572 5292 628
rect 5348 572 5452 628
rect 5508 572 5612 628
rect 5668 572 5772 628
rect 5828 572 5932 628
rect 5988 572 6092 628
rect 6148 572 6252 628
rect 6308 572 6412 628
rect 6468 572 6572 628
rect 6628 572 6732 628
rect 6788 572 6892 628
rect 6948 572 7212 628
rect 7268 572 7372 628
rect 7428 572 7532 628
rect 7588 572 7692 628
rect 7748 572 7852 628
rect 7908 572 8012 628
rect 8068 572 8172 628
rect 8228 572 8400 628
rect 0 560 8400 572
rect 320 328 400 360
rect 320 272 332 328
rect 388 272 400 328
rect 320 266 334 272
rect 386 266 400 272
rect 320 254 400 266
rect 320 248 334 254
rect 386 248 400 254
rect 320 192 332 248
rect 388 192 400 248
rect 320 160 400 192
rect 8000 328 8080 360
rect 8000 272 8012 328
rect 8068 272 8080 328
rect 8000 266 8014 272
rect 8066 266 8080 272
rect 8000 254 8080 266
rect 8000 248 8014 254
rect 8066 248 8080 254
rect 8000 192 8012 248
rect 8068 192 8080 248
rect 8000 160 8080 192
<< via2 >>
rect 4172 3582 4174 3628
rect 4174 3582 4226 3628
rect 4226 3582 4228 3628
rect 4172 3572 4228 3582
rect 4172 3518 4174 3548
rect 4174 3518 4226 3548
rect 4226 3518 4228 3548
rect 4172 3506 4228 3518
rect 4172 3492 4174 3506
rect 4174 3492 4226 3506
rect 4226 3492 4228 3506
rect 4172 3454 4174 3468
rect 4174 3454 4226 3468
rect 4226 3454 4228 3468
rect 4172 3442 4228 3454
rect 4172 3412 4174 3442
rect 4174 3412 4226 3442
rect 4226 3412 4228 3442
rect 4172 3378 4228 3388
rect 4172 3332 4174 3378
rect 4174 3332 4226 3378
rect 4226 3332 4228 3378
rect 12 2786 68 2788
rect 12 2734 14 2786
rect 14 2734 66 2786
rect 66 2734 68 2786
rect 12 2732 68 2734
rect 172 2786 228 2788
rect 172 2734 174 2786
rect 174 2734 226 2786
rect 226 2734 228 2786
rect 172 2732 228 2734
rect 332 2786 388 2788
rect 332 2734 334 2786
rect 334 2734 386 2786
rect 386 2734 388 2786
rect 332 2732 388 2734
rect 492 2786 548 2788
rect 492 2734 494 2786
rect 494 2734 546 2786
rect 546 2734 548 2786
rect 492 2732 548 2734
rect 652 2786 708 2788
rect 652 2734 654 2786
rect 654 2734 706 2786
rect 706 2734 708 2786
rect 652 2732 708 2734
rect 812 2786 868 2788
rect 812 2734 814 2786
rect 814 2734 866 2786
rect 866 2734 868 2786
rect 812 2732 868 2734
rect 972 2786 1028 2788
rect 972 2734 974 2786
rect 974 2734 1026 2786
rect 1026 2734 1028 2786
rect 972 2732 1028 2734
rect 1132 2786 1188 2788
rect 1132 2734 1134 2786
rect 1134 2734 1186 2786
rect 1186 2734 1188 2786
rect 1132 2732 1188 2734
rect 1452 2786 1508 2788
rect 1452 2734 1454 2786
rect 1454 2734 1506 2786
rect 1506 2734 1508 2786
rect 1452 2732 1508 2734
rect 1612 2786 1668 2788
rect 1612 2734 1614 2786
rect 1614 2734 1666 2786
rect 1666 2734 1668 2786
rect 1612 2732 1668 2734
rect 1772 2786 1828 2788
rect 1772 2734 1774 2786
rect 1774 2734 1826 2786
rect 1826 2734 1828 2786
rect 1772 2732 1828 2734
rect 1932 2786 1988 2788
rect 1932 2734 1934 2786
rect 1934 2734 1986 2786
rect 1986 2734 1988 2786
rect 1932 2732 1988 2734
rect 2092 2786 2148 2788
rect 2092 2734 2094 2786
rect 2094 2734 2146 2786
rect 2146 2734 2148 2786
rect 2092 2732 2148 2734
rect 2252 2786 2308 2788
rect 2252 2734 2254 2786
rect 2254 2734 2306 2786
rect 2306 2734 2308 2786
rect 2252 2732 2308 2734
rect 2412 2786 2468 2788
rect 2412 2734 2414 2786
rect 2414 2734 2466 2786
rect 2466 2734 2468 2786
rect 2412 2732 2468 2734
rect 2572 2786 2628 2788
rect 2572 2734 2574 2786
rect 2574 2734 2626 2786
rect 2626 2734 2628 2786
rect 2572 2732 2628 2734
rect 2732 2786 2788 2788
rect 2732 2734 2734 2786
rect 2734 2734 2786 2786
rect 2786 2734 2788 2786
rect 2732 2732 2788 2734
rect 2892 2786 2948 2788
rect 2892 2734 2894 2786
rect 2894 2734 2946 2786
rect 2946 2734 2948 2786
rect 2892 2732 2948 2734
rect 3052 2786 3108 2788
rect 3052 2734 3054 2786
rect 3054 2734 3106 2786
rect 3106 2734 3108 2786
rect 3052 2732 3108 2734
rect 3372 2786 3428 2788
rect 3372 2734 3374 2786
rect 3374 2734 3426 2786
rect 3426 2734 3428 2786
rect 3372 2732 3428 2734
rect 3532 2786 3588 2788
rect 3532 2734 3534 2786
rect 3534 2734 3586 2786
rect 3586 2734 3588 2786
rect 3532 2732 3588 2734
rect 3692 2786 3748 2788
rect 3692 2734 3694 2786
rect 3694 2734 3746 2786
rect 3746 2734 3748 2786
rect 3692 2732 3748 2734
rect 3852 2786 3908 2788
rect 3852 2734 3854 2786
rect 3854 2734 3906 2786
rect 3906 2734 3908 2786
rect 3852 2732 3908 2734
rect 4012 2786 4068 2788
rect 4012 2734 4014 2786
rect 4014 2734 4066 2786
rect 4066 2734 4068 2786
rect 4012 2732 4068 2734
rect 4172 2786 4228 2788
rect 4172 2734 4174 2786
rect 4174 2734 4226 2786
rect 4226 2734 4228 2786
rect 4172 2732 4228 2734
rect 4332 2786 4388 2788
rect 4332 2734 4334 2786
rect 4334 2734 4386 2786
rect 4386 2734 4388 2786
rect 4332 2732 4388 2734
rect 4492 2786 4548 2788
rect 4492 2734 4494 2786
rect 4494 2734 4546 2786
rect 4546 2734 4548 2786
rect 4492 2732 4548 2734
rect 4652 2786 4708 2788
rect 4652 2734 4654 2786
rect 4654 2734 4706 2786
rect 4706 2734 4708 2786
rect 4652 2732 4708 2734
rect 4812 2786 4868 2788
rect 4812 2734 4814 2786
rect 4814 2734 4866 2786
rect 4866 2734 4868 2786
rect 4812 2732 4868 2734
rect 4972 2786 5028 2788
rect 4972 2734 4974 2786
rect 4974 2734 5026 2786
rect 5026 2734 5028 2786
rect 4972 2732 5028 2734
rect 5292 2786 5348 2788
rect 5292 2734 5294 2786
rect 5294 2734 5346 2786
rect 5346 2734 5348 2786
rect 5292 2732 5348 2734
rect 5452 2786 5508 2788
rect 5452 2734 5454 2786
rect 5454 2734 5506 2786
rect 5506 2734 5508 2786
rect 5452 2732 5508 2734
rect 5612 2786 5668 2788
rect 5612 2734 5614 2786
rect 5614 2734 5666 2786
rect 5666 2734 5668 2786
rect 5612 2732 5668 2734
rect 5772 2786 5828 2788
rect 5772 2734 5774 2786
rect 5774 2734 5826 2786
rect 5826 2734 5828 2786
rect 5772 2732 5828 2734
rect 5932 2786 5988 2788
rect 5932 2734 5934 2786
rect 5934 2734 5986 2786
rect 5986 2734 5988 2786
rect 5932 2732 5988 2734
rect 6092 2786 6148 2788
rect 6092 2734 6094 2786
rect 6094 2734 6146 2786
rect 6146 2734 6148 2786
rect 6092 2732 6148 2734
rect 6252 2786 6308 2788
rect 6252 2734 6254 2786
rect 6254 2734 6306 2786
rect 6306 2734 6308 2786
rect 6252 2732 6308 2734
rect 6412 2786 6468 2788
rect 6412 2734 6414 2786
rect 6414 2734 6466 2786
rect 6466 2734 6468 2786
rect 6412 2732 6468 2734
rect 6572 2786 6628 2788
rect 6572 2734 6574 2786
rect 6574 2734 6626 2786
rect 6626 2734 6628 2786
rect 6572 2732 6628 2734
rect 6732 2786 6788 2788
rect 6732 2734 6734 2786
rect 6734 2734 6786 2786
rect 6786 2734 6788 2786
rect 6732 2732 6788 2734
rect 6892 2786 6948 2788
rect 6892 2734 6894 2786
rect 6894 2734 6946 2786
rect 6946 2734 6948 2786
rect 6892 2732 6948 2734
rect 7212 2786 7268 2788
rect 7212 2734 7214 2786
rect 7214 2734 7266 2786
rect 7266 2734 7268 2786
rect 7212 2732 7268 2734
rect 7372 2786 7428 2788
rect 7372 2734 7374 2786
rect 7374 2734 7426 2786
rect 7426 2734 7428 2786
rect 7372 2732 7428 2734
rect 7532 2786 7588 2788
rect 7532 2734 7534 2786
rect 7534 2734 7586 2786
rect 7586 2734 7588 2786
rect 7532 2732 7588 2734
rect 7692 2786 7748 2788
rect 7692 2734 7694 2786
rect 7694 2734 7746 2786
rect 7746 2734 7748 2786
rect 7692 2732 7748 2734
rect 7852 2786 7908 2788
rect 7852 2734 7854 2786
rect 7854 2734 7906 2786
rect 7906 2734 7908 2786
rect 7852 2732 7908 2734
rect 8012 2786 8068 2788
rect 8012 2734 8014 2786
rect 8014 2734 8066 2786
rect 8066 2734 8068 2786
rect 8012 2732 8068 2734
rect 8172 2786 8228 2788
rect 8172 2734 8174 2786
rect 8174 2734 8226 2786
rect 8226 2734 8228 2786
rect 8172 2732 8228 2734
rect 8332 2786 8388 2788
rect 8332 2734 8334 2786
rect 8334 2734 8386 2786
rect 8386 2734 8388 2786
rect 8332 2732 8388 2734
rect 12 2466 68 2468
rect 12 2414 14 2466
rect 14 2414 66 2466
rect 66 2414 68 2466
rect 12 2412 68 2414
rect 172 2466 228 2468
rect 172 2414 174 2466
rect 174 2414 226 2466
rect 226 2414 228 2466
rect 172 2412 228 2414
rect 332 2466 388 2468
rect 332 2414 334 2466
rect 334 2414 386 2466
rect 386 2414 388 2466
rect 332 2412 388 2414
rect 492 2466 548 2468
rect 492 2414 494 2466
rect 494 2414 546 2466
rect 546 2414 548 2466
rect 492 2412 548 2414
rect 652 2466 708 2468
rect 652 2414 654 2466
rect 654 2414 706 2466
rect 706 2414 708 2466
rect 652 2412 708 2414
rect 812 2466 868 2468
rect 812 2414 814 2466
rect 814 2414 866 2466
rect 866 2414 868 2466
rect 812 2412 868 2414
rect 972 2466 1028 2468
rect 972 2414 974 2466
rect 974 2414 1026 2466
rect 1026 2414 1028 2466
rect 972 2412 1028 2414
rect 1132 2466 1188 2468
rect 1132 2414 1134 2466
rect 1134 2414 1186 2466
rect 1186 2414 1188 2466
rect 1132 2412 1188 2414
rect 1452 2466 1508 2468
rect 1452 2414 1454 2466
rect 1454 2414 1506 2466
rect 1506 2414 1508 2466
rect 1452 2412 1508 2414
rect 1612 2466 1668 2468
rect 1612 2414 1614 2466
rect 1614 2414 1666 2466
rect 1666 2414 1668 2466
rect 1612 2412 1668 2414
rect 1772 2466 1828 2468
rect 1772 2414 1774 2466
rect 1774 2414 1826 2466
rect 1826 2414 1828 2466
rect 1772 2412 1828 2414
rect 1932 2466 1988 2468
rect 1932 2414 1934 2466
rect 1934 2414 1986 2466
rect 1986 2414 1988 2466
rect 1932 2412 1988 2414
rect 2092 2466 2148 2468
rect 2092 2414 2094 2466
rect 2094 2414 2146 2466
rect 2146 2414 2148 2466
rect 2092 2412 2148 2414
rect 2252 2466 2308 2468
rect 2252 2414 2254 2466
rect 2254 2414 2306 2466
rect 2306 2414 2308 2466
rect 2252 2412 2308 2414
rect 2412 2466 2468 2468
rect 2412 2414 2414 2466
rect 2414 2414 2466 2466
rect 2466 2414 2468 2466
rect 2412 2412 2468 2414
rect 2572 2466 2628 2468
rect 2572 2414 2574 2466
rect 2574 2414 2626 2466
rect 2626 2414 2628 2466
rect 2572 2412 2628 2414
rect 2732 2466 2788 2468
rect 2732 2414 2734 2466
rect 2734 2414 2786 2466
rect 2786 2414 2788 2466
rect 2732 2412 2788 2414
rect 2892 2466 2948 2468
rect 2892 2414 2894 2466
rect 2894 2414 2946 2466
rect 2946 2414 2948 2466
rect 2892 2412 2948 2414
rect 3052 2466 3108 2468
rect 3052 2414 3054 2466
rect 3054 2414 3106 2466
rect 3106 2414 3108 2466
rect 3052 2412 3108 2414
rect 3372 2466 3428 2468
rect 3372 2414 3374 2466
rect 3374 2414 3426 2466
rect 3426 2414 3428 2466
rect 3372 2412 3428 2414
rect 3532 2466 3588 2468
rect 3532 2414 3534 2466
rect 3534 2414 3586 2466
rect 3586 2414 3588 2466
rect 3532 2412 3588 2414
rect 3692 2466 3748 2468
rect 3692 2414 3694 2466
rect 3694 2414 3746 2466
rect 3746 2414 3748 2466
rect 3692 2412 3748 2414
rect 3852 2466 3908 2468
rect 3852 2414 3854 2466
rect 3854 2414 3906 2466
rect 3906 2414 3908 2466
rect 3852 2412 3908 2414
rect 4012 2466 4068 2468
rect 4012 2414 4014 2466
rect 4014 2414 4066 2466
rect 4066 2414 4068 2466
rect 4012 2412 4068 2414
rect 4172 2466 4228 2468
rect 4172 2414 4174 2466
rect 4174 2414 4226 2466
rect 4226 2414 4228 2466
rect 4172 2412 4228 2414
rect 4332 2466 4388 2468
rect 4332 2414 4334 2466
rect 4334 2414 4386 2466
rect 4386 2414 4388 2466
rect 4332 2412 4388 2414
rect 4492 2466 4548 2468
rect 4492 2414 4494 2466
rect 4494 2414 4546 2466
rect 4546 2414 4548 2466
rect 4492 2412 4548 2414
rect 4652 2466 4708 2468
rect 4652 2414 4654 2466
rect 4654 2414 4706 2466
rect 4706 2414 4708 2466
rect 4652 2412 4708 2414
rect 4812 2466 4868 2468
rect 4812 2414 4814 2466
rect 4814 2414 4866 2466
rect 4866 2414 4868 2466
rect 4812 2412 4868 2414
rect 4972 2466 5028 2468
rect 4972 2414 4974 2466
rect 4974 2414 5026 2466
rect 5026 2414 5028 2466
rect 4972 2412 5028 2414
rect 5292 2466 5348 2468
rect 5292 2414 5294 2466
rect 5294 2414 5346 2466
rect 5346 2414 5348 2466
rect 5292 2412 5348 2414
rect 5452 2466 5508 2468
rect 5452 2414 5454 2466
rect 5454 2414 5506 2466
rect 5506 2414 5508 2466
rect 5452 2412 5508 2414
rect 5612 2466 5668 2468
rect 5612 2414 5614 2466
rect 5614 2414 5666 2466
rect 5666 2414 5668 2466
rect 5612 2412 5668 2414
rect 5772 2466 5828 2468
rect 5772 2414 5774 2466
rect 5774 2414 5826 2466
rect 5826 2414 5828 2466
rect 5772 2412 5828 2414
rect 5932 2466 5988 2468
rect 5932 2414 5934 2466
rect 5934 2414 5986 2466
rect 5986 2414 5988 2466
rect 5932 2412 5988 2414
rect 6092 2466 6148 2468
rect 6092 2414 6094 2466
rect 6094 2414 6146 2466
rect 6146 2414 6148 2466
rect 6092 2412 6148 2414
rect 6252 2466 6308 2468
rect 6252 2414 6254 2466
rect 6254 2414 6306 2466
rect 6306 2414 6308 2466
rect 6252 2412 6308 2414
rect 6412 2466 6468 2468
rect 6412 2414 6414 2466
rect 6414 2414 6466 2466
rect 6466 2414 6468 2466
rect 6412 2412 6468 2414
rect 6572 2466 6628 2468
rect 6572 2414 6574 2466
rect 6574 2414 6626 2466
rect 6626 2414 6628 2466
rect 6572 2412 6628 2414
rect 6732 2466 6788 2468
rect 6732 2414 6734 2466
rect 6734 2414 6786 2466
rect 6786 2414 6788 2466
rect 6732 2412 6788 2414
rect 6892 2466 6948 2468
rect 6892 2414 6894 2466
rect 6894 2414 6946 2466
rect 6946 2414 6948 2466
rect 6892 2412 6948 2414
rect 7212 2466 7268 2468
rect 7212 2414 7214 2466
rect 7214 2414 7266 2466
rect 7266 2414 7268 2466
rect 7212 2412 7268 2414
rect 7372 2466 7428 2468
rect 7372 2414 7374 2466
rect 7374 2414 7426 2466
rect 7426 2414 7428 2466
rect 7372 2412 7428 2414
rect 7532 2466 7588 2468
rect 7532 2414 7534 2466
rect 7534 2414 7586 2466
rect 7586 2414 7588 2466
rect 7532 2412 7588 2414
rect 7692 2466 7748 2468
rect 7692 2414 7694 2466
rect 7694 2414 7746 2466
rect 7746 2414 7748 2466
rect 7692 2412 7748 2414
rect 7852 2466 7908 2468
rect 7852 2414 7854 2466
rect 7854 2414 7906 2466
rect 7906 2414 7908 2466
rect 7852 2412 7908 2414
rect 8012 2466 8068 2468
rect 8012 2414 8014 2466
rect 8014 2414 8066 2466
rect 8066 2414 8068 2466
rect 8012 2412 8068 2414
rect 8172 2466 8228 2468
rect 8172 2414 8174 2466
rect 8174 2414 8226 2466
rect 8226 2414 8228 2466
rect 8172 2412 8228 2414
rect 8332 2466 8388 2468
rect 8332 2414 8334 2466
rect 8334 2414 8386 2466
rect 8386 2414 8388 2466
rect 8332 2412 8388 2414
rect 172 1212 228 1268
rect 332 1212 388 1268
rect 492 1212 548 1268
rect 652 1212 708 1268
rect 812 1212 868 1268
rect 972 1212 1028 1268
rect 1132 1212 1188 1268
rect 1452 1212 1508 1268
rect 1612 1212 1668 1268
rect 1772 1212 1828 1268
rect 1932 1212 1988 1268
rect 2092 1212 2148 1268
rect 2252 1212 2308 1268
rect 2412 1212 2468 1268
rect 2572 1212 2628 1268
rect 2732 1212 2788 1268
rect 2892 1212 2948 1268
rect 3052 1212 3108 1268
rect 3372 1212 3428 1268
rect 3532 1212 3588 1268
rect 3692 1212 3748 1268
rect 3852 1212 3908 1268
rect 4012 1212 4068 1268
rect 4332 1212 4388 1268
rect 4492 1212 4548 1268
rect 4652 1212 4708 1268
rect 4812 1212 4868 1268
rect 4972 1212 5028 1268
rect 5292 1212 5348 1268
rect 5452 1212 5508 1268
rect 5612 1212 5668 1268
rect 5772 1212 5828 1268
rect 5932 1212 5988 1268
rect 6092 1212 6148 1268
rect 6252 1212 6308 1268
rect 6412 1212 6468 1268
rect 6572 1212 6628 1268
rect 6732 1212 6788 1268
rect 6892 1212 6948 1268
rect 7212 1212 7268 1268
rect 7372 1212 7428 1268
rect 7532 1212 7588 1268
rect 7692 1212 7748 1268
rect 7852 1212 7908 1268
rect 8012 1212 8068 1268
rect 8172 1212 8228 1268
rect 172 946 228 948
rect 172 894 174 946
rect 174 894 226 946
rect 226 894 228 946
rect 172 892 228 894
rect 332 892 388 948
rect 492 892 548 948
rect 652 892 708 948
rect 812 892 868 948
rect 972 892 1028 948
rect 1132 892 1188 948
rect 1452 892 1508 948
rect 1612 892 1668 948
rect 1772 892 1828 948
rect 1932 892 1988 948
rect 2092 892 2148 948
rect 2252 892 2308 948
rect 2412 892 2468 948
rect 2572 892 2628 948
rect 2732 892 2788 948
rect 2892 892 2948 948
rect 3052 892 3108 948
rect 3372 892 3428 948
rect 3532 892 3588 948
rect 3692 892 3748 948
rect 3852 892 3908 948
rect 4012 892 4068 948
rect 4332 892 4388 948
rect 4492 892 4548 948
rect 4652 892 4708 948
rect 4812 892 4868 948
rect 4972 892 5028 948
rect 5292 892 5348 948
rect 5452 892 5508 948
rect 5612 892 5668 948
rect 5772 892 5828 948
rect 5932 892 5988 948
rect 6092 892 6148 948
rect 6252 892 6308 948
rect 6412 892 6468 948
rect 6572 892 6628 948
rect 6732 892 6788 948
rect 6892 892 6948 948
rect 7212 892 7268 948
rect 7372 892 7428 948
rect 7532 892 7588 948
rect 7692 892 7748 948
rect 7852 892 7908 948
rect 8012 892 8068 948
rect 8172 892 8228 948
rect 172 572 228 628
rect 332 572 388 628
rect 492 572 548 628
rect 652 572 708 628
rect 812 572 868 628
rect 972 572 1028 628
rect 1132 572 1188 628
rect 1452 572 1508 628
rect 1612 572 1668 628
rect 1772 572 1828 628
rect 1932 572 1988 628
rect 2092 572 2148 628
rect 2252 572 2308 628
rect 2412 572 2468 628
rect 2572 572 2628 628
rect 2732 572 2788 628
rect 2892 572 2948 628
rect 3052 572 3108 628
rect 3372 572 3428 628
rect 3532 572 3588 628
rect 3692 572 3748 628
rect 3852 572 3908 628
rect 4012 572 4068 628
rect 4332 572 4388 628
rect 4492 572 4548 628
rect 4652 572 4708 628
rect 4812 572 4868 628
rect 4972 572 5028 628
rect 5292 572 5348 628
rect 5452 572 5508 628
rect 5612 572 5668 628
rect 5772 572 5828 628
rect 5932 572 5988 628
rect 6092 572 6148 628
rect 6252 572 6308 628
rect 6412 572 6468 628
rect 6572 572 6628 628
rect 6732 572 6788 628
rect 6892 572 6948 628
rect 7212 572 7268 628
rect 7372 572 7428 628
rect 7532 572 7588 628
rect 7692 572 7748 628
rect 7852 572 7908 628
rect 8012 572 8068 628
rect 8172 572 8228 628
rect 332 318 388 328
rect 332 272 334 318
rect 334 272 386 318
rect 386 272 388 318
rect 332 202 334 248
rect 334 202 386 248
rect 386 202 388 248
rect 332 192 388 202
rect 8012 318 8068 328
rect 8012 272 8014 318
rect 8014 272 8066 318
rect 8066 272 8068 318
rect 8012 202 8014 248
rect 8014 202 8066 248
rect 8066 202 8068 248
rect 8012 192 8068 202
<< metal3 >>
rect 4160 3632 4240 3680
rect 4160 3568 4168 3632
rect 4232 3568 4240 3632
rect 4160 3552 4240 3568
rect 4160 3488 4168 3552
rect 4232 3488 4240 3552
rect 4160 3472 4240 3488
rect 4160 3408 4168 3472
rect 4232 3408 4240 3472
rect 4160 3392 4240 3408
rect 4160 3328 4168 3392
rect 4232 3328 4240 3392
rect 4160 3280 4240 3328
rect 0 2792 80 2800
rect 0 2728 8 2792
rect 72 2728 80 2792
rect 0 2472 80 2728
rect 0 2408 8 2472
rect 72 2408 80 2472
rect 0 2400 80 2408
rect 160 2792 240 2800
rect 160 2728 168 2792
rect 232 2728 240 2792
rect 160 2472 240 2728
rect 160 2408 168 2472
rect 232 2408 240 2472
rect 160 2400 240 2408
rect 320 2792 400 2800
rect 320 2728 328 2792
rect 392 2728 400 2792
rect 320 2472 400 2728
rect 320 2408 328 2472
rect 392 2408 400 2472
rect 320 2400 400 2408
rect 480 2792 560 2800
rect 480 2728 488 2792
rect 552 2728 560 2792
rect 480 2472 560 2728
rect 480 2408 488 2472
rect 552 2408 560 2472
rect 480 2400 560 2408
rect 640 2792 720 2800
rect 640 2728 648 2792
rect 712 2728 720 2792
rect 640 2472 720 2728
rect 640 2408 648 2472
rect 712 2408 720 2472
rect 640 2400 720 2408
rect 800 2792 880 2800
rect 800 2728 808 2792
rect 872 2728 880 2792
rect 800 2472 880 2728
rect 800 2408 808 2472
rect 872 2408 880 2472
rect 800 2400 880 2408
rect 960 2792 1040 2800
rect 960 2728 968 2792
rect 1032 2728 1040 2792
rect 960 2472 1040 2728
rect 960 2408 968 2472
rect 1032 2408 1040 2472
rect 960 2400 1040 2408
rect 1120 2792 1200 2800
rect 1120 2728 1128 2792
rect 1192 2728 1200 2792
rect 1120 2472 1200 2728
rect 1120 2408 1128 2472
rect 1192 2408 1200 2472
rect 1120 2400 1200 2408
rect 1440 2792 1520 2800
rect 1440 2728 1448 2792
rect 1512 2728 1520 2792
rect 1440 2472 1520 2728
rect 1440 2408 1448 2472
rect 1512 2408 1520 2472
rect 1440 2400 1520 2408
rect 1600 2792 1680 2800
rect 1600 2728 1608 2792
rect 1672 2728 1680 2792
rect 1600 2472 1680 2728
rect 1600 2408 1608 2472
rect 1672 2408 1680 2472
rect 1600 2400 1680 2408
rect 1760 2792 1840 2800
rect 1760 2728 1768 2792
rect 1832 2728 1840 2792
rect 1760 2472 1840 2728
rect 1760 2408 1768 2472
rect 1832 2408 1840 2472
rect 1760 2400 1840 2408
rect 1920 2792 2000 2800
rect 1920 2728 1928 2792
rect 1992 2728 2000 2792
rect 1920 2472 2000 2728
rect 1920 2408 1928 2472
rect 1992 2408 2000 2472
rect 1920 2400 2000 2408
rect 2080 2792 2160 2800
rect 2080 2728 2088 2792
rect 2152 2728 2160 2792
rect 2080 2472 2160 2728
rect 2080 2408 2088 2472
rect 2152 2408 2160 2472
rect 2080 2400 2160 2408
rect 2240 2792 2320 2800
rect 2240 2728 2248 2792
rect 2312 2728 2320 2792
rect 2240 2472 2320 2728
rect 2240 2408 2248 2472
rect 2312 2408 2320 2472
rect 2240 2400 2320 2408
rect 2400 2792 2480 2800
rect 2400 2728 2408 2792
rect 2472 2728 2480 2792
rect 2400 2472 2480 2728
rect 2400 2408 2408 2472
rect 2472 2408 2480 2472
rect 2400 2400 2480 2408
rect 2560 2792 2640 2800
rect 2560 2728 2568 2792
rect 2632 2728 2640 2792
rect 2560 2472 2640 2728
rect 2560 2408 2568 2472
rect 2632 2408 2640 2472
rect 2560 2400 2640 2408
rect 2720 2792 2800 2800
rect 2720 2728 2728 2792
rect 2792 2728 2800 2792
rect 2720 2472 2800 2728
rect 2720 2408 2728 2472
rect 2792 2408 2800 2472
rect 2720 2400 2800 2408
rect 2880 2792 2960 2800
rect 2880 2728 2888 2792
rect 2952 2728 2960 2792
rect 2880 2472 2960 2728
rect 2880 2408 2888 2472
rect 2952 2408 2960 2472
rect 2880 2400 2960 2408
rect 3040 2792 3120 2800
rect 3040 2728 3048 2792
rect 3112 2728 3120 2792
rect 3040 2472 3120 2728
rect 3040 2408 3048 2472
rect 3112 2408 3120 2472
rect 3040 2400 3120 2408
rect 3360 2792 3440 2800
rect 3360 2728 3368 2792
rect 3432 2728 3440 2792
rect 3360 2472 3440 2728
rect 3360 2408 3368 2472
rect 3432 2408 3440 2472
rect 3360 2400 3440 2408
rect 3520 2792 3600 2800
rect 3520 2728 3528 2792
rect 3592 2728 3600 2792
rect 3520 2472 3600 2728
rect 3520 2408 3528 2472
rect 3592 2408 3600 2472
rect 3520 2400 3600 2408
rect 3680 2792 3760 2800
rect 3680 2728 3688 2792
rect 3752 2728 3760 2792
rect 3680 2472 3760 2728
rect 3680 2408 3688 2472
rect 3752 2408 3760 2472
rect 3680 2400 3760 2408
rect 3840 2792 3920 2800
rect 3840 2728 3848 2792
rect 3912 2728 3920 2792
rect 3840 2472 3920 2728
rect 3840 2408 3848 2472
rect 3912 2408 3920 2472
rect 3840 2400 3920 2408
rect 4000 2792 4080 2800
rect 4000 2728 4008 2792
rect 4072 2728 4080 2792
rect 4000 2472 4080 2728
rect 4000 2408 4008 2472
rect 4072 2408 4080 2472
rect 4000 2400 4080 2408
rect 4160 2792 4240 2800
rect 4160 2728 4168 2792
rect 4232 2728 4240 2792
rect 4160 2472 4240 2728
rect 4160 2408 4168 2472
rect 4232 2408 4240 2472
rect 4160 2400 4240 2408
rect 4320 2792 4400 2800
rect 4320 2728 4328 2792
rect 4392 2728 4400 2792
rect 4320 2472 4400 2728
rect 4320 2408 4328 2472
rect 4392 2408 4400 2472
rect 4320 2400 4400 2408
rect 4480 2792 4560 2800
rect 4480 2728 4488 2792
rect 4552 2728 4560 2792
rect 4480 2472 4560 2728
rect 4480 2408 4488 2472
rect 4552 2408 4560 2472
rect 4480 2400 4560 2408
rect 4640 2792 4720 2800
rect 4640 2728 4648 2792
rect 4712 2728 4720 2792
rect 4640 2472 4720 2728
rect 4640 2408 4648 2472
rect 4712 2408 4720 2472
rect 4640 2400 4720 2408
rect 4800 2792 4880 2800
rect 4800 2728 4808 2792
rect 4872 2728 4880 2792
rect 4800 2472 4880 2728
rect 4800 2408 4808 2472
rect 4872 2408 4880 2472
rect 4800 2400 4880 2408
rect 4960 2792 5040 2800
rect 4960 2728 4968 2792
rect 5032 2728 5040 2792
rect 4960 2472 5040 2728
rect 4960 2408 4968 2472
rect 5032 2408 5040 2472
rect 4960 2400 5040 2408
rect 5280 2792 5360 2800
rect 5280 2728 5288 2792
rect 5352 2728 5360 2792
rect 5280 2472 5360 2728
rect 5280 2408 5288 2472
rect 5352 2408 5360 2472
rect 5280 2400 5360 2408
rect 5440 2792 5520 2800
rect 5440 2728 5448 2792
rect 5512 2728 5520 2792
rect 5440 2472 5520 2728
rect 5440 2408 5448 2472
rect 5512 2408 5520 2472
rect 5440 2400 5520 2408
rect 5600 2792 5680 2800
rect 5600 2728 5608 2792
rect 5672 2728 5680 2792
rect 5600 2472 5680 2728
rect 5600 2408 5608 2472
rect 5672 2408 5680 2472
rect 5600 2400 5680 2408
rect 5760 2792 5840 2800
rect 5760 2728 5768 2792
rect 5832 2728 5840 2792
rect 5760 2472 5840 2728
rect 5760 2408 5768 2472
rect 5832 2408 5840 2472
rect 5760 2400 5840 2408
rect 5920 2792 6000 2800
rect 5920 2728 5928 2792
rect 5992 2728 6000 2792
rect 5920 2472 6000 2728
rect 5920 2408 5928 2472
rect 5992 2408 6000 2472
rect 5920 2400 6000 2408
rect 6080 2792 6160 2800
rect 6080 2728 6088 2792
rect 6152 2728 6160 2792
rect 6080 2472 6160 2728
rect 6080 2408 6088 2472
rect 6152 2408 6160 2472
rect 6080 2400 6160 2408
rect 6240 2792 6320 2800
rect 6240 2728 6248 2792
rect 6312 2728 6320 2792
rect 6240 2472 6320 2728
rect 6240 2408 6248 2472
rect 6312 2408 6320 2472
rect 6240 2400 6320 2408
rect 6400 2792 6480 2800
rect 6400 2728 6408 2792
rect 6472 2728 6480 2792
rect 6400 2472 6480 2728
rect 6400 2408 6408 2472
rect 6472 2408 6480 2472
rect 6400 2400 6480 2408
rect 6560 2792 6640 2800
rect 6560 2728 6568 2792
rect 6632 2728 6640 2792
rect 6560 2472 6640 2728
rect 6560 2408 6568 2472
rect 6632 2408 6640 2472
rect 6560 2400 6640 2408
rect 6720 2792 6800 2800
rect 6720 2728 6728 2792
rect 6792 2728 6800 2792
rect 6720 2472 6800 2728
rect 6720 2408 6728 2472
rect 6792 2408 6800 2472
rect 6720 2400 6800 2408
rect 6880 2792 6960 2800
rect 6880 2728 6888 2792
rect 6952 2728 6960 2792
rect 6880 2472 6960 2728
rect 6880 2408 6888 2472
rect 6952 2408 6960 2472
rect 6880 2400 6960 2408
rect 7200 2792 7280 2800
rect 7200 2728 7208 2792
rect 7272 2728 7280 2792
rect 7200 2472 7280 2728
rect 7200 2408 7208 2472
rect 7272 2408 7280 2472
rect 7200 2400 7280 2408
rect 7360 2792 7440 2800
rect 7360 2728 7368 2792
rect 7432 2728 7440 2792
rect 7360 2472 7440 2728
rect 7360 2408 7368 2472
rect 7432 2408 7440 2472
rect 7360 2400 7440 2408
rect 7520 2792 7600 2800
rect 7520 2728 7528 2792
rect 7592 2728 7600 2792
rect 7520 2472 7600 2728
rect 7520 2408 7528 2472
rect 7592 2408 7600 2472
rect 7520 2400 7600 2408
rect 7680 2792 7760 2800
rect 7680 2728 7688 2792
rect 7752 2728 7760 2792
rect 7680 2472 7760 2728
rect 7680 2408 7688 2472
rect 7752 2408 7760 2472
rect 7680 2400 7760 2408
rect 7840 2792 7920 2800
rect 7840 2728 7848 2792
rect 7912 2728 7920 2792
rect 7840 2472 7920 2728
rect 7840 2408 7848 2472
rect 7912 2408 7920 2472
rect 7840 2400 7920 2408
rect 8000 2792 8080 2800
rect 8000 2728 8008 2792
rect 8072 2728 8080 2792
rect 8000 2472 8080 2728
rect 8000 2408 8008 2472
rect 8072 2408 8080 2472
rect 8000 2400 8080 2408
rect 8160 2792 8240 2800
rect 8160 2728 8168 2792
rect 8232 2728 8240 2792
rect 8160 2472 8240 2728
rect 8160 2408 8168 2472
rect 8232 2408 8240 2472
rect 8160 2400 8240 2408
rect 8320 2792 8400 2800
rect 8320 2728 8328 2792
rect 8392 2728 8400 2792
rect 8320 2472 8400 2728
rect 8320 2408 8328 2472
rect 8392 2408 8400 2472
rect 8320 2400 8400 2408
rect 160 1268 240 1280
rect 160 1212 172 1268
rect 228 1212 240 1268
rect 160 1112 240 1212
rect 160 1048 168 1112
rect 232 1048 240 1112
rect 160 952 240 1048
rect 160 888 168 952
rect 232 888 240 952
rect 160 792 240 888
rect 160 728 168 792
rect 232 728 240 792
rect 160 628 240 728
rect 160 572 172 628
rect 228 572 240 628
rect 160 560 240 572
rect 320 1268 400 1280
rect 320 1212 332 1268
rect 388 1212 400 1268
rect 320 1112 400 1212
rect 320 1048 328 1112
rect 392 1048 400 1112
rect 320 952 400 1048
rect 320 888 328 952
rect 392 888 400 952
rect 320 792 400 888
rect 320 728 328 792
rect 392 728 400 792
rect 320 628 400 728
rect 320 572 332 628
rect 388 572 400 628
rect 320 560 400 572
rect 480 1268 560 1280
rect 480 1212 492 1268
rect 548 1212 560 1268
rect 480 1112 560 1212
rect 480 1048 488 1112
rect 552 1048 560 1112
rect 480 952 560 1048
rect 480 888 488 952
rect 552 888 560 952
rect 480 792 560 888
rect 480 728 488 792
rect 552 728 560 792
rect 480 628 560 728
rect 480 572 492 628
rect 548 572 560 628
rect 480 560 560 572
rect 640 1268 720 1280
rect 640 1212 652 1268
rect 708 1212 720 1268
rect 640 1112 720 1212
rect 640 1048 648 1112
rect 712 1048 720 1112
rect 640 952 720 1048
rect 640 888 648 952
rect 712 888 720 952
rect 640 792 720 888
rect 640 728 648 792
rect 712 728 720 792
rect 640 628 720 728
rect 640 572 652 628
rect 708 572 720 628
rect 640 560 720 572
rect 800 1268 880 1280
rect 800 1212 812 1268
rect 868 1212 880 1268
rect 800 1112 880 1212
rect 800 1048 808 1112
rect 872 1048 880 1112
rect 800 952 880 1048
rect 800 888 808 952
rect 872 888 880 952
rect 800 792 880 888
rect 800 728 808 792
rect 872 728 880 792
rect 800 628 880 728
rect 800 572 812 628
rect 868 572 880 628
rect 800 560 880 572
rect 960 1268 1040 1280
rect 960 1212 972 1268
rect 1028 1212 1040 1268
rect 960 1112 1040 1212
rect 960 1048 968 1112
rect 1032 1048 1040 1112
rect 960 952 1040 1048
rect 960 888 968 952
rect 1032 888 1040 952
rect 960 792 1040 888
rect 960 728 968 792
rect 1032 728 1040 792
rect 960 628 1040 728
rect 960 572 972 628
rect 1028 572 1040 628
rect 960 560 1040 572
rect 1120 1268 1200 1280
rect 1120 1212 1132 1268
rect 1188 1212 1200 1268
rect 1120 1112 1200 1212
rect 1120 1048 1128 1112
rect 1192 1048 1200 1112
rect 1120 952 1200 1048
rect 1120 888 1128 952
rect 1192 888 1200 952
rect 1120 792 1200 888
rect 1120 728 1128 792
rect 1192 728 1200 792
rect 1120 628 1200 728
rect 1120 572 1132 628
rect 1188 572 1200 628
rect 1120 560 1200 572
rect 1440 1268 1520 1280
rect 1440 1212 1452 1268
rect 1508 1212 1520 1268
rect 1440 1112 1520 1212
rect 1440 1048 1448 1112
rect 1512 1048 1520 1112
rect 1440 952 1520 1048
rect 1440 888 1448 952
rect 1512 888 1520 952
rect 1440 792 1520 888
rect 1440 728 1448 792
rect 1512 728 1520 792
rect 1440 628 1520 728
rect 1440 572 1452 628
rect 1508 572 1520 628
rect 1440 560 1520 572
rect 1600 1268 1680 1280
rect 1600 1212 1612 1268
rect 1668 1212 1680 1268
rect 1600 1112 1680 1212
rect 1600 1048 1608 1112
rect 1672 1048 1680 1112
rect 1600 952 1680 1048
rect 1600 888 1608 952
rect 1672 888 1680 952
rect 1600 792 1680 888
rect 1600 728 1608 792
rect 1672 728 1680 792
rect 1600 628 1680 728
rect 1600 572 1612 628
rect 1668 572 1680 628
rect 1600 560 1680 572
rect 1760 1268 1840 1280
rect 1760 1212 1772 1268
rect 1828 1212 1840 1268
rect 1760 1112 1840 1212
rect 1760 1048 1768 1112
rect 1832 1048 1840 1112
rect 1760 952 1840 1048
rect 1760 888 1768 952
rect 1832 888 1840 952
rect 1760 792 1840 888
rect 1760 728 1768 792
rect 1832 728 1840 792
rect 1760 628 1840 728
rect 1760 572 1772 628
rect 1828 572 1840 628
rect 1760 560 1840 572
rect 1920 1268 2000 1280
rect 1920 1212 1932 1268
rect 1988 1212 2000 1268
rect 1920 1112 2000 1212
rect 1920 1048 1928 1112
rect 1992 1048 2000 1112
rect 1920 952 2000 1048
rect 1920 888 1928 952
rect 1992 888 2000 952
rect 1920 792 2000 888
rect 1920 728 1928 792
rect 1992 728 2000 792
rect 1920 628 2000 728
rect 1920 572 1932 628
rect 1988 572 2000 628
rect 1920 560 2000 572
rect 2080 1268 2160 1280
rect 2080 1212 2092 1268
rect 2148 1212 2160 1268
rect 2080 1112 2160 1212
rect 2080 1048 2088 1112
rect 2152 1048 2160 1112
rect 2080 952 2160 1048
rect 2080 888 2088 952
rect 2152 888 2160 952
rect 2080 792 2160 888
rect 2080 728 2088 792
rect 2152 728 2160 792
rect 2080 628 2160 728
rect 2080 572 2092 628
rect 2148 572 2160 628
rect 2080 560 2160 572
rect 2240 1268 2320 1280
rect 2240 1212 2252 1268
rect 2308 1212 2320 1268
rect 2240 1112 2320 1212
rect 2240 1048 2248 1112
rect 2312 1048 2320 1112
rect 2240 952 2320 1048
rect 2240 888 2248 952
rect 2312 888 2320 952
rect 2240 792 2320 888
rect 2240 728 2248 792
rect 2312 728 2320 792
rect 2240 628 2320 728
rect 2240 572 2252 628
rect 2308 572 2320 628
rect 2240 560 2320 572
rect 2400 1268 2480 1280
rect 2400 1212 2412 1268
rect 2468 1212 2480 1268
rect 2400 1112 2480 1212
rect 2400 1048 2408 1112
rect 2472 1048 2480 1112
rect 2400 952 2480 1048
rect 2400 888 2408 952
rect 2472 888 2480 952
rect 2400 792 2480 888
rect 2400 728 2408 792
rect 2472 728 2480 792
rect 2400 628 2480 728
rect 2400 572 2412 628
rect 2468 572 2480 628
rect 2400 560 2480 572
rect 2560 1268 2640 1280
rect 2560 1212 2572 1268
rect 2628 1212 2640 1268
rect 2560 1112 2640 1212
rect 2560 1048 2568 1112
rect 2632 1048 2640 1112
rect 2560 952 2640 1048
rect 2560 888 2568 952
rect 2632 888 2640 952
rect 2560 792 2640 888
rect 2560 728 2568 792
rect 2632 728 2640 792
rect 2560 628 2640 728
rect 2560 572 2572 628
rect 2628 572 2640 628
rect 2560 560 2640 572
rect 2720 1268 2800 1280
rect 2720 1212 2732 1268
rect 2788 1212 2800 1268
rect 2720 1112 2800 1212
rect 2720 1048 2728 1112
rect 2792 1048 2800 1112
rect 2720 952 2800 1048
rect 2720 888 2728 952
rect 2792 888 2800 952
rect 2720 792 2800 888
rect 2720 728 2728 792
rect 2792 728 2800 792
rect 2720 628 2800 728
rect 2720 572 2732 628
rect 2788 572 2800 628
rect 2720 560 2800 572
rect 2880 1268 2960 1280
rect 2880 1212 2892 1268
rect 2948 1212 2960 1268
rect 2880 1112 2960 1212
rect 2880 1048 2888 1112
rect 2952 1048 2960 1112
rect 2880 952 2960 1048
rect 2880 888 2888 952
rect 2952 888 2960 952
rect 2880 792 2960 888
rect 2880 728 2888 792
rect 2952 728 2960 792
rect 2880 628 2960 728
rect 2880 572 2892 628
rect 2948 572 2960 628
rect 2880 560 2960 572
rect 3040 1268 3120 1280
rect 3040 1212 3052 1268
rect 3108 1212 3120 1268
rect 3040 1112 3120 1212
rect 3040 1048 3048 1112
rect 3112 1048 3120 1112
rect 3040 952 3120 1048
rect 3040 888 3048 952
rect 3112 888 3120 952
rect 3040 792 3120 888
rect 3040 728 3048 792
rect 3112 728 3120 792
rect 3040 628 3120 728
rect 3040 572 3052 628
rect 3108 572 3120 628
rect 3040 560 3120 572
rect 3360 1268 3440 1280
rect 3360 1212 3372 1268
rect 3428 1212 3440 1268
rect 3360 1112 3440 1212
rect 3360 1048 3368 1112
rect 3432 1048 3440 1112
rect 3360 952 3440 1048
rect 3360 888 3368 952
rect 3432 888 3440 952
rect 3360 792 3440 888
rect 3360 728 3368 792
rect 3432 728 3440 792
rect 3360 628 3440 728
rect 3360 572 3372 628
rect 3428 572 3440 628
rect 3360 560 3440 572
rect 3520 1268 3600 1280
rect 3520 1212 3532 1268
rect 3588 1212 3600 1268
rect 3520 1112 3600 1212
rect 3520 1048 3528 1112
rect 3592 1048 3600 1112
rect 3520 952 3600 1048
rect 3520 888 3528 952
rect 3592 888 3600 952
rect 3520 792 3600 888
rect 3520 728 3528 792
rect 3592 728 3600 792
rect 3520 628 3600 728
rect 3520 572 3532 628
rect 3588 572 3600 628
rect 3520 560 3600 572
rect 3680 1268 3760 1280
rect 3680 1212 3692 1268
rect 3748 1212 3760 1268
rect 3680 1112 3760 1212
rect 3680 1048 3688 1112
rect 3752 1048 3760 1112
rect 3680 952 3760 1048
rect 3680 888 3688 952
rect 3752 888 3760 952
rect 3680 792 3760 888
rect 3680 728 3688 792
rect 3752 728 3760 792
rect 3680 628 3760 728
rect 3680 572 3692 628
rect 3748 572 3760 628
rect 3680 560 3760 572
rect 3840 1268 3920 1280
rect 3840 1212 3852 1268
rect 3908 1212 3920 1268
rect 3840 1112 3920 1212
rect 3840 1048 3848 1112
rect 3912 1048 3920 1112
rect 3840 952 3920 1048
rect 3840 888 3848 952
rect 3912 888 3920 952
rect 3840 792 3920 888
rect 3840 728 3848 792
rect 3912 728 3920 792
rect 3840 628 3920 728
rect 3840 572 3852 628
rect 3908 572 3920 628
rect 3840 560 3920 572
rect 4000 1268 4080 1280
rect 4000 1212 4012 1268
rect 4068 1212 4080 1268
rect 4000 1112 4080 1212
rect 4000 1048 4008 1112
rect 4072 1048 4080 1112
rect 4000 952 4080 1048
rect 4000 888 4008 952
rect 4072 888 4080 952
rect 4000 792 4080 888
rect 4000 728 4008 792
rect 4072 728 4080 792
rect 4000 628 4080 728
rect 4000 572 4012 628
rect 4068 572 4080 628
rect 4000 560 4080 572
rect 4320 1268 4400 1280
rect 4320 1212 4332 1268
rect 4388 1212 4400 1268
rect 4320 1112 4400 1212
rect 4320 1048 4328 1112
rect 4392 1048 4400 1112
rect 4320 952 4400 1048
rect 4320 888 4328 952
rect 4392 888 4400 952
rect 4320 792 4400 888
rect 4320 728 4328 792
rect 4392 728 4400 792
rect 4320 628 4400 728
rect 4320 572 4332 628
rect 4388 572 4400 628
rect 4320 560 4400 572
rect 4480 1268 4560 1280
rect 4480 1212 4492 1268
rect 4548 1212 4560 1268
rect 4480 1112 4560 1212
rect 4480 1048 4488 1112
rect 4552 1048 4560 1112
rect 4480 952 4560 1048
rect 4480 888 4488 952
rect 4552 888 4560 952
rect 4480 792 4560 888
rect 4480 728 4488 792
rect 4552 728 4560 792
rect 4480 628 4560 728
rect 4480 572 4492 628
rect 4548 572 4560 628
rect 4480 560 4560 572
rect 4640 1268 4720 1280
rect 4640 1212 4652 1268
rect 4708 1212 4720 1268
rect 4640 1112 4720 1212
rect 4640 1048 4648 1112
rect 4712 1048 4720 1112
rect 4640 952 4720 1048
rect 4640 888 4648 952
rect 4712 888 4720 952
rect 4640 792 4720 888
rect 4640 728 4648 792
rect 4712 728 4720 792
rect 4640 628 4720 728
rect 4640 572 4652 628
rect 4708 572 4720 628
rect 4640 560 4720 572
rect 4800 1268 4880 1280
rect 4800 1212 4812 1268
rect 4868 1212 4880 1268
rect 4800 1112 4880 1212
rect 4800 1048 4808 1112
rect 4872 1048 4880 1112
rect 4800 952 4880 1048
rect 4800 888 4808 952
rect 4872 888 4880 952
rect 4800 792 4880 888
rect 4800 728 4808 792
rect 4872 728 4880 792
rect 4800 628 4880 728
rect 4800 572 4812 628
rect 4868 572 4880 628
rect 4800 560 4880 572
rect 4960 1268 5040 1280
rect 4960 1212 4972 1268
rect 5028 1212 5040 1268
rect 4960 1112 5040 1212
rect 4960 1048 4968 1112
rect 5032 1048 5040 1112
rect 4960 952 5040 1048
rect 4960 888 4968 952
rect 5032 888 5040 952
rect 4960 792 5040 888
rect 4960 728 4968 792
rect 5032 728 5040 792
rect 4960 628 5040 728
rect 4960 572 4972 628
rect 5028 572 5040 628
rect 4960 560 5040 572
rect 5280 1268 5360 1280
rect 5280 1212 5292 1268
rect 5348 1212 5360 1268
rect 5280 1112 5360 1212
rect 5280 1048 5288 1112
rect 5352 1048 5360 1112
rect 5280 952 5360 1048
rect 5280 888 5288 952
rect 5352 888 5360 952
rect 5280 792 5360 888
rect 5280 728 5288 792
rect 5352 728 5360 792
rect 5280 628 5360 728
rect 5280 572 5292 628
rect 5348 572 5360 628
rect 5280 560 5360 572
rect 5440 1268 5520 1280
rect 5440 1212 5452 1268
rect 5508 1212 5520 1268
rect 5440 1112 5520 1212
rect 5440 1048 5448 1112
rect 5512 1048 5520 1112
rect 5440 952 5520 1048
rect 5440 888 5448 952
rect 5512 888 5520 952
rect 5440 792 5520 888
rect 5440 728 5448 792
rect 5512 728 5520 792
rect 5440 628 5520 728
rect 5440 572 5452 628
rect 5508 572 5520 628
rect 5440 560 5520 572
rect 5600 1268 5680 1280
rect 5600 1212 5612 1268
rect 5668 1212 5680 1268
rect 5600 1112 5680 1212
rect 5600 1048 5608 1112
rect 5672 1048 5680 1112
rect 5600 952 5680 1048
rect 5600 888 5608 952
rect 5672 888 5680 952
rect 5600 792 5680 888
rect 5600 728 5608 792
rect 5672 728 5680 792
rect 5600 628 5680 728
rect 5600 572 5612 628
rect 5668 572 5680 628
rect 5600 560 5680 572
rect 5760 1268 5840 1280
rect 5760 1212 5772 1268
rect 5828 1212 5840 1268
rect 5760 1112 5840 1212
rect 5760 1048 5768 1112
rect 5832 1048 5840 1112
rect 5760 952 5840 1048
rect 5760 888 5768 952
rect 5832 888 5840 952
rect 5760 792 5840 888
rect 5760 728 5768 792
rect 5832 728 5840 792
rect 5760 628 5840 728
rect 5760 572 5772 628
rect 5828 572 5840 628
rect 5760 560 5840 572
rect 5920 1268 6000 1280
rect 5920 1212 5932 1268
rect 5988 1212 6000 1268
rect 5920 1112 6000 1212
rect 5920 1048 5928 1112
rect 5992 1048 6000 1112
rect 5920 952 6000 1048
rect 5920 888 5928 952
rect 5992 888 6000 952
rect 5920 792 6000 888
rect 5920 728 5928 792
rect 5992 728 6000 792
rect 5920 628 6000 728
rect 5920 572 5932 628
rect 5988 572 6000 628
rect 5920 560 6000 572
rect 6080 1268 6160 1280
rect 6080 1212 6092 1268
rect 6148 1212 6160 1268
rect 6080 1112 6160 1212
rect 6080 1048 6088 1112
rect 6152 1048 6160 1112
rect 6080 952 6160 1048
rect 6080 888 6088 952
rect 6152 888 6160 952
rect 6080 792 6160 888
rect 6080 728 6088 792
rect 6152 728 6160 792
rect 6080 628 6160 728
rect 6080 572 6092 628
rect 6148 572 6160 628
rect 6080 560 6160 572
rect 6240 1268 6320 1280
rect 6240 1212 6252 1268
rect 6308 1212 6320 1268
rect 6240 1112 6320 1212
rect 6240 1048 6248 1112
rect 6312 1048 6320 1112
rect 6240 952 6320 1048
rect 6240 888 6248 952
rect 6312 888 6320 952
rect 6240 792 6320 888
rect 6240 728 6248 792
rect 6312 728 6320 792
rect 6240 628 6320 728
rect 6240 572 6252 628
rect 6308 572 6320 628
rect 6240 560 6320 572
rect 6400 1268 6480 1280
rect 6400 1212 6412 1268
rect 6468 1212 6480 1268
rect 6400 1112 6480 1212
rect 6400 1048 6408 1112
rect 6472 1048 6480 1112
rect 6400 952 6480 1048
rect 6400 888 6408 952
rect 6472 888 6480 952
rect 6400 792 6480 888
rect 6400 728 6408 792
rect 6472 728 6480 792
rect 6400 628 6480 728
rect 6400 572 6412 628
rect 6468 572 6480 628
rect 6400 560 6480 572
rect 6560 1268 6640 1280
rect 6560 1212 6572 1268
rect 6628 1212 6640 1268
rect 6560 1112 6640 1212
rect 6560 1048 6568 1112
rect 6632 1048 6640 1112
rect 6560 952 6640 1048
rect 6560 888 6568 952
rect 6632 888 6640 952
rect 6560 792 6640 888
rect 6560 728 6568 792
rect 6632 728 6640 792
rect 6560 628 6640 728
rect 6560 572 6572 628
rect 6628 572 6640 628
rect 6560 560 6640 572
rect 6720 1268 6800 1280
rect 6720 1212 6732 1268
rect 6788 1212 6800 1268
rect 6720 1112 6800 1212
rect 6720 1048 6728 1112
rect 6792 1048 6800 1112
rect 6720 952 6800 1048
rect 6720 888 6728 952
rect 6792 888 6800 952
rect 6720 792 6800 888
rect 6720 728 6728 792
rect 6792 728 6800 792
rect 6720 628 6800 728
rect 6720 572 6732 628
rect 6788 572 6800 628
rect 6720 560 6800 572
rect 6880 1268 6960 1280
rect 6880 1212 6892 1268
rect 6948 1212 6960 1268
rect 6880 1112 6960 1212
rect 6880 1048 6888 1112
rect 6952 1048 6960 1112
rect 6880 952 6960 1048
rect 6880 888 6888 952
rect 6952 888 6960 952
rect 6880 792 6960 888
rect 6880 728 6888 792
rect 6952 728 6960 792
rect 6880 628 6960 728
rect 6880 572 6892 628
rect 6948 572 6960 628
rect 6880 560 6960 572
rect 7200 1268 7280 1280
rect 7200 1212 7212 1268
rect 7268 1212 7280 1268
rect 7200 1112 7280 1212
rect 7200 1048 7208 1112
rect 7272 1048 7280 1112
rect 7200 952 7280 1048
rect 7200 888 7208 952
rect 7272 888 7280 952
rect 7200 792 7280 888
rect 7200 728 7208 792
rect 7272 728 7280 792
rect 7200 628 7280 728
rect 7200 572 7212 628
rect 7268 572 7280 628
rect 7200 560 7280 572
rect 7360 1268 7440 1280
rect 7360 1212 7372 1268
rect 7428 1212 7440 1268
rect 7360 1112 7440 1212
rect 7360 1048 7368 1112
rect 7432 1048 7440 1112
rect 7360 952 7440 1048
rect 7360 888 7368 952
rect 7432 888 7440 952
rect 7360 792 7440 888
rect 7360 728 7368 792
rect 7432 728 7440 792
rect 7360 628 7440 728
rect 7360 572 7372 628
rect 7428 572 7440 628
rect 7360 560 7440 572
rect 7520 1268 7600 1280
rect 7520 1212 7532 1268
rect 7588 1212 7600 1268
rect 7520 1112 7600 1212
rect 7520 1048 7528 1112
rect 7592 1048 7600 1112
rect 7520 952 7600 1048
rect 7520 888 7528 952
rect 7592 888 7600 952
rect 7520 792 7600 888
rect 7520 728 7528 792
rect 7592 728 7600 792
rect 7520 628 7600 728
rect 7520 572 7532 628
rect 7588 572 7600 628
rect 7520 560 7600 572
rect 7680 1268 7760 1280
rect 7680 1212 7692 1268
rect 7748 1212 7760 1268
rect 7680 1112 7760 1212
rect 7680 1048 7688 1112
rect 7752 1048 7760 1112
rect 7680 952 7760 1048
rect 7680 888 7688 952
rect 7752 888 7760 952
rect 7680 792 7760 888
rect 7680 728 7688 792
rect 7752 728 7760 792
rect 7680 628 7760 728
rect 7680 572 7692 628
rect 7748 572 7760 628
rect 7680 560 7760 572
rect 7840 1268 7920 1280
rect 7840 1212 7852 1268
rect 7908 1212 7920 1268
rect 7840 1112 7920 1212
rect 7840 1048 7848 1112
rect 7912 1048 7920 1112
rect 7840 952 7920 1048
rect 7840 888 7848 952
rect 7912 888 7920 952
rect 7840 792 7920 888
rect 7840 728 7848 792
rect 7912 728 7920 792
rect 7840 628 7920 728
rect 7840 572 7852 628
rect 7908 572 7920 628
rect 7840 560 7920 572
rect 8000 1268 8080 1280
rect 8000 1212 8012 1268
rect 8068 1212 8080 1268
rect 8000 1112 8080 1212
rect 8000 1048 8008 1112
rect 8072 1048 8080 1112
rect 8000 952 8080 1048
rect 8000 888 8008 952
rect 8072 888 8080 952
rect 8000 792 8080 888
rect 8000 728 8008 792
rect 8072 728 8080 792
rect 8000 628 8080 728
rect 8000 572 8012 628
rect 8068 572 8080 628
rect 8000 560 8080 572
rect 8160 1268 8240 1280
rect 8160 1212 8172 1268
rect 8228 1212 8240 1268
rect 8160 1112 8240 1212
rect 8160 1048 8168 1112
rect 8232 1048 8240 1112
rect 8160 952 8240 1048
rect 8160 888 8168 952
rect 8232 888 8240 952
rect 8160 792 8240 888
rect 8160 728 8168 792
rect 8232 728 8240 792
rect 8160 628 8240 728
rect 8160 572 8172 628
rect 8228 572 8240 628
rect 8160 560 8240 572
rect 320 332 400 360
rect 320 268 328 332
rect 392 268 400 332
rect 320 252 400 268
rect 320 188 328 252
rect 392 188 400 252
rect 320 160 400 188
rect 8000 332 8080 360
rect 8000 268 8008 332
rect 8072 268 8080 332
rect 8000 252 8080 268
rect 8000 188 8008 252
rect 8072 188 8080 252
rect 8000 160 8080 188
<< via3 >>
rect 4168 3628 4232 3632
rect 4168 3572 4172 3628
rect 4172 3572 4228 3628
rect 4228 3572 4232 3628
rect 4168 3568 4232 3572
rect 4168 3548 4232 3552
rect 4168 3492 4172 3548
rect 4172 3492 4228 3548
rect 4228 3492 4232 3548
rect 4168 3488 4232 3492
rect 4168 3468 4232 3472
rect 4168 3412 4172 3468
rect 4172 3412 4228 3468
rect 4228 3412 4232 3468
rect 4168 3408 4232 3412
rect 4168 3388 4232 3392
rect 4168 3332 4172 3388
rect 4172 3332 4228 3388
rect 4228 3332 4232 3388
rect 4168 3328 4232 3332
rect 8 2788 72 2792
rect 8 2732 12 2788
rect 12 2732 68 2788
rect 68 2732 72 2788
rect 8 2728 72 2732
rect 8 2468 72 2472
rect 8 2412 12 2468
rect 12 2412 68 2468
rect 68 2412 72 2468
rect 8 2408 72 2412
rect 168 2788 232 2792
rect 168 2732 172 2788
rect 172 2732 228 2788
rect 228 2732 232 2788
rect 168 2728 232 2732
rect 168 2468 232 2472
rect 168 2412 172 2468
rect 172 2412 228 2468
rect 228 2412 232 2468
rect 168 2408 232 2412
rect 328 2788 392 2792
rect 328 2732 332 2788
rect 332 2732 388 2788
rect 388 2732 392 2788
rect 328 2728 392 2732
rect 328 2468 392 2472
rect 328 2412 332 2468
rect 332 2412 388 2468
rect 388 2412 392 2468
rect 328 2408 392 2412
rect 488 2788 552 2792
rect 488 2732 492 2788
rect 492 2732 548 2788
rect 548 2732 552 2788
rect 488 2728 552 2732
rect 488 2468 552 2472
rect 488 2412 492 2468
rect 492 2412 548 2468
rect 548 2412 552 2468
rect 488 2408 552 2412
rect 648 2788 712 2792
rect 648 2732 652 2788
rect 652 2732 708 2788
rect 708 2732 712 2788
rect 648 2728 712 2732
rect 648 2468 712 2472
rect 648 2412 652 2468
rect 652 2412 708 2468
rect 708 2412 712 2468
rect 648 2408 712 2412
rect 808 2788 872 2792
rect 808 2732 812 2788
rect 812 2732 868 2788
rect 868 2732 872 2788
rect 808 2728 872 2732
rect 808 2468 872 2472
rect 808 2412 812 2468
rect 812 2412 868 2468
rect 868 2412 872 2468
rect 808 2408 872 2412
rect 968 2788 1032 2792
rect 968 2732 972 2788
rect 972 2732 1028 2788
rect 1028 2732 1032 2788
rect 968 2728 1032 2732
rect 968 2468 1032 2472
rect 968 2412 972 2468
rect 972 2412 1028 2468
rect 1028 2412 1032 2468
rect 968 2408 1032 2412
rect 1128 2788 1192 2792
rect 1128 2732 1132 2788
rect 1132 2732 1188 2788
rect 1188 2732 1192 2788
rect 1128 2728 1192 2732
rect 1128 2468 1192 2472
rect 1128 2412 1132 2468
rect 1132 2412 1188 2468
rect 1188 2412 1192 2468
rect 1128 2408 1192 2412
rect 1448 2788 1512 2792
rect 1448 2732 1452 2788
rect 1452 2732 1508 2788
rect 1508 2732 1512 2788
rect 1448 2728 1512 2732
rect 1448 2468 1512 2472
rect 1448 2412 1452 2468
rect 1452 2412 1508 2468
rect 1508 2412 1512 2468
rect 1448 2408 1512 2412
rect 1608 2788 1672 2792
rect 1608 2732 1612 2788
rect 1612 2732 1668 2788
rect 1668 2732 1672 2788
rect 1608 2728 1672 2732
rect 1608 2468 1672 2472
rect 1608 2412 1612 2468
rect 1612 2412 1668 2468
rect 1668 2412 1672 2468
rect 1608 2408 1672 2412
rect 1768 2788 1832 2792
rect 1768 2732 1772 2788
rect 1772 2732 1828 2788
rect 1828 2732 1832 2788
rect 1768 2728 1832 2732
rect 1768 2468 1832 2472
rect 1768 2412 1772 2468
rect 1772 2412 1828 2468
rect 1828 2412 1832 2468
rect 1768 2408 1832 2412
rect 1928 2788 1992 2792
rect 1928 2732 1932 2788
rect 1932 2732 1988 2788
rect 1988 2732 1992 2788
rect 1928 2728 1992 2732
rect 1928 2468 1992 2472
rect 1928 2412 1932 2468
rect 1932 2412 1988 2468
rect 1988 2412 1992 2468
rect 1928 2408 1992 2412
rect 2088 2788 2152 2792
rect 2088 2732 2092 2788
rect 2092 2732 2148 2788
rect 2148 2732 2152 2788
rect 2088 2728 2152 2732
rect 2088 2468 2152 2472
rect 2088 2412 2092 2468
rect 2092 2412 2148 2468
rect 2148 2412 2152 2468
rect 2088 2408 2152 2412
rect 2248 2788 2312 2792
rect 2248 2732 2252 2788
rect 2252 2732 2308 2788
rect 2308 2732 2312 2788
rect 2248 2728 2312 2732
rect 2248 2468 2312 2472
rect 2248 2412 2252 2468
rect 2252 2412 2308 2468
rect 2308 2412 2312 2468
rect 2248 2408 2312 2412
rect 2408 2788 2472 2792
rect 2408 2732 2412 2788
rect 2412 2732 2468 2788
rect 2468 2732 2472 2788
rect 2408 2728 2472 2732
rect 2408 2468 2472 2472
rect 2408 2412 2412 2468
rect 2412 2412 2468 2468
rect 2468 2412 2472 2468
rect 2408 2408 2472 2412
rect 2568 2788 2632 2792
rect 2568 2732 2572 2788
rect 2572 2732 2628 2788
rect 2628 2732 2632 2788
rect 2568 2728 2632 2732
rect 2568 2468 2632 2472
rect 2568 2412 2572 2468
rect 2572 2412 2628 2468
rect 2628 2412 2632 2468
rect 2568 2408 2632 2412
rect 2728 2788 2792 2792
rect 2728 2732 2732 2788
rect 2732 2732 2788 2788
rect 2788 2732 2792 2788
rect 2728 2728 2792 2732
rect 2728 2468 2792 2472
rect 2728 2412 2732 2468
rect 2732 2412 2788 2468
rect 2788 2412 2792 2468
rect 2728 2408 2792 2412
rect 2888 2788 2952 2792
rect 2888 2732 2892 2788
rect 2892 2732 2948 2788
rect 2948 2732 2952 2788
rect 2888 2728 2952 2732
rect 2888 2468 2952 2472
rect 2888 2412 2892 2468
rect 2892 2412 2948 2468
rect 2948 2412 2952 2468
rect 2888 2408 2952 2412
rect 3048 2788 3112 2792
rect 3048 2732 3052 2788
rect 3052 2732 3108 2788
rect 3108 2732 3112 2788
rect 3048 2728 3112 2732
rect 3048 2468 3112 2472
rect 3048 2412 3052 2468
rect 3052 2412 3108 2468
rect 3108 2412 3112 2468
rect 3048 2408 3112 2412
rect 3368 2788 3432 2792
rect 3368 2732 3372 2788
rect 3372 2732 3428 2788
rect 3428 2732 3432 2788
rect 3368 2728 3432 2732
rect 3368 2468 3432 2472
rect 3368 2412 3372 2468
rect 3372 2412 3428 2468
rect 3428 2412 3432 2468
rect 3368 2408 3432 2412
rect 3528 2788 3592 2792
rect 3528 2732 3532 2788
rect 3532 2732 3588 2788
rect 3588 2732 3592 2788
rect 3528 2728 3592 2732
rect 3528 2468 3592 2472
rect 3528 2412 3532 2468
rect 3532 2412 3588 2468
rect 3588 2412 3592 2468
rect 3528 2408 3592 2412
rect 3688 2788 3752 2792
rect 3688 2732 3692 2788
rect 3692 2732 3748 2788
rect 3748 2732 3752 2788
rect 3688 2728 3752 2732
rect 3688 2468 3752 2472
rect 3688 2412 3692 2468
rect 3692 2412 3748 2468
rect 3748 2412 3752 2468
rect 3688 2408 3752 2412
rect 3848 2788 3912 2792
rect 3848 2732 3852 2788
rect 3852 2732 3908 2788
rect 3908 2732 3912 2788
rect 3848 2728 3912 2732
rect 3848 2468 3912 2472
rect 3848 2412 3852 2468
rect 3852 2412 3908 2468
rect 3908 2412 3912 2468
rect 3848 2408 3912 2412
rect 4008 2788 4072 2792
rect 4008 2732 4012 2788
rect 4012 2732 4068 2788
rect 4068 2732 4072 2788
rect 4008 2728 4072 2732
rect 4008 2468 4072 2472
rect 4008 2412 4012 2468
rect 4012 2412 4068 2468
rect 4068 2412 4072 2468
rect 4008 2408 4072 2412
rect 4168 2788 4232 2792
rect 4168 2732 4172 2788
rect 4172 2732 4228 2788
rect 4228 2732 4232 2788
rect 4168 2728 4232 2732
rect 4168 2468 4232 2472
rect 4168 2412 4172 2468
rect 4172 2412 4228 2468
rect 4228 2412 4232 2468
rect 4168 2408 4232 2412
rect 4328 2788 4392 2792
rect 4328 2732 4332 2788
rect 4332 2732 4388 2788
rect 4388 2732 4392 2788
rect 4328 2728 4392 2732
rect 4328 2468 4392 2472
rect 4328 2412 4332 2468
rect 4332 2412 4388 2468
rect 4388 2412 4392 2468
rect 4328 2408 4392 2412
rect 4488 2788 4552 2792
rect 4488 2732 4492 2788
rect 4492 2732 4548 2788
rect 4548 2732 4552 2788
rect 4488 2728 4552 2732
rect 4488 2468 4552 2472
rect 4488 2412 4492 2468
rect 4492 2412 4548 2468
rect 4548 2412 4552 2468
rect 4488 2408 4552 2412
rect 4648 2788 4712 2792
rect 4648 2732 4652 2788
rect 4652 2732 4708 2788
rect 4708 2732 4712 2788
rect 4648 2728 4712 2732
rect 4648 2468 4712 2472
rect 4648 2412 4652 2468
rect 4652 2412 4708 2468
rect 4708 2412 4712 2468
rect 4648 2408 4712 2412
rect 4808 2788 4872 2792
rect 4808 2732 4812 2788
rect 4812 2732 4868 2788
rect 4868 2732 4872 2788
rect 4808 2728 4872 2732
rect 4808 2468 4872 2472
rect 4808 2412 4812 2468
rect 4812 2412 4868 2468
rect 4868 2412 4872 2468
rect 4808 2408 4872 2412
rect 4968 2788 5032 2792
rect 4968 2732 4972 2788
rect 4972 2732 5028 2788
rect 5028 2732 5032 2788
rect 4968 2728 5032 2732
rect 4968 2468 5032 2472
rect 4968 2412 4972 2468
rect 4972 2412 5028 2468
rect 5028 2412 5032 2468
rect 4968 2408 5032 2412
rect 5288 2788 5352 2792
rect 5288 2732 5292 2788
rect 5292 2732 5348 2788
rect 5348 2732 5352 2788
rect 5288 2728 5352 2732
rect 5288 2468 5352 2472
rect 5288 2412 5292 2468
rect 5292 2412 5348 2468
rect 5348 2412 5352 2468
rect 5288 2408 5352 2412
rect 5448 2788 5512 2792
rect 5448 2732 5452 2788
rect 5452 2732 5508 2788
rect 5508 2732 5512 2788
rect 5448 2728 5512 2732
rect 5448 2468 5512 2472
rect 5448 2412 5452 2468
rect 5452 2412 5508 2468
rect 5508 2412 5512 2468
rect 5448 2408 5512 2412
rect 5608 2788 5672 2792
rect 5608 2732 5612 2788
rect 5612 2732 5668 2788
rect 5668 2732 5672 2788
rect 5608 2728 5672 2732
rect 5608 2468 5672 2472
rect 5608 2412 5612 2468
rect 5612 2412 5668 2468
rect 5668 2412 5672 2468
rect 5608 2408 5672 2412
rect 5768 2788 5832 2792
rect 5768 2732 5772 2788
rect 5772 2732 5828 2788
rect 5828 2732 5832 2788
rect 5768 2728 5832 2732
rect 5768 2468 5832 2472
rect 5768 2412 5772 2468
rect 5772 2412 5828 2468
rect 5828 2412 5832 2468
rect 5768 2408 5832 2412
rect 5928 2788 5992 2792
rect 5928 2732 5932 2788
rect 5932 2732 5988 2788
rect 5988 2732 5992 2788
rect 5928 2728 5992 2732
rect 5928 2468 5992 2472
rect 5928 2412 5932 2468
rect 5932 2412 5988 2468
rect 5988 2412 5992 2468
rect 5928 2408 5992 2412
rect 6088 2788 6152 2792
rect 6088 2732 6092 2788
rect 6092 2732 6148 2788
rect 6148 2732 6152 2788
rect 6088 2728 6152 2732
rect 6088 2468 6152 2472
rect 6088 2412 6092 2468
rect 6092 2412 6148 2468
rect 6148 2412 6152 2468
rect 6088 2408 6152 2412
rect 6248 2788 6312 2792
rect 6248 2732 6252 2788
rect 6252 2732 6308 2788
rect 6308 2732 6312 2788
rect 6248 2728 6312 2732
rect 6248 2468 6312 2472
rect 6248 2412 6252 2468
rect 6252 2412 6308 2468
rect 6308 2412 6312 2468
rect 6248 2408 6312 2412
rect 6408 2788 6472 2792
rect 6408 2732 6412 2788
rect 6412 2732 6468 2788
rect 6468 2732 6472 2788
rect 6408 2728 6472 2732
rect 6408 2468 6472 2472
rect 6408 2412 6412 2468
rect 6412 2412 6468 2468
rect 6468 2412 6472 2468
rect 6408 2408 6472 2412
rect 6568 2788 6632 2792
rect 6568 2732 6572 2788
rect 6572 2732 6628 2788
rect 6628 2732 6632 2788
rect 6568 2728 6632 2732
rect 6568 2468 6632 2472
rect 6568 2412 6572 2468
rect 6572 2412 6628 2468
rect 6628 2412 6632 2468
rect 6568 2408 6632 2412
rect 6728 2788 6792 2792
rect 6728 2732 6732 2788
rect 6732 2732 6788 2788
rect 6788 2732 6792 2788
rect 6728 2728 6792 2732
rect 6728 2468 6792 2472
rect 6728 2412 6732 2468
rect 6732 2412 6788 2468
rect 6788 2412 6792 2468
rect 6728 2408 6792 2412
rect 6888 2788 6952 2792
rect 6888 2732 6892 2788
rect 6892 2732 6948 2788
rect 6948 2732 6952 2788
rect 6888 2728 6952 2732
rect 6888 2468 6952 2472
rect 6888 2412 6892 2468
rect 6892 2412 6948 2468
rect 6948 2412 6952 2468
rect 6888 2408 6952 2412
rect 7208 2788 7272 2792
rect 7208 2732 7212 2788
rect 7212 2732 7268 2788
rect 7268 2732 7272 2788
rect 7208 2728 7272 2732
rect 7208 2468 7272 2472
rect 7208 2412 7212 2468
rect 7212 2412 7268 2468
rect 7268 2412 7272 2468
rect 7208 2408 7272 2412
rect 7368 2788 7432 2792
rect 7368 2732 7372 2788
rect 7372 2732 7428 2788
rect 7428 2732 7432 2788
rect 7368 2728 7432 2732
rect 7368 2468 7432 2472
rect 7368 2412 7372 2468
rect 7372 2412 7428 2468
rect 7428 2412 7432 2468
rect 7368 2408 7432 2412
rect 7528 2788 7592 2792
rect 7528 2732 7532 2788
rect 7532 2732 7588 2788
rect 7588 2732 7592 2788
rect 7528 2728 7592 2732
rect 7528 2468 7592 2472
rect 7528 2412 7532 2468
rect 7532 2412 7588 2468
rect 7588 2412 7592 2468
rect 7528 2408 7592 2412
rect 7688 2788 7752 2792
rect 7688 2732 7692 2788
rect 7692 2732 7748 2788
rect 7748 2732 7752 2788
rect 7688 2728 7752 2732
rect 7688 2468 7752 2472
rect 7688 2412 7692 2468
rect 7692 2412 7748 2468
rect 7748 2412 7752 2468
rect 7688 2408 7752 2412
rect 7848 2788 7912 2792
rect 7848 2732 7852 2788
rect 7852 2732 7908 2788
rect 7908 2732 7912 2788
rect 7848 2728 7912 2732
rect 7848 2468 7912 2472
rect 7848 2412 7852 2468
rect 7852 2412 7908 2468
rect 7908 2412 7912 2468
rect 7848 2408 7912 2412
rect 8008 2788 8072 2792
rect 8008 2732 8012 2788
rect 8012 2732 8068 2788
rect 8068 2732 8072 2788
rect 8008 2728 8072 2732
rect 8008 2468 8072 2472
rect 8008 2412 8012 2468
rect 8012 2412 8068 2468
rect 8068 2412 8072 2468
rect 8008 2408 8072 2412
rect 8168 2788 8232 2792
rect 8168 2732 8172 2788
rect 8172 2732 8228 2788
rect 8228 2732 8232 2788
rect 8168 2728 8232 2732
rect 8168 2468 8232 2472
rect 8168 2412 8172 2468
rect 8172 2412 8228 2468
rect 8228 2412 8232 2468
rect 8168 2408 8232 2412
rect 8328 2788 8392 2792
rect 8328 2732 8332 2788
rect 8332 2732 8388 2788
rect 8388 2732 8392 2788
rect 8328 2728 8392 2732
rect 8328 2468 8392 2472
rect 8328 2412 8332 2468
rect 8332 2412 8388 2468
rect 8388 2412 8392 2468
rect 8328 2408 8392 2412
rect 168 1048 232 1112
rect 168 948 232 952
rect 168 892 172 948
rect 172 892 228 948
rect 228 892 232 948
rect 168 888 232 892
rect 168 728 232 792
rect 328 1048 392 1112
rect 328 948 392 952
rect 328 892 332 948
rect 332 892 388 948
rect 388 892 392 948
rect 328 888 392 892
rect 328 728 392 792
rect 488 1048 552 1112
rect 488 948 552 952
rect 488 892 492 948
rect 492 892 548 948
rect 548 892 552 948
rect 488 888 552 892
rect 488 728 552 792
rect 648 1048 712 1112
rect 648 948 712 952
rect 648 892 652 948
rect 652 892 708 948
rect 708 892 712 948
rect 648 888 712 892
rect 648 728 712 792
rect 808 1048 872 1112
rect 808 948 872 952
rect 808 892 812 948
rect 812 892 868 948
rect 868 892 872 948
rect 808 888 872 892
rect 808 728 872 792
rect 968 1048 1032 1112
rect 968 948 1032 952
rect 968 892 972 948
rect 972 892 1028 948
rect 1028 892 1032 948
rect 968 888 1032 892
rect 968 728 1032 792
rect 1128 1048 1192 1112
rect 1128 948 1192 952
rect 1128 892 1132 948
rect 1132 892 1188 948
rect 1188 892 1192 948
rect 1128 888 1192 892
rect 1128 728 1192 792
rect 1448 1048 1512 1112
rect 1448 948 1512 952
rect 1448 892 1452 948
rect 1452 892 1508 948
rect 1508 892 1512 948
rect 1448 888 1512 892
rect 1448 728 1512 792
rect 1608 1048 1672 1112
rect 1608 948 1672 952
rect 1608 892 1612 948
rect 1612 892 1668 948
rect 1668 892 1672 948
rect 1608 888 1672 892
rect 1608 728 1672 792
rect 1768 1048 1832 1112
rect 1768 948 1832 952
rect 1768 892 1772 948
rect 1772 892 1828 948
rect 1828 892 1832 948
rect 1768 888 1832 892
rect 1768 728 1832 792
rect 1928 1048 1992 1112
rect 1928 948 1992 952
rect 1928 892 1932 948
rect 1932 892 1988 948
rect 1988 892 1992 948
rect 1928 888 1992 892
rect 1928 728 1992 792
rect 2088 1048 2152 1112
rect 2088 948 2152 952
rect 2088 892 2092 948
rect 2092 892 2148 948
rect 2148 892 2152 948
rect 2088 888 2152 892
rect 2088 728 2152 792
rect 2248 1048 2312 1112
rect 2248 948 2312 952
rect 2248 892 2252 948
rect 2252 892 2308 948
rect 2308 892 2312 948
rect 2248 888 2312 892
rect 2248 728 2312 792
rect 2408 1048 2472 1112
rect 2408 948 2472 952
rect 2408 892 2412 948
rect 2412 892 2468 948
rect 2468 892 2472 948
rect 2408 888 2472 892
rect 2408 728 2472 792
rect 2568 1048 2632 1112
rect 2568 948 2632 952
rect 2568 892 2572 948
rect 2572 892 2628 948
rect 2628 892 2632 948
rect 2568 888 2632 892
rect 2568 728 2632 792
rect 2728 1048 2792 1112
rect 2728 948 2792 952
rect 2728 892 2732 948
rect 2732 892 2788 948
rect 2788 892 2792 948
rect 2728 888 2792 892
rect 2728 728 2792 792
rect 2888 1048 2952 1112
rect 2888 948 2952 952
rect 2888 892 2892 948
rect 2892 892 2948 948
rect 2948 892 2952 948
rect 2888 888 2952 892
rect 2888 728 2952 792
rect 3048 1048 3112 1112
rect 3048 948 3112 952
rect 3048 892 3052 948
rect 3052 892 3108 948
rect 3108 892 3112 948
rect 3048 888 3112 892
rect 3048 728 3112 792
rect 3368 1048 3432 1112
rect 3368 948 3432 952
rect 3368 892 3372 948
rect 3372 892 3428 948
rect 3428 892 3432 948
rect 3368 888 3432 892
rect 3368 728 3432 792
rect 3528 1048 3592 1112
rect 3528 948 3592 952
rect 3528 892 3532 948
rect 3532 892 3588 948
rect 3588 892 3592 948
rect 3528 888 3592 892
rect 3528 728 3592 792
rect 3688 1048 3752 1112
rect 3688 948 3752 952
rect 3688 892 3692 948
rect 3692 892 3748 948
rect 3748 892 3752 948
rect 3688 888 3752 892
rect 3688 728 3752 792
rect 3848 1048 3912 1112
rect 3848 948 3912 952
rect 3848 892 3852 948
rect 3852 892 3908 948
rect 3908 892 3912 948
rect 3848 888 3912 892
rect 3848 728 3912 792
rect 4008 1048 4072 1112
rect 4008 948 4072 952
rect 4008 892 4012 948
rect 4012 892 4068 948
rect 4068 892 4072 948
rect 4008 888 4072 892
rect 4008 728 4072 792
rect 4328 1048 4392 1112
rect 4328 948 4392 952
rect 4328 892 4332 948
rect 4332 892 4388 948
rect 4388 892 4392 948
rect 4328 888 4392 892
rect 4328 728 4392 792
rect 4488 1048 4552 1112
rect 4488 948 4552 952
rect 4488 892 4492 948
rect 4492 892 4548 948
rect 4548 892 4552 948
rect 4488 888 4552 892
rect 4488 728 4552 792
rect 4648 1048 4712 1112
rect 4648 948 4712 952
rect 4648 892 4652 948
rect 4652 892 4708 948
rect 4708 892 4712 948
rect 4648 888 4712 892
rect 4648 728 4712 792
rect 4808 1048 4872 1112
rect 4808 948 4872 952
rect 4808 892 4812 948
rect 4812 892 4868 948
rect 4868 892 4872 948
rect 4808 888 4872 892
rect 4808 728 4872 792
rect 4968 1048 5032 1112
rect 4968 948 5032 952
rect 4968 892 4972 948
rect 4972 892 5028 948
rect 5028 892 5032 948
rect 4968 888 5032 892
rect 4968 728 5032 792
rect 5288 1048 5352 1112
rect 5288 948 5352 952
rect 5288 892 5292 948
rect 5292 892 5348 948
rect 5348 892 5352 948
rect 5288 888 5352 892
rect 5288 728 5352 792
rect 5448 1048 5512 1112
rect 5448 948 5512 952
rect 5448 892 5452 948
rect 5452 892 5508 948
rect 5508 892 5512 948
rect 5448 888 5512 892
rect 5448 728 5512 792
rect 5608 1048 5672 1112
rect 5608 948 5672 952
rect 5608 892 5612 948
rect 5612 892 5668 948
rect 5668 892 5672 948
rect 5608 888 5672 892
rect 5608 728 5672 792
rect 5768 1048 5832 1112
rect 5768 948 5832 952
rect 5768 892 5772 948
rect 5772 892 5828 948
rect 5828 892 5832 948
rect 5768 888 5832 892
rect 5768 728 5832 792
rect 5928 1048 5992 1112
rect 5928 948 5992 952
rect 5928 892 5932 948
rect 5932 892 5988 948
rect 5988 892 5992 948
rect 5928 888 5992 892
rect 5928 728 5992 792
rect 6088 1048 6152 1112
rect 6088 948 6152 952
rect 6088 892 6092 948
rect 6092 892 6148 948
rect 6148 892 6152 948
rect 6088 888 6152 892
rect 6088 728 6152 792
rect 6248 1048 6312 1112
rect 6248 948 6312 952
rect 6248 892 6252 948
rect 6252 892 6308 948
rect 6308 892 6312 948
rect 6248 888 6312 892
rect 6248 728 6312 792
rect 6408 1048 6472 1112
rect 6408 948 6472 952
rect 6408 892 6412 948
rect 6412 892 6468 948
rect 6468 892 6472 948
rect 6408 888 6472 892
rect 6408 728 6472 792
rect 6568 1048 6632 1112
rect 6568 948 6632 952
rect 6568 892 6572 948
rect 6572 892 6628 948
rect 6628 892 6632 948
rect 6568 888 6632 892
rect 6568 728 6632 792
rect 6728 1048 6792 1112
rect 6728 948 6792 952
rect 6728 892 6732 948
rect 6732 892 6788 948
rect 6788 892 6792 948
rect 6728 888 6792 892
rect 6728 728 6792 792
rect 6888 1048 6952 1112
rect 6888 948 6952 952
rect 6888 892 6892 948
rect 6892 892 6948 948
rect 6948 892 6952 948
rect 6888 888 6952 892
rect 6888 728 6952 792
rect 7208 1048 7272 1112
rect 7208 948 7272 952
rect 7208 892 7212 948
rect 7212 892 7268 948
rect 7268 892 7272 948
rect 7208 888 7272 892
rect 7208 728 7272 792
rect 7368 1048 7432 1112
rect 7368 948 7432 952
rect 7368 892 7372 948
rect 7372 892 7428 948
rect 7428 892 7432 948
rect 7368 888 7432 892
rect 7368 728 7432 792
rect 7528 1048 7592 1112
rect 7528 948 7592 952
rect 7528 892 7532 948
rect 7532 892 7588 948
rect 7588 892 7592 948
rect 7528 888 7592 892
rect 7528 728 7592 792
rect 7688 1048 7752 1112
rect 7688 948 7752 952
rect 7688 892 7692 948
rect 7692 892 7748 948
rect 7748 892 7752 948
rect 7688 888 7752 892
rect 7688 728 7752 792
rect 7848 1048 7912 1112
rect 7848 948 7912 952
rect 7848 892 7852 948
rect 7852 892 7908 948
rect 7908 892 7912 948
rect 7848 888 7912 892
rect 7848 728 7912 792
rect 8008 1048 8072 1112
rect 8008 948 8072 952
rect 8008 892 8012 948
rect 8012 892 8068 948
rect 8068 892 8072 948
rect 8008 888 8072 892
rect 8008 728 8072 792
rect 8168 1048 8232 1112
rect 8168 948 8232 952
rect 8168 892 8172 948
rect 8172 892 8228 948
rect 8228 892 8232 948
rect 8168 888 8232 892
rect 8168 728 8232 792
rect 328 328 392 332
rect 328 272 332 328
rect 332 272 388 328
rect 388 272 392 328
rect 328 268 392 272
rect 328 248 392 252
rect 328 192 332 248
rect 332 192 388 248
rect 388 192 392 248
rect 328 188 392 192
rect 8008 328 8072 332
rect 8008 272 8012 328
rect 8012 272 8068 328
rect 8068 272 8072 328
rect 8008 268 8072 272
rect 8008 248 8072 252
rect 8008 192 8012 248
rect 8012 192 8068 248
rect 8068 192 8072 248
rect 8008 188 8072 192
<< metal4 >>
rect 0 3632 8400 3680
rect 0 3598 4168 3632
rect 0 3362 242 3598
rect 478 3568 4168 3598
rect 4232 3598 8400 3632
rect 4232 3568 7922 3598
rect 478 3552 7922 3568
rect 478 3488 4168 3552
rect 4232 3488 7922 3552
rect 478 3472 7922 3488
rect 478 3408 4168 3472
rect 4232 3408 7922 3472
rect 478 3392 7922 3408
rect 478 3362 4168 3392
rect 0 3328 4168 3362
rect 4232 3362 7922 3392
rect 8158 3362 8400 3598
rect 4232 3328 8400 3362
rect 0 3280 8400 3328
rect 0 2792 8400 2800
rect 0 2728 8 2792
rect 72 2728 168 2792
rect 232 2728 328 2792
rect 392 2728 488 2792
rect 552 2728 648 2792
rect 712 2728 808 2792
rect 872 2728 968 2792
rect 1032 2728 1128 2792
rect 1192 2728 1448 2792
rect 1512 2728 1608 2792
rect 1672 2728 1768 2792
rect 1832 2728 1928 2792
rect 1992 2728 2088 2792
rect 2152 2728 2248 2792
rect 2312 2728 2408 2792
rect 2472 2728 2568 2792
rect 2632 2728 2728 2792
rect 2792 2728 2888 2792
rect 2952 2728 3048 2792
rect 3112 2728 3368 2792
rect 3432 2728 3528 2792
rect 3592 2728 3688 2792
rect 3752 2728 3848 2792
rect 3912 2728 4008 2792
rect 4072 2728 4168 2792
rect 4232 2728 4328 2792
rect 4392 2728 4488 2792
rect 4552 2728 4648 2792
rect 4712 2728 4808 2792
rect 4872 2728 4968 2792
rect 5032 2728 5288 2792
rect 5352 2728 5448 2792
rect 5512 2728 5608 2792
rect 5672 2728 5768 2792
rect 5832 2728 5928 2792
rect 5992 2728 6088 2792
rect 6152 2728 6248 2792
rect 6312 2728 6408 2792
rect 6472 2728 6568 2792
rect 6632 2728 6728 2792
rect 6792 2728 6888 2792
rect 6952 2728 7208 2792
rect 7272 2728 7368 2792
rect 7432 2728 7528 2792
rect 7592 2728 7688 2792
rect 7752 2728 7848 2792
rect 7912 2728 8008 2792
rect 8072 2728 8168 2792
rect 8232 2728 8328 2792
rect 8392 2728 8400 2792
rect 0 2718 8400 2728
rect 0 2482 1202 2718
rect 1438 2482 6962 2718
rect 7198 2482 8400 2718
rect 0 2472 8400 2482
rect 0 2408 8 2472
rect 72 2408 168 2472
rect 232 2408 328 2472
rect 392 2408 488 2472
rect 552 2408 648 2472
rect 712 2408 808 2472
rect 872 2408 968 2472
rect 1032 2408 1128 2472
rect 1192 2408 1448 2472
rect 1512 2408 1608 2472
rect 1672 2408 1768 2472
rect 1832 2408 1928 2472
rect 1992 2408 2088 2472
rect 2152 2408 2248 2472
rect 2312 2408 2408 2472
rect 2472 2408 2568 2472
rect 2632 2408 2728 2472
rect 2792 2408 2888 2472
rect 2952 2408 3048 2472
rect 3112 2408 3368 2472
rect 3432 2408 3528 2472
rect 3592 2408 3688 2472
rect 3752 2408 3848 2472
rect 3912 2408 4008 2472
rect 4072 2408 4168 2472
rect 4232 2408 4328 2472
rect 4392 2408 4488 2472
rect 4552 2408 4648 2472
rect 4712 2408 4808 2472
rect 4872 2408 4968 2472
rect 5032 2408 5288 2472
rect 5352 2408 5448 2472
rect 5512 2408 5608 2472
rect 5672 2408 5768 2472
rect 5832 2408 5928 2472
rect 5992 2408 6088 2472
rect 6152 2408 6248 2472
rect 6312 2408 6408 2472
rect 6472 2408 6568 2472
rect 6632 2408 6728 2472
rect 6792 2408 6888 2472
rect 6952 2408 7208 2472
rect 7272 2408 7368 2472
rect 7432 2408 7528 2472
rect 7592 2408 7688 2472
rect 7752 2408 7848 2472
rect 7912 2408 8008 2472
rect 8072 2408 8168 2472
rect 8232 2408 8328 2472
rect 8392 2408 8400 2472
rect 0 2400 8400 2408
rect 0 1112 8400 1120
rect 0 1048 168 1112
rect 232 1048 328 1112
rect 392 1048 488 1112
rect 552 1048 648 1112
rect 712 1048 808 1112
rect 872 1048 968 1112
rect 1032 1048 1128 1112
rect 1192 1048 1448 1112
rect 1512 1048 1608 1112
rect 1672 1048 1768 1112
rect 1832 1048 1928 1112
rect 1992 1048 2088 1112
rect 2152 1048 2248 1112
rect 2312 1048 2408 1112
rect 2472 1048 2568 1112
rect 2632 1048 2728 1112
rect 2792 1048 2888 1112
rect 2952 1048 3048 1112
rect 3112 1048 3368 1112
rect 3432 1048 3528 1112
rect 3592 1048 3688 1112
rect 3752 1048 3848 1112
rect 3912 1048 4008 1112
rect 4072 1048 4328 1112
rect 4392 1048 4488 1112
rect 4552 1048 4648 1112
rect 4712 1048 4808 1112
rect 4872 1048 4968 1112
rect 5032 1048 5288 1112
rect 5352 1048 5448 1112
rect 5512 1048 5608 1112
rect 5672 1048 5768 1112
rect 5832 1048 5928 1112
rect 5992 1048 6088 1112
rect 6152 1048 6248 1112
rect 6312 1048 6408 1112
rect 6472 1048 6568 1112
rect 6632 1048 6728 1112
rect 6792 1048 6888 1112
rect 6952 1048 7208 1112
rect 7272 1048 7368 1112
rect 7432 1048 7528 1112
rect 7592 1048 7688 1112
rect 7752 1048 7848 1112
rect 7912 1048 8008 1112
rect 8072 1048 8168 1112
rect 8232 1048 8400 1112
rect 0 1038 8400 1048
rect 0 952 2162 1038
rect 2398 952 4082 1038
rect 0 888 168 952
rect 232 888 328 952
rect 392 888 488 952
rect 552 888 648 952
rect 712 888 808 952
rect 872 888 968 952
rect 1032 888 1128 952
rect 1192 888 1448 952
rect 1512 888 1608 952
rect 1672 888 1768 952
rect 1832 888 1928 952
rect 1992 888 2088 952
rect 2152 888 2162 952
rect 2398 888 2408 952
rect 2472 888 2568 952
rect 2632 888 2728 952
rect 2792 888 2888 952
rect 2952 888 3048 952
rect 3112 888 3368 952
rect 3432 888 3528 952
rect 3592 888 3688 952
rect 3752 888 3848 952
rect 3912 888 4008 952
rect 4072 888 4082 952
rect 0 802 2162 888
rect 2398 802 4082 888
rect 4318 952 6002 1038
rect 6238 952 8400 1038
rect 4318 888 4328 952
rect 4392 888 4488 952
rect 4552 888 4648 952
rect 4712 888 4808 952
rect 4872 888 4968 952
rect 5032 888 5288 952
rect 5352 888 5448 952
rect 5512 888 5608 952
rect 5672 888 5768 952
rect 5832 888 5928 952
rect 5992 888 6002 952
rect 6238 888 6248 952
rect 6312 888 6408 952
rect 6472 888 6568 952
rect 6632 888 6728 952
rect 6792 888 6888 952
rect 6952 888 7208 952
rect 7272 888 7368 952
rect 7432 888 7528 952
rect 7592 888 7688 952
rect 7752 888 7848 952
rect 7912 888 8008 952
rect 8072 888 8168 952
rect 8232 888 8400 952
rect 4318 802 6002 888
rect 6238 802 8400 888
rect 0 792 8400 802
rect 0 728 168 792
rect 232 728 328 792
rect 392 728 488 792
rect 552 728 648 792
rect 712 728 808 792
rect 872 728 968 792
rect 1032 728 1128 792
rect 1192 728 1448 792
rect 1512 728 1608 792
rect 1672 728 1768 792
rect 1832 728 1928 792
rect 1992 728 2088 792
rect 2152 728 2248 792
rect 2312 728 2408 792
rect 2472 728 2568 792
rect 2632 728 2728 792
rect 2792 728 2888 792
rect 2952 728 3048 792
rect 3112 728 3368 792
rect 3432 728 3528 792
rect 3592 728 3688 792
rect 3752 728 3848 792
rect 3912 728 4008 792
rect 4072 728 4328 792
rect 4392 728 4488 792
rect 4552 728 4648 792
rect 4712 728 4808 792
rect 4872 728 4968 792
rect 5032 728 5288 792
rect 5352 728 5448 792
rect 5512 728 5608 792
rect 5672 728 5768 792
rect 5832 728 5928 792
rect 5992 728 6088 792
rect 6152 728 6248 792
rect 6312 728 6408 792
rect 6472 728 6568 792
rect 6632 728 6728 792
rect 6792 728 6888 792
rect 6952 728 7208 792
rect 7272 728 7368 792
rect 7432 728 7528 792
rect 7592 728 7688 792
rect 7752 728 7848 792
rect 7912 728 8008 792
rect 8072 728 8168 792
rect 8232 728 8400 792
rect 0 720 8400 728
rect 0 332 8400 400
rect 0 268 328 332
rect 392 318 8008 332
rect 392 268 3122 318
rect 0 252 3122 268
rect 0 188 328 252
rect 392 188 3122 252
rect 0 82 3122 188
rect 3358 82 5042 318
rect 5278 268 8008 318
rect 8072 268 8400 332
rect 5278 252 8400 268
rect 5278 188 8008 252
rect 8072 188 8400 252
rect 5278 82 8400 188
rect 0 0 8400 82
<< via4 >>
rect 242 3362 478 3598
rect 7922 3362 8158 3598
rect 1202 2482 1438 2718
rect 6962 2482 7198 2718
rect 2162 952 2398 1038
rect 2162 888 2248 952
rect 2248 888 2312 952
rect 2312 888 2398 952
rect 2162 802 2398 888
rect 4082 802 4318 1038
rect 6002 952 6238 1038
rect 6002 888 6088 952
rect 6088 888 6152 952
rect 6152 888 6238 952
rect 6002 802 6238 888
rect 3122 82 3358 318
rect 5042 82 5278 318
<< metal5 >>
rect 160 3598 560 4000
rect 160 3362 242 3598
rect 478 3362 560 3598
rect 160 0 560 3362
rect 1120 2718 1520 4000
rect 1120 2482 1202 2718
rect 1438 2482 1520 2718
rect 1120 0 1520 2482
rect 2080 1038 2480 4000
rect 2080 802 2162 1038
rect 2398 802 2480 1038
rect 2080 0 2480 802
rect 3040 318 3440 4000
rect 3040 82 3122 318
rect 3358 82 3440 318
rect 3040 0 3440 82
rect 4000 1038 4400 4000
rect 4000 802 4082 1038
rect 4318 802 4400 1038
rect 4000 0 4400 802
rect 4960 318 5360 4000
rect 4960 82 5042 318
rect 5278 82 5360 318
rect 4960 0 5360 82
rect 5920 1038 6320 4000
rect 5920 802 6002 1038
rect 6238 802 6320 1038
rect 5920 0 6320 802
rect 6880 2718 7280 4000
rect 6880 2482 6962 2718
rect 7198 2482 7280 2718
rect 6880 0 7280 2482
rect 7840 3598 8240 4000
rect 7840 3362 7922 3598
rect 8158 3362 8240 3598
rect 7840 0 8240 3362
<< labels >>
rlabel metal1 s 2240 3080 2320 3680 4 pa1
rlabel metal1 s 2240 1640 2320 2240 4 pb1
rlabel metal1 s 6080 1640 6160 2240 4 pb2
rlabel metal1 s 2240 160 2320 360 4 n1
rlabel metal1 s 6080 160 6160 360 4 n2
rlabel metal1 s 6080 3080 6160 3680 4 pa2
rlabel metal2 s 0 1040 8400 1120 4 in
port 1 nsew
rlabel metal2 s 0 720 8400 800 4 out
port 2 nsew
rlabel metal5 s 160 0 560 4000 4 vdda
port 3 nsew
rlabel metal2 s 0 2560 8400 2640 4 bp
port 4 nsew
rlabel metal5 s 1120 0 1520 4000 4 vddx
port 5 nsew
rlabel metal5 s 2080 0 2480 4000 4 gnda
port 6 nsew
rlabel metal5 s 3040 0 3440 4000 4 vssa
port 7 nsew
<< end >>
