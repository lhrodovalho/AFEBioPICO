magic
tech sky130A
timestamp 1637516460
<< nwell >>
rect -180 1620 2220 2100
rect 4060 1620 6460 2100
rect -180 980 2220 1460
rect 4060 980 6460 1460
rect -180 340 2220 820
rect 4060 340 6460 820
rect -180 -300 2220 180
rect 4060 -300 6460 180
<< mvpmos >>
rect 20 1958 2020 2000
rect 20 1798 2020 1840
rect 4260 1958 6260 2000
rect 4260 1798 6260 1840
rect 20 1240 2020 1282
rect 20 1080 2020 1122
rect 4260 1240 6260 1282
rect 4260 1080 6260 1122
rect 20 678 2020 720
rect 20 518 2020 560
rect 4260 678 6260 720
rect 4260 518 6260 560
rect 20 -40 2020 2
rect 20 -200 2020 -158
rect 4260 -40 6260 2
rect 4260 -200 6260 -158
<< mvpdiff >>
rect -80 1990 20 2000
rect -80 1970 -70 1990
rect -50 1970 20 1990
rect -80 1958 20 1970
rect 2020 1990 2120 2000
rect 2020 1970 2090 1990
rect 2110 1970 2120 1990
rect 2020 1958 2120 1970
rect -80 1830 20 1840
rect -80 1810 -70 1830
rect -50 1810 20 1830
rect -80 1798 20 1810
rect 2020 1830 2120 1840
rect 2020 1810 2090 1830
rect 2110 1810 2120 1830
rect 2020 1798 2120 1810
rect 4160 1990 4260 2000
rect 4160 1970 4170 1990
rect 4190 1970 4260 1990
rect 4160 1958 4260 1970
rect 6260 1990 6360 2000
rect 6260 1970 6330 1990
rect 6350 1970 6360 1990
rect 6260 1958 6360 1970
rect 4160 1830 4260 1840
rect 4160 1810 4170 1830
rect 4190 1810 4260 1830
rect 4160 1798 4260 1810
rect 6260 1830 6360 1840
rect 6260 1810 6330 1830
rect 6350 1810 6360 1830
rect 6260 1798 6360 1810
rect -80 1270 20 1282
rect -80 1250 -70 1270
rect -50 1250 20 1270
rect -80 1240 20 1250
rect 2020 1270 2120 1282
rect 2020 1250 2090 1270
rect 2110 1250 2120 1270
rect 2020 1240 2120 1250
rect -80 1110 20 1122
rect -80 1090 -70 1110
rect -50 1090 20 1110
rect -80 1080 20 1090
rect 2020 1110 2120 1122
rect 2020 1090 2090 1110
rect 2110 1090 2120 1110
rect 2020 1080 2120 1090
rect 4160 1270 4260 1282
rect 4160 1250 4170 1270
rect 4190 1250 4260 1270
rect 4160 1240 4260 1250
rect 6260 1270 6360 1282
rect 6260 1250 6330 1270
rect 6350 1250 6360 1270
rect 6260 1240 6360 1250
rect 4160 1110 4260 1122
rect 4160 1090 4170 1110
rect 4190 1090 4260 1110
rect 4160 1080 4260 1090
rect 6260 1110 6360 1122
rect 6260 1090 6330 1110
rect 6350 1090 6360 1110
rect 6260 1080 6360 1090
rect -80 710 20 720
rect -80 690 -70 710
rect -50 690 20 710
rect -80 678 20 690
rect 2020 710 2120 720
rect 2020 690 2090 710
rect 2110 690 2120 710
rect 2020 678 2120 690
rect -80 550 20 560
rect -80 530 -70 550
rect -50 530 20 550
rect -80 518 20 530
rect 2020 550 2120 560
rect 2020 530 2090 550
rect 2110 530 2120 550
rect 2020 518 2120 530
rect 4160 710 4260 720
rect 4160 690 4170 710
rect 4190 690 4260 710
rect 4160 678 4260 690
rect 6260 710 6360 720
rect 6260 690 6330 710
rect 6350 690 6360 710
rect 6260 678 6360 690
rect 4160 550 4260 560
rect 4160 530 4170 550
rect 4190 530 4260 550
rect 4160 518 4260 530
rect 6260 550 6360 560
rect 6260 530 6330 550
rect 6350 530 6360 550
rect 6260 518 6360 530
rect -80 -10 20 2
rect -80 -30 -70 -10
rect -50 -30 20 -10
rect -80 -40 20 -30
rect 2020 -10 2120 2
rect 2020 -30 2090 -10
rect 2110 -30 2120 -10
rect 2020 -40 2120 -30
rect -80 -170 20 -158
rect -80 -190 -70 -170
rect -50 -190 20 -170
rect -80 -200 20 -190
rect 2020 -170 2120 -158
rect 2020 -190 2090 -170
rect 2110 -190 2120 -170
rect 2020 -200 2120 -190
rect 4160 -10 4260 2
rect 4160 -30 4170 -10
rect 4190 -30 4260 -10
rect 4160 -40 4260 -30
rect 6260 -10 6360 2
rect 6260 -30 6330 -10
rect 6350 -30 6360 -10
rect 6260 -40 6360 -30
rect 4160 -170 4260 -158
rect 4160 -190 4170 -170
rect 4190 -190 4260 -170
rect 4160 -200 4260 -190
rect 6260 -170 6360 -158
rect 6260 -190 6330 -170
rect 6350 -190 6360 -170
rect 6260 -200 6360 -190
<< mvpdiffc >>
rect -70 1970 -50 1990
rect 2090 1970 2110 1990
rect -70 1810 -50 1830
rect 2090 1810 2110 1830
rect 4170 1970 4190 1990
rect 6330 1970 6350 1990
rect 4170 1810 4190 1830
rect 6330 1810 6350 1830
rect -70 1250 -50 1270
rect 2090 1250 2110 1270
rect -70 1090 -50 1110
rect 2090 1090 2110 1110
rect 4170 1250 4190 1270
rect 6330 1250 6350 1270
rect 4170 1090 4190 1110
rect 6330 1090 6350 1110
rect -70 690 -50 710
rect 2090 690 2110 710
rect -70 530 -50 550
rect 2090 530 2110 550
rect 4170 690 4190 710
rect 6330 690 6350 710
rect 4170 530 4190 550
rect 6330 530 6350 550
rect -70 -30 -50 -10
rect 2090 -30 2110 -10
rect -70 -190 -50 -170
rect 2090 -190 2110 -170
rect 4170 -30 4190 -10
rect 6330 -30 6350 -10
rect 4170 -190 4190 -170
rect 6330 -190 6350 -170
<< psubdiff >>
rect -240 2120 -180 2160
rect 2220 2120 2280 2160
rect -240 2100 -200 2120
rect 2240 2100 2280 2120
rect -240 1600 -200 1640
rect 2240 1600 2280 1640
rect -240 1560 -180 1600
rect 2220 1560 2280 1600
rect 4000 2120 4060 2160
rect 6460 2120 6520 2160
rect 4000 2100 4040 2120
rect 6480 2100 6520 2120
rect 4000 1600 4040 1640
rect 6480 1600 6520 1640
rect 4000 1560 4060 1600
rect 6460 1560 6520 1600
rect -240 1480 -180 1520
rect 2220 1480 2280 1520
rect -240 1440 -200 1480
rect 2240 1440 2280 1480
rect -240 960 -200 980
rect 2240 960 2280 980
rect -240 920 -180 960
rect 2220 920 2280 960
rect 4000 1480 4060 1520
rect 6460 1480 6520 1520
rect 4000 1440 4040 1480
rect 6480 1440 6520 1480
rect 4000 960 4040 980
rect 6480 960 6520 980
rect 4000 920 4060 960
rect 6460 920 6520 960
rect -240 840 -180 880
rect 2220 840 2280 880
rect -240 820 -200 840
rect 2240 820 2280 840
rect -240 320 -200 360
rect 2240 320 2280 360
rect -240 280 -180 320
rect 2220 280 2280 320
rect 4000 840 4060 880
rect 6460 840 6520 880
rect 4000 820 4040 840
rect 6480 820 6520 840
rect 4000 320 4040 360
rect 6480 320 6520 360
rect 4000 280 4060 320
rect 6460 280 6520 320
rect -240 200 -180 240
rect 2220 200 2280 240
rect -240 160 -200 200
rect 2240 160 2280 200
rect -240 -320 -200 -300
rect 2240 -320 2280 -300
rect -240 -360 -180 -320
rect 2220 -360 2280 -320
rect 4000 200 4060 240
rect 6460 200 6520 240
rect 4000 160 4040 200
rect 6480 160 6520 200
rect 4000 -320 4040 -300
rect 6480 -320 6520 -300
rect 4000 -360 4060 -320
rect 6460 -360 6520 -320
<< nsubdiff >>
rect -160 2040 -100 2080
rect 2140 2040 2200 2080
rect -160 2020 -120 2040
rect 2160 2020 2200 2040
rect -160 1640 -100 1680
rect 2140 1640 2200 1680
rect 4080 2040 4140 2080
rect 6380 2040 6440 2080
rect 4080 2020 4120 2040
rect 6400 2020 6440 2040
rect 4080 1640 4140 1680
rect 6380 1640 6440 1680
rect -160 1400 -100 1440
rect 2140 1400 2200 1440
rect -160 1040 -120 1060
rect 2160 1040 2200 1060
rect -160 1000 -100 1040
rect 2140 1000 2200 1040
rect 4080 1400 4140 1440
rect 6380 1400 6440 1440
rect 4080 1040 4120 1060
rect 6400 1040 6440 1060
rect 4080 1000 4140 1040
rect 6380 1000 6440 1040
rect -160 760 -100 800
rect 2140 760 2200 800
rect -160 740 -120 760
rect 2160 740 2200 760
rect -160 360 -100 400
rect 2140 360 2200 400
rect 4080 760 4140 800
rect 6380 760 6440 800
rect 4080 740 4120 760
rect 6400 740 6440 760
rect 4080 360 4140 400
rect 6380 360 6440 400
rect -160 120 -100 160
rect 2140 120 2200 160
rect -160 -240 -120 -220
rect 2160 -240 2200 -220
rect -160 -280 -100 -240
rect 2140 -280 2200 -240
rect 4080 120 4140 160
rect 6380 120 6440 160
rect 4080 -240 4120 -220
rect 6400 -240 6440 -220
rect 4080 -280 4140 -240
rect 6380 -280 6440 -240
<< psubdiffcont >>
rect -180 2120 2220 2160
rect -240 1640 -200 2100
rect 2240 1640 2280 2100
rect -180 1560 2220 1600
rect 4060 2120 6460 2160
rect 4000 1640 4040 2100
rect 6480 1640 6520 2100
rect 4060 1560 6460 1600
rect -180 1480 2220 1520
rect -240 980 -200 1440
rect 2240 980 2280 1440
rect -180 920 2220 960
rect 4060 1480 6460 1520
rect 4000 980 4040 1440
rect 6480 980 6520 1440
rect 4060 920 6460 960
rect -180 840 2220 880
rect -240 360 -200 820
rect 2240 360 2280 820
rect -180 280 2220 320
rect 4060 840 6460 880
rect 4000 360 4040 820
rect 6480 360 6520 820
rect 4060 280 6460 320
rect -180 200 2220 240
rect -240 -300 -200 160
rect 2240 -300 2280 160
rect -180 -360 2220 -320
rect 4060 200 6460 240
rect 4000 -300 4040 160
rect 6480 -300 6520 160
rect 4060 -360 6460 -320
<< nsubdiffcont >>
rect -100 2040 2140 2080
rect -160 1680 -120 2020
rect 2160 1680 2200 2020
rect -100 1640 2140 1680
rect 4140 2040 6380 2080
rect 4080 1680 4120 2020
rect 6400 1680 6440 2020
rect 4140 1640 6380 1680
rect -100 1400 2140 1440
rect -160 1060 -120 1400
rect 2160 1060 2200 1400
rect -100 1000 2140 1040
rect 4140 1400 6380 1440
rect 4080 1060 4120 1400
rect 6400 1060 6440 1400
rect 4140 1000 6380 1040
rect -100 760 2140 800
rect -160 400 -120 740
rect 2160 400 2200 740
rect -100 360 2140 400
rect 4140 760 6380 800
rect 4080 400 4120 740
rect 6400 400 6440 740
rect 4140 360 6380 400
rect -100 120 2140 160
rect -160 -220 -120 120
rect 2160 -220 2200 120
rect -100 -280 2140 -240
rect 4140 120 6380 160
rect 4080 -220 4120 120
rect 6400 -220 6440 120
rect 4140 -280 6380 -240
<< poly >>
rect 20 2000 2020 2020
rect 20 1915 2020 1958
rect 20 1885 30 1915
rect 2010 1885 2020 1915
rect 20 1880 2020 1885
rect 20 1840 2020 1855
rect 20 1755 2020 1798
rect 20 1725 30 1755
rect 2010 1725 2020 1755
rect 20 1720 2020 1725
rect 4260 2000 6260 2020
rect 4260 1915 6260 1958
rect 4260 1885 4270 1915
rect 6250 1885 6260 1915
rect 4260 1880 6260 1885
rect 4260 1840 6260 1855
rect 4260 1755 6260 1798
rect 4260 1725 4270 1755
rect 6250 1725 6260 1755
rect 4260 1720 6260 1725
rect 20 1355 2020 1360
rect 20 1325 30 1355
rect 2010 1325 2020 1355
rect 20 1282 2020 1325
rect 20 1225 2020 1240
rect 20 1195 2020 1200
rect 20 1165 30 1195
rect 2010 1165 2020 1195
rect 20 1122 2020 1165
rect 20 1060 2020 1080
rect 4260 1355 6260 1360
rect 4260 1325 4270 1355
rect 6250 1325 6260 1355
rect 4260 1282 6260 1325
rect 4260 1225 6260 1240
rect 4260 1195 6260 1200
rect 4260 1165 4270 1195
rect 6250 1165 6260 1195
rect 4260 1122 6260 1165
rect 4260 1060 6260 1080
rect 20 720 2020 740
rect 20 635 2020 678
rect 20 605 30 635
rect 2010 605 2020 635
rect 20 600 2020 605
rect 20 560 2020 575
rect 20 475 2020 518
rect 20 445 30 475
rect 2010 445 2020 475
rect 20 440 2020 445
rect 4260 720 6260 740
rect 4260 635 6260 678
rect 4260 605 4270 635
rect 6250 605 6260 635
rect 4260 600 6260 605
rect 4260 560 6260 575
rect 4260 475 6260 518
rect 4260 445 4270 475
rect 6250 445 6260 475
rect 4260 440 6260 445
rect 20 75 2020 80
rect 20 45 30 75
rect 2010 45 2020 75
rect 20 2 2020 45
rect 20 -55 2020 -40
rect 20 -85 2020 -80
rect 20 -115 30 -85
rect 2010 -115 2020 -85
rect 20 -158 2020 -115
rect 20 -220 2020 -200
rect 4260 75 6260 80
rect 4260 45 4270 75
rect 6250 45 6260 75
rect 4260 2 6260 45
rect 4260 -55 6260 -40
rect 4260 -85 6260 -80
rect 4260 -115 4270 -85
rect 6250 -115 6260 -85
rect 4260 -158 6260 -115
rect 4260 -220 6260 -200
<< polycont >>
rect 30 1885 2010 1915
rect 30 1725 2010 1755
rect 4270 1885 6250 1915
rect 4270 1725 6250 1755
rect 30 1325 2010 1355
rect 30 1165 2010 1195
rect 4270 1325 6250 1355
rect 4270 1165 6250 1195
rect 30 605 2010 635
rect 30 445 2010 475
rect 4270 605 6250 635
rect 4270 445 6250 475
rect 30 45 2010 75
rect 30 -115 2010 -85
rect 4270 45 6250 75
rect 4270 -115 6250 -85
<< locali >>
rect -240 2120 -180 2160
rect 2220 2120 4060 2160
rect 6460 2120 6520 2160
rect -240 2100 -200 2120
rect 2240 2100 2280 2120
rect -160 2070 -100 2080
rect -160 2050 -150 2070
rect -130 2050 -100 2070
rect -160 2040 -100 2050
rect 2140 2040 2200 2080
rect -160 2020 -120 2040
rect 2160 2020 2200 2040
rect -80 1990 -40 2000
rect -80 1970 -70 1990
rect -50 1970 -40 1990
rect -80 1958 -40 1970
rect 2080 1990 2120 2000
rect 2080 1970 2090 1990
rect 2110 1970 2120 1990
rect 2080 1958 2120 1970
rect 20 1915 2020 1920
rect 20 1885 30 1915
rect 2010 1885 2020 1915
rect 20 1880 2020 1885
rect -80 1830 -40 1840
rect -80 1810 -70 1830
rect -50 1810 -40 1830
rect -80 1798 -40 1810
rect 2080 1830 2120 1840
rect 2080 1810 2090 1830
rect 2110 1810 2120 1830
rect 2080 1798 2120 1810
rect 20 1755 2020 1760
rect 20 1725 30 1755
rect 2010 1725 2020 1755
rect 20 1720 2020 1725
rect -160 1640 -100 1680
rect 2140 1640 2200 1680
rect -240 1600 -200 1640
rect 2240 1600 2280 1640
rect -240 1560 -180 1600
rect 2220 1560 2280 1600
rect -240 1520 -200 1560
rect 2240 1520 2280 1560
rect -240 1480 -180 1520
rect 2220 1480 2280 1520
rect -240 1440 -200 1480
rect 2240 1440 2280 1480
rect -160 1400 -100 1440
rect 2140 1400 2200 1440
rect 20 1355 2020 1360
rect 20 1325 30 1355
rect 2010 1325 2020 1355
rect 20 1320 2020 1325
rect -80 1270 -40 1282
rect -80 1250 -70 1270
rect -50 1250 -40 1270
rect -80 1240 -40 1250
rect 2080 1270 2120 1282
rect 2080 1250 2090 1270
rect 2110 1250 2120 1270
rect 2080 1240 2120 1250
rect 20 1195 2020 1200
rect 20 1165 30 1195
rect 2010 1165 2020 1195
rect 20 1160 2020 1165
rect -80 1110 -40 1122
rect -80 1090 -70 1110
rect -50 1090 -40 1110
rect -80 1080 -40 1090
rect 2080 1110 2120 1122
rect 2080 1090 2090 1110
rect 2110 1090 2120 1110
rect 2080 1080 2120 1090
rect -160 1040 -120 1060
rect 2160 1040 2200 1060
rect -160 1000 -100 1040
rect 2140 1000 2200 1040
rect -240 960 -200 980
rect 2240 960 2280 980
rect -240 920 -180 960
rect 2220 920 2280 960
rect -240 880 -160 920
rect -120 880 -80 920
rect 2240 880 2280 920
rect -240 840 -180 880
rect 2220 840 2280 880
rect -240 820 -200 840
rect 2240 820 2280 840
rect -160 760 -100 800
rect 2140 760 2200 800
rect -160 740 -120 760
rect 2160 740 2200 760
rect -80 710 -40 720
rect -80 690 -70 710
rect -50 690 -40 710
rect -80 678 -40 690
rect 2080 710 2120 720
rect 2080 690 2090 710
rect 2110 690 2120 710
rect 2080 678 2120 690
rect 20 635 2020 640
rect 20 605 30 635
rect 2010 605 2020 635
rect 20 600 2020 605
rect -80 550 -40 560
rect -80 530 -70 550
rect -50 530 -40 550
rect -80 518 -40 530
rect 2080 550 2120 560
rect 2080 530 2090 550
rect 2110 530 2120 550
rect 2080 518 2120 530
rect 20 475 2020 480
rect 20 445 30 475
rect 2010 445 2020 475
rect 20 440 2020 445
rect -160 360 -100 400
rect 2140 360 2200 400
rect -240 320 -200 360
rect 2240 320 2280 360
rect -240 280 -180 320
rect 2220 280 2280 320
rect -240 240 -200 280
rect 2240 240 2280 280
rect -240 200 -180 240
rect 2220 200 2280 240
rect -240 160 -200 200
rect 2240 160 2280 200
rect -160 120 -100 160
rect 2140 120 2200 160
rect 20 75 2020 80
rect 20 45 30 75
rect 2010 45 2020 75
rect 20 40 2020 45
rect -80 -10 -40 2
rect -80 -30 -70 -10
rect -50 -30 -40 -10
rect -80 -40 -40 -30
rect 2080 -10 2120 2
rect 2080 -30 2090 -10
rect 2110 -30 2120 -10
rect 2080 -40 2120 -30
rect 20 -85 2020 -80
rect 20 -115 30 -85
rect 2010 -115 2020 -85
rect 20 -120 2020 -115
rect -80 -170 -40 -158
rect -80 -190 -70 -170
rect -50 -190 -40 -170
rect -80 -200 -40 -190
rect 2080 -170 2120 -158
rect 2080 -190 2090 -170
rect 2110 -190 2120 -170
rect 2080 -200 2120 -190
rect -160 -240 -120 -220
rect 2160 -240 2200 -220
rect -160 -250 -100 -240
rect -160 -270 -150 -250
rect -130 -270 -100 -250
rect -160 -280 -100 -270
rect 2140 -280 2200 -240
rect -240 -320 -200 -300
rect 2240 -320 2280 -300
rect 4000 2100 4040 2120
rect 6480 2100 6520 2120
rect 4080 2040 4140 2080
rect 6380 2070 6440 2080
rect 6380 2050 6410 2070
rect 6430 2050 6440 2070
rect 6380 2040 6440 2050
rect 4080 2020 4120 2040
rect 6400 2020 6440 2040
rect 4160 1990 4200 2000
rect 4160 1970 4170 1990
rect 4190 1970 4200 1990
rect 4160 1958 4200 1970
rect 6320 1990 6360 2000
rect 6320 1970 6330 1990
rect 6350 1970 6360 1990
rect 6320 1958 6360 1970
rect 4260 1915 6260 1920
rect 4260 1885 4270 1915
rect 6250 1885 6260 1915
rect 4260 1880 6260 1885
rect 4160 1830 4200 1840
rect 4160 1810 4170 1830
rect 4190 1810 4200 1830
rect 4160 1798 4200 1810
rect 6320 1830 6360 1840
rect 6320 1810 6330 1830
rect 6350 1810 6360 1830
rect 6320 1798 6360 1810
rect 4260 1755 6260 1760
rect 4260 1725 4270 1755
rect 6250 1725 6260 1755
rect 4260 1720 6260 1725
rect 4080 1640 4140 1680
rect 6380 1640 6440 1680
rect 4000 1600 4040 1640
rect 6480 1600 6520 1640
rect 4000 1560 4060 1600
rect 6460 1560 6520 1600
rect 4000 1520 4040 1560
rect 6480 1520 6520 1560
rect 4000 1480 4060 1520
rect 6460 1480 6520 1520
rect 4000 1440 4040 1480
rect 6480 1440 6520 1480
rect 4080 1400 4140 1440
rect 6380 1400 6440 1440
rect 4260 1355 6260 1360
rect 4260 1325 4270 1355
rect 6250 1325 6260 1355
rect 4260 1320 6260 1325
rect 4160 1270 4200 1282
rect 4160 1250 4170 1270
rect 4190 1250 4200 1270
rect 4160 1240 4200 1250
rect 6320 1270 6360 1282
rect 6320 1250 6330 1270
rect 6350 1250 6360 1270
rect 6320 1240 6360 1250
rect 4260 1195 6260 1200
rect 4260 1165 4270 1195
rect 6250 1165 6260 1195
rect 4260 1160 6260 1165
rect 4160 1110 4200 1122
rect 4160 1090 4170 1110
rect 4190 1090 4200 1110
rect 4160 1080 4200 1090
rect 6320 1110 6360 1122
rect 6320 1090 6330 1110
rect 6350 1090 6360 1110
rect 6320 1080 6360 1090
rect 4080 1040 4120 1060
rect 6400 1040 6440 1060
rect 4080 1000 4140 1040
rect 6380 1000 6440 1040
rect 4000 960 4040 980
rect 6480 960 6520 980
rect 4000 920 4060 960
rect 6460 920 6520 960
rect 4000 880 4040 920
rect 6360 880 6400 920
rect 6440 880 6520 920
rect 4000 840 4060 880
rect 6460 840 6520 880
rect 4000 820 4040 840
rect 6480 820 6520 840
rect 4080 760 4140 800
rect 6380 760 6440 800
rect 4080 740 4120 760
rect 6400 740 6440 760
rect 4160 710 4200 720
rect 4160 690 4170 710
rect 4190 690 4200 710
rect 4160 678 4200 690
rect 6320 710 6360 720
rect 6320 690 6330 710
rect 6350 690 6360 710
rect 6320 678 6360 690
rect 4260 635 6260 640
rect 4260 605 4270 635
rect 6250 605 6260 635
rect 4260 600 6260 605
rect 4160 550 4200 560
rect 4160 530 4170 550
rect 4190 530 4200 550
rect 4160 518 4200 530
rect 6320 550 6360 560
rect 6320 530 6330 550
rect 6350 530 6360 550
rect 6320 518 6360 530
rect 4260 475 6260 480
rect 4260 445 4270 475
rect 6250 445 6260 475
rect 4260 440 6260 445
rect 4080 360 4140 400
rect 6380 360 6440 400
rect 4000 320 4040 360
rect 6480 320 6520 360
rect 4000 280 4060 320
rect 6460 280 6520 320
rect 4000 240 4040 280
rect 6480 240 6520 280
rect 4000 200 4060 240
rect 6460 200 6520 240
rect 4000 160 4040 200
rect 6480 160 6520 200
rect 4080 120 4140 160
rect 6380 120 6440 160
rect 4260 75 6260 80
rect 4260 45 4270 75
rect 6250 45 6260 75
rect 4260 40 6260 45
rect 4160 -10 4200 2
rect 4160 -30 4170 -10
rect 4190 -30 4200 -10
rect 4160 -40 4200 -30
rect 6320 -10 6360 2
rect 6320 -30 6330 -10
rect 6350 -30 6360 -10
rect 6320 -40 6360 -30
rect 4260 -85 6260 -80
rect 4260 -115 4270 -85
rect 6250 -115 6260 -85
rect 4260 -120 6260 -115
rect 4160 -170 4200 -158
rect 4160 -190 4170 -170
rect 4190 -190 4200 -170
rect 4160 -200 4200 -190
rect 6320 -170 6360 -158
rect 6320 -190 6330 -170
rect 6350 -190 6360 -170
rect 6320 -200 6360 -190
rect 4080 -240 4120 -220
rect 6400 -240 6440 -220
rect 4080 -280 4140 -240
rect 6380 -250 6440 -240
rect 6380 -270 6410 -250
rect 6430 -270 6440 -250
rect 6380 -280 6440 -270
rect 4000 -320 4040 -300
rect 6480 -320 6520 -300
rect -240 -360 -180 -320
rect 2220 -360 4060 -320
rect 6460 -360 6520 -320
<< viali >>
rect -150 2050 -130 2070
rect -70 1970 -50 1990
rect 2090 1970 2110 1990
rect 30 1885 2010 1915
rect -70 1810 -50 1830
rect 2090 1810 2110 1830
rect 30 1725 2010 1755
rect 2090 1410 2110 1430
rect 30 1325 2010 1355
rect -70 1250 -50 1270
rect 2090 1250 2110 1270
rect 30 1165 2010 1195
rect -70 1090 -50 1110
rect 2090 1090 2110 1110
rect -160 880 -120 920
rect -70 690 -50 710
rect 2090 690 2110 710
rect 30 605 2010 635
rect -70 530 -50 550
rect 2090 530 2110 550
rect 30 445 2010 475
rect 2090 370 2110 390
rect 30 45 2010 75
rect -70 -30 -50 -10
rect 2090 -30 2110 -10
rect 30 -115 2010 -85
rect -70 -190 -50 -170
rect 2090 -190 2110 -170
rect -150 -270 -130 -250
rect 6410 2050 6430 2070
rect 4170 1970 4190 1990
rect 6330 1970 6350 1990
rect 4270 1885 6250 1915
rect 4170 1810 4190 1830
rect 6330 1810 6350 1830
rect 4270 1725 6250 1755
rect 4170 1410 4190 1430
rect 4270 1325 6250 1355
rect 4170 1250 4190 1270
rect 6330 1250 6350 1270
rect 4270 1165 6250 1195
rect 4170 1090 4190 1110
rect 6330 1090 6350 1110
rect 6400 880 6440 920
rect 4170 690 4190 710
rect 6330 690 6350 710
rect 4270 605 6250 635
rect 4170 530 4190 550
rect 6330 530 6350 550
rect 4270 445 6250 475
rect 4170 370 4190 390
rect 4270 45 6250 75
rect 4170 -30 4190 -10
rect 6330 -30 6350 -10
rect 4270 -115 6250 -85
rect 4170 -190 4190 -170
rect 6330 -190 6350 -170
rect 6410 -270 6430 -250
<< metal1 >>
rect -160 2075 -120 2080
rect -160 2045 -155 2075
rect -125 2045 -120 2075
rect -160 2040 -120 2045
rect 6400 2075 6440 2080
rect 6400 2045 6405 2075
rect 6435 2045 6440 2075
rect 6400 2040 6440 2045
rect -80 1990 -40 2000
rect -80 1970 -70 1990
rect -50 1970 -40 1990
rect -80 1830 -40 1970
rect 2080 1990 2120 2000
rect 2080 1970 2090 1990
rect 2110 1970 2120 1990
rect 20 1915 2020 1920
rect 20 1885 30 1915
rect 2010 1885 2020 1915
rect 20 1880 2020 1885
rect -80 1810 -70 1830
rect -50 1810 -40 1830
rect -80 1755 -40 1810
rect 2080 1830 2120 1970
rect 2080 1810 2090 1830
rect 2110 1810 2120 1830
rect -80 1725 -75 1755
rect -45 1725 -40 1755
rect -80 1270 -40 1725
rect 20 1755 2020 1760
rect 20 1725 30 1755
rect 2010 1725 2020 1755
rect 20 1720 2020 1725
rect 2080 1430 2120 1810
rect 2080 1410 2090 1430
rect 2110 1410 2120 1430
rect 20 1355 2020 1360
rect 20 1325 30 1355
rect 2010 1325 2020 1355
rect 20 1320 2020 1325
rect 2080 1355 2120 1410
rect 2080 1325 2085 1355
rect 2115 1325 2120 1355
rect -80 1250 -70 1270
rect -50 1250 -40 1270
rect -80 1110 -40 1250
rect 2080 1270 2120 1325
rect 2080 1250 2090 1270
rect 2110 1250 2120 1270
rect 20 1195 2020 1200
rect 20 1165 30 1195
rect 2010 1165 2020 1195
rect 20 1160 2020 1165
rect -80 1090 -70 1110
rect -50 1090 -40 1110
rect -80 1080 -40 1090
rect 2080 1110 2120 1250
rect 2080 1090 2090 1110
rect 2110 1090 2120 1110
rect 2080 1080 2120 1090
rect 4160 1990 4200 2000
rect 4160 1970 4170 1990
rect 4190 1970 4200 1990
rect 4160 1830 4200 1970
rect 6320 1990 6360 2000
rect 6320 1970 6330 1990
rect 6350 1970 6360 1990
rect 4260 1915 6260 1920
rect 4260 1885 4270 1915
rect 6250 1885 6260 1915
rect 4260 1880 6260 1885
rect 4160 1810 4170 1830
rect 4190 1810 4200 1830
rect 4160 1430 4200 1810
rect 6320 1830 6360 1970
rect 6320 1810 6330 1830
rect 6350 1810 6360 1830
rect 4260 1755 6260 1760
rect 4260 1725 4270 1755
rect 6250 1725 6260 1755
rect 4260 1720 6260 1725
rect 6320 1755 6360 1810
rect 6320 1725 6325 1755
rect 6355 1725 6360 1755
rect 4160 1410 4170 1430
rect 4190 1410 4200 1430
rect 4160 1355 4200 1410
rect 4160 1325 4165 1355
rect 4195 1325 4200 1355
rect 4160 1270 4200 1325
rect 4260 1355 6260 1360
rect 4260 1325 4270 1355
rect 6250 1325 6260 1355
rect 4260 1320 6260 1325
rect 4160 1250 4170 1270
rect 4190 1250 4200 1270
rect 4160 1110 4200 1250
rect 6320 1270 6360 1725
rect 6320 1250 6330 1270
rect 6350 1250 6360 1270
rect 4260 1195 6260 1200
rect 4260 1165 4270 1195
rect 6250 1165 6260 1195
rect 4260 1160 6260 1165
rect 4160 1090 4170 1110
rect 4190 1090 4200 1110
rect 4160 1080 4200 1090
rect 6320 1110 6360 1250
rect 6320 1090 6330 1110
rect 6350 1090 6360 1110
rect 6320 1080 6360 1090
rect -200 920 -80 960
rect -200 880 -160 920
rect -120 880 -80 920
rect -200 840 -80 880
rect 6360 920 6480 960
rect 6360 880 6400 920
rect 6440 880 6480 920
rect 6360 840 6480 880
rect -80 710 -40 720
rect -80 690 -70 710
rect -50 690 -40 710
rect -80 550 -40 690
rect 2080 710 2120 720
rect 2080 690 2090 710
rect 2110 690 2120 710
rect 20 635 2020 640
rect 20 605 30 635
rect 2010 605 2020 635
rect 20 600 2020 605
rect -80 530 -70 550
rect -50 530 -40 550
rect -80 75 -40 530
rect 2080 550 2120 690
rect 2080 530 2090 550
rect 2110 530 2120 550
rect 20 475 2020 480
rect 20 445 30 475
rect 2010 445 2020 475
rect 20 440 2020 445
rect 2080 475 2120 530
rect 2080 445 2085 475
rect 2115 445 2120 475
rect 2080 390 2120 445
rect 2080 370 2090 390
rect 2110 370 2120 390
rect -80 45 -75 75
rect -45 45 -40 75
rect -80 -10 -40 45
rect 20 75 2020 80
rect 20 45 30 75
rect 2010 45 2020 75
rect 20 40 2020 45
rect -80 -30 -70 -10
rect -50 -30 -40 -10
rect -80 -170 -40 -30
rect 2080 -10 2120 370
rect 2080 -30 2090 -10
rect 2110 -30 2120 -10
rect 20 -85 2020 -80
rect 20 -115 30 -85
rect 2010 -115 2020 -85
rect 20 -120 2020 -115
rect -80 -190 -70 -170
rect -50 -190 -40 -170
rect -80 -200 -40 -190
rect 2080 -170 2120 -30
rect 2080 -190 2090 -170
rect 2110 -190 2120 -170
rect 2080 -200 2120 -190
rect 4160 710 4200 720
rect 4160 690 4170 710
rect 4190 690 4200 710
rect 4160 550 4200 690
rect 6320 710 6360 720
rect 6320 690 6330 710
rect 6350 690 6360 710
rect 4260 635 6260 640
rect 4260 605 4270 635
rect 6250 605 6260 635
rect 4260 600 6260 605
rect 4160 530 4170 550
rect 4190 530 4200 550
rect 4160 475 4200 530
rect 6320 550 6360 690
rect 6320 530 6330 550
rect 6350 530 6360 550
rect 4160 445 4165 475
rect 4195 445 4200 475
rect 4160 390 4200 445
rect 4260 475 6260 480
rect 4260 445 4270 475
rect 6250 445 6260 475
rect 4260 440 6260 445
rect 4160 370 4170 390
rect 4190 370 4200 390
rect 4160 -10 4200 370
rect 4260 75 6260 80
rect 4260 45 4270 75
rect 6250 45 6260 75
rect 4260 40 6260 45
rect 6320 75 6360 530
rect 6320 45 6325 75
rect 6355 45 6360 75
rect 4160 -30 4170 -10
rect 4190 -30 4200 -10
rect 4160 -170 4200 -30
rect 6320 -10 6360 45
rect 6320 -30 6330 -10
rect 6350 -30 6360 -10
rect 4260 -85 6260 -80
rect 4260 -115 4270 -85
rect 6250 -115 6260 -85
rect 4260 -120 6260 -115
rect 4160 -190 4170 -170
rect 4190 -190 4200 -170
rect 4160 -200 4200 -190
rect 6320 -170 6360 -30
rect 6320 -190 6330 -170
rect 6350 -190 6360 -170
rect 6320 -200 6360 -190
rect -160 -245 -120 -240
rect -160 -275 -155 -245
rect -125 -275 -120 -245
rect -160 -280 -120 -275
rect 6400 -245 6440 -240
rect 6400 -275 6405 -245
rect 6435 -275 6440 -245
rect 6400 -280 6440 -275
<< via1 >>
rect -155 2070 -125 2075
rect -155 2050 -150 2070
rect -150 2050 -130 2070
rect -130 2050 -125 2070
rect -155 2045 -125 2050
rect 6405 2070 6435 2075
rect 6405 2050 6410 2070
rect 6410 2050 6430 2070
rect 6430 2050 6435 2070
rect 6405 2045 6435 2050
rect 30 1885 2010 1915
rect -75 1725 -45 1755
rect 30 1725 2010 1755
rect 30 1325 2010 1355
rect 2085 1325 2115 1355
rect 30 1165 2010 1195
rect 4270 1885 6250 1915
rect 4270 1725 6250 1755
rect 6325 1725 6355 1755
rect 4165 1325 4195 1355
rect 4270 1325 6250 1355
rect 4270 1165 6250 1195
rect -160 880 -120 920
rect 6400 880 6440 920
rect 30 605 2010 635
rect 30 445 2010 475
rect 2085 445 2115 475
rect -75 45 -45 75
rect 30 45 2010 75
rect 30 -115 2010 -85
rect 4270 605 6250 635
rect 4165 445 4195 475
rect 4270 445 6250 475
rect 4270 45 6250 75
rect 6325 45 6355 75
rect 4270 -115 6250 -85
rect -155 -250 -125 -245
rect -155 -270 -150 -250
rect -150 -270 -130 -250
rect -130 -270 -125 -250
rect -155 -275 -125 -270
rect 6405 -250 6435 -245
rect 6405 -270 6410 -250
rect 6410 -270 6430 -250
rect 6430 -270 6435 -250
rect 6405 -275 6435 -270
<< metal2 >>
rect 2320 2155 3960 2160
rect 2320 2125 2325 2155
rect 2355 2125 2485 2155
rect 2515 2125 2645 2155
rect 2675 2125 2805 2155
rect 2835 2125 2965 2155
rect 2995 2125 3125 2155
rect 3155 2125 3285 2155
rect 3315 2125 3445 2155
rect 3475 2125 3605 2155
rect 3635 2125 3765 2155
rect 3795 2125 3925 2155
rect 3955 2125 3960 2155
rect 2320 2120 3960 2125
rect -240 2075 6520 2080
rect -240 2045 -155 2075
rect -125 2045 3205 2075
rect 3235 2045 6405 2075
rect 6435 2045 6520 2075
rect -240 2040 6520 2045
rect 2320 1995 3960 2000
rect 2320 1965 2325 1995
rect 2355 1965 2485 1995
rect 2515 1965 2645 1995
rect 2675 1965 2805 1995
rect 2835 1965 2965 1995
rect 2995 1965 3125 1995
rect 3155 1965 3285 1995
rect 3315 1965 3445 1995
rect 3475 1965 3605 1995
rect 3635 1965 3765 1995
rect 3795 1965 3925 1995
rect 3955 1965 3960 1995
rect 2320 1960 3960 1965
rect -240 1915 6520 1920
rect -240 1885 30 1915
rect 2010 1885 3045 1915
rect 3075 1885 4270 1915
rect 6250 1885 6520 1915
rect -240 1880 6520 1885
rect 2320 1835 3960 1840
rect 2320 1805 2325 1835
rect 2355 1805 2485 1835
rect 2515 1805 2645 1835
rect 2675 1805 2805 1835
rect 2835 1805 2965 1835
rect 2995 1805 3125 1835
rect 3155 1805 3285 1835
rect 3315 1805 3445 1835
rect 3475 1805 3605 1835
rect 3635 1805 3765 1835
rect 3795 1805 3925 1835
rect 3955 1805 3960 1835
rect 2320 1800 3960 1805
rect -240 1755 2920 1760
rect -240 1725 -75 1755
rect -45 1725 30 1755
rect 2010 1725 2725 1755
rect 2755 1725 2920 1755
rect -240 1720 2920 1725
rect 2960 1755 3320 1760
rect 2960 1725 2965 1755
rect 2995 1725 3125 1755
rect 3155 1725 3285 1755
rect 3315 1725 3320 1755
rect 2960 1720 3320 1725
rect 3360 1755 6520 1760
rect 3360 1725 3845 1755
rect 3875 1725 4270 1755
rect 6250 1725 6325 1755
rect 6355 1725 6520 1755
rect 3360 1720 6520 1725
rect 2320 1675 3960 1680
rect 2320 1645 2325 1675
rect 2355 1645 2485 1675
rect 2515 1645 2645 1675
rect 2675 1645 2805 1675
rect 2835 1645 2965 1675
rect 2995 1645 3125 1675
rect 3155 1645 3285 1675
rect 3315 1645 3445 1675
rect 3475 1645 3605 1675
rect 3635 1645 3765 1675
rect 3795 1645 3925 1675
rect 3955 1645 3960 1675
rect 2320 1640 3960 1645
rect 2320 1595 3960 1600
rect 2320 1565 2325 1595
rect 2355 1565 2485 1595
rect 2515 1565 2645 1595
rect 2675 1565 2805 1595
rect 2835 1565 2965 1595
rect 2995 1565 3125 1595
rect 3155 1565 3285 1595
rect 3315 1565 3445 1595
rect 3475 1565 3605 1595
rect 3635 1565 3765 1595
rect 3795 1565 3925 1595
rect 3955 1565 3960 1595
rect 2320 1560 3960 1565
rect 2320 1515 3960 1520
rect 2320 1485 2885 1515
rect 2915 1485 3365 1515
rect 3395 1485 3960 1515
rect 2320 1480 3960 1485
rect 2320 1435 3960 1440
rect 2320 1405 2325 1435
rect 2355 1405 2485 1435
rect 2515 1405 2645 1435
rect 2675 1405 2805 1435
rect 2835 1405 2965 1435
rect 2995 1405 3125 1435
rect 3155 1405 3285 1435
rect 3315 1405 3445 1435
rect 3475 1405 3605 1435
rect 3635 1405 3765 1435
rect 3795 1405 3925 1435
rect 3955 1405 3960 1435
rect 2320 1400 3960 1405
rect -240 1355 2920 1360
rect -240 1325 30 1355
rect 2010 1325 2085 1355
rect 2115 1325 2885 1355
rect 2915 1325 2920 1355
rect -240 1320 2920 1325
rect 2960 1355 3320 1360
rect 2960 1325 2965 1355
rect 2995 1325 3125 1355
rect 3155 1325 3285 1355
rect 3315 1325 3320 1355
rect 2960 1320 3320 1325
rect 3360 1355 6520 1360
rect 3360 1325 3685 1355
rect 3715 1325 4165 1355
rect 4195 1325 4270 1355
rect 6250 1325 6520 1355
rect 3360 1320 6520 1325
rect 2320 1275 3960 1280
rect 2320 1245 2325 1275
rect 2355 1245 2485 1275
rect 2515 1245 2645 1275
rect 2675 1245 2805 1275
rect 2835 1245 2965 1275
rect 2995 1245 3125 1275
rect 3155 1245 3285 1275
rect 3315 1245 3445 1275
rect 3475 1245 3605 1275
rect 3635 1245 3765 1275
rect 3795 1245 3925 1275
rect 3955 1245 3960 1275
rect 2320 1240 3960 1245
rect -240 1195 6520 1200
rect -240 1165 30 1195
rect 2010 1165 3045 1195
rect 3075 1165 4270 1195
rect 6250 1165 6520 1195
rect -240 1160 6520 1165
rect 2320 1115 3960 1120
rect 2320 1085 2325 1115
rect 2355 1085 2485 1115
rect 2515 1085 2645 1115
rect 2675 1085 2805 1115
rect 2835 1085 2965 1115
rect 2995 1085 3125 1115
rect 3155 1085 3285 1115
rect 3315 1085 3445 1115
rect 3475 1085 3605 1115
rect 3635 1085 3765 1115
rect 3795 1085 3925 1115
rect 3955 1085 3960 1115
rect 2320 1080 3960 1085
rect -240 1000 2280 1040
rect 2320 1035 3960 1040
rect 2320 1005 2725 1035
rect 2755 1005 3525 1035
rect 3555 1005 3960 1035
rect 2320 1000 3960 1005
rect 4000 1000 6520 1040
rect -200 920 -80 960
rect 2320 955 3960 960
rect 2320 925 2325 955
rect 2355 925 2485 955
rect 2515 925 2645 955
rect 2675 925 2805 955
rect 2835 925 2965 955
rect 2995 925 3125 955
rect 3155 925 3285 955
rect 3315 925 3445 955
rect 3475 925 3605 955
rect 3635 925 3765 955
rect 3795 925 3925 955
rect 3955 925 3960 955
rect 2320 920 3960 925
rect 6360 920 6480 960
rect -200 880 -160 920
rect -120 880 -80 920
rect 6360 880 6400 920
rect 6440 880 6480 920
rect -200 840 -80 880
rect 2320 875 3960 880
rect 2320 845 2325 875
rect 2355 845 2485 875
rect 2515 845 2645 875
rect 2675 845 2805 875
rect 2835 845 2965 875
rect 2995 845 3125 875
rect 3155 845 3285 875
rect 3315 845 3445 875
rect 3475 845 3605 875
rect 3635 845 3765 875
rect 3795 845 3925 875
rect 3955 845 3960 875
rect 2320 840 3960 845
rect 6360 840 6480 880
rect -240 760 2280 800
rect 2320 795 3960 800
rect 2320 765 2405 795
rect 2435 765 3845 795
rect 3875 765 3960 795
rect 2320 760 3960 765
rect 4000 760 6520 800
rect 2320 715 3960 720
rect 2320 685 2325 715
rect 2355 685 2485 715
rect 2515 685 2645 715
rect 2675 685 2805 715
rect 2835 685 2965 715
rect 2995 685 3125 715
rect 3155 685 3285 715
rect 3315 685 3445 715
rect 3475 685 3605 715
rect 3635 685 3765 715
rect 3795 685 3925 715
rect 3955 685 3960 715
rect 2320 680 3960 685
rect -240 635 6520 640
rect -240 605 30 635
rect 2010 605 3045 635
rect 3075 605 4270 635
rect 6250 605 6520 635
rect -240 600 6520 605
rect 2320 555 3960 560
rect 2320 525 2325 555
rect 2355 525 2485 555
rect 2515 525 2645 555
rect 2675 525 2805 555
rect 2835 525 2965 555
rect 2995 525 3125 555
rect 3155 525 3285 555
rect 3315 525 3445 555
rect 3475 525 3605 555
rect 3635 525 3765 555
rect 3795 525 3925 555
rect 3955 525 3960 555
rect 2320 520 3960 525
rect -240 475 2920 480
rect -240 445 30 475
rect 2010 445 2085 475
rect 2115 445 2565 475
rect 2595 445 2920 475
rect -240 440 2920 445
rect 2960 475 3320 480
rect 2960 445 2965 475
rect 2995 445 3125 475
rect 3155 445 3285 475
rect 3315 445 3320 475
rect 2960 440 3320 445
rect 3360 475 6520 480
rect 3360 445 3365 475
rect 3395 445 4165 475
rect 4195 445 4270 475
rect 6250 445 6520 475
rect 3360 440 6520 445
rect 2320 395 3960 400
rect 2320 365 2325 395
rect 2355 365 2485 395
rect 2515 365 2645 395
rect 2675 365 2805 395
rect 2835 365 2965 395
rect 2995 365 3125 395
rect 3155 365 3285 395
rect 3315 365 3445 395
rect 3475 365 3605 395
rect 3635 365 3765 395
rect 3795 365 3925 395
rect 3955 365 3960 395
rect 2320 360 3960 365
rect 2320 315 3960 320
rect 2320 285 2565 315
rect 2595 285 3685 315
rect 3715 285 3960 315
rect 2320 280 3960 285
rect 2320 235 3960 240
rect 2320 205 2325 235
rect 2355 205 2485 235
rect 2515 205 2645 235
rect 2675 205 2805 235
rect 2835 205 2965 235
rect 2995 205 3125 235
rect 3155 205 3285 235
rect 3315 205 3445 235
rect 3475 205 3605 235
rect 3635 205 3765 235
rect 3795 205 3925 235
rect 3955 205 3960 235
rect 2320 200 3960 205
rect 2320 155 3960 160
rect 2320 125 2325 155
rect 2355 125 2485 155
rect 2515 125 2645 155
rect 2675 125 2805 155
rect 2835 125 2965 155
rect 2995 125 3125 155
rect 3155 125 3285 155
rect 3315 125 3445 155
rect 3475 125 3605 155
rect 3635 125 3765 155
rect 3795 125 3925 155
rect 3955 125 3960 155
rect 2320 120 3960 125
rect -240 75 2920 80
rect -240 45 -75 75
rect -45 45 30 75
rect 2010 45 2405 75
rect 2435 45 2920 75
rect -240 40 2920 45
rect 2960 75 3320 80
rect 2960 45 2965 75
rect 2995 45 3125 75
rect 3155 45 3285 75
rect 3315 45 3320 75
rect 2960 40 3320 45
rect 3360 75 6520 80
rect 3360 45 3525 75
rect 3555 45 4270 75
rect 6250 45 6325 75
rect 6355 45 6520 75
rect 3360 40 6520 45
rect 2320 -5 3960 0
rect 2320 -35 2325 -5
rect 2355 -35 2485 -5
rect 2515 -35 2645 -5
rect 2675 -35 2805 -5
rect 2835 -35 2965 -5
rect 2995 -35 3125 -5
rect 3155 -35 3285 -5
rect 3315 -35 3445 -5
rect 3475 -35 3605 -5
rect 3635 -35 3765 -5
rect 3795 -35 3925 -5
rect 3955 -35 3960 -5
rect 2320 -40 3960 -35
rect -240 -85 6520 -80
rect -240 -115 30 -85
rect 2010 -115 3045 -85
rect 3075 -115 4270 -85
rect 6250 -115 6520 -85
rect -240 -120 6520 -115
rect 2320 -165 3960 -160
rect 2320 -195 2325 -165
rect 2355 -195 2485 -165
rect 2515 -195 2645 -165
rect 2675 -195 2805 -165
rect 2835 -195 2965 -165
rect 2995 -195 3125 -165
rect 3155 -195 3285 -165
rect 3315 -195 3445 -165
rect 3475 -195 3605 -165
rect 3635 -195 3765 -165
rect 3795 -195 3925 -165
rect 3955 -195 3960 -165
rect 2320 -200 3960 -195
rect -240 -245 6520 -240
rect -240 -275 -155 -245
rect -125 -275 3205 -245
rect 3235 -275 6405 -245
rect 6435 -275 6520 -245
rect -240 -280 6520 -275
rect 2320 -325 3960 -320
rect 2320 -355 2325 -325
rect 2355 -355 2485 -325
rect 2515 -355 2645 -325
rect 2675 -355 2805 -325
rect 2835 -355 2965 -325
rect 2995 -355 3125 -325
rect 3155 -355 3285 -325
rect 3315 -355 3445 -325
rect 3475 -355 3605 -325
rect 3635 -355 3765 -325
rect 3795 -355 3925 -325
rect 3955 -355 3960 -325
rect 2320 -360 3960 -355
<< via2 >>
rect 2325 2125 2355 2155
rect 2485 2125 2515 2155
rect 2645 2125 2675 2155
rect 2805 2125 2835 2155
rect 2965 2125 2995 2155
rect 3125 2125 3155 2155
rect 3285 2125 3315 2155
rect 3445 2125 3475 2155
rect 3605 2125 3635 2155
rect 3765 2125 3795 2155
rect 3925 2125 3955 2155
rect 3205 2045 3235 2075
rect 2325 1965 2355 1995
rect 2485 1965 2515 1995
rect 2645 1965 2675 1995
rect 2805 1965 2835 1995
rect 2965 1965 2995 1995
rect 3125 1965 3155 1995
rect 3285 1965 3315 1995
rect 3445 1965 3475 1995
rect 3605 1965 3635 1995
rect 3765 1965 3795 1995
rect 3925 1965 3955 1995
rect 3045 1885 3075 1915
rect 2325 1805 2355 1835
rect 2485 1805 2515 1835
rect 2645 1805 2675 1835
rect 2805 1805 2835 1835
rect 2965 1805 2995 1835
rect 3125 1805 3155 1835
rect 3285 1805 3315 1835
rect 3445 1805 3475 1835
rect 3605 1805 3635 1835
rect 3765 1805 3795 1835
rect 3925 1805 3955 1835
rect 2725 1725 2755 1755
rect 2965 1725 2995 1755
rect 3125 1725 3155 1755
rect 3285 1725 3315 1755
rect 3845 1725 3875 1755
rect 2325 1645 2355 1675
rect 2485 1645 2515 1675
rect 2645 1645 2675 1675
rect 2805 1645 2835 1675
rect 2965 1645 2995 1675
rect 3125 1645 3155 1675
rect 3285 1645 3315 1675
rect 3445 1645 3475 1675
rect 3605 1645 3635 1675
rect 3765 1645 3795 1675
rect 3925 1645 3955 1675
rect 2325 1565 2355 1595
rect 2485 1565 2515 1595
rect 2645 1565 2675 1595
rect 2805 1565 2835 1595
rect 2965 1565 2995 1595
rect 3125 1565 3155 1595
rect 3285 1565 3315 1595
rect 3445 1565 3475 1595
rect 3605 1565 3635 1595
rect 3765 1565 3795 1595
rect 3925 1565 3955 1595
rect 2885 1485 2915 1515
rect 3365 1485 3395 1515
rect 2325 1405 2355 1435
rect 2485 1405 2515 1435
rect 2645 1405 2675 1435
rect 2805 1405 2835 1435
rect 2965 1405 2995 1435
rect 3125 1405 3155 1435
rect 3285 1405 3315 1435
rect 3445 1405 3475 1435
rect 3605 1405 3635 1435
rect 3765 1405 3795 1435
rect 3925 1405 3955 1435
rect 2885 1325 2915 1355
rect 2965 1325 2995 1355
rect 3125 1325 3155 1355
rect 3285 1325 3315 1355
rect 3685 1325 3715 1355
rect 2325 1245 2355 1275
rect 2485 1245 2515 1275
rect 2645 1245 2675 1275
rect 2805 1245 2835 1275
rect 2965 1245 2995 1275
rect 3125 1245 3155 1275
rect 3285 1245 3315 1275
rect 3445 1245 3475 1275
rect 3605 1245 3635 1275
rect 3765 1245 3795 1275
rect 3925 1245 3955 1275
rect 3045 1165 3075 1195
rect 2325 1085 2355 1115
rect 2485 1085 2515 1115
rect 2645 1085 2675 1115
rect 2805 1085 2835 1115
rect 2965 1085 2995 1115
rect 3125 1085 3155 1115
rect 3285 1085 3315 1115
rect 3445 1085 3475 1115
rect 3605 1085 3635 1115
rect 3765 1085 3795 1115
rect 3925 1085 3955 1115
rect 2725 1005 2755 1035
rect 3525 1005 3555 1035
rect 2325 925 2355 955
rect 2485 925 2515 955
rect 2645 925 2675 955
rect 2805 925 2835 955
rect 2965 925 2995 955
rect 3125 925 3155 955
rect 3285 925 3315 955
rect 3445 925 3475 955
rect 3605 925 3635 955
rect 3765 925 3795 955
rect 3925 925 3955 955
rect -160 880 -120 920
rect 6400 880 6440 920
rect 2325 845 2355 875
rect 2485 845 2515 875
rect 2645 845 2675 875
rect 2805 845 2835 875
rect 2965 845 2995 875
rect 3125 845 3155 875
rect 3285 845 3315 875
rect 3445 845 3475 875
rect 3605 845 3635 875
rect 3765 845 3795 875
rect 3925 845 3955 875
rect 2405 765 2435 795
rect 3845 765 3875 795
rect 2325 685 2355 715
rect 2485 685 2515 715
rect 2645 685 2675 715
rect 2805 685 2835 715
rect 2965 685 2995 715
rect 3125 685 3155 715
rect 3285 685 3315 715
rect 3445 685 3475 715
rect 3605 685 3635 715
rect 3765 685 3795 715
rect 3925 685 3955 715
rect 3045 605 3075 635
rect 2325 525 2355 555
rect 2485 525 2515 555
rect 2645 525 2675 555
rect 2805 525 2835 555
rect 2965 525 2995 555
rect 3125 525 3155 555
rect 3285 525 3315 555
rect 3445 525 3475 555
rect 3605 525 3635 555
rect 3765 525 3795 555
rect 3925 525 3955 555
rect 2565 445 2595 475
rect 2965 445 2995 475
rect 3125 445 3155 475
rect 3285 445 3315 475
rect 3365 445 3395 475
rect 2325 365 2355 395
rect 2485 365 2515 395
rect 2645 365 2675 395
rect 2805 365 2835 395
rect 2965 365 2995 395
rect 3125 365 3155 395
rect 3285 365 3315 395
rect 3445 365 3475 395
rect 3605 365 3635 395
rect 3765 365 3795 395
rect 3925 365 3955 395
rect 2565 285 2595 315
rect 3685 285 3715 315
rect 2325 205 2355 235
rect 2485 205 2515 235
rect 2645 205 2675 235
rect 2805 205 2835 235
rect 2965 205 2995 235
rect 3125 205 3155 235
rect 3285 205 3315 235
rect 3445 205 3475 235
rect 3605 205 3635 235
rect 3765 205 3795 235
rect 3925 205 3955 235
rect 2325 125 2355 155
rect 2485 125 2515 155
rect 2645 125 2675 155
rect 2805 125 2835 155
rect 2965 125 2995 155
rect 3125 125 3155 155
rect 3285 125 3315 155
rect 3445 125 3475 155
rect 3605 125 3635 155
rect 3765 125 3795 155
rect 3925 125 3955 155
rect 2405 45 2435 75
rect 2965 45 2995 75
rect 3125 45 3155 75
rect 3285 45 3315 75
rect 3525 45 3555 75
rect 2325 -35 2355 -5
rect 2485 -35 2515 -5
rect 2645 -35 2675 -5
rect 2805 -35 2835 -5
rect 2965 -35 2995 -5
rect 3125 -35 3155 -5
rect 3285 -35 3315 -5
rect 3445 -35 3475 -5
rect 3605 -35 3635 -5
rect 3765 -35 3795 -5
rect 3925 -35 3955 -5
rect 3045 -115 3075 -85
rect 2325 -195 2355 -165
rect 2485 -195 2515 -165
rect 2645 -195 2675 -165
rect 2805 -195 2835 -165
rect 2965 -195 2995 -165
rect 3125 -195 3155 -165
rect 3285 -195 3315 -165
rect 3445 -195 3475 -165
rect 3605 -195 3635 -165
rect 3765 -195 3795 -165
rect 3925 -195 3955 -165
rect 3205 -275 3235 -245
rect 2325 -355 2355 -325
rect 2485 -355 2515 -325
rect 2645 -355 2675 -325
rect 2805 -355 2835 -325
rect 2965 -355 2995 -325
rect 3125 -355 3155 -325
rect 3285 -355 3315 -325
rect 3445 -355 3475 -325
rect 3605 -355 3635 -325
rect 3765 -355 3795 -325
rect 3925 -355 3955 -325
<< metal3 >>
rect 2320 2156 2360 2160
rect 2320 2124 2324 2156
rect 2356 2124 2360 2156
rect 2320 1996 2360 2124
rect 2320 1964 2324 1996
rect 2356 1964 2360 1996
rect 2320 1836 2360 1964
rect 2320 1804 2324 1836
rect 2356 1804 2360 1836
rect 2320 1676 2360 1804
rect 2320 1644 2324 1676
rect 2356 1644 2360 1676
rect 2320 1596 2360 1644
rect 2320 1564 2324 1596
rect 2356 1564 2360 1596
rect 2320 1436 2360 1564
rect 2320 1404 2324 1436
rect 2356 1404 2360 1436
rect 2320 1276 2360 1404
rect 2320 1244 2324 1276
rect 2356 1244 2360 1276
rect 2320 1116 2360 1244
rect 2320 1084 2324 1116
rect 2356 1084 2360 1116
rect -200 920 -80 960
rect -200 880 -160 920
rect -120 880 -80 920
rect -200 840 -80 880
rect 2320 956 2360 1084
rect 2320 924 2324 956
rect 2356 924 2360 956
rect 2320 876 2360 924
rect 2320 844 2324 876
rect 2356 844 2360 876
rect 2320 716 2360 844
rect 2320 684 2324 716
rect 2356 684 2360 716
rect 2320 556 2360 684
rect 2320 524 2324 556
rect 2356 524 2360 556
rect 2320 396 2360 524
rect 2320 364 2324 396
rect 2356 364 2360 396
rect 2320 236 2360 364
rect 2320 204 2324 236
rect 2356 204 2360 236
rect 2320 156 2360 204
rect 2320 124 2324 156
rect 2356 124 2360 156
rect 2320 -4 2360 124
rect 2320 -36 2324 -4
rect 2356 -36 2360 -4
rect 2320 -164 2360 -36
rect 2320 -196 2324 -164
rect 2356 -196 2360 -164
rect 2320 -324 2360 -196
rect 2320 -356 2324 -324
rect 2356 -356 2360 -324
rect 2320 -360 2360 -356
rect 2400 795 2440 2160
rect 2400 765 2405 795
rect 2435 765 2440 795
rect 2400 75 2440 765
rect 2400 45 2405 75
rect 2435 45 2440 75
rect 2400 -360 2440 45
rect 2480 2156 2520 2160
rect 2480 2124 2484 2156
rect 2516 2124 2520 2156
rect 2480 1996 2520 2124
rect 2480 1964 2484 1996
rect 2516 1964 2520 1996
rect 2480 1836 2520 1964
rect 2480 1804 2484 1836
rect 2516 1804 2520 1836
rect 2480 1676 2520 1804
rect 2480 1644 2484 1676
rect 2516 1644 2520 1676
rect 2480 1596 2520 1644
rect 2480 1564 2484 1596
rect 2516 1564 2520 1596
rect 2480 1436 2520 1564
rect 2480 1404 2484 1436
rect 2516 1404 2520 1436
rect 2480 1276 2520 1404
rect 2480 1244 2484 1276
rect 2516 1244 2520 1276
rect 2480 1116 2520 1244
rect 2480 1084 2484 1116
rect 2516 1084 2520 1116
rect 2480 956 2520 1084
rect 2480 924 2484 956
rect 2516 924 2520 956
rect 2480 876 2520 924
rect 2480 844 2484 876
rect 2516 844 2520 876
rect 2480 716 2520 844
rect 2480 684 2484 716
rect 2516 684 2520 716
rect 2480 556 2520 684
rect 2480 524 2484 556
rect 2516 524 2520 556
rect 2480 396 2520 524
rect 2480 364 2484 396
rect 2516 364 2520 396
rect 2480 236 2520 364
rect 2480 204 2484 236
rect 2516 204 2520 236
rect 2480 156 2520 204
rect 2480 124 2484 156
rect 2516 124 2520 156
rect 2480 -4 2520 124
rect 2480 -36 2484 -4
rect 2516 -36 2520 -4
rect 2480 -164 2520 -36
rect 2480 -196 2484 -164
rect 2516 -196 2520 -164
rect 2480 -324 2520 -196
rect 2480 -356 2484 -324
rect 2516 -356 2520 -324
rect 2480 -360 2520 -356
rect 2560 475 2600 2160
rect 2560 445 2565 475
rect 2595 445 2600 475
rect 2560 315 2600 445
rect 2560 285 2565 315
rect 2595 285 2600 315
rect 2560 -360 2600 285
rect 2640 2156 2680 2160
rect 2640 2124 2644 2156
rect 2676 2124 2680 2156
rect 2640 1996 2680 2124
rect 2640 1964 2644 1996
rect 2676 1964 2680 1996
rect 2640 1836 2680 1964
rect 2640 1804 2644 1836
rect 2676 1804 2680 1836
rect 2640 1676 2680 1804
rect 2640 1644 2644 1676
rect 2676 1644 2680 1676
rect 2640 1596 2680 1644
rect 2640 1564 2644 1596
rect 2676 1564 2680 1596
rect 2640 1436 2680 1564
rect 2640 1404 2644 1436
rect 2676 1404 2680 1436
rect 2640 1276 2680 1404
rect 2640 1244 2644 1276
rect 2676 1244 2680 1276
rect 2640 1116 2680 1244
rect 2640 1084 2644 1116
rect 2676 1084 2680 1116
rect 2640 956 2680 1084
rect 2640 924 2644 956
rect 2676 924 2680 956
rect 2640 876 2680 924
rect 2640 844 2644 876
rect 2676 844 2680 876
rect 2640 716 2680 844
rect 2640 684 2644 716
rect 2676 684 2680 716
rect 2640 556 2680 684
rect 2640 524 2644 556
rect 2676 524 2680 556
rect 2640 396 2680 524
rect 2640 364 2644 396
rect 2676 364 2680 396
rect 2640 236 2680 364
rect 2640 204 2644 236
rect 2676 204 2680 236
rect 2640 156 2680 204
rect 2640 124 2644 156
rect 2676 124 2680 156
rect 2640 -4 2680 124
rect 2640 -36 2644 -4
rect 2676 -36 2680 -4
rect 2640 -164 2680 -36
rect 2640 -196 2644 -164
rect 2676 -196 2680 -164
rect 2640 -324 2680 -196
rect 2640 -356 2644 -324
rect 2676 -356 2680 -324
rect 2640 -360 2680 -356
rect 2720 1755 2760 2160
rect 2720 1725 2725 1755
rect 2755 1725 2760 1755
rect 2720 1035 2760 1725
rect 2720 1005 2725 1035
rect 2755 1005 2760 1035
rect 2720 -360 2760 1005
rect 2800 2156 2840 2160
rect 2800 2124 2804 2156
rect 2836 2124 2840 2156
rect 2800 1996 2840 2124
rect 2800 1964 2804 1996
rect 2836 1964 2840 1996
rect 2800 1836 2840 1964
rect 2800 1804 2804 1836
rect 2836 1804 2840 1836
rect 2800 1676 2840 1804
rect 2800 1644 2804 1676
rect 2836 1644 2840 1676
rect 2800 1596 2840 1644
rect 2800 1564 2804 1596
rect 2836 1564 2840 1596
rect 2800 1436 2840 1564
rect 2800 1404 2804 1436
rect 2836 1404 2840 1436
rect 2800 1276 2840 1404
rect 2800 1244 2804 1276
rect 2836 1244 2840 1276
rect 2800 1116 2840 1244
rect 2800 1084 2804 1116
rect 2836 1084 2840 1116
rect 2800 956 2840 1084
rect 2800 924 2804 956
rect 2836 924 2840 956
rect 2800 876 2840 924
rect 2800 844 2804 876
rect 2836 844 2840 876
rect 2800 716 2840 844
rect 2800 684 2804 716
rect 2836 684 2840 716
rect 2800 556 2840 684
rect 2800 524 2804 556
rect 2836 524 2840 556
rect 2800 396 2840 524
rect 2800 364 2804 396
rect 2836 364 2840 396
rect 2800 236 2840 364
rect 2800 204 2804 236
rect 2836 204 2840 236
rect 2800 156 2840 204
rect 2800 124 2804 156
rect 2836 124 2840 156
rect 2800 -4 2840 124
rect 2800 -36 2804 -4
rect 2836 -36 2840 -4
rect 2800 -164 2840 -36
rect 2800 -196 2804 -164
rect 2836 -196 2840 -164
rect 2800 -324 2840 -196
rect 2800 -356 2804 -324
rect 2836 -356 2840 -324
rect 2800 -360 2840 -356
rect 2880 1515 2920 2160
rect 2880 1485 2885 1515
rect 2915 1485 2920 1515
rect 2880 1355 2920 1485
rect 2880 1325 2885 1355
rect 2915 1325 2920 1355
rect 2880 -360 2920 1325
rect 2960 2156 3000 2160
rect 2960 2124 2964 2156
rect 2996 2124 3000 2156
rect 2960 1996 3000 2124
rect 2960 1964 2964 1996
rect 2996 1964 3000 1996
rect 2960 1836 3000 1964
rect 2960 1804 2964 1836
rect 2996 1804 3000 1836
rect 2960 1756 3000 1804
rect 2960 1724 2964 1756
rect 2996 1724 3000 1756
rect 2960 1676 3000 1724
rect 2960 1644 2964 1676
rect 2996 1644 3000 1676
rect 2960 1596 3000 1644
rect 2960 1564 2964 1596
rect 2996 1564 3000 1596
rect 2960 1436 3000 1564
rect 2960 1404 2964 1436
rect 2996 1404 3000 1436
rect 2960 1356 3000 1404
rect 2960 1324 2964 1356
rect 2996 1324 3000 1356
rect 2960 1276 3000 1324
rect 2960 1244 2964 1276
rect 2996 1244 3000 1276
rect 2960 1116 3000 1244
rect 2960 1084 2964 1116
rect 2996 1084 3000 1116
rect 2960 956 3000 1084
rect 2960 924 2964 956
rect 2996 924 3000 956
rect 2960 876 3000 924
rect 2960 844 2964 876
rect 2996 844 3000 876
rect 2960 716 3000 844
rect 2960 684 2964 716
rect 2996 684 3000 716
rect 2960 556 3000 684
rect 2960 524 2964 556
rect 2996 524 3000 556
rect 2960 476 3000 524
rect 2960 444 2964 476
rect 2996 444 3000 476
rect 2960 396 3000 444
rect 2960 364 2964 396
rect 2996 364 3000 396
rect 2960 236 3000 364
rect 2960 204 2964 236
rect 2996 204 3000 236
rect 2960 156 3000 204
rect 2960 124 2964 156
rect 2996 124 3000 156
rect 2960 76 3000 124
rect 2960 44 2964 76
rect 2996 44 3000 76
rect 2960 -4 3000 44
rect 2960 -36 2964 -4
rect 2996 -36 3000 -4
rect 2960 -164 3000 -36
rect 2960 -196 2964 -164
rect 2996 -196 3000 -164
rect 2960 -324 3000 -196
rect 2960 -356 2964 -324
rect 2996 -356 3000 -324
rect 2960 -360 3000 -356
rect 3040 1915 3080 2160
rect 3040 1885 3045 1915
rect 3075 1885 3080 1915
rect 3040 1195 3080 1885
rect 3040 1165 3045 1195
rect 3075 1165 3080 1195
rect 3040 635 3080 1165
rect 3040 605 3045 635
rect 3075 605 3080 635
rect 3040 -85 3080 605
rect 3040 -115 3045 -85
rect 3075 -115 3080 -85
rect 3040 -360 3080 -115
rect 3120 2156 3160 2160
rect 3120 2124 3124 2156
rect 3156 2124 3160 2156
rect 3120 1996 3160 2124
rect 3120 1964 3124 1996
rect 3156 1964 3160 1996
rect 3120 1836 3160 1964
rect 3120 1804 3124 1836
rect 3156 1804 3160 1836
rect 3120 1756 3160 1804
rect 3120 1724 3124 1756
rect 3156 1724 3160 1756
rect 3120 1676 3160 1724
rect 3120 1644 3124 1676
rect 3156 1644 3160 1676
rect 3120 1596 3160 1644
rect 3120 1564 3124 1596
rect 3156 1564 3160 1596
rect 3120 1436 3160 1564
rect 3120 1404 3124 1436
rect 3156 1404 3160 1436
rect 3120 1356 3160 1404
rect 3120 1324 3124 1356
rect 3156 1324 3160 1356
rect 3120 1276 3160 1324
rect 3120 1244 3124 1276
rect 3156 1244 3160 1276
rect 3120 1116 3160 1244
rect 3120 1084 3124 1116
rect 3156 1084 3160 1116
rect 3120 956 3160 1084
rect 3120 924 3124 956
rect 3156 924 3160 956
rect 3120 876 3160 924
rect 3120 844 3124 876
rect 3156 844 3160 876
rect 3120 716 3160 844
rect 3120 684 3124 716
rect 3156 684 3160 716
rect 3120 556 3160 684
rect 3120 524 3124 556
rect 3156 524 3160 556
rect 3120 476 3160 524
rect 3120 444 3124 476
rect 3156 444 3160 476
rect 3120 396 3160 444
rect 3120 364 3124 396
rect 3156 364 3160 396
rect 3120 236 3160 364
rect 3120 204 3124 236
rect 3156 204 3160 236
rect 3120 156 3160 204
rect 3120 124 3124 156
rect 3156 124 3160 156
rect 3120 76 3160 124
rect 3120 44 3124 76
rect 3156 44 3160 76
rect 3120 -4 3160 44
rect 3120 -36 3124 -4
rect 3156 -36 3160 -4
rect 3120 -164 3160 -36
rect 3120 -196 3124 -164
rect 3156 -196 3160 -164
rect 3120 -324 3160 -196
rect 3120 -356 3124 -324
rect 3156 -356 3160 -324
rect 3120 -360 3160 -356
rect 3200 2075 3240 2160
rect 3200 2045 3205 2075
rect 3235 2045 3240 2075
rect 3200 -245 3240 2045
rect 3200 -275 3205 -245
rect 3235 -275 3240 -245
rect 3200 -360 3240 -275
rect 3280 2156 3320 2160
rect 3280 2124 3284 2156
rect 3316 2124 3320 2156
rect 3280 1996 3320 2124
rect 3280 1964 3284 1996
rect 3316 1964 3320 1996
rect 3280 1836 3320 1964
rect 3280 1804 3284 1836
rect 3316 1804 3320 1836
rect 3280 1756 3320 1804
rect 3280 1724 3284 1756
rect 3316 1724 3320 1756
rect 3280 1676 3320 1724
rect 3280 1644 3284 1676
rect 3316 1644 3320 1676
rect 3280 1596 3320 1644
rect 3280 1564 3284 1596
rect 3316 1564 3320 1596
rect 3280 1436 3320 1564
rect 3280 1404 3284 1436
rect 3316 1404 3320 1436
rect 3280 1356 3320 1404
rect 3280 1324 3284 1356
rect 3316 1324 3320 1356
rect 3280 1276 3320 1324
rect 3280 1244 3284 1276
rect 3316 1244 3320 1276
rect 3280 1116 3320 1244
rect 3280 1084 3284 1116
rect 3316 1084 3320 1116
rect 3280 956 3320 1084
rect 3280 924 3284 956
rect 3316 924 3320 956
rect 3280 876 3320 924
rect 3280 844 3284 876
rect 3316 844 3320 876
rect 3280 716 3320 844
rect 3280 684 3284 716
rect 3316 684 3320 716
rect 3280 556 3320 684
rect 3280 524 3284 556
rect 3316 524 3320 556
rect 3280 476 3320 524
rect 3280 444 3284 476
rect 3316 444 3320 476
rect 3280 396 3320 444
rect 3280 364 3284 396
rect 3316 364 3320 396
rect 3280 236 3320 364
rect 3280 204 3284 236
rect 3316 204 3320 236
rect 3280 156 3320 204
rect 3280 124 3284 156
rect 3316 124 3320 156
rect 3280 76 3320 124
rect 3280 44 3284 76
rect 3316 44 3320 76
rect 3280 -4 3320 44
rect 3280 -36 3284 -4
rect 3316 -36 3320 -4
rect 3280 -164 3320 -36
rect 3280 -196 3284 -164
rect 3316 -196 3320 -164
rect 3280 -324 3320 -196
rect 3280 -356 3284 -324
rect 3316 -356 3320 -324
rect 3280 -360 3320 -356
rect 3360 1515 3400 2160
rect 3360 1485 3365 1515
rect 3395 1485 3400 1515
rect 3360 475 3400 1485
rect 3360 445 3365 475
rect 3395 445 3400 475
rect 3360 -360 3400 445
rect 3440 2156 3480 2160
rect 3440 2124 3444 2156
rect 3476 2124 3480 2156
rect 3440 1996 3480 2124
rect 3440 1964 3444 1996
rect 3476 1964 3480 1996
rect 3440 1836 3480 1964
rect 3440 1804 3444 1836
rect 3476 1804 3480 1836
rect 3440 1676 3480 1804
rect 3440 1644 3444 1676
rect 3476 1644 3480 1676
rect 3440 1596 3480 1644
rect 3440 1564 3444 1596
rect 3476 1564 3480 1596
rect 3440 1436 3480 1564
rect 3440 1404 3444 1436
rect 3476 1404 3480 1436
rect 3440 1276 3480 1404
rect 3440 1244 3444 1276
rect 3476 1244 3480 1276
rect 3440 1116 3480 1244
rect 3440 1084 3444 1116
rect 3476 1084 3480 1116
rect 3440 956 3480 1084
rect 3440 924 3444 956
rect 3476 924 3480 956
rect 3440 876 3480 924
rect 3440 844 3444 876
rect 3476 844 3480 876
rect 3440 716 3480 844
rect 3440 684 3444 716
rect 3476 684 3480 716
rect 3440 556 3480 684
rect 3440 524 3444 556
rect 3476 524 3480 556
rect 3440 396 3480 524
rect 3440 364 3444 396
rect 3476 364 3480 396
rect 3440 236 3480 364
rect 3440 204 3444 236
rect 3476 204 3480 236
rect 3440 156 3480 204
rect 3440 124 3444 156
rect 3476 124 3480 156
rect 3440 -4 3480 124
rect 3440 -36 3444 -4
rect 3476 -36 3480 -4
rect 3440 -164 3480 -36
rect 3440 -196 3444 -164
rect 3476 -196 3480 -164
rect 3440 -324 3480 -196
rect 3440 -356 3444 -324
rect 3476 -356 3480 -324
rect 3440 -360 3480 -356
rect 3520 1035 3560 2160
rect 3520 1005 3525 1035
rect 3555 1005 3560 1035
rect 3520 75 3560 1005
rect 3520 45 3525 75
rect 3555 45 3560 75
rect 3520 -360 3560 45
rect 3600 2156 3640 2160
rect 3600 2124 3604 2156
rect 3636 2124 3640 2156
rect 3600 1996 3640 2124
rect 3600 1964 3604 1996
rect 3636 1964 3640 1996
rect 3600 1836 3640 1964
rect 3600 1804 3604 1836
rect 3636 1804 3640 1836
rect 3600 1676 3640 1804
rect 3600 1644 3604 1676
rect 3636 1644 3640 1676
rect 3600 1596 3640 1644
rect 3600 1564 3604 1596
rect 3636 1564 3640 1596
rect 3600 1436 3640 1564
rect 3600 1404 3604 1436
rect 3636 1404 3640 1436
rect 3600 1276 3640 1404
rect 3600 1244 3604 1276
rect 3636 1244 3640 1276
rect 3600 1116 3640 1244
rect 3600 1084 3604 1116
rect 3636 1084 3640 1116
rect 3600 956 3640 1084
rect 3600 924 3604 956
rect 3636 924 3640 956
rect 3600 876 3640 924
rect 3600 844 3604 876
rect 3636 844 3640 876
rect 3600 716 3640 844
rect 3600 684 3604 716
rect 3636 684 3640 716
rect 3600 556 3640 684
rect 3600 524 3604 556
rect 3636 524 3640 556
rect 3600 396 3640 524
rect 3600 364 3604 396
rect 3636 364 3640 396
rect 3600 236 3640 364
rect 3600 204 3604 236
rect 3636 204 3640 236
rect 3600 156 3640 204
rect 3600 124 3604 156
rect 3636 124 3640 156
rect 3600 -4 3640 124
rect 3600 -36 3604 -4
rect 3636 -36 3640 -4
rect 3600 -164 3640 -36
rect 3600 -196 3604 -164
rect 3636 -196 3640 -164
rect 3600 -324 3640 -196
rect 3600 -356 3604 -324
rect 3636 -356 3640 -324
rect 3600 -360 3640 -356
rect 3680 1355 3720 2160
rect 3680 1325 3685 1355
rect 3715 1325 3720 1355
rect 3680 315 3720 1325
rect 3680 285 3685 315
rect 3715 285 3720 315
rect 3680 -360 3720 285
rect 3760 2156 3800 2160
rect 3760 2124 3764 2156
rect 3796 2124 3800 2156
rect 3760 1996 3800 2124
rect 3760 1964 3764 1996
rect 3796 1964 3800 1996
rect 3760 1836 3800 1964
rect 3760 1804 3764 1836
rect 3796 1804 3800 1836
rect 3760 1676 3800 1804
rect 3760 1644 3764 1676
rect 3796 1644 3800 1676
rect 3760 1596 3800 1644
rect 3760 1564 3764 1596
rect 3796 1564 3800 1596
rect 3760 1436 3800 1564
rect 3760 1404 3764 1436
rect 3796 1404 3800 1436
rect 3760 1276 3800 1404
rect 3760 1244 3764 1276
rect 3796 1244 3800 1276
rect 3760 1116 3800 1244
rect 3760 1084 3764 1116
rect 3796 1084 3800 1116
rect 3760 956 3800 1084
rect 3760 924 3764 956
rect 3796 924 3800 956
rect 3760 876 3800 924
rect 3760 844 3764 876
rect 3796 844 3800 876
rect 3760 716 3800 844
rect 3760 684 3764 716
rect 3796 684 3800 716
rect 3760 556 3800 684
rect 3760 524 3764 556
rect 3796 524 3800 556
rect 3760 396 3800 524
rect 3760 364 3764 396
rect 3796 364 3800 396
rect 3760 236 3800 364
rect 3760 204 3764 236
rect 3796 204 3800 236
rect 3760 156 3800 204
rect 3760 124 3764 156
rect 3796 124 3800 156
rect 3760 -4 3800 124
rect 3760 -36 3764 -4
rect 3796 -36 3800 -4
rect 3760 -164 3800 -36
rect 3760 -196 3764 -164
rect 3796 -196 3800 -164
rect 3760 -324 3800 -196
rect 3760 -356 3764 -324
rect 3796 -356 3800 -324
rect 3760 -360 3800 -356
rect 3840 1755 3880 2160
rect 3840 1725 3845 1755
rect 3875 1725 3880 1755
rect 3840 795 3880 1725
rect 3840 765 3845 795
rect 3875 765 3880 795
rect 3840 -360 3880 765
rect 3920 2156 3960 2160
rect 3920 2124 3924 2156
rect 3956 2124 3960 2156
rect 3920 1996 3960 2124
rect 3920 1964 3924 1996
rect 3956 1964 3960 1996
rect 3920 1836 3960 1964
rect 3920 1804 3924 1836
rect 3956 1804 3960 1836
rect 3920 1676 3960 1804
rect 3920 1644 3924 1676
rect 3956 1644 3960 1676
rect 3920 1596 3960 1644
rect 3920 1564 3924 1596
rect 3956 1564 3960 1596
rect 3920 1436 3960 1564
rect 3920 1404 3924 1436
rect 3956 1404 3960 1436
rect 3920 1276 3960 1404
rect 3920 1244 3924 1276
rect 3956 1244 3960 1276
rect 3920 1116 3960 1244
rect 3920 1084 3924 1116
rect 3956 1084 3960 1116
rect 3920 956 3960 1084
rect 3920 924 3924 956
rect 3956 924 3960 956
rect 3920 876 3960 924
rect 3920 844 3924 876
rect 3956 844 3960 876
rect 3920 716 3960 844
rect 6360 920 6480 960
rect 6360 880 6400 920
rect 6440 880 6480 920
rect 6360 840 6480 880
rect 3920 684 3924 716
rect 3956 684 3960 716
rect 3920 556 3960 684
rect 3920 524 3924 556
rect 3956 524 3960 556
rect 3920 396 3960 524
rect 3920 364 3924 396
rect 3956 364 3960 396
rect 3920 236 3960 364
rect 3920 204 3924 236
rect 3956 204 3960 236
rect 3920 156 3960 204
rect 3920 124 3924 156
rect 3956 124 3960 156
rect 3920 -4 3960 124
rect 3920 -36 3924 -4
rect 3956 -36 3960 -4
rect 3920 -164 3960 -36
rect 3920 -196 3924 -164
rect 3956 -196 3960 -164
rect 3920 -324 3960 -196
rect 3920 -356 3924 -324
rect 3956 -356 3960 -324
rect 3920 -360 3960 -356
<< via3 >>
rect 2324 2155 2356 2156
rect 2324 2125 2325 2155
rect 2325 2125 2355 2155
rect 2355 2125 2356 2155
rect 2324 2124 2356 2125
rect 2324 1995 2356 1996
rect 2324 1965 2325 1995
rect 2325 1965 2355 1995
rect 2355 1965 2356 1995
rect 2324 1964 2356 1965
rect 2324 1835 2356 1836
rect 2324 1805 2325 1835
rect 2325 1805 2355 1835
rect 2355 1805 2356 1835
rect 2324 1804 2356 1805
rect 2324 1675 2356 1676
rect 2324 1645 2325 1675
rect 2325 1645 2355 1675
rect 2355 1645 2356 1675
rect 2324 1644 2356 1645
rect 2324 1595 2356 1596
rect 2324 1565 2325 1595
rect 2325 1565 2355 1595
rect 2355 1565 2356 1595
rect 2324 1564 2356 1565
rect 2324 1435 2356 1436
rect 2324 1405 2325 1435
rect 2325 1405 2355 1435
rect 2355 1405 2356 1435
rect 2324 1404 2356 1405
rect 2324 1275 2356 1276
rect 2324 1245 2325 1275
rect 2325 1245 2355 1275
rect 2355 1245 2356 1275
rect 2324 1244 2356 1245
rect 2324 1115 2356 1116
rect 2324 1085 2325 1115
rect 2325 1085 2355 1115
rect 2355 1085 2356 1115
rect 2324 1084 2356 1085
rect -160 880 -120 920
rect 2324 955 2356 956
rect 2324 925 2325 955
rect 2325 925 2355 955
rect 2355 925 2356 955
rect 2324 924 2356 925
rect 2324 875 2356 876
rect 2324 845 2325 875
rect 2325 845 2355 875
rect 2355 845 2356 875
rect 2324 844 2356 845
rect 2324 715 2356 716
rect 2324 685 2325 715
rect 2325 685 2355 715
rect 2355 685 2356 715
rect 2324 684 2356 685
rect 2324 555 2356 556
rect 2324 525 2325 555
rect 2325 525 2355 555
rect 2355 525 2356 555
rect 2324 524 2356 525
rect 2324 395 2356 396
rect 2324 365 2325 395
rect 2325 365 2355 395
rect 2355 365 2356 395
rect 2324 364 2356 365
rect 2324 235 2356 236
rect 2324 205 2325 235
rect 2325 205 2355 235
rect 2355 205 2356 235
rect 2324 204 2356 205
rect 2324 155 2356 156
rect 2324 125 2325 155
rect 2325 125 2355 155
rect 2355 125 2356 155
rect 2324 124 2356 125
rect 2324 -5 2356 -4
rect 2324 -35 2325 -5
rect 2325 -35 2355 -5
rect 2355 -35 2356 -5
rect 2324 -36 2356 -35
rect 2324 -165 2356 -164
rect 2324 -195 2325 -165
rect 2325 -195 2355 -165
rect 2355 -195 2356 -165
rect 2324 -196 2356 -195
rect 2324 -325 2356 -324
rect 2324 -355 2325 -325
rect 2325 -355 2355 -325
rect 2355 -355 2356 -325
rect 2324 -356 2356 -355
rect 2484 2155 2516 2156
rect 2484 2125 2485 2155
rect 2485 2125 2515 2155
rect 2515 2125 2516 2155
rect 2484 2124 2516 2125
rect 2484 1995 2516 1996
rect 2484 1965 2485 1995
rect 2485 1965 2515 1995
rect 2515 1965 2516 1995
rect 2484 1964 2516 1965
rect 2484 1835 2516 1836
rect 2484 1805 2485 1835
rect 2485 1805 2515 1835
rect 2515 1805 2516 1835
rect 2484 1804 2516 1805
rect 2484 1675 2516 1676
rect 2484 1645 2485 1675
rect 2485 1645 2515 1675
rect 2515 1645 2516 1675
rect 2484 1644 2516 1645
rect 2484 1595 2516 1596
rect 2484 1565 2485 1595
rect 2485 1565 2515 1595
rect 2515 1565 2516 1595
rect 2484 1564 2516 1565
rect 2484 1435 2516 1436
rect 2484 1405 2485 1435
rect 2485 1405 2515 1435
rect 2515 1405 2516 1435
rect 2484 1404 2516 1405
rect 2484 1275 2516 1276
rect 2484 1245 2485 1275
rect 2485 1245 2515 1275
rect 2515 1245 2516 1275
rect 2484 1244 2516 1245
rect 2484 1115 2516 1116
rect 2484 1085 2485 1115
rect 2485 1085 2515 1115
rect 2515 1085 2516 1115
rect 2484 1084 2516 1085
rect 2484 955 2516 956
rect 2484 925 2485 955
rect 2485 925 2515 955
rect 2515 925 2516 955
rect 2484 924 2516 925
rect 2484 875 2516 876
rect 2484 845 2485 875
rect 2485 845 2515 875
rect 2515 845 2516 875
rect 2484 844 2516 845
rect 2484 715 2516 716
rect 2484 685 2485 715
rect 2485 685 2515 715
rect 2515 685 2516 715
rect 2484 684 2516 685
rect 2484 555 2516 556
rect 2484 525 2485 555
rect 2485 525 2515 555
rect 2515 525 2516 555
rect 2484 524 2516 525
rect 2484 395 2516 396
rect 2484 365 2485 395
rect 2485 365 2515 395
rect 2515 365 2516 395
rect 2484 364 2516 365
rect 2484 235 2516 236
rect 2484 205 2485 235
rect 2485 205 2515 235
rect 2515 205 2516 235
rect 2484 204 2516 205
rect 2484 155 2516 156
rect 2484 125 2485 155
rect 2485 125 2515 155
rect 2515 125 2516 155
rect 2484 124 2516 125
rect 2484 -5 2516 -4
rect 2484 -35 2485 -5
rect 2485 -35 2515 -5
rect 2515 -35 2516 -5
rect 2484 -36 2516 -35
rect 2484 -165 2516 -164
rect 2484 -195 2485 -165
rect 2485 -195 2515 -165
rect 2515 -195 2516 -165
rect 2484 -196 2516 -195
rect 2484 -325 2516 -324
rect 2484 -355 2485 -325
rect 2485 -355 2515 -325
rect 2515 -355 2516 -325
rect 2484 -356 2516 -355
rect 2644 2155 2676 2156
rect 2644 2125 2645 2155
rect 2645 2125 2675 2155
rect 2675 2125 2676 2155
rect 2644 2124 2676 2125
rect 2644 1995 2676 1996
rect 2644 1965 2645 1995
rect 2645 1965 2675 1995
rect 2675 1965 2676 1995
rect 2644 1964 2676 1965
rect 2644 1835 2676 1836
rect 2644 1805 2645 1835
rect 2645 1805 2675 1835
rect 2675 1805 2676 1835
rect 2644 1804 2676 1805
rect 2644 1675 2676 1676
rect 2644 1645 2645 1675
rect 2645 1645 2675 1675
rect 2675 1645 2676 1675
rect 2644 1644 2676 1645
rect 2644 1595 2676 1596
rect 2644 1565 2645 1595
rect 2645 1565 2675 1595
rect 2675 1565 2676 1595
rect 2644 1564 2676 1565
rect 2644 1435 2676 1436
rect 2644 1405 2645 1435
rect 2645 1405 2675 1435
rect 2675 1405 2676 1435
rect 2644 1404 2676 1405
rect 2644 1275 2676 1276
rect 2644 1245 2645 1275
rect 2645 1245 2675 1275
rect 2675 1245 2676 1275
rect 2644 1244 2676 1245
rect 2644 1115 2676 1116
rect 2644 1085 2645 1115
rect 2645 1085 2675 1115
rect 2675 1085 2676 1115
rect 2644 1084 2676 1085
rect 2644 955 2676 956
rect 2644 925 2645 955
rect 2645 925 2675 955
rect 2675 925 2676 955
rect 2644 924 2676 925
rect 2644 875 2676 876
rect 2644 845 2645 875
rect 2645 845 2675 875
rect 2675 845 2676 875
rect 2644 844 2676 845
rect 2644 715 2676 716
rect 2644 685 2645 715
rect 2645 685 2675 715
rect 2675 685 2676 715
rect 2644 684 2676 685
rect 2644 555 2676 556
rect 2644 525 2645 555
rect 2645 525 2675 555
rect 2675 525 2676 555
rect 2644 524 2676 525
rect 2644 395 2676 396
rect 2644 365 2645 395
rect 2645 365 2675 395
rect 2675 365 2676 395
rect 2644 364 2676 365
rect 2644 235 2676 236
rect 2644 205 2645 235
rect 2645 205 2675 235
rect 2675 205 2676 235
rect 2644 204 2676 205
rect 2644 155 2676 156
rect 2644 125 2645 155
rect 2645 125 2675 155
rect 2675 125 2676 155
rect 2644 124 2676 125
rect 2644 -5 2676 -4
rect 2644 -35 2645 -5
rect 2645 -35 2675 -5
rect 2675 -35 2676 -5
rect 2644 -36 2676 -35
rect 2644 -165 2676 -164
rect 2644 -195 2645 -165
rect 2645 -195 2675 -165
rect 2675 -195 2676 -165
rect 2644 -196 2676 -195
rect 2644 -325 2676 -324
rect 2644 -355 2645 -325
rect 2645 -355 2675 -325
rect 2675 -355 2676 -325
rect 2644 -356 2676 -355
rect 2804 2155 2836 2156
rect 2804 2125 2805 2155
rect 2805 2125 2835 2155
rect 2835 2125 2836 2155
rect 2804 2124 2836 2125
rect 2804 1995 2836 1996
rect 2804 1965 2805 1995
rect 2805 1965 2835 1995
rect 2835 1965 2836 1995
rect 2804 1964 2836 1965
rect 2804 1835 2836 1836
rect 2804 1805 2805 1835
rect 2805 1805 2835 1835
rect 2835 1805 2836 1835
rect 2804 1804 2836 1805
rect 2804 1675 2836 1676
rect 2804 1645 2805 1675
rect 2805 1645 2835 1675
rect 2835 1645 2836 1675
rect 2804 1644 2836 1645
rect 2804 1595 2836 1596
rect 2804 1565 2805 1595
rect 2805 1565 2835 1595
rect 2835 1565 2836 1595
rect 2804 1564 2836 1565
rect 2804 1435 2836 1436
rect 2804 1405 2805 1435
rect 2805 1405 2835 1435
rect 2835 1405 2836 1435
rect 2804 1404 2836 1405
rect 2804 1275 2836 1276
rect 2804 1245 2805 1275
rect 2805 1245 2835 1275
rect 2835 1245 2836 1275
rect 2804 1244 2836 1245
rect 2804 1115 2836 1116
rect 2804 1085 2805 1115
rect 2805 1085 2835 1115
rect 2835 1085 2836 1115
rect 2804 1084 2836 1085
rect 2804 955 2836 956
rect 2804 925 2805 955
rect 2805 925 2835 955
rect 2835 925 2836 955
rect 2804 924 2836 925
rect 2804 875 2836 876
rect 2804 845 2805 875
rect 2805 845 2835 875
rect 2835 845 2836 875
rect 2804 844 2836 845
rect 2804 715 2836 716
rect 2804 685 2805 715
rect 2805 685 2835 715
rect 2835 685 2836 715
rect 2804 684 2836 685
rect 2804 555 2836 556
rect 2804 525 2805 555
rect 2805 525 2835 555
rect 2835 525 2836 555
rect 2804 524 2836 525
rect 2804 395 2836 396
rect 2804 365 2805 395
rect 2805 365 2835 395
rect 2835 365 2836 395
rect 2804 364 2836 365
rect 2804 235 2836 236
rect 2804 205 2805 235
rect 2805 205 2835 235
rect 2835 205 2836 235
rect 2804 204 2836 205
rect 2804 155 2836 156
rect 2804 125 2805 155
rect 2805 125 2835 155
rect 2835 125 2836 155
rect 2804 124 2836 125
rect 2804 -5 2836 -4
rect 2804 -35 2805 -5
rect 2805 -35 2835 -5
rect 2835 -35 2836 -5
rect 2804 -36 2836 -35
rect 2804 -165 2836 -164
rect 2804 -195 2805 -165
rect 2805 -195 2835 -165
rect 2835 -195 2836 -165
rect 2804 -196 2836 -195
rect 2804 -325 2836 -324
rect 2804 -355 2805 -325
rect 2805 -355 2835 -325
rect 2835 -355 2836 -325
rect 2804 -356 2836 -355
rect 2964 2155 2996 2156
rect 2964 2125 2965 2155
rect 2965 2125 2995 2155
rect 2995 2125 2996 2155
rect 2964 2124 2996 2125
rect 2964 1995 2996 1996
rect 2964 1965 2965 1995
rect 2965 1965 2995 1995
rect 2995 1965 2996 1995
rect 2964 1964 2996 1965
rect 2964 1835 2996 1836
rect 2964 1805 2965 1835
rect 2965 1805 2995 1835
rect 2995 1805 2996 1835
rect 2964 1804 2996 1805
rect 2964 1755 2996 1756
rect 2964 1725 2965 1755
rect 2965 1725 2995 1755
rect 2995 1725 2996 1755
rect 2964 1724 2996 1725
rect 2964 1675 2996 1676
rect 2964 1645 2965 1675
rect 2965 1645 2995 1675
rect 2995 1645 2996 1675
rect 2964 1644 2996 1645
rect 2964 1595 2996 1596
rect 2964 1565 2965 1595
rect 2965 1565 2995 1595
rect 2995 1565 2996 1595
rect 2964 1564 2996 1565
rect 2964 1435 2996 1436
rect 2964 1405 2965 1435
rect 2965 1405 2995 1435
rect 2995 1405 2996 1435
rect 2964 1404 2996 1405
rect 2964 1355 2996 1356
rect 2964 1325 2965 1355
rect 2965 1325 2995 1355
rect 2995 1325 2996 1355
rect 2964 1324 2996 1325
rect 2964 1275 2996 1276
rect 2964 1245 2965 1275
rect 2965 1245 2995 1275
rect 2995 1245 2996 1275
rect 2964 1244 2996 1245
rect 2964 1115 2996 1116
rect 2964 1085 2965 1115
rect 2965 1085 2995 1115
rect 2995 1085 2996 1115
rect 2964 1084 2996 1085
rect 2964 955 2996 956
rect 2964 925 2965 955
rect 2965 925 2995 955
rect 2995 925 2996 955
rect 2964 924 2996 925
rect 2964 875 2996 876
rect 2964 845 2965 875
rect 2965 845 2995 875
rect 2995 845 2996 875
rect 2964 844 2996 845
rect 2964 715 2996 716
rect 2964 685 2965 715
rect 2965 685 2995 715
rect 2995 685 2996 715
rect 2964 684 2996 685
rect 2964 555 2996 556
rect 2964 525 2965 555
rect 2965 525 2995 555
rect 2995 525 2996 555
rect 2964 524 2996 525
rect 2964 475 2996 476
rect 2964 445 2965 475
rect 2965 445 2995 475
rect 2995 445 2996 475
rect 2964 444 2996 445
rect 2964 395 2996 396
rect 2964 365 2965 395
rect 2965 365 2995 395
rect 2995 365 2996 395
rect 2964 364 2996 365
rect 2964 235 2996 236
rect 2964 205 2965 235
rect 2965 205 2995 235
rect 2995 205 2996 235
rect 2964 204 2996 205
rect 2964 155 2996 156
rect 2964 125 2965 155
rect 2965 125 2995 155
rect 2995 125 2996 155
rect 2964 124 2996 125
rect 2964 75 2996 76
rect 2964 45 2965 75
rect 2965 45 2995 75
rect 2995 45 2996 75
rect 2964 44 2996 45
rect 2964 -5 2996 -4
rect 2964 -35 2965 -5
rect 2965 -35 2995 -5
rect 2995 -35 2996 -5
rect 2964 -36 2996 -35
rect 2964 -165 2996 -164
rect 2964 -195 2965 -165
rect 2965 -195 2995 -165
rect 2995 -195 2996 -165
rect 2964 -196 2996 -195
rect 2964 -325 2996 -324
rect 2964 -355 2965 -325
rect 2965 -355 2995 -325
rect 2995 -355 2996 -325
rect 2964 -356 2996 -355
rect 3124 2155 3156 2156
rect 3124 2125 3125 2155
rect 3125 2125 3155 2155
rect 3155 2125 3156 2155
rect 3124 2124 3156 2125
rect 3124 1995 3156 1996
rect 3124 1965 3125 1995
rect 3125 1965 3155 1995
rect 3155 1965 3156 1995
rect 3124 1964 3156 1965
rect 3124 1835 3156 1836
rect 3124 1805 3125 1835
rect 3125 1805 3155 1835
rect 3155 1805 3156 1835
rect 3124 1804 3156 1805
rect 3124 1755 3156 1756
rect 3124 1725 3125 1755
rect 3125 1725 3155 1755
rect 3155 1725 3156 1755
rect 3124 1724 3156 1725
rect 3124 1675 3156 1676
rect 3124 1645 3125 1675
rect 3125 1645 3155 1675
rect 3155 1645 3156 1675
rect 3124 1644 3156 1645
rect 3124 1595 3156 1596
rect 3124 1565 3125 1595
rect 3125 1565 3155 1595
rect 3155 1565 3156 1595
rect 3124 1564 3156 1565
rect 3124 1435 3156 1436
rect 3124 1405 3125 1435
rect 3125 1405 3155 1435
rect 3155 1405 3156 1435
rect 3124 1404 3156 1405
rect 3124 1355 3156 1356
rect 3124 1325 3125 1355
rect 3125 1325 3155 1355
rect 3155 1325 3156 1355
rect 3124 1324 3156 1325
rect 3124 1275 3156 1276
rect 3124 1245 3125 1275
rect 3125 1245 3155 1275
rect 3155 1245 3156 1275
rect 3124 1244 3156 1245
rect 3124 1115 3156 1116
rect 3124 1085 3125 1115
rect 3125 1085 3155 1115
rect 3155 1085 3156 1115
rect 3124 1084 3156 1085
rect 3124 955 3156 956
rect 3124 925 3125 955
rect 3125 925 3155 955
rect 3155 925 3156 955
rect 3124 924 3156 925
rect 3124 875 3156 876
rect 3124 845 3125 875
rect 3125 845 3155 875
rect 3155 845 3156 875
rect 3124 844 3156 845
rect 3124 715 3156 716
rect 3124 685 3125 715
rect 3125 685 3155 715
rect 3155 685 3156 715
rect 3124 684 3156 685
rect 3124 555 3156 556
rect 3124 525 3125 555
rect 3125 525 3155 555
rect 3155 525 3156 555
rect 3124 524 3156 525
rect 3124 475 3156 476
rect 3124 445 3125 475
rect 3125 445 3155 475
rect 3155 445 3156 475
rect 3124 444 3156 445
rect 3124 395 3156 396
rect 3124 365 3125 395
rect 3125 365 3155 395
rect 3155 365 3156 395
rect 3124 364 3156 365
rect 3124 235 3156 236
rect 3124 205 3125 235
rect 3125 205 3155 235
rect 3155 205 3156 235
rect 3124 204 3156 205
rect 3124 155 3156 156
rect 3124 125 3125 155
rect 3125 125 3155 155
rect 3155 125 3156 155
rect 3124 124 3156 125
rect 3124 75 3156 76
rect 3124 45 3125 75
rect 3125 45 3155 75
rect 3155 45 3156 75
rect 3124 44 3156 45
rect 3124 -5 3156 -4
rect 3124 -35 3125 -5
rect 3125 -35 3155 -5
rect 3155 -35 3156 -5
rect 3124 -36 3156 -35
rect 3124 -165 3156 -164
rect 3124 -195 3125 -165
rect 3125 -195 3155 -165
rect 3155 -195 3156 -165
rect 3124 -196 3156 -195
rect 3124 -325 3156 -324
rect 3124 -355 3125 -325
rect 3125 -355 3155 -325
rect 3155 -355 3156 -325
rect 3124 -356 3156 -355
rect 3284 2155 3316 2156
rect 3284 2125 3285 2155
rect 3285 2125 3315 2155
rect 3315 2125 3316 2155
rect 3284 2124 3316 2125
rect 3284 1995 3316 1996
rect 3284 1965 3285 1995
rect 3285 1965 3315 1995
rect 3315 1965 3316 1995
rect 3284 1964 3316 1965
rect 3284 1835 3316 1836
rect 3284 1805 3285 1835
rect 3285 1805 3315 1835
rect 3315 1805 3316 1835
rect 3284 1804 3316 1805
rect 3284 1755 3316 1756
rect 3284 1725 3285 1755
rect 3285 1725 3315 1755
rect 3315 1725 3316 1755
rect 3284 1724 3316 1725
rect 3284 1675 3316 1676
rect 3284 1645 3285 1675
rect 3285 1645 3315 1675
rect 3315 1645 3316 1675
rect 3284 1644 3316 1645
rect 3284 1595 3316 1596
rect 3284 1565 3285 1595
rect 3285 1565 3315 1595
rect 3315 1565 3316 1595
rect 3284 1564 3316 1565
rect 3284 1435 3316 1436
rect 3284 1405 3285 1435
rect 3285 1405 3315 1435
rect 3315 1405 3316 1435
rect 3284 1404 3316 1405
rect 3284 1355 3316 1356
rect 3284 1325 3285 1355
rect 3285 1325 3315 1355
rect 3315 1325 3316 1355
rect 3284 1324 3316 1325
rect 3284 1275 3316 1276
rect 3284 1245 3285 1275
rect 3285 1245 3315 1275
rect 3315 1245 3316 1275
rect 3284 1244 3316 1245
rect 3284 1115 3316 1116
rect 3284 1085 3285 1115
rect 3285 1085 3315 1115
rect 3315 1085 3316 1115
rect 3284 1084 3316 1085
rect 3284 955 3316 956
rect 3284 925 3285 955
rect 3285 925 3315 955
rect 3315 925 3316 955
rect 3284 924 3316 925
rect 3284 875 3316 876
rect 3284 845 3285 875
rect 3285 845 3315 875
rect 3315 845 3316 875
rect 3284 844 3316 845
rect 3284 715 3316 716
rect 3284 685 3285 715
rect 3285 685 3315 715
rect 3315 685 3316 715
rect 3284 684 3316 685
rect 3284 555 3316 556
rect 3284 525 3285 555
rect 3285 525 3315 555
rect 3315 525 3316 555
rect 3284 524 3316 525
rect 3284 475 3316 476
rect 3284 445 3285 475
rect 3285 445 3315 475
rect 3315 445 3316 475
rect 3284 444 3316 445
rect 3284 395 3316 396
rect 3284 365 3285 395
rect 3285 365 3315 395
rect 3315 365 3316 395
rect 3284 364 3316 365
rect 3284 235 3316 236
rect 3284 205 3285 235
rect 3285 205 3315 235
rect 3315 205 3316 235
rect 3284 204 3316 205
rect 3284 155 3316 156
rect 3284 125 3285 155
rect 3285 125 3315 155
rect 3315 125 3316 155
rect 3284 124 3316 125
rect 3284 75 3316 76
rect 3284 45 3285 75
rect 3285 45 3315 75
rect 3315 45 3316 75
rect 3284 44 3316 45
rect 3284 -5 3316 -4
rect 3284 -35 3285 -5
rect 3285 -35 3315 -5
rect 3315 -35 3316 -5
rect 3284 -36 3316 -35
rect 3284 -165 3316 -164
rect 3284 -195 3285 -165
rect 3285 -195 3315 -165
rect 3315 -195 3316 -165
rect 3284 -196 3316 -195
rect 3284 -325 3316 -324
rect 3284 -355 3285 -325
rect 3285 -355 3315 -325
rect 3315 -355 3316 -325
rect 3284 -356 3316 -355
rect 3444 2155 3476 2156
rect 3444 2125 3445 2155
rect 3445 2125 3475 2155
rect 3475 2125 3476 2155
rect 3444 2124 3476 2125
rect 3444 1995 3476 1996
rect 3444 1965 3445 1995
rect 3445 1965 3475 1995
rect 3475 1965 3476 1995
rect 3444 1964 3476 1965
rect 3444 1835 3476 1836
rect 3444 1805 3445 1835
rect 3445 1805 3475 1835
rect 3475 1805 3476 1835
rect 3444 1804 3476 1805
rect 3444 1675 3476 1676
rect 3444 1645 3445 1675
rect 3445 1645 3475 1675
rect 3475 1645 3476 1675
rect 3444 1644 3476 1645
rect 3444 1595 3476 1596
rect 3444 1565 3445 1595
rect 3445 1565 3475 1595
rect 3475 1565 3476 1595
rect 3444 1564 3476 1565
rect 3444 1435 3476 1436
rect 3444 1405 3445 1435
rect 3445 1405 3475 1435
rect 3475 1405 3476 1435
rect 3444 1404 3476 1405
rect 3444 1275 3476 1276
rect 3444 1245 3445 1275
rect 3445 1245 3475 1275
rect 3475 1245 3476 1275
rect 3444 1244 3476 1245
rect 3444 1115 3476 1116
rect 3444 1085 3445 1115
rect 3445 1085 3475 1115
rect 3475 1085 3476 1115
rect 3444 1084 3476 1085
rect 3444 955 3476 956
rect 3444 925 3445 955
rect 3445 925 3475 955
rect 3475 925 3476 955
rect 3444 924 3476 925
rect 3444 875 3476 876
rect 3444 845 3445 875
rect 3445 845 3475 875
rect 3475 845 3476 875
rect 3444 844 3476 845
rect 3444 715 3476 716
rect 3444 685 3445 715
rect 3445 685 3475 715
rect 3475 685 3476 715
rect 3444 684 3476 685
rect 3444 555 3476 556
rect 3444 525 3445 555
rect 3445 525 3475 555
rect 3475 525 3476 555
rect 3444 524 3476 525
rect 3444 395 3476 396
rect 3444 365 3445 395
rect 3445 365 3475 395
rect 3475 365 3476 395
rect 3444 364 3476 365
rect 3444 235 3476 236
rect 3444 205 3445 235
rect 3445 205 3475 235
rect 3475 205 3476 235
rect 3444 204 3476 205
rect 3444 155 3476 156
rect 3444 125 3445 155
rect 3445 125 3475 155
rect 3475 125 3476 155
rect 3444 124 3476 125
rect 3444 -5 3476 -4
rect 3444 -35 3445 -5
rect 3445 -35 3475 -5
rect 3475 -35 3476 -5
rect 3444 -36 3476 -35
rect 3444 -165 3476 -164
rect 3444 -195 3445 -165
rect 3445 -195 3475 -165
rect 3475 -195 3476 -165
rect 3444 -196 3476 -195
rect 3444 -325 3476 -324
rect 3444 -355 3445 -325
rect 3445 -355 3475 -325
rect 3475 -355 3476 -325
rect 3444 -356 3476 -355
rect 3604 2155 3636 2156
rect 3604 2125 3605 2155
rect 3605 2125 3635 2155
rect 3635 2125 3636 2155
rect 3604 2124 3636 2125
rect 3604 1995 3636 1996
rect 3604 1965 3605 1995
rect 3605 1965 3635 1995
rect 3635 1965 3636 1995
rect 3604 1964 3636 1965
rect 3604 1835 3636 1836
rect 3604 1805 3605 1835
rect 3605 1805 3635 1835
rect 3635 1805 3636 1835
rect 3604 1804 3636 1805
rect 3604 1675 3636 1676
rect 3604 1645 3605 1675
rect 3605 1645 3635 1675
rect 3635 1645 3636 1675
rect 3604 1644 3636 1645
rect 3604 1595 3636 1596
rect 3604 1565 3605 1595
rect 3605 1565 3635 1595
rect 3635 1565 3636 1595
rect 3604 1564 3636 1565
rect 3604 1435 3636 1436
rect 3604 1405 3605 1435
rect 3605 1405 3635 1435
rect 3635 1405 3636 1435
rect 3604 1404 3636 1405
rect 3604 1275 3636 1276
rect 3604 1245 3605 1275
rect 3605 1245 3635 1275
rect 3635 1245 3636 1275
rect 3604 1244 3636 1245
rect 3604 1115 3636 1116
rect 3604 1085 3605 1115
rect 3605 1085 3635 1115
rect 3635 1085 3636 1115
rect 3604 1084 3636 1085
rect 3604 955 3636 956
rect 3604 925 3605 955
rect 3605 925 3635 955
rect 3635 925 3636 955
rect 3604 924 3636 925
rect 3604 875 3636 876
rect 3604 845 3605 875
rect 3605 845 3635 875
rect 3635 845 3636 875
rect 3604 844 3636 845
rect 3604 715 3636 716
rect 3604 685 3605 715
rect 3605 685 3635 715
rect 3635 685 3636 715
rect 3604 684 3636 685
rect 3604 555 3636 556
rect 3604 525 3605 555
rect 3605 525 3635 555
rect 3635 525 3636 555
rect 3604 524 3636 525
rect 3604 395 3636 396
rect 3604 365 3605 395
rect 3605 365 3635 395
rect 3635 365 3636 395
rect 3604 364 3636 365
rect 3604 235 3636 236
rect 3604 205 3605 235
rect 3605 205 3635 235
rect 3635 205 3636 235
rect 3604 204 3636 205
rect 3604 155 3636 156
rect 3604 125 3605 155
rect 3605 125 3635 155
rect 3635 125 3636 155
rect 3604 124 3636 125
rect 3604 -5 3636 -4
rect 3604 -35 3605 -5
rect 3605 -35 3635 -5
rect 3635 -35 3636 -5
rect 3604 -36 3636 -35
rect 3604 -165 3636 -164
rect 3604 -195 3605 -165
rect 3605 -195 3635 -165
rect 3635 -195 3636 -165
rect 3604 -196 3636 -195
rect 3604 -325 3636 -324
rect 3604 -355 3605 -325
rect 3605 -355 3635 -325
rect 3635 -355 3636 -325
rect 3604 -356 3636 -355
rect 3764 2155 3796 2156
rect 3764 2125 3765 2155
rect 3765 2125 3795 2155
rect 3795 2125 3796 2155
rect 3764 2124 3796 2125
rect 3764 1995 3796 1996
rect 3764 1965 3765 1995
rect 3765 1965 3795 1995
rect 3795 1965 3796 1995
rect 3764 1964 3796 1965
rect 3764 1835 3796 1836
rect 3764 1805 3765 1835
rect 3765 1805 3795 1835
rect 3795 1805 3796 1835
rect 3764 1804 3796 1805
rect 3764 1675 3796 1676
rect 3764 1645 3765 1675
rect 3765 1645 3795 1675
rect 3795 1645 3796 1675
rect 3764 1644 3796 1645
rect 3764 1595 3796 1596
rect 3764 1565 3765 1595
rect 3765 1565 3795 1595
rect 3795 1565 3796 1595
rect 3764 1564 3796 1565
rect 3764 1435 3796 1436
rect 3764 1405 3765 1435
rect 3765 1405 3795 1435
rect 3795 1405 3796 1435
rect 3764 1404 3796 1405
rect 3764 1275 3796 1276
rect 3764 1245 3765 1275
rect 3765 1245 3795 1275
rect 3795 1245 3796 1275
rect 3764 1244 3796 1245
rect 3764 1115 3796 1116
rect 3764 1085 3765 1115
rect 3765 1085 3795 1115
rect 3795 1085 3796 1115
rect 3764 1084 3796 1085
rect 3764 955 3796 956
rect 3764 925 3765 955
rect 3765 925 3795 955
rect 3795 925 3796 955
rect 3764 924 3796 925
rect 3764 875 3796 876
rect 3764 845 3765 875
rect 3765 845 3795 875
rect 3795 845 3796 875
rect 3764 844 3796 845
rect 3764 715 3796 716
rect 3764 685 3765 715
rect 3765 685 3795 715
rect 3795 685 3796 715
rect 3764 684 3796 685
rect 3764 555 3796 556
rect 3764 525 3765 555
rect 3765 525 3795 555
rect 3795 525 3796 555
rect 3764 524 3796 525
rect 3764 395 3796 396
rect 3764 365 3765 395
rect 3765 365 3795 395
rect 3795 365 3796 395
rect 3764 364 3796 365
rect 3764 235 3796 236
rect 3764 205 3765 235
rect 3765 205 3795 235
rect 3795 205 3796 235
rect 3764 204 3796 205
rect 3764 155 3796 156
rect 3764 125 3765 155
rect 3765 125 3795 155
rect 3795 125 3796 155
rect 3764 124 3796 125
rect 3764 -5 3796 -4
rect 3764 -35 3765 -5
rect 3765 -35 3795 -5
rect 3795 -35 3796 -5
rect 3764 -36 3796 -35
rect 3764 -165 3796 -164
rect 3764 -195 3765 -165
rect 3765 -195 3795 -165
rect 3795 -195 3796 -165
rect 3764 -196 3796 -195
rect 3764 -325 3796 -324
rect 3764 -355 3765 -325
rect 3765 -355 3795 -325
rect 3795 -355 3796 -325
rect 3764 -356 3796 -355
rect 3924 2155 3956 2156
rect 3924 2125 3925 2155
rect 3925 2125 3955 2155
rect 3955 2125 3956 2155
rect 3924 2124 3956 2125
rect 3924 1995 3956 1996
rect 3924 1965 3925 1995
rect 3925 1965 3955 1995
rect 3955 1965 3956 1995
rect 3924 1964 3956 1965
rect 3924 1835 3956 1836
rect 3924 1805 3925 1835
rect 3925 1805 3955 1835
rect 3955 1805 3956 1835
rect 3924 1804 3956 1805
rect 3924 1675 3956 1676
rect 3924 1645 3925 1675
rect 3925 1645 3955 1675
rect 3955 1645 3956 1675
rect 3924 1644 3956 1645
rect 3924 1595 3956 1596
rect 3924 1565 3925 1595
rect 3925 1565 3955 1595
rect 3955 1565 3956 1595
rect 3924 1564 3956 1565
rect 3924 1435 3956 1436
rect 3924 1405 3925 1435
rect 3925 1405 3955 1435
rect 3955 1405 3956 1435
rect 3924 1404 3956 1405
rect 3924 1275 3956 1276
rect 3924 1245 3925 1275
rect 3925 1245 3955 1275
rect 3955 1245 3956 1275
rect 3924 1244 3956 1245
rect 3924 1115 3956 1116
rect 3924 1085 3925 1115
rect 3925 1085 3955 1115
rect 3955 1085 3956 1115
rect 3924 1084 3956 1085
rect 3924 955 3956 956
rect 3924 925 3925 955
rect 3925 925 3955 955
rect 3955 925 3956 955
rect 3924 924 3956 925
rect 3924 875 3956 876
rect 3924 845 3925 875
rect 3925 845 3955 875
rect 3955 845 3956 875
rect 3924 844 3956 845
rect 6400 880 6440 920
rect 3924 715 3956 716
rect 3924 685 3925 715
rect 3925 685 3955 715
rect 3955 685 3956 715
rect 3924 684 3956 685
rect 3924 555 3956 556
rect 3924 525 3925 555
rect 3925 525 3955 555
rect 3955 525 3956 555
rect 3924 524 3956 525
rect 3924 395 3956 396
rect 3924 365 3925 395
rect 3925 365 3955 395
rect 3955 365 3956 395
rect 3924 364 3956 365
rect 3924 235 3956 236
rect 3924 205 3925 235
rect 3925 205 3955 235
rect 3955 205 3956 235
rect 3924 204 3956 205
rect 3924 155 3956 156
rect 3924 125 3925 155
rect 3925 125 3955 155
rect 3955 125 3956 155
rect 3924 124 3956 125
rect 3924 -5 3956 -4
rect 3924 -35 3925 -5
rect 3925 -35 3955 -5
rect 3955 -35 3956 -5
rect 3924 -36 3956 -35
rect 3924 -165 3956 -164
rect 3924 -195 3925 -165
rect 3925 -195 3955 -165
rect 3955 -195 3956 -165
rect 3924 -196 3956 -195
rect 3924 -325 3956 -324
rect 3924 -355 3925 -325
rect 3925 -355 3955 -325
rect 3955 -355 3956 -325
rect 3924 -356 3956 -355
<< metal4 >>
rect 2320 2156 3960 2160
rect 2320 2124 2324 2156
rect 2356 2124 2484 2156
rect 2516 2124 2644 2156
rect 2676 2124 2804 2156
rect 2836 2124 2964 2156
rect 2996 2124 3124 2156
rect 3156 2124 3284 2156
rect 3316 2124 3444 2156
rect 3476 2124 3604 2156
rect 3636 2124 3764 2156
rect 3796 2124 3924 2156
rect 3956 2124 3960 2156
rect 2320 2120 3960 2124
rect 2320 1996 3960 2000
rect 2320 1964 2324 1996
rect 2356 1964 2484 1996
rect 2516 1964 2644 1996
rect 2676 1964 2804 1996
rect 2836 1964 2964 1996
rect 2996 1964 3124 1996
rect 3156 1964 3284 1996
rect 3316 1964 3444 1996
rect 3476 1964 3604 1996
rect 3636 1964 3764 1996
rect 3796 1964 3924 1996
rect 3956 1964 3960 1996
rect 2320 1960 3960 1964
rect 2320 1836 3960 1840
rect 2320 1804 2324 1836
rect 2356 1804 2484 1836
rect 2516 1804 2644 1836
rect 2676 1804 2804 1836
rect 2836 1804 2964 1836
rect 2996 1804 3124 1836
rect 3156 1804 3284 1836
rect 3316 1804 3444 1836
rect 3476 1804 3604 1836
rect 3636 1804 3764 1836
rect 3796 1804 3924 1836
rect 3956 1804 3960 1836
rect 2320 1800 3960 1804
rect 2960 1756 3320 1760
rect 2960 1724 2964 1756
rect 2996 1724 3124 1756
rect 3156 1724 3284 1756
rect 3316 1724 3320 1756
rect 2960 1720 3320 1724
rect 2320 1676 3960 1680
rect 2320 1644 2324 1676
rect 2356 1644 2484 1676
rect 2516 1644 2644 1676
rect 2676 1644 2804 1676
rect 2836 1644 2964 1676
rect 2996 1644 3124 1676
rect 3156 1644 3284 1676
rect 3316 1644 3444 1676
rect 3476 1644 3604 1676
rect 3636 1644 3764 1676
rect 3796 1644 3924 1676
rect 3956 1644 3960 1676
rect 2320 1640 3960 1644
rect 2320 1596 3960 1600
rect 2320 1564 2324 1596
rect 2356 1564 2484 1596
rect 2516 1564 2644 1596
rect 2676 1564 2804 1596
rect 2836 1564 2964 1596
rect 2996 1564 3124 1596
rect 3156 1564 3284 1596
rect 3316 1564 3444 1596
rect 3476 1564 3604 1596
rect 3636 1564 3764 1596
rect 3796 1564 3924 1596
rect 3956 1564 3960 1596
rect 2320 1560 3960 1564
rect 2320 1436 3960 1440
rect 2320 1404 2324 1436
rect 2356 1404 2484 1436
rect 2516 1404 2644 1436
rect 2676 1404 2804 1436
rect 2836 1404 2964 1436
rect 2996 1404 3124 1436
rect 3156 1404 3284 1436
rect 3316 1404 3444 1436
rect 3476 1404 3604 1436
rect 3636 1404 3764 1436
rect 3796 1404 3924 1436
rect 3956 1404 3960 1436
rect 2320 1400 3960 1404
rect 2960 1356 3320 1360
rect 2960 1324 2964 1356
rect 2996 1324 3124 1356
rect 3156 1324 3284 1356
rect 3316 1324 3320 1356
rect 2960 1320 3320 1324
rect 2320 1276 3960 1280
rect 2320 1244 2324 1276
rect 2356 1244 2484 1276
rect 2516 1244 2644 1276
rect 2676 1244 2804 1276
rect 2836 1244 2964 1276
rect 2996 1244 3124 1276
rect 3156 1244 3284 1276
rect 3316 1244 3444 1276
rect 3476 1244 3604 1276
rect 3636 1244 3764 1276
rect 3796 1244 3924 1276
rect 3956 1244 3960 1276
rect 2320 1240 3960 1244
rect 2320 1116 3960 1120
rect 2320 1084 2324 1116
rect 2356 1084 2484 1116
rect 2516 1084 2644 1116
rect 2676 1084 2804 1116
rect 2836 1084 2964 1116
rect 2996 1084 3124 1116
rect 3156 1084 3284 1116
rect 3316 1084 3444 1116
rect 3476 1084 3604 1116
rect 3636 1084 3764 1116
rect 3796 1084 3924 1116
rect 3956 1084 3960 1116
rect 2320 1080 3960 1084
rect -240 960 -40 1000
rect 6320 960 6520 1000
rect -240 840 -200 960
rect -80 840 -40 960
rect 2320 956 3960 960
rect 2320 924 2324 956
rect 2356 924 2484 956
rect 2516 924 2644 956
rect 2676 924 2804 956
rect 2836 924 2964 956
rect 2996 924 3124 956
rect 3156 924 3284 956
rect 3316 924 3444 956
rect 3476 924 3604 956
rect 3636 924 3764 956
rect 3796 924 3924 956
rect 3956 924 3960 956
rect 2320 920 3960 924
rect 2320 876 3960 880
rect 2320 844 2324 876
rect 2356 844 2484 876
rect 2516 844 2644 876
rect 2676 844 2804 876
rect 2836 844 2964 876
rect 2996 844 3124 876
rect 3156 844 3284 876
rect 3316 844 3444 876
rect 3476 844 3604 876
rect 3636 844 3764 876
rect 3796 844 3924 876
rect 3956 844 3960 876
rect 2320 840 3960 844
rect 6320 840 6360 960
rect 6480 840 6520 960
rect -240 800 -40 840
rect 6320 800 6520 840
rect 2320 716 3960 720
rect 2320 684 2324 716
rect 2356 684 2484 716
rect 2516 684 2644 716
rect 2676 684 2804 716
rect 2836 684 2964 716
rect 2996 684 3124 716
rect 3156 684 3284 716
rect 3316 684 3444 716
rect 3476 684 3604 716
rect 3636 684 3764 716
rect 3796 684 3924 716
rect 3956 684 3960 716
rect 2320 680 3960 684
rect 2320 556 3960 560
rect 2320 524 2324 556
rect 2356 524 2484 556
rect 2516 524 2644 556
rect 2676 524 2804 556
rect 2836 524 2964 556
rect 2996 524 3124 556
rect 3156 524 3284 556
rect 3316 524 3444 556
rect 3476 524 3604 556
rect 3636 524 3764 556
rect 3796 524 3924 556
rect 3956 524 3960 556
rect 2320 520 3960 524
rect 2960 476 3320 480
rect 2960 444 2964 476
rect 2996 444 3124 476
rect 3156 444 3284 476
rect 3316 444 3320 476
rect 2960 440 3320 444
rect 2320 396 3960 400
rect 2320 364 2324 396
rect 2356 364 2484 396
rect 2516 364 2644 396
rect 2676 364 2804 396
rect 2836 364 2964 396
rect 2996 364 3124 396
rect 3156 364 3284 396
rect 3316 364 3444 396
rect 3476 364 3604 396
rect 3636 364 3764 396
rect 3796 364 3924 396
rect 3956 364 3960 396
rect 2320 360 3960 364
rect 2320 236 3960 240
rect 2320 204 2324 236
rect 2356 204 2484 236
rect 2516 204 2644 236
rect 2676 204 2804 236
rect 2836 204 2964 236
rect 2996 204 3124 236
rect 3156 204 3284 236
rect 3316 204 3444 236
rect 3476 204 3604 236
rect 3636 204 3764 236
rect 3796 204 3924 236
rect 3956 204 3960 236
rect 2320 200 3960 204
rect 2320 156 3960 160
rect 2320 124 2324 156
rect 2356 124 2484 156
rect 2516 124 2644 156
rect 2676 124 2804 156
rect 2836 124 2964 156
rect 2996 124 3124 156
rect 3156 124 3284 156
rect 3316 124 3444 156
rect 3476 124 3604 156
rect 3636 124 3764 156
rect 3796 124 3924 156
rect 3956 124 3960 156
rect 2320 120 3960 124
rect 2960 76 3320 80
rect 2960 44 2964 76
rect 2996 44 3124 76
rect 3156 44 3284 76
rect 3316 44 3320 76
rect 2960 40 3320 44
rect 2320 -4 3960 0
rect 2320 -36 2324 -4
rect 2356 -36 2484 -4
rect 2516 -36 2644 -4
rect 2676 -36 2804 -4
rect 2836 -36 2964 -4
rect 2996 -36 3124 -4
rect 3156 -36 3284 -4
rect 3316 -36 3444 -4
rect 3476 -36 3604 -4
rect 3636 -36 3764 -4
rect 3796 -36 3924 -4
rect 3956 -36 3960 -4
rect 2320 -40 3960 -36
rect 2320 -164 3960 -160
rect 2320 -196 2324 -164
rect 2356 -196 2484 -164
rect 2516 -196 2644 -164
rect 2676 -196 2804 -164
rect 2836 -196 2964 -164
rect 2996 -196 3124 -164
rect 3156 -196 3284 -164
rect 3316 -196 3444 -164
rect 3476 -196 3604 -164
rect 3636 -196 3764 -164
rect 3796 -196 3924 -164
rect 3956 -196 3960 -164
rect 2320 -200 3960 -196
rect 2320 -324 3960 -320
rect 2320 -356 2324 -324
rect 2356 -356 2484 -324
rect 2516 -356 2644 -324
rect 2676 -356 2804 -324
rect 2836 -356 2964 -324
rect 2996 -356 3124 -324
rect 3156 -356 3284 -324
rect 3316 -356 3444 -324
rect 3476 -356 3604 -324
rect 3636 -356 3764 -324
rect 3796 -356 3924 -324
rect 3956 -356 3960 -324
rect 2320 -360 3960 -356
<< via4 >>
rect -200 920 -80 960
rect -200 880 -160 920
rect -160 880 -120 920
rect -120 880 -80 920
rect -200 840 -80 880
rect 6360 920 6480 960
rect 6360 880 6400 920
rect 6400 880 6440 920
rect 6440 880 6480 920
rect 6360 840 6480 880
<< metal5 >>
rect -240 960 -40 2160
rect -240 840 -200 960
rect -80 840 -40 960
rect -240 -360 -40 840
rect 6320 960 6520 2160
rect 6320 840 6360 960
rect 6480 840 6520 960
rect 6320 -360 6520 840
<< labels >>
rlabel metal3 2400 -360 2440 2160 0 xp
port 1 nsew
rlabel metal3 2560 -360 2600 2160 0 om
port 2 nsew
rlabel metal3 2720 -360 2760 2160 0 xm
port 3 nsew
rlabel metal3 2880 -360 2920 2160 0 op
port 4 nsew
rlabel metal3 3040 -360 3080 2160 0 fsb
port 5 nsew
rlabel metal3 3200 -360 3240 2160 0 q
port 6 nsew
rlabel metal3 2320 -320 2360 -280 0 gnda
port 7 nsew
rlabel metal5 -240 -360 -40 -320 0 vssa
port 8 nsew
<< end >>
