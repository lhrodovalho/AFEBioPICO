**.subckt pseudo_tb
XM1 X X B B sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 X X A A sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
VA A GND 0
VB B GND 0
**** begin user architecture code


.include ~/git/open_pdks/sources/sky130-pdk/libraries/sky130_fd_pr/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include ~/git/open_pdks/sources/sky130-pdk/libraries/sky130_fd_pr/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/git/open_pdks/sources/sky130-pdk/libraries/sky130_fd_pr/latest/models/all.spice

* All models
*.include /usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice




.options gmin=1e-13
.options rshunt = 1.0e13

.control
  dc VA -0.9 0.9 0.011
  let r=abs(deriv(v(a))/deriv(i(va)))
  plot r ylog
.endc


**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
