**.subckt iref_tb
VDD vdd GND 1.8
VSS vss GND 0.0
x1 vdd io vss iref
VO io GND 0.0
**** begin user architecture code



.include /usr/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_g5v0d10v5__ss.corner.spice
.include /usr/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include /usr/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include /usr/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice

.include /usr/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include /usr/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include /usr/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include /usr/share/pdk/sky130A/libs.ref/spi/sky130_fd_pr/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice

.include /usr/share/pdk/sky130A/libs.tech/ngspice/all.spice





.param mc_mm_switch=0

.options gmin=1e-12
.options reltol=1e-5
.options abstol=1e-15
*.options rshunt = 1.0e15

.control
  op
  print i(VO)

  dc VDD 0.3 1.8 1m

  let io = i(VO)
  wrdata ../../SIM_DATA/iref_io.txt io
  plot io

  let psrr = deriv(io)/io
  wrdata ../../SIM_DATA/iref_psrr.txt io
  plot ylog abs(psrr)

.endc


**** end user architecture code
**.ends

* expanding   symbol:  iref.sym # of pins=3
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/IREF/iref.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/IREF/iref.sch
.subckt iref  vdd io vss
*.iopin vdd
*.iopin vss
*.iopin io
x12 net4 p1 vdd vdd p1_2
x25 net11 net12 vss vss n1_2
x31 net14 lo vdd vdd p2_1
x32 vdd lo net14 vdd p2_1
x7 x p2 net2 vdd p2_1
x8 net2 p1 vdd vdd p2_1
x9 net3 p1 vdd vdd p1_2
x10 net8 p0 vdd vdd p1_2
x11 net6 p2 vdd vdd p1_2
x15 net13 p1 vdd vdd p1_2
x16 net10 p0 vdd vdd p1_2
x19 n1 p2 net4 vdd p1_2
x20 y p2 net3 vdd p1_2
x23 p0 p2 net8 vdd p1_2
x24 p2 p2 net6 vdd p1_2
x27 io p2 net13 vdd p1_2
x33 p1 p2 net10 vdd p1_2
x1 net12 net12 net11 vss n1_2
x2 net9 n1 vss vss n1_2
x3 p1 n1 net9 vss n1_2
x4 net7 y vss vss n1_2
x5 p0 y net7 vss n1_2
x6 net5 n1 vss vss n2_1
x13 p2 n1 net5 vss n2_1
x14 net1 n1 vss vss n1_2
x17 n1 n1 net1 vss n1_2
x18 z x vss vss n1_2
x21 y y z vss n1_2
x22 z x vss vss n1_2
x26 x x z vss n1_2
x29 lo n1 vss vss n1_2
x30 p1 lo n1 vss n1_2
.ends


* expanding   symbol:  ../ARRAY/p1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_2.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_2.sch
.subckt p1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_1
xd D G X B p1_1
.ends


* expanding   symbol:  ../ARRAY/n1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_2.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_2.sch
.subckt n1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_1
xs X G S B n1_1
.ends


* expanding   symbol:  ../ARRAY/p2_1.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p2_1.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p2_1.sch
.subckt p2_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xl D G S B p1_1
xr D G S B p1_1
.ends


* expanding   symbol:  ../ARRAY/n2_1.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n2_1.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n2_1.sch
.subckt n2_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xr D G S B n1_1
xl D G S B n1_1
.ends


* expanding   symbol:  p1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_1.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_1.sch
.subckt p1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8_lvt L=8 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
.ends


* expanding   symbol:  n1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_1.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_1.sch
.subckt n1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8_lvt L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
.ends

.GLOBAL GND
** flattened .save nodes
.end
