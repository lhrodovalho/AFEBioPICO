.subckt load ip im ib vdda gnda vssa
xpa1 ib ib vdda vdda vssa p1_8

xpd1 ip ib vdda vdda vssa p1_8
xnd3 ip n  vssa vssa n1_8

xpe1 im  ib vdda vdda vssa p1_8
xne3 im n  vssa vssa n1_8

xpf1 y  ib   vdda vdda vssa p1_8
xpf2 n  gnda y    vdda vssa p1_8
xnf3 n  n    vssa vssa n1_8

xpg1 y  ib   vdda vdda vssa p1_8
xpg2 n  gnda y    vdda vssa p1_8
xng3 n  n    vssa vssa n1_8

xph1 y  ib   vdda vdda vssa p1_8
xph2 z  ip   y    vdda vssa p1_8
xnh3 z  z    vssa vssa n1_8

xpi1 y  ib   vdda vdda vssa p1_8
xpi2 z  im   y    vdda vssa p1_8
xni3 z  z    vssa vssa n1_8

.ends

.subckt load2 ip im ib vdda gnda vssa
xpa1 ib ib vdda vdda vssa p8_1

xpb1 x  ib vdda vdda vssa p1_8
xpb2 y  ip x    vdda vssa p1_8
xnb3 y  n  vssa vssa      n1_8

xpc1 x  ib vdda vdda vssa p1_8
xpc2 y  im x    vdda vssa p1_8
xnc3 y  n  vssa vssa      n1_8

xpd1 x  ib vdda vdda vssa p1_8
xpd2 y  y  x    vdda vssa p1_8
xnd3 y  n  vssa vssa	  n1_8

xpe1 x  ib vdda vdda vssa p1_8
xpe2 y  y  x    vdda vssa p1_8
xne3 y  n  vssa vssa	  n1_8

xpf1 x  ib vdda vdda vssa p1_8
xpf2 z  y  x    vdda vssa p1_8
xnf3 z  n  vssa vssa	  n1_8

xpg1 x  ib vdda vdda vssa p1_8
xpg2 z  z  x    vdda vssa p1_8
xng3 z  n  vssa vssa	  n1_8

xph1 x  ib vdda vdda vssa p1_8
xph2 im z  x    vdda vssa p1_8
xnh3 im n  vssa vssa	  n1_8

xpi1 x  ib vdda vdda vssa p1_8
xpi2 ip z  x    vdda vssa p1_8
xni3 ip n  vssa vssa	  n1_8

xpj1 x ib   vdda vdda vssa p1_8
xpj2 n gnda x    vdda vssa p1_8
xnj3 n n    vssa vssa	  n1_8

.ends

.subckt load3 ip im ib vdda gnda vssa
xpa1 ib ib vdda vdda vssa p8_1

xpb1 x  ib vdda vdda vssa p1_8
xpb2 im ip x    vdda vssa p1_8
xnb3 im n  vssa vssa      n1_8

xpc1 x  ib vdda vdda vssa p1_8
xpc2 ip im x    vdda vssa p1_8
xnc3 ip n  vssa vssa      n1_8

xpd1 x  ib vdda vdda vssa p1_8
xpd2 ip ip x    vdda vssa p1_8
xnd3 ip n  vssa vssa      n1_8

xpe1 x  ib vdda vdda vssa p1_8
xpe2 im im x    vdda vssa p1_8
xne3 im n  vssa vssa      n1_8

xpj1 x ib   vdda vdda vssa p1_8
xpj2 n gnda x    vdda vssa p1_8
xnj3 n n    vssa vssa	   n1_8

.ends
