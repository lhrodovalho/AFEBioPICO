magic
tech sky130A
timestamp 1637779139
<< nwell >>
rect -180 -500 5180 460
<< mvnmos >>
rect 0 -1240 200 -1140
rect 320 -1240 520 -1140
rect 640 -1240 840 -1140
rect 960 -1240 1160 -1140
rect 1280 -1240 1480 -1140
rect 1600 -1240 1800 -1140
rect 1920 -1240 2120 -1140
rect 2240 -1240 2440 -1140
rect 2560 -1240 2760 -1140
rect 2880 -1240 3080 -1140
rect 3200 -1240 3400 -1140
rect 3520 -1240 3720 -1140
rect 3840 -1240 4040 -1140
rect 4160 -1240 4360 -1140
rect 4480 -1240 4680 -1140
rect 4800 -1240 5000 -1140
rect 0 -1440 200 -1340
rect 320 -1440 520 -1340
rect 640 -1440 840 -1340
rect 960 -1440 1160 -1340
rect 1280 -1440 1480 -1340
rect 1600 -1440 1800 -1340
rect 1920 -1440 2120 -1340
rect 2240 -1440 2440 -1340
rect 2560 -1440 2760 -1340
rect 2880 -1440 3080 -1340
rect 3200 -1440 3400 -1340
rect 3520 -1440 3720 -1340
rect 3840 -1440 4040 -1340
rect 4160 -1440 4360 -1340
rect 4480 -1440 4680 -1340
rect 4800 -1440 5000 -1340
<< mvpmos >>
rect 0 60 200 360
rect 320 60 520 360
rect 640 60 840 360
rect 960 60 1160 360
rect 1280 60 1480 360
rect 1600 60 1800 360
rect 1920 60 2120 360
rect 2240 60 2440 360
rect 2560 60 2760 360
rect 2880 60 3080 360
rect 3200 60 3400 360
rect 3520 60 3720 360
rect 3840 60 4040 360
rect 4160 60 4360 360
rect 4480 60 4680 360
rect 4800 60 5000 360
rect 0 -340 200 -40
rect 320 -340 520 -40
rect 640 -340 840 -40
rect 960 -340 1160 -40
rect 1280 -340 1480 -40
rect 1600 -340 1800 -40
rect 1920 -340 2120 -40
rect 2240 -340 2440 -40
rect 2560 -340 2760 -40
rect 2880 -340 3080 -40
rect 3200 -340 3400 -40
rect 3520 -340 3720 -40
rect 3840 -340 4040 -40
rect 4160 -340 4360 -40
rect 4480 -340 4680 -40
rect 4800 -340 5000 -40
<< mvndiff >>
rect -80 -1150 0 -1140
rect -80 -1230 -75 -1150
rect -45 -1230 0 -1150
rect -80 -1240 0 -1230
rect 200 -1150 320 -1140
rect 200 -1230 245 -1150
rect 275 -1230 320 -1150
rect 200 -1240 320 -1230
rect 520 -1150 640 -1140
rect 520 -1230 565 -1150
rect 595 -1230 640 -1150
rect 520 -1240 640 -1230
rect 840 -1150 960 -1140
rect 840 -1230 885 -1150
rect 915 -1230 960 -1150
rect 840 -1240 960 -1230
rect 1160 -1150 1280 -1140
rect 1160 -1230 1205 -1150
rect 1235 -1230 1280 -1150
rect 1160 -1240 1280 -1230
rect 1480 -1150 1600 -1140
rect 1480 -1230 1525 -1150
rect 1555 -1230 1600 -1150
rect 1480 -1240 1600 -1230
rect 1800 -1150 1920 -1140
rect 1800 -1230 1845 -1150
rect 1875 -1230 1920 -1150
rect 1800 -1240 1920 -1230
rect 2120 -1150 2240 -1140
rect 2120 -1230 2165 -1150
rect 2195 -1230 2240 -1150
rect 2120 -1240 2240 -1230
rect 2440 -1150 2560 -1140
rect 2440 -1230 2485 -1150
rect 2515 -1230 2560 -1150
rect 2440 -1240 2560 -1230
rect 2760 -1150 2880 -1140
rect 2760 -1230 2805 -1150
rect 2835 -1230 2880 -1150
rect 2760 -1240 2880 -1230
rect 3080 -1150 3200 -1140
rect 3080 -1230 3125 -1150
rect 3155 -1230 3200 -1150
rect 3080 -1240 3200 -1230
rect 3400 -1150 3520 -1140
rect 3400 -1230 3445 -1150
rect 3475 -1230 3520 -1150
rect 3400 -1240 3520 -1230
rect 3720 -1150 3840 -1140
rect 3720 -1230 3765 -1150
rect 3795 -1230 3840 -1150
rect 3720 -1240 3840 -1230
rect 4040 -1150 4160 -1140
rect 4040 -1230 4085 -1150
rect 4115 -1230 4160 -1150
rect 4040 -1240 4160 -1230
rect 4360 -1150 4480 -1140
rect 4360 -1230 4405 -1150
rect 4435 -1230 4480 -1150
rect 4360 -1240 4480 -1230
rect 4680 -1150 4800 -1140
rect 4680 -1230 4725 -1150
rect 4755 -1230 4800 -1150
rect 4680 -1240 4800 -1230
rect 5000 -1150 5080 -1140
rect 5000 -1230 5045 -1150
rect 5075 -1230 5080 -1150
rect 5000 -1240 5080 -1230
rect -80 -1350 0 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 0 -1350
rect -80 -1440 0 -1430
rect 200 -1350 320 -1340
rect 200 -1430 245 -1350
rect 275 -1430 320 -1350
rect 200 -1440 320 -1430
rect 520 -1350 640 -1340
rect 520 -1430 565 -1350
rect 595 -1430 640 -1350
rect 520 -1440 640 -1430
rect 840 -1350 960 -1340
rect 840 -1430 885 -1350
rect 915 -1430 960 -1350
rect 840 -1440 960 -1430
rect 1160 -1350 1280 -1340
rect 1160 -1430 1205 -1350
rect 1235 -1430 1280 -1350
rect 1160 -1440 1280 -1430
rect 1480 -1350 1600 -1340
rect 1480 -1430 1525 -1350
rect 1555 -1430 1600 -1350
rect 1480 -1440 1600 -1430
rect 1800 -1350 1920 -1340
rect 1800 -1430 1845 -1350
rect 1875 -1430 1920 -1350
rect 1800 -1440 1920 -1430
rect 2120 -1350 2240 -1340
rect 2120 -1430 2165 -1350
rect 2195 -1430 2240 -1350
rect 2120 -1440 2240 -1430
rect 2440 -1350 2560 -1340
rect 2440 -1430 2485 -1350
rect 2515 -1430 2560 -1350
rect 2440 -1440 2560 -1430
rect 2760 -1350 2880 -1340
rect 2760 -1430 2805 -1350
rect 2835 -1430 2880 -1350
rect 2760 -1440 2880 -1430
rect 3080 -1350 3200 -1340
rect 3080 -1430 3125 -1350
rect 3155 -1430 3200 -1350
rect 3080 -1440 3200 -1430
rect 3400 -1350 3520 -1340
rect 3400 -1430 3445 -1350
rect 3475 -1430 3520 -1350
rect 3400 -1440 3520 -1430
rect 3720 -1350 3840 -1340
rect 3720 -1430 3765 -1350
rect 3795 -1430 3840 -1350
rect 3720 -1440 3840 -1430
rect 4040 -1350 4160 -1340
rect 4040 -1430 4085 -1350
rect 4115 -1430 4160 -1350
rect 4040 -1440 4160 -1430
rect 4360 -1350 4480 -1340
rect 4360 -1430 4405 -1350
rect 4435 -1430 4480 -1350
rect 4360 -1440 4480 -1430
rect 4680 -1350 4800 -1340
rect 4680 -1430 4725 -1350
rect 4755 -1430 4800 -1350
rect 4680 -1440 4800 -1430
rect 5000 -1350 5080 -1340
rect 5000 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5000 -1440 5080 -1430
<< mvpdiff >>
rect -80 350 0 360
rect -80 70 -75 350
rect -45 70 0 350
rect -80 60 0 70
rect 200 350 320 360
rect 200 70 245 350
rect 275 70 320 350
rect 200 60 320 70
rect 520 350 640 360
rect 520 70 565 350
rect 595 70 640 350
rect 520 60 640 70
rect 840 350 960 360
rect 840 70 885 350
rect 915 70 960 350
rect 840 60 960 70
rect 1160 350 1280 360
rect 1160 70 1205 350
rect 1235 70 1280 350
rect 1160 60 1280 70
rect 1480 350 1600 360
rect 1480 70 1525 350
rect 1555 70 1600 350
rect 1480 60 1600 70
rect 1800 350 1920 360
rect 1800 70 1845 350
rect 1875 70 1920 350
rect 1800 60 1920 70
rect 2120 350 2240 360
rect 2120 70 2165 350
rect 2195 70 2240 350
rect 2120 60 2240 70
rect 2440 350 2560 360
rect 2440 70 2485 350
rect 2515 70 2560 350
rect 2440 60 2560 70
rect 2760 350 2880 360
rect 2760 70 2805 350
rect 2835 70 2880 350
rect 2760 60 2880 70
rect 3080 350 3200 360
rect 3080 70 3125 350
rect 3155 70 3200 350
rect 3080 60 3200 70
rect 3400 350 3520 360
rect 3400 70 3445 350
rect 3475 70 3520 350
rect 3400 60 3520 70
rect 3720 350 3840 360
rect 3720 70 3765 350
rect 3795 70 3840 350
rect 3720 60 3840 70
rect 4040 350 4160 360
rect 4040 70 4085 350
rect 4115 70 4160 350
rect 4040 60 4160 70
rect 4360 350 4480 360
rect 4360 70 4405 350
rect 4435 70 4480 350
rect 4360 60 4480 70
rect 4680 350 4800 360
rect 4680 70 4725 350
rect 4755 70 4800 350
rect 4680 60 4800 70
rect 5000 350 5080 360
rect 5000 70 5045 350
rect 5075 70 5080 350
rect 5000 60 5080 70
rect -80 -50 0 -40
rect -80 -330 -75 -50
rect -45 -330 0 -50
rect -80 -340 0 -330
rect 200 -50 320 -40
rect 200 -330 245 -50
rect 275 -330 320 -50
rect 200 -340 320 -330
rect 520 -50 640 -40
rect 520 -330 565 -50
rect 595 -330 640 -50
rect 520 -340 640 -330
rect 840 -50 960 -40
rect 840 -330 885 -50
rect 915 -330 960 -50
rect 840 -340 960 -330
rect 1160 -50 1280 -40
rect 1160 -330 1205 -50
rect 1235 -330 1280 -50
rect 1160 -340 1280 -330
rect 1480 -50 1600 -40
rect 1480 -330 1525 -50
rect 1555 -330 1600 -50
rect 1480 -340 1600 -330
rect 1800 -50 1920 -40
rect 1800 -330 1845 -50
rect 1875 -330 1920 -50
rect 1800 -340 1920 -330
rect 2120 -50 2240 -40
rect 2120 -330 2165 -50
rect 2195 -330 2240 -50
rect 2120 -340 2240 -330
rect 2440 -50 2560 -40
rect 2440 -330 2485 -50
rect 2515 -330 2560 -50
rect 2440 -340 2560 -330
rect 2760 -50 2880 -40
rect 2760 -330 2805 -50
rect 2835 -330 2880 -50
rect 2760 -340 2880 -330
rect 3080 -50 3200 -40
rect 3080 -330 3125 -50
rect 3155 -330 3200 -50
rect 3080 -340 3200 -330
rect 3400 -50 3520 -40
rect 3400 -330 3445 -50
rect 3475 -330 3520 -50
rect 3400 -340 3520 -330
rect 3720 -50 3840 -40
rect 3720 -330 3765 -50
rect 3795 -330 3840 -50
rect 3720 -340 3840 -330
rect 4040 -50 4160 -40
rect 4040 -330 4085 -50
rect 4115 -330 4160 -50
rect 4040 -340 4160 -330
rect 4360 -50 4480 -40
rect 4360 -330 4405 -50
rect 4435 -330 4480 -50
rect 4360 -340 4480 -330
rect 4680 -50 4800 -40
rect 4680 -330 4725 -50
rect 4755 -330 4800 -50
rect 4680 -340 4800 -330
rect 5000 -50 5080 -40
rect 5000 -330 5045 -50
rect 5075 -330 5080 -50
rect 5000 -340 5080 -330
<< mvndiffc >>
rect -75 -1230 -45 -1150
rect 245 -1230 275 -1150
rect 565 -1230 595 -1150
rect 885 -1230 915 -1150
rect 1205 -1230 1235 -1150
rect 1525 -1230 1555 -1150
rect 1845 -1230 1875 -1150
rect 2165 -1230 2195 -1150
rect 2485 -1230 2515 -1150
rect 2805 -1230 2835 -1150
rect 3125 -1230 3155 -1150
rect 3445 -1230 3475 -1150
rect 3765 -1230 3795 -1150
rect 4085 -1230 4115 -1150
rect 4405 -1230 4435 -1150
rect 4725 -1230 4755 -1150
rect 5045 -1230 5075 -1150
rect -75 -1430 -45 -1350
rect 245 -1430 275 -1350
rect 565 -1430 595 -1350
rect 885 -1430 915 -1350
rect 1205 -1430 1235 -1350
rect 1525 -1430 1555 -1350
rect 1845 -1430 1875 -1350
rect 2165 -1430 2195 -1350
rect 2485 -1430 2515 -1350
rect 2805 -1430 2835 -1350
rect 3125 -1430 3155 -1350
rect 3445 -1430 3475 -1350
rect 3765 -1430 3795 -1350
rect 4085 -1430 4115 -1350
rect 4405 -1430 4435 -1350
rect 4725 -1430 4755 -1350
rect 5045 -1430 5075 -1350
<< mvpdiffc >>
rect -75 70 -45 350
rect 245 70 275 350
rect 565 70 595 350
rect 885 70 915 350
rect 1205 70 1235 350
rect 1525 70 1555 350
rect 1845 70 1875 350
rect 2165 70 2195 350
rect 2485 70 2515 350
rect 2805 70 2835 350
rect 3125 70 3155 350
rect 3445 70 3475 350
rect 3765 70 3795 350
rect 4085 70 4115 350
rect 4405 70 4435 350
rect 4725 70 4755 350
rect 5045 70 5075 350
rect -75 -330 -45 -50
rect 245 -330 275 -50
rect 565 -330 595 -50
rect 885 -330 915 -50
rect 1205 -330 1235 -50
rect 1525 -330 1555 -50
rect 1845 -330 1875 -50
rect 2165 -330 2195 -50
rect 2485 -330 2515 -50
rect 2805 -330 2835 -50
rect 3125 -330 3155 -50
rect 3445 -330 3475 -50
rect 3765 -330 3795 -50
rect 4085 -330 4115 -50
rect 4405 -330 4435 -50
rect 4725 -330 4755 -50
rect 5045 -330 5075 -50
<< psubdiff >>
rect -240 480 -180 520
rect 5180 480 5240 520
rect -240 460 -200 480
rect 5200 460 5240 480
rect -200 -1040 -180 -1000
rect 5180 -1040 5200 -1000
rect -240 -1480 -200 -1460
rect 5200 -1480 5240 -1460
rect -240 -1520 -180 -1480
rect 5180 -1520 5240 -1480
<< nsubdiff >>
rect -160 400 -100 440
rect 5100 400 5160 440
rect -160 380 -120 400
rect 5120 380 5160 400
rect -160 -440 -120 -420
rect 5120 -440 5160 -420
rect -160 -480 -100 -440
rect 5100 -480 5160 -440
<< psubdiffcont >>
rect -180 480 5180 520
rect -240 -1460 -200 460
rect -180 -1040 5180 -1000
rect 5200 -1460 5240 460
rect -180 -1520 5180 -1480
<< nsubdiffcont >>
rect -100 400 5100 440
rect -160 -420 -120 380
rect 5120 -420 5160 380
rect -100 -480 5100 -440
<< poly >>
rect 0 360 200 380
rect 320 360 520 380
rect 640 360 840 380
rect 960 360 1160 380
rect 1280 360 1480 380
rect 1600 360 1800 380
rect 1920 360 2120 380
rect 2240 360 2440 380
rect 2560 360 2760 380
rect 2880 360 3080 380
rect 3200 360 3400 380
rect 3520 360 3720 380
rect 3840 360 4040 380
rect 4160 360 4360 380
rect 4480 360 4680 380
rect 4800 360 5000 380
rect 0 -40 200 60
rect 320 -40 520 60
rect 640 -40 840 60
rect 960 -40 1160 60
rect 1280 -40 1480 60
rect 1600 -40 1800 60
rect 1920 -40 2120 60
rect 2240 -40 2440 60
rect 2560 -40 2760 60
rect 2880 -40 3080 60
rect 3200 -40 3400 60
rect 3520 -40 3720 60
rect 3840 -40 4040 60
rect 4160 -40 4360 60
rect 4480 -40 4680 60
rect 4800 -40 5000 60
rect 0 -365 200 -340
rect 0 -395 10 -365
rect 190 -395 200 -365
rect 0 -400 200 -395
rect 320 -365 520 -340
rect 320 -395 330 -365
rect 510 -395 520 -365
rect 320 -400 520 -395
rect 640 -365 840 -340
rect 640 -395 650 -365
rect 830 -395 840 -365
rect 640 -400 840 -395
rect 960 -365 1160 -340
rect 960 -395 970 -365
rect 1150 -395 1160 -365
rect 960 -400 1160 -395
rect 1280 -365 1480 -340
rect 1280 -395 1290 -365
rect 1470 -395 1480 -365
rect 1280 -400 1480 -395
rect 1600 -365 1800 -340
rect 1600 -395 1610 -365
rect 1790 -395 1800 -365
rect 1600 -400 1800 -395
rect 1920 -365 2120 -340
rect 1920 -395 1930 -365
rect 2110 -395 2120 -365
rect 1920 -400 2120 -395
rect 2240 -365 2440 -340
rect 2240 -395 2250 -365
rect 2430 -395 2440 -365
rect 2240 -400 2440 -395
rect 2560 -365 2760 -340
rect 2560 -395 2570 -365
rect 2750 -395 2760 -365
rect 2560 -400 2760 -395
rect 2880 -365 3080 -340
rect 2880 -395 2890 -365
rect 3070 -395 3080 -365
rect 2880 -400 3080 -395
rect 3200 -365 3400 -340
rect 3200 -395 3210 -365
rect 3390 -395 3400 -365
rect 3200 -400 3400 -395
rect 3520 -365 3720 -340
rect 3520 -395 3530 -365
rect 3710 -395 3720 -365
rect 3520 -400 3720 -395
rect 3840 -365 4040 -340
rect 3840 -395 3850 -365
rect 4030 -395 4040 -365
rect 3840 -400 4040 -395
rect 4160 -365 4360 -340
rect 4160 -395 4170 -365
rect 4350 -395 4360 -365
rect 4160 -400 4360 -395
rect 4480 -365 4680 -340
rect 4480 -395 4490 -365
rect 4670 -395 4680 -365
rect 4480 -400 4680 -395
rect 4800 -365 5000 -340
rect 4800 -395 4810 -365
rect 4990 -395 5000 -365
rect 4800 -400 5000 -395
rect 0 -1085 200 -1080
rect 0 -1115 10 -1085
rect 190 -1115 200 -1085
rect 0 -1140 200 -1115
rect 320 -1085 520 -1080
rect 320 -1115 330 -1085
rect 510 -1115 520 -1085
rect 320 -1140 520 -1115
rect 640 -1085 840 -1080
rect 640 -1115 650 -1085
rect 830 -1115 840 -1085
rect 640 -1140 840 -1115
rect 960 -1085 1160 -1080
rect 960 -1115 970 -1085
rect 1150 -1115 1160 -1085
rect 960 -1140 1160 -1115
rect 1280 -1085 1480 -1080
rect 1280 -1115 1290 -1085
rect 1470 -1115 1480 -1085
rect 1280 -1140 1480 -1115
rect 1600 -1085 1800 -1080
rect 1600 -1115 1610 -1085
rect 1790 -1115 1800 -1085
rect 1600 -1140 1800 -1115
rect 1920 -1085 2120 -1080
rect 1920 -1115 1930 -1085
rect 2110 -1115 2120 -1085
rect 1920 -1140 2120 -1115
rect 2240 -1085 2440 -1080
rect 2240 -1115 2250 -1085
rect 2430 -1115 2440 -1085
rect 2240 -1140 2440 -1115
rect 2560 -1085 2760 -1080
rect 2560 -1115 2570 -1085
rect 2750 -1115 2760 -1085
rect 2560 -1140 2760 -1115
rect 2880 -1085 3080 -1080
rect 2880 -1115 2890 -1085
rect 3070 -1115 3080 -1085
rect 2880 -1140 3080 -1115
rect 3200 -1085 3400 -1080
rect 3200 -1115 3210 -1085
rect 3390 -1115 3400 -1085
rect 3200 -1140 3400 -1115
rect 3520 -1085 3720 -1080
rect 3520 -1115 3530 -1085
rect 3710 -1115 3720 -1085
rect 3520 -1140 3720 -1115
rect 3840 -1085 4040 -1080
rect 3840 -1115 3850 -1085
rect 4030 -1115 4040 -1085
rect 3840 -1140 4040 -1115
rect 4160 -1085 4360 -1080
rect 4160 -1115 4170 -1085
rect 4350 -1115 4360 -1085
rect 4160 -1140 4360 -1115
rect 4480 -1085 4680 -1080
rect 4480 -1115 4490 -1085
rect 4670 -1115 4680 -1085
rect 4480 -1140 4680 -1115
rect 4800 -1085 5000 -1080
rect 4800 -1115 4810 -1085
rect 4990 -1115 5000 -1085
rect 4800 -1140 5000 -1115
rect 0 -1340 200 -1240
rect 320 -1340 520 -1240
rect 640 -1340 840 -1240
rect 960 -1340 1160 -1240
rect 1280 -1340 1480 -1240
rect 1600 -1340 1800 -1240
rect 1920 -1340 2120 -1240
rect 2240 -1340 2440 -1240
rect 2560 -1340 2760 -1240
rect 2880 -1340 3080 -1240
rect 3200 -1340 3400 -1240
rect 3520 -1340 3720 -1240
rect 3840 -1340 4040 -1240
rect 4160 -1340 4360 -1240
rect 4480 -1340 4680 -1240
rect 4800 -1340 5000 -1240
rect 0 -1460 200 -1440
rect 320 -1460 520 -1440
rect 640 -1460 840 -1440
rect 960 -1460 1160 -1440
rect 1280 -1460 1480 -1440
rect 1600 -1460 1800 -1440
rect 1920 -1460 2120 -1440
rect 2240 -1460 2440 -1440
rect 2560 -1460 2760 -1440
rect 2880 -1460 3080 -1440
rect 3200 -1460 3400 -1440
rect 3520 -1460 3720 -1440
rect 3840 -1460 4040 -1440
rect 4160 -1460 4360 -1440
rect 4480 -1460 4680 -1440
rect 4800 -1460 5000 -1440
<< polycont >>
rect 10 -395 190 -365
rect 330 -395 510 -365
rect 650 -395 830 -365
rect 970 -395 1150 -365
rect 1290 -395 1470 -365
rect 1610 -395 1790 -365
rect 1930 -395 2110 -365
rect 2250 -395 2430 -365
rect 2570 -395 2750 -365
rect 2890 -395 3070 -365
rect 3210 -395 3390 -365
rect 3530 -395 3710 -365
rect 3850 -395 4030 -365
rect 4170 -395 4350 -365
rect 4490 -395 4670 -365
rect 4810 -395 4990 -365
rect 10 -1115 190 -1085
rect 330 -1115 510 -1085
rect 650 -1115 830 -1085
rect 970 -1115 1150 -1085
rect 1290 -1115 1470 -1085
rect 1610 -1115 1790 -1085
rect 1930 -1115 2110 -1085
rect 2250 -1115 2430 -1085
rect 2570 -1115 2750 -1085
rect 2890 -1115 3070 -1085
rect 3210 -1115 3390 -1085
rect 3530 -1115 3710 -1085
rect 3850 -1115 4030 -1085
rect 4170 -1115 4350 -1085
rect 4490 -1115 4670 -1085
rect 4810 -1115 4990 -1085
<< locali >>
rect -240 480 -180 520
rect 5180 480 5240 520
rect -240 460 -200 480
rect 5200 460 5240 480
rect -160 400 -100 440
rect 5100 400 5160 440
rect -160 380 -120 400
rect -80 350 -40 400
rect -80 70 -75 350
rect -45 70 -40 350
rect -80 60 -40 70
rect 240 350 280 360
rect 240 70 245 350
rect 275 70 280 350
rect 240 60 280 70
rect 560 350 600 360
rect 560 70 565 350
rect 595 70 600 350
rect 560 40 600 70
rect 880 350 920 360
rect 880 70 885 350
rect 915 70 920 350
rect 880 60 920 70
rect 1200 350 1240 400
rect 1200 70 1205 350
rect 1235 70 1240 350
rect 1200 60 1240 70
rect 1520 350 1560 360
rect 1520 70 1525 350
rect 1555 70 1560 350
rect 1520 60 1560 70
rect 1840 350 1880 360
rect 1840 70 1845 350
rect 1875 70 1880 350
rect 1840 40 1880 70
rect 2160 350 2200 360
rect 2160 70 2165 350
rect 2195 70 2200 350
rect 2160 60 2200 70
rect 2480 350 2520 400
rect 2480 70 2485 350
rect 2515 70 2520 350
rect 2480 60 2520 70
rect 2800 350 2840 360
rect 2800 70 2805 350
rect 2835 70 2840 350
rect 2800 60 2840 70
rect 3120 350 3160 360
rect 3120 70 3125 350
rect 3155 70 3160 350
rect 3120 40 3160 70
rect 3440 350 3480 360
rect 3440 70 3445 350
rect 3475 70 3480 350
rect 3440 60 3480 70
rect 3760 350 3800 400
rect 3760 70 3765 350
rect 3795 70 3800 350
rect 3760 60 3800 70
rect 4080 350 4120 360
rect 4080 70 4085 350
rect 4115 70 4120 350
rect 4080 60 4120 70
rect 4400 350 4440 360
rect 4400 70 4405 350
rect 4435 70 4440 350
rect 4400 40 4440 70
rect 4720 350 4760 360
rect 4720 70 4725 350
rect 4755 70 4760 350
rect 4720 60 4760 70
rect 5040 350 5080 400
rect 5040 70 5045 350
rect 5075 70 5080 350
rect 5040 60 5080 70
rect 5120 380 5160 400
rect -80 0 5080 40
rect -80 -50 -40 0
rect -80 -330 -75 -50
rect -45 -330 -40 -50
rect -80 -340 -40 -330
rect 240 -50 280 -40
rect 240 -330 245 -50
rect 275 -330 280 -50
rect 240 -340 280 -330
rect 560 -50 600 0
rect 560 -330 565 -50
rect 595 -330 600 -50
rect 560 -340 600 -330
rect 880 -50 920 -40
rect 880 -330 885 -50
rect 915 -330 920 -50
rect 880 -340 920 -330
rect 1200 -50 1240 0
rect 1200 -330 1205 -50
rect 1235 -330 1240 -50
rect 1200 -340 1240 -330
rect 1520 -50 1560 -40
rect 1520 -330 1525 -50
rect 1555 -330 1560 -50
rect 1520 -340 1560 -330
rect 1840 -50 1880 0
rect 1840 -330 1845 -50
rect 1875 -330 1880 -50
rect 1840 -340 1880 -330
rect 2160 -50 2200 -40
rect 2160 -330 2165 -50
rect 2195 -330 2200 -50
rect 2160 -340 2200 -330
rect 2480 -50 2520 0
rect 2480 -330 2485 -50
rect 2515 -330 2520 -50
rect 2480 -340 2520 -330
rect 2800 -50 2840 -40
rect 2800 -330 2805 -50
rect 2835 -330 2840 -50
rect 2800 -340 2840 -330
rect 3120 -50 3160 0
rect 3120 -330 3125 -50
rect 3155 -330 3160 -50
rect 3120 -340 3160 -330
rect 3440 -50 3480 -40
rect 3440 -330 3445 -50
rect 3475 -330 3480 -50
rect 3440 -340 3480 -330
rect 3760 -50 3800 0
rect 3760 -330 3765 -50
rect 3795 -330 3800 -50
rect 3760 -340 3800 -330
rect 4080 -50 4120 -40
rect 4080 -330 4085 -50
rect 4115 -330 4120 -50
rect 4080 -340 4120 -330
rect 4400 -50 4440 0
rect 4400 -330 4405 -50
rect 4435 -330 4440 -50
rect 4400 -340 4440 -330
rect 4720 -50 4760 -40
rect 4720 -330 4725 -50
rect 4755 -330 4760 -50
rect 4720 -340 4760 -330
rect 5040 -50 5080 0
rect 5040 -330 5045 -50
rect 5075 -330 5080 -50
rect 5040 -340 5080 -330
rect 0 -365 200 -360
rect 0 -395 10 -365
rect 190 -395 200 -365
rect 0 -400 200 -395
rect 320 -365 520 -360
rect 320 -395 330 -365
rect 510 -395 520 -365
rect 320 -400 520 -395
rect 640 -365 840 -360
rect 640 -395 650 -365
rect 830 -395 840 -365
rect 640 -400 840 -395
rect 960 -365 1160 -360
rect 960 -395 970 -365
rect 1150 -395 1160 -365
rect 960 -400 1160 -395
rect 1280 -365 1480 -360
rect 1280 -395 1290 -365
rect 1470 -395 1480 -365
rect 1280 -400 1480 -395
rect 1600 -365 1800 -360
rect 1600 -395 1610 -365
rect 1790 -395 1800 -365
rect 1600 -400 1800 -395
rect 1920 -365 2120 -360
rect 1920 -395 1930 -365
rect 2110 -395 2120 -365
rect 1920 -400 2120 -395
rect 2240 -365 2440 -360
rect 2240 -395 2250 -365
rect 2430 -395 2440 -365
rect 2240 -400 2440 -395
rect 2560 -365 2760 -360
rect 2560 -395 2570 -365
rect 2750 -395 2760 -365
rect 2560 -400 2760 -395
rect 2880 -365 3080 -360
rect 2880 -395 2890 -365
rect 3070 -395 3080 -365
rect 2880 -400 3080 -395
rect 3200 -365 3400 -360
rect 3200 -395 3210 -365
rect 3390 -395 3400 -365
rect 3200 -400 3400 -395
rect 3520 -365 3720 -360
rect 3520 -395 3530 -365
rect 3710 -395 3720 -365
rect 3520 -400 3720 -395
rect 3840 -365 4040 -360
rect 3840 -395 3850 -365
rect 4030 -395 4040 -365
rect 3840 -400 4040 -395
rect 4160 -365 4360 -360
rect 4160 -395 4170 -365
rect 4350 -395 4360 -365
rect 4160 -400 4360 -395
rect 4480 -365 4680 -360
rect 4480 -395 4490 -365
rect 4670 -395 4680 -365
rect 4480 -400 4680 -395
rect 4800 -365 5000 -360
rect 4800 -395 4810 -365
rect 4990 -395 5000 -365
rect 4800 -400 5000 -395
rect -160 -440 -120 -420
rect 5120 -440 5160 -420
rect -160 -480 -100 -440
rect 5100 -480 5160 -440
rect -200 -1040 -180 -1000
rect 5180 -1040 5200 -1000
rect 0 -1085 200 -1080
rect 0 -1115 10 -1085
rect 190 -1115 200 -1085
rect 0 -1120 200 -1115
rect 320 -1085 520 -1080
rect 320 -1115 330 -1085
rect 510 -1115 520 -1085
rect 320 -1120 520 -1115
rect 640 -1085 840 -1080
rect 640 -1115 650 -1085
rect 830 -1115 840 -1085
rect 640 -1120 840 -1115
rect 960 -1085 1160 -1080
rect 960 -1115 970 -1085
rect 1150 -1115 1160 -1085
rect 960 -1120 1160 -1115
rect 1280 -1085 1480 -1080
rect 1280 -1115 1290 -1085
rect 1470 -1115 1480 -1085
rect 1280 -1120 1480 -1115
rect 1600 -1085 1800 -1080
rect 1600 -1115 1610 -1085
rect 1790 -1115 1800 -1085
rect 1600 -1120 1800 -1115
rect 1920 -1085 2120 -1080
rect 1920 -1115 1930 -1085
rect 2110 -1115 2120 -1085
rect 1920 -1120 2120 -1115
rect 2240 -1085 2440 -1080
rect 2240 -1115 2250 -1085
rect 2430 -1115 2440 -1085
rect 2240 -1120 2440 -1115
rect 2560 -1085 2760 -1080
rect 2560 -1115 2570 -1085
rect 2750 -1115 2760 -1085
rect 2560 -1120 2760 -1115
rect 2880 -1085 3080 -1080
rect 2880 -1115 2890 -1085
rect 3070 -1115 3080 -1085
rect 2880 -1120 3080 -1115
rect 3200 -1085 3400 -1080
rect 3200 -1115 3210 -1085
rect 3390 -1115 3400 -1085
rect 3200 -1120 3400 -1115
rect 3520 -1085 3720 -1080
rect 3520 -1115 3530 -1085
rect 3710 -1115 3720 -1085
rect 3520 -1120 3720 -1115
rect 3840 -1085 4040 -1080
rect 3840 -1115 3850 -1085
rect 4030 -1115 4040 -1085
rect 3840 -1120 4040 -1115
rect 4160 -1085 4360 -1080
rect 4160 -1115 4170 -1085
rect 4350 -1115 4360 -1085
rect 4160 -1120 4360 -1115
rect 4480 -1085 4680 -1080
rect 4480 -1115 4490 -1085
rect 4670 -1115 4680 -1085
rect 4480 -1120 4680 -1115
rect 4800 -1085 5000 -1080
rect 4800 -1115 4810 -1085
rect 4990 -1115 5000 -1085
rect 4800 -1120 5000 -1115
rect -80 -1150 -40 -1140
rect -80 -1230 -75 -1150
rect -45 -1230 -40 -1150
rect -80 -1240 -40 -1230
rect 240 -1150 280 -1140
rect 240 -1230 245 -1150
rect 275 -1230 280 -1150
rect 240 -1280 280 -1230
rect 560 -1150 600 -1140
rect 560 -1230 565 -1150
rect 595 -1230 600 -1150
rect 560 -1240 600 -1230
rect 880 -1150 920 -1140
rect 880 -1230 885 -1150
rect 915 -1230 920 -1150
rect 880 -1280 920 -1230
rect 1200 -1150 1240 -1140
rect 1200 -1230 1205 -1150
rect 1235 -1230 1240 -1150
rect 1200 -1240 1240 -1230
rect 1520 -1150 1560 -1140
rect 1520 -1230 1525 -1150
rect 1555 -1230 1560 -1150
rect 1520 -1280 1560 -1230
rect 1840 -1150 1880 -1140
rect 1840 -1230 1845 -1150
rect 1875 -1230 1880 -1150
rect 1840 -1240 1880 -1230
rect 2160 -1150 2200 -1140
rect 2160 -1230 2165 -1150
rect 2195 -1230 2200 -1150
rect 2160 -1280 2200 -1230
rect 2480 -1150 2520 -1140
rect 2480 -1230 2485 -1150
rect 2515 -1230 2520 -1150
rect 2480 -1240 2520 -1230
rect 2800 -1150 2840 -1140
rect 2800 -1230 2805 -1150
rect 2835 -1230 2840 -1150
rect 2800 -1280 2840 -1230
rect 3120 -1150 3160 -1140
rect 3120 -1230 3125 -1150
rect 3155 -1230 3160 -1150
rect 3120 -1240 3160 -1230
rect 3440 -1150 3480 -1140
rect 3440 -1230 3445 -1150
rect 3475 -1230 3480 -1150
rect 3440 -1280 3480 -1230
rect 3760 -1150 3800 -1140
rect 3760 -1230 3765 -1150
rect 3795 -1230 3800 -1150
rect 3760 -1240 3800 -1230
rect 4080 -1150 4120 -1140
rect 4080 -1230 4085 -1150
rect 4115 -1230 4120 -1150
rect 4080 -1280 4120 -1230
rect 4400 -1150 4440 -1140
rect 4400 -1230 4405 -1150
rect 4435 -1230 4440 -1150
rect 4400 -1240 4440 -1230
rect 4720 -1150 4760 -1140
rect 4720 -1230 4725 -1150
rect 4755 -1230 4760 -1150
rect 4720 -1280 4760 -1230
rect 5040 -1150 5080 -1140
rect 5040 -1230 5045 -1150
rect 5075 -1230 5080 -1150
rect 5040 -1240 5080 -1230
rect -80 -1320 5080 -1280
rect -240 -1480 -200 -1460
rect -80 -1350 -40 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 -40 -1350
rect -80 -1480 -40 -1430
rect 240 -1350 280 -1340
rect 240 -1430 245 -1350
rect 275 -1430 280 -1350
rect 240 -1440 280 -1430
rect 560 -1350 600 -1320
rect 560 -1430 565 -1350
rect 595 -1430 600 -1350
rect 560 -1440 600 -1430
rect 880 -1350 920 -1340
rect 880 -1430 885 -1350
rect 915 -1430 920 -1350
rect 880 -1440 920 -1430
rect 1200 -1350 1240 -1340
rect 1200 -1430 1205 -1350
rect 1235 -1430 1240 -1350
rect 1200 -1480 1240 -1430
rect 1520 -1350 1560 -1340
rect 1520 -1430 1525 -1350
rect 1555 -1430 1560 -1350
rect 1520 -1440 1560 -1430
rect 1840 -1350 1880 -1320
rect 1840 -1430 1845 -1350
rect 1875 -1430 1880 -1350
rect 1840 -1440 1880 -1430
rect 2160 -1350 2200 -1340
rect 2160 -1430 2165 -1350
rect 2195 -1430 2200 -1350
rect 2160 -1440 2200 -1430
rect 2480 -1350 2520 -1340
rect 2480 -1430 2485 -1350
rect 2515 -1430 2520 -1350
rect 2480 -1480 2520 -1430
rect 2800 -1350 2840 -1340
rect 2800 -1430 2805 -1350
rect 2835 -1430 2840 -1350
rect 2800 -1440 2840 -1430
rect 3120 -1350 3160 -1320
rect 3120 -1430 3125 -1350
rect 3155 -1430 3160 -1350
rect 3120 -1440 3160 -1430
rect 3440 -1350 3480 -1340
rect 3440 -1430 3445 -1350
rect 3475 -1430 3480 -1350
rect 3440 -1440 3480 -1430
rect 3760 -1350 3800 -1340
rect 3760 -1430 3765 -1350
rect 3795 -1430 3800 -1350
rect 3760 -1480 3800 -1430
rect 4080 -1350 4120 -1340
rect 4080 -1430 4085 -1350
rect 4115 -1430 4120 -1350
rect 4080 -1440 4120 -1430
rect 4400 -1350 4440 -1320
rect 4400 -1430 4405 -1350
rect 4435 -1430 4440 -1350
rect 4400 -1440 4440 -1430
rect 4720 -1350 4760 -1340
rect 4720 -1430 4725 -1350
rect 4755 -1430 4760 -1350
rect 4720 -1440 4760 -1430
rect 5040 -1350 5080 -1340
rect 5040 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5040 -1480 5080 -1430
rect 5200 -1480 5240 -1460
rect -240 -1520 -180 -1480
rect 5180 -1520 5240 -1480
<< viali >>
rect -75 70 -45 350
rect 245 70 275 350
rect 565 70 595 350
rect 885 70 915 350
rect 1205 70 1235 350
rect 1525 70 1555 350
rect 1845 70 1875 350
rect 2165 70 2195 350
rect 2485 70 2515 350
rect 2805 70 2835 350
rect 3125 70 3155 350
rect 3445 70 3475 350
rect 3765 70 3795 350
rect 4085 70 4115 350
rect 4405 70 4435 350
rect 4725 70 4755 350
rect 5045 70 5075 350
rect -75 -330 -45 -50
rect 245 -330 275 -50
rect 565 -330 595 -50
rect 885 -330 915 -50
rect 1205 -330 1235 -50
rect 1525 -330 1555 -50
rect 1845 -330 1875 -50
rect 2165 -330 2195 -50
rect 2485 -330 2515 -50
rect 2805 -330 2835 -50
rect 3125 -330 3155 -50
rect 3445 -330 3475 -50
rect 3765 -330 3795 -50
rect 4085 -330 4115 -50
rect 4405 -330 4435 -50
rect 4725 -330 4755 -50
rect 5045 -330 5075 -50
rect 10 -395 190 -365
rect 330 -395 510 -365
rect 650 -395 830 -365
rect 970 -395 1150 -365
rect 1290 -395 1470 -365
rect 1610 -395 1790 -365
rect 1930 -395 2110 -365
rect 2250 -395 2430 -365
rect 2570 -395 2750 -365
rect 2890 -395 3070 -365
rect 3210 -395 3390 -365
rect 3530 -395 3710 -365
rect 3850 -395 4030 -365
rect 4170 -395 4350 -365
rect 4490 -395 4670 -365
rect 4810 -395 4990 -365
rect 10 -1115 190 -1085
rect 330 -1115 510 -1085
rect 650 -1115 830 -1085
rect 970 -1115 1150 -1085
rect 1290 -1115 1470 -1085
rect 1610 -1115 1790 -1085
rect 1930 -1115 2110 -1085
rect 2250 -1115 2430 -1085
rect 2570 -1115 2750 -1085
rect 2890 -1115 3070 -1085
rect 3210 -1115 3390 -1085
rect 3530 -1115 3710 -1085
rect 3850 -1115 4030 -1085
rect 4170 -1115 4350 -1085
rect 4490 -1115 4670 -1085
rect 4810 -1115 4990 -1085
rect -75 -1230 -45 -1150
rect 245 -1230 275 -1150
rect 565 -1230 595 -1150
rect 885 -1230 915 -1150
rect 1205 -1230 1235 -1150
rect 1525 -1230 1555 -1150
rect 1845 -1230 1875 -1150
rect 2165 -1230 2195 -1150
rect 2485 -1230 2515 -1150
rect 2805 -1230 2835 -1150
rect 3125 -1230 3155 -1150
rect 3445 -1230 3475 -1150
rect 3765 -1230 3795 -1150
rect 4085 -1230 4115 -1150
rect 4405 -1230 4435 -1150
rect 4725 -1230 4755 -1150
rect 5045 -1230 5075 -1150
rect -75 -1430 -45 -1350
rect 245 -1430 275 -1350
rect 565 -1430 595 -1350
rect 885 -1430 915 -1350
rect 1205 -1430 1235 -1350
rect 1525 -1430 1555 -1350
rect 1845 -1430 1875 -1350
rect 2165 -1430 2195 -1350
rect 2485 -1430 2515 -1350
rect 2805 -1430 2835 -1350
rect 3125 -1430 3155 -1350
rect 3445 -1430 3475 -1350
rect 3765 -1430 3795 -1350
rect 4085 -1430 4115 -1350
rect 4405 -1430 4435 -1350
rect 4725 -1430 4755 -1350
rect 5045 -1430 5075 -1350
<< metal1 >>
rect -80 350 -40 360
rect -80 70 -75 350
rect -45 70 -40 350
rect -80 60 -40 70
rect 240 350 280 360
rect 240 70 245 350
rect 275 70 280 350
rect 240 60 280 70
rect 560 350 600 360
rect 560 70 565 350
rect 595 70 600 350
rect 560 60 600 70
rect 880 350 920 360
rect 880 70 885 350
rect 915 70 920 350
rect 880 60 920 70
rect 1200 350 1240 360
rect 1200 70 1205 350
rect 1235 70 1240 350
rect 1200 60 1240 70
rect 1520 350 1560 360
rect 1520 70 1525 350
rect 1555 70 1560 350
rect 1520 60 1560 70
rect 1840 350 1880 360
rect 1840 70 1845 350
rect 1875 70 1880 350
rect 1840 60 1880 70
rect 2160 350 2200 360
rect 2160 70 2165 350
rect 2195 70 2200 350
rect 2160 60 2200 70
rect 2480 350 2520 360
rect 2480 70 2485 350
rect 2515 70 2520 350
rect 2480 60 2520 70
rect 2800 350 2840 360
rect 2800 70 2805 350
rect 2835 70 2840 350
rect 2800 60 2840 70
rect 3120 350 3160 360
rect 3120 70 3125 350
rect 3155 70 3160 350
rect 3120 60 3160 70
rect 3440 350 3480 360
rect 3440 70 3445 350
rect 3475 70 3480 350
rect 3440 60 3480 70
rect 3760 350 3800 360
rect 3760 70 3765 350
rect 3795 70 3800 350
rect 3760 60 3800 70
rect 4080 350 4120 360
rect 4080 70 4085 350
rect 4115 70 4120 350
rect 4080 60 4120 70
rect 4400 350 4440 360
rect 4400 70 4405 350
rect 4435 70 4440 350
rect 4400 60 4440 70
rect 4720 350 4760 360
rect 4720 70 4725 350
rect 4755 70 4760 350
rect 4720 60 4760 70
rect 5040 350 5080 360
rect 5040 70 5045 350
rect 5075 70 5080 350
rect 5040 60 5080 70
rect -80 -50 -40 -40
rect -80 -330 -75 -50
rect -45 -330 -40 -50
rect -80 -340 -40 -330
rect 240 -50 280 -40
rect 240 -330 245 -50
rect 275 -330 280 -50
rect 0 -365 200 -360
rect 0 -395 10 -365
rect 190 -395 200 -365
rect 0 -400 200 -395
rect 240 -685 280 -330
rect 560 -50 600 -40
rect 560 -330 565 -50
rect 595 -330 600 -50
rect 560 -340 600 -330
rect 880 -50 920 -40
rect 880 -330 885 -50
rect 915 -330 920 -50
rect 320 -365 520 -360
rect 320 -395 330 -365
rect 510 -395 520 -365
rect 320 -400 520 -395
rect 640 -365 840 -360
rect 640 -395 650 -365
rect 830 -395 840 -365
rect 640 -400 840 -395
rect 240 -715 245 -685
rect 275 -715 280 -685
rect 240 -720 280 -715
rect 880 -685 920 -330
rect 1200 -50 1240 -40
rect 1200 -330 1205 -50
rect 1235 -330 1240 -50
rect 1200 -340 1240 -330
rect 1520 -50 1560 -40
rect 1520 -330 1525 -50
rect 1555 -330 1560 -50
rect 960 -365 1160 -360
rect 960 -395 970 -365
rect 1150 -395 1160 -365
rect 960 -400 1160 -395
rect 1280 -365 1480 -360
rect 1280 -395 1290 -365
rect 1470 -395 1480 -365
rect 1280 -400 1480 -395
rect 880 -715 885 -685
rect 915 -715 920 -685
rect 880 -720 920 -715
rect 1520 -685 1560 -330
rect 1840 -50 1880 -40
rect 1840 -330 1845 -50
rect 1875 -330 1880 -50
rect 1840 -340 1880 -330
rect 2160 -50 2200 -40
rect 2160 -330 2165 -50
rect 2195 -330 2200 -50
rect 1600 -365 1800 -360
rect 1600 -395 1610 -365
rect 1790 -395 1800 -365
rect 1600 -400 1800 -395
rect 1920 -365 2120 -360
rect 1920 -395 1930 -365
rect 2110 -395 2120 -365
rect 1920 -400 2120 -395
rect 1520 -715 1525 -685
rect 1555 -715 1560 -685
rect 1520 -720 1560 -715
rect 2160 -685 2200 -330
rect 2480 -50 2520 -40
rect 2480 -330 2485 -50
rect 2515 -330 2520 -50
rect 2480 -340 2520 -330
rect 2800 -50 2840 -40
rect 2800 -330 2805 -50
rect 2835 -330 2840 -50
rect 2240 -365 2440 -360
rect 2240 -395 2250 -365
rect 2430 -395 2440 -365
rect 2240 -400 2440 -395
rect 2560 -365 2760 -360
rect 2560 -395 2570 -365
rect 2750 -395 2760 -365
rect 2560 -400 2760 -395
rect 2160 -715 2165 -685
rect 2195 -715 2200 -685
rect 2160 -720 2200 -715
rect 2800 -685 2840 -330
rect 3120 -50 3160 -40
rect 3120 -330 3125 -50
rect 3155 -330 3160 -50
rect 3120 -340 3160 -330
rect 3440 -50 3480 -40
rect 3440 -330 3445 -50
rect 3475 -330 3480 -50
rect 2880 -365 3080 -360
rect 2880 -395 2890 -365
rect 3070 -395 3080 -365
rect 2880 -400 3080 -395
rect 3200 -365 3400 -360
rect 3200 -395 3210 -365
rect 3390 -395 3400 -365
rect 3200 -400 3400 -395
rect 2800 -715 2805 -685
rect 2835 -715 2840 -685
rect 2800 -720 2840 -715
rect 3440 -685 3480 -330
rect 3760 -50 3800 -40
rect 3760 -330 3765 -50
rect 3795 -330 3800 -50
rect 3760 -340 3800 -330
rect 4080 -50 4120 -40
rect 4080 -330 4085 -50
rect 4115 -330 4120 -50
rect 3520 -365 3720 -360
rect 3520 -395 3530 -365
rect 3710 -395 3720 -365
rect 3520 -400 3720 -395
rect 3840 -365 4040 -360
rect 3840 -395 3850 -365
rect 4030 -395 4040 -365
rect 3840 -400 4040 -395
rect 3440 -715 3445 -685
rect 3475 -715 3480 -685
rect 3440 -720 3480 -715
rect 4080 -685 4120 -330
rect 4400 -50 4440 -40
rect 4400 -330 4405 -50
rect 4435 -330 4440 -50
rect 4400 -340 4440 -330
rect 4720 -50 4760 -40
rect 4720 -330 4725 -50
rect 4755 -330 4760 -50
rect 4160 -365 4360 -360
rect 4160 -395 4170 -365
rect 4350 -395 4360 -365
rect 4160 -400 4360 -395
rect 4480 -365 4680 -360
rect 4480 -395 4490 -365
rect 4670 -395 4680 -365
rect 4480 -400 4680 -395
rect 4080 -715 4085 -685
rect 4115 -715 4120 -685
rect 4080 -720 4120 -715
rect 4720 -685 4760 -330
rect 5040 -50 5080 -40
rect 5040 -330 5045 -50
rect 5075 -330 5080 -50
rect 5040 -340 5080 -330
rect 4800 -365 5000 -360
rect 4800 -395 4810 -365
rect 4990 -395 5000 -365
rect 4800 -400 5000 -395
rect 4720 -715 4725 -685
rect 4755 -715 4760 -685
rect 4720 -720 4760 -715
rect -80 -845 -40 -840
rect -80 -875 -75 -845
rect -45 -875 -40 -845
rect -80 -1150 -40 -875
rect 560 -845 600 -840
rect 560 -875 565 -845
rect 595 -875 600 -845
rect 0 -1085 200 -1080
rect 0 -1115 10 -1085
rect 190 -1115 200 -1085
rect 0 -1120 200 -1115
rect 320 -1085 520 -1080
rect 320 -1115 330 -1085
rect 510 -1115 520 -1085
rect 320 -1120 520 -1115
rect -80 -1230 -75 -1150
rect -45 -1230 -40 -1150
rect -80 -1240 -40 -1230
rect 240 -1150 280 -1140
rect 240 -1230 245 -1150
rect 275 -1230 280 -1150
rect 240 -1245 280 -1230
rect 560 -1150 600 -875
rect 1200 -845 1240 -840
rect 1200 -875 1205 -845
rect 1235 -875 1240 -845
rect 640 -1085 840 -1080
rect 640 -1115 650 -1085
rect 830 -1115 840 -1085
rect 640 -1120 840 -1115
rect 960 -1085 1160 -1080
rect 960 -1115 970 -1085
rect 1150 -1115 1160 -1085
rect 960 -1120 1160 -1115
rect 560 -1230 565 -1150
rect 595 -1230 600 -1150
rect 560 -1240 600 -1230
rect 880 -1150 920 -1140
rect 880 -1230 885 -1150
rect 915 -1230 920 -1150
rect 240 -1275 245 -1245
rect 275 -1275 280 -1245
rect 240 -1280 280 -1275
rect 880 -1245 920 -1230
rect 1200 -1150 1240 -875
rect 1840 -845 1880 -840
rect 1840 -875 1845 -845
rect 1875 -875 1880 -845
rect 1280 -1085 1480 -1080
rect 1280 -1115 1290 -1085
rect 1470 -1115 1480 -1085
rect 1280 -1120 1480 -1115
rect 1600 -1085 1800 -1080
rect 1600 -1115 1610 -1085
rect 1790 -1115 1800 -1085
rect 1600 -1120 1800 -1115
rect 1200 -1230 1205 -1150
rect 1235 -1230 1240 -1150
rect 1200 -1240 1240 -1230
rect 1520 -1150 1560 -1140
rect 1520 -1230 1525 -1150
rect 1555 -1230 1560 -1150
rect 880 -1275 885 -1245
rect 915 -1275 920 -1245
rect 880 -1280 920 -1275
rect 1520 -1245 1560 -1230
rect 1840 -1150 1880 -875
rect 2480 -845 2520 -840
rect 2480 -875 2485 -845
rect 2515 -875 2520 -845
rect 1920 -1085 2120 -1080
rect 1920 -1115 1930 -1085
rect 2110 -1115 2120 -1085
rect 1920 -1120 2120 -1115
rect 2240 -1085 2440 -1080
rect 2240 -1115 2250 -1085
rect 2430 -1115 2440 -1085
rect 2240 -1120 2440 -1115
rect 1840 -1230 1845 -1150
rect 1875 -1230 1880 -1150
rect 1840 -1240 1880 -1230
rect 2160 -1150 2200 -1140
rect 2160 -1230 2165 -1150
rect 2195 -1230 2200 -1150
rect 1520 -1275 1525 -1245
rect 1555 -1275 1560 -1245
rect 1520 -1280 1560 -1275
rect 2160 -1245 2200 -1230
rect 2480 -1150 2520 -875
rect 3120 -845 3160 -840
rect 3120 -875 3125 -845
rect 3155 -875 3160 -845
rect 2560 -1085 2760 -1080
rect 2560 -1115 2570 -1085
rect 2750 -1115 2760 -1085
rect 2560 -1120 2760 -1115
rect 2880 -1085 3080 -1080
rect 2880 -1115 2890 -1085
rect 3070 -1115 3080 -1085
rect 2880 -1120 3080 -1115
rect 2480 -1230 2485 -1150
rect 2515 -1230 2520 -1150
rect 2480 -1240 2520 -1230
rect 2800 -1150 2840 -1140
rect 2800 -1230 2805 -1150
rect 2835 -1230 2840 -1150
rect 2160 -1275 2165 -1245
rect 2195 -1275 2200 -1245
rect 2160 -1280 2200 -1275
rect 2800 -1245 2840 -1230
rect 3120 -1150 3160 -875
rect 3760 -845 3800 -840
rect 3760 -875 3765 -845
rect 3795 -875 3800 -845
rect 3200 -1085 3400 -1080
rect 3200 -1115 3210 -1085
rect 3390 -1115 3400 -1085
rect 3200 -1120 3400 -1115
rect 3520 -1085 3720 -1080
rect 3520 -1115 3530 -1085
rect 3710 -1115 3720 -1085
rect 3520 -1120 3720 -1115
rect 3120 -1230 3125 -1150
rect 3155 -1230 3160 -1150
rect 3120 -1240 3160 -1230
rect 3440 -1150 3480 -1140
rect 3440 -1230 3445 -1150
rect 3475 -1230 3480 -1150
rect 2800 -1275 2805 -1245
rect 2835 -1275 2840 -1245
rect 2800 -1280 2840 -1275
rect 3440 -1245 3480 -1230
rect 3760 -1150 3800 -875
rect 4400 -845 4440 -840
rect 4400 -875 4405 -845
rect 4435 -875 4440 -845
rect 3840 -1085 4040 -1080
rect 3840 -1115 3850 -1085
rect 4030 -1115 4040 -1085
rect 3840 -1120 4040 -1115
rect 4160 -1085 4360 -1080
rect 4160 -1115 4170 -1085
rect 4350 -1115 4360 -1085
rect 4160 -1120 4360 -1115
rect 3760 -1230 3765 -1150
rect 3795 -1230 3800 -1150
rect 3760 -1240 3800 -1230
rect 4080 -1150 4120 -1140
rect 4080 -1230 4085 -1150
rect 4115 -1230 4120 -1150
rect 3440 -1275 3445 -1245
rect 3475 -1275 3480 -1245
rect 3440 -1280 3480 -1275
rect 4080 -1245 4120 -1230
rect 4400 -1150 4440 -875
rect 5040 -845 5080 -840
rect 5040 -875 5045 -845
rect 5075 -875 5080 -845
rect 4480 -1085 4680 -1080
rect 4480 -1115 4490 -1085
rect 4670 -1115 4680 -1085
rect 4480 -1120 4680 -1115
rect 4800 -1085 5000 -1080
rect 4800 -1115 4810 -1085
rect 4990 -1115 5000 -1085
rect 4800 -1120 5000 -1115
rect 4400 -1230 4405 -1150
rect 4435 -1230 4440 -1150
rect 4400 -1240 4440 -1230
rect 4720 -1150 4760 -1140
rect 4720 -1230 4725 -1150
rect 4755 -1230 4760 -1150
rect 4080 -1275 4085 -1245
rect 4115 -1275 4120 -1245
rect 4080 -1280 4120 -1275
rect 4720 -1245 4760 -1230
rect 5040 -1150 5080 -875
rect 5040 -1230 5045 -1150
rect 5075 -1230 5080 -1150
rect 5040 -1240 5080 -1230
rect 4720 -1275 4725 -1245
rect 4755 -1275 4760 -1245
rect 4720 -1280 4760 -1275
rect -80 -1350 -40 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 -40 -1350
rect -80 -1440 -40 -1430
rect 240 -1350 280 -1340
rect 240 -1430 245 -1350
rect 275 -1430 280 -1350
rect 240 -1440 280 -1430
rect 560 -1350 600 -1340
rect 560 -1430 565 -1350
rect 595 -1430 600 -1350
rect 560 -1440 600 -1430
rect 880 -1350 920 -1340
rect 880 -1430 885 -1350
rect 915 -1430 920 -1350
rect 880 -1440 920 -1430
rect 1200 -1350 1240 -1340
rect 1200 -1430 1205 -1350
rect 1235 -1430 1240 -1350
rect 1200 -1440 1240 -1430
rect 1520 -1350 1560 -1340
rect 1520 -1430 1525 -1350
rect 1555 -1430 1560 -1350
rect 1520 -1440 1560 -1430
rect 1840 -1350 1880 -1340
rect 1840 -1430 1845 -1350
rect 1875 -1430 1880 -1350
rect 1840 -1440 1880 -1430
rect 2160 -1350 2200 -1340
rect 2160 -1430 2165 -1350
rect 2195 -1430 2200 -1350
rect 2160 -1440 2200 -1430
rect 2480 -1350 2520 -1340
rect 2480 -1430 2485 -1350
rect 2515 -1430 2520 -1350
rect 2480 -1440 2520 -1430
rect 2800 -1350 2840 -1340
rect 2800 -1430 2805 -1350
rect 2835 -1430 2840 -1350
rect 2800 -1440 2840 -1430
rect 3120 -1350 3160 -1340
rect 3120 -1430 3125 -1350
rect 3155 -1430 3160 -1350
rect 3120 -1440 3160 -1430
rect 3440 -1350 3480 -1340
rect 3440 -1430 3445 -1350
rect 3475 -1430 3480 -1350
rect 3440 -1440 3480 -1430
rect 3760 -1350 3800 -1340
rect 3760 -1430 3765 -1350
rect 3795 -1430 3800 -1350
rect 3760 -1440 3800 -1430
rect 4080 -1350 4120 -1340
rect 4080 -1430 4085 -1350
rect 4115 -1430 4120 -1350
rect 4080 -1440 4120 -1430
rect 4400 -1350 4440 -1340
rect 4400 -1430 4405 -1350
rect 4435 -1430 4440 -1350
rect 4400 -1440 4440 -1430
rect 4720 -1350 4760 -1340
rect 4720 -1430 4725 -1350
rect 4755 -1430 4760 -1350
rect 4720 -1440 4760 -1430
rect 5040 -1350 5080 -1340
rect 5040 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5040 -1440 5080 -1430
<< via1 >>
rect -75 130 -45 310
rect 1205 130 1235 310
rect 2485 130 2515 310
rect 3765 130 3795 310
rect 5045 130 5075 310
rect 10 -395 190 -365
rect 330 -395 510 -365
rect 650 -395 830 -365
rect 245 -715 275 -685
rect 970 -395 1150 -365
rect 1290 -395 1470 -365
rect 885 -715 915 -685
rect 1610 -395 1790 -365
rect 1930 -395 2110 -365
rect 1525 -715 1555 -685
rect 2250 -395 2430 -365
rect 2570 -395 2750 -365
rect 2165 -715 2195 -685
rect 2890 -395 3070 -365
rect 3210 -395 3390 -365
rect 2805 -715 2835 -685
rect 3530 -395 3710 -365
rect 3850 -395 4030 -365
rect 3445 -715 3475 -685
rect 4170 -395 4350 -365
rect 4490 -395 4670 -365
rect 4085 -715 4115 -685
rect 4810 -395 4990 -365
rect 4725 -715 4755 -685
rect -75 -875 -45 -845
rect 565 -875 595 -845
rect 10 -1115 190 -1085
rect 330 -1115 510 -1085
rect 1205 -875 1235 -845
rect 650 -1115 830 -1085
rect 970 -1115 1150 -1085
rect 245 -1275 275 -1245
rect 1845 -875 1875 -845
rect 1290 -1115 1470 -1085
rect 1610 -1115 1790 -1085
rect 885 -1275 915 -1245
rect 2485 -875 2515 -845
rect 1930 -1115 2110 -1085
rect 2250 -1115 2430 -1085
rect 1525 -1275 1555 -1245
rect 3125 -875 3155 -845
rect 2570 -1115 2750 -1085
rect 2890 -1115 3070 -1085
rect 2165 -1275 2195 -1245
rect 3765 -875 3795 -845
rect 3210 -1115 3390 -1085
rect 3530 -1115 3710 -1085
rect 2805 -1275 2835 -1245
rect 4405 -875 4435 -845
rect 3850 -1115 4030 -1085
rect 4170 -1115 4350 -1085
rect 3445 -1275 3475 -1245
rect 5045 -875 5075 -845
rect 4490 -1115 4670 -1085
rect 4810 -1115 4990 -1085
rect 4085 -1275 4115 -1245
rect 4725 -1275 4755 -1245
rect -75 -1430 -45 -1350
rect 1205 -1430 1235 -1350
rect 2485 -1430 2515 -1350
rect 3765 -1430 3795 -1350
rect 5045 -1430 5075 -1350
<< metal2 >>
rect -80 310 -40 320
rect -80 130 -75 310
rect -45 130 -40 310
rect -80 120 -40 130
rect 1200 310 1240 320
rect 1200 130 1205 310
rect 1235 130 1240 310
rect 1200 120 1240 130
rect 2480 310 2520 320
rect 2480 130 2485 310
rect 2515 130 2520 310
rect 2480 120 2520 130
rect 3760 310 3800 320
rect 3760 130 3765 310
rect 3795 130 3800 310
rect 3760 120 3800 130
rect 5040 310 5080 320
rect 5040 130 5045 310
rect 5075 130 5080 310
rect 5040 120 5080 130
rect -240 -320 5240 -280
rect -240 -365 5240 -360
rect -240 -395 10 -365
rect 190 -395 330 -365
rect 510 -395 650 -365
rect 830 -395 970 -365
rect 1150 -395 1290 -365
rect 1470 -395 1610 -365
rect 1790 -395 1930 -365
rect 2110 -395 2250 -365
rect 2430 -395 2570 -365
rect 2750 -395 2890 -365
rect 3070 -395 3210 -365
rect 3390 -395 3530 -365
rect 3710 -395 3850 -365
rect 4030 -395 4170 -365
rect 4350 -395 4490 -365
rect 4670 -395 4810 -365
rect 4990 -395 5240 -365
rect -240 -400 5240 -395
rect -240 -480 5240 -440
rect -240 -560 5240 -520
rect -240 -640 5240 -600
rect -240 -685 5240 -680
rect -240 -715 245 -685
rect 275 -715 885 -685
rect 915 -715 1525 -685
rect 1555 -715 2165 -685
rect 2195 -715 2805 -685
rect 2835 -715 3445 -685
rect 3475 -715 4085 -685
rect 4115 -715 4725 -685
rect 4755 -715 5240 -685
rect -240 -720 5240 -715
rect -240 -800 5240 -760
rect -240 -845 5240 -840
rect -240 -875 -75 -845
rect -45 -875 565 -845
rect 595 -875 1205 -845
rect 1235 -875 1845 -845
rect 1875 -875 2485 -845
rect 2515 -875 3125 -845
rect 3155 -875 3765 -845
rect 3795 -875 4405 -845
rect 4435 -875 5045 -845
rect 5075 -875 5240 -845
rect -240 -880 5240 -875
rect -240 -960 5240 -920
rect -240 -1005 5240 -1000
rect -240 -1035 -235 -1005
rect -205 -1035 -155 -1005
rect -125 -1035 -75 -1005
rect -45 -1035 5 -1005
rect 35 -1035 85 -1005
rect 115 -1035 165 -1005
rect 195 -1035 245 -1005
rect 275 -1035 325 -1005
rect 355 -1035 405 -1005
rect 435 -1035 485 -1005
rect 515 -1035 565 -1005
rect 595 -1035 645 -1005
rect 675 -1035 725 -1005
rect 755 -1035 805 -1005
rect 835 -1035 885 -1005
rect 915 -1035 965 -1005
rect 995 -1035 1045 -1005
rect 1075 -1035 1125 -1005
rect 1155 -1035 1205 -1005
rect 1235 -1035 1285 -1005
rect 1315 -1035 1365 -1005
rect 1395 -1035 1445 -1005
rect 1475 -1035 1525 -1005
rect 1555 -1035 1605 -1005
rect 1635 -1035 1685 -1005
rect 1715 -1035 1765 -1005
rect 1795 -1035 1845 -1005
rect 1875 -1035 1925 -1005
rect 1955 -1035 2005 -1005
rect 2035 -1035 2085 -1005
rect 2115 -1035 2165 -1005
rect 2195 -1035 2245 -1005
rect 2275 -1035 2325 -1005
rect 2355 -1035 2405 -1005
rect 2435 -1035 2485 -1005
rect 2515 -1035 2565 -1005
rect 2595 -1035 2645 -1005
rect 2675 -1035 2725 -1005
rect 2755 -1035 2805 -1005
rect 2835 -1035 2885 -1005
rect 2915 -1035 2965 -1005
rect 2995 -1035 3045 -1005
rect 3075 -1035 3125 -1005
rect 3155 -1035 3205 -1005
rect 3235 -1035 3285 -1005
rect 3315 -1035 3365 -1005
rect 3395 -1035 3445 -1005
rect 3475 -1035 3525 -1005
rect 3555 -1035 3605 -1005
rect 3635 -1035 3685 -1005
rect 3715 -1035 3765 -1005
rect 3795 -1035 3845 -1005
rect 3875 -1035 3925 -1005
rect 3955 -1035 4005 -1005
rect 4035 -1035 4085 -1005
rect 4115 -1035 4165 -1005
rect 4195 -1035 4245 -1005
rect 4275 -1035 4325 -1005
rect 4355 -1035 4405 -1005
rect 4435 -1035 4485 -1005
rect 4515 -1035 4565 -1005
rect 4595 -1035 4645 -1005
rect 4675 -1035 4725 -1005
rect 4755 -1035 4805 -1005
rect 4835 -1035 4885 -1005
rect 4915 -1035 4965 -1005
rect 4995 -1035 5045 -1005
rect 5075 -1035 5125 -1005
rect 5155 -1035 5205 -1005
rect 5235 -1035 5240 -1005
rect -240 -1040 5240 -1035
rect -240 -1085 5240 -1080
rect -240 -1115 10 -1085
rect 190 -1115 330 -1085
rect 510 -1115 650 -1085
rect 830 -1115 970 -1085
rect 1150 -1115 1290 -1085
rect 1470 -1115 1610 -1085
rect 1790 -1115 1930 -1085
rect 2110 -1115 2250 -1085
rect 2430 -1115 2570 -1085
rect 2750 -1115 2890 -1085
rect 3070 -1115 3210 -1085
rect 3390 -1115 3530 -1085
rect 3710 -1115 3850 -1085
rect 4030 -1115 4170 -1085
rect 4350 -1115 4490 -1085
rect 4670 -1115 4810 -1085
rect 4990 -1115 5240 -1085
rect -240 -1120 5240 -1115
rect -240 -1165 5240 -1160
rect -240 -1195 -235 -1165
rect -205 -1195 -155 -1165
rect -125 -1195 -75 -1165
rect -45 -1195 5 -1165
rect 35 -1195 85 -1165
rect 115 -1195 165 -1165
rect 195 -1195 245 -1165
rect 275 -1195 325 -1165
rect 355 -1195 405 -1165
rect 435 -1195 485 -1165
rect 515 -1195 565 -1165
rect 595 -1195 645 -1165
rect 675 -1195 725 -1165
rect 755 -1195 805 -1165
rect 835 -1195 885 -1165
rect 915 -1195 965 -1165
rect 995 -1195 1045 -1165
rect 1075 -1195 1125 -1165
rect 1155 -1195 1205 -1165
rect 1235 -1195 1285 -1165
rect 1315 -1195 1365 -1165
rect 1395 -1195 1445 -1165
rect 1475 -1195 1525 -1165
rect 1555 -1195 1605 -1165
rect 1635 -1195 1685 -1165
rect 1715 -1195 1765 -1165
rect 1795 -1195 1845 -1165
rect 1875 -1195 1925 -1165
rect 1955 -1195 2005 -1165
rect 2035 -1195 2085 -1165
rect 2115 -1195 2165 -1165
rect 2195 -1195 2245 -1165
rect 2275 -1195 2325 -1165
rect 2355 -1195 2405 -1165
rect 2435 -1195 2485 -1165
rect 2515 -1195 2565 -1165
rect 2595 -1195 2645 -1165
rect 2675 -1195 2725 -1165
rect 2755 -1195 2805 -1165
rect 2835 -1195 2885 -1165
rect 2915 -1195 2965 -1165
rect 2995 -1195 3045 -1165
rect 3075 -1195 3125 -1165
rect 3155 -1195 3205 -1165
rect 3235 -1195 3285 -1165
rect 3315 -1195 3365 -1165
rect 3395 -1195 3445 -1165
rect 3475 -1195 3525 -1165
rect 3555 -1195 3605 -1165
rect 3635 -1195 3685 -1165
rect 3715 -1195 3765 -1165
rect 3795 -1195 3845 -1165
rect 3875 -1195 3925 -1165
rect 3955 -1195 4005 -1165
rect 4035 -1195 4085 -1165
rect 4115 -1195 4165 -1165
rect 4195 -1195 4245 -1165
rect 4275 -1195 4325 -1165
rect 4355 -1195 4405 -1165
rect 4435 -1195 4485 -1165
rect 4515 -1195 4565 -1165
rect 4595 -1195 4645 -1165
rect 4675 -1195 4725 -1165
rect 4755 -1195 4805 -1165
rect 4835 -1195 4885 -1165
rect 4915 -1195 4965 -1165
rect 4995 -1195 5045 -1165
rect 5075 -1195 5125 -1165
rect 5155 -1195 5205 -1165
rect 5235 -1195 5240 -1165
rect -240 -1200 5240 -1195
rect -240 -1245 5240 -1240
rect -240 -1275 245 -1245
rect 275 -1275 885 -1245
rect 915 -1275 1525 -1245
rect 1555 -1275 2165 -1245
rect 2195 -1275 2805 -1245
rect 2835 -1275 3445 -1245
rect 3475 -1275 4085 -1245
rect 4115 -1275 4725 -1245
rect 4755 -1275 5240 -1245
rect -240 -1280 5240 -1275
rect -240 -1325 5080 -1320
rect -240 -1355 -235 -1325
rect -205 -1355 -155 -1325
rect -125 -1355 -75 -1325
rect -240 -1360 -75 -1355
rect -80 -1430 -75 -1360
rect -45 -1355 5 -1325
rect 35 -1355 85 -1325
rect 115 -1355 165 -1325
rect 195 -1355 245 -1325
rect 275 -1355 325 -1325
rect 355 -1355 405 -1325
rect 435 -1355 485 -1325
rect 515 -1355 645 -1325
rect 675 -1355 725 -1325
rect 755 -1355 805 -1325
rect 835 -1355 885 -1325
rect 915 -1355 965 -1325
rect 995 -1355 1045 -1325
rect 1075 -1355 1125 -1325
rect 1155 -1355 1205 -1325
rect -45 -1360 1205 -1355
rect -45 -1430 -40 -1360
rect -80 -1440 -40 -1430
rect 1200 -1430 1205 -1360
rect 1235 -1355 1285 -1325
rect 1315 -1355 1365 -1325
rect 1395 -1355 1445 -1325
rect 1475 -1355 1525 -1325
rect 1555 -1355 1605 -1325
rect 1635 -1355 1685 -1325
rect 1715 -1355 1765 -1325
rect 1795 -1355 1925 -1325
rect 1955 -1355 2005 -1325
rect 2035 -1355 2085 -1325
rect 2115 -1355 2165 -1325
rect 2195 -1355 2245 -1325
rect 2275 -1355 2325 -1325
rect 2355 -1355 2405 -1325
rect 2435 -1355 2485 -1325
rect 1235 -1360 2485 -1355
rect 1235 -1430 1240 -1360
rect 1200 -1440 1240 -1430
rect 2480 -1430 2485 -1360
rect 2515 -1355 2565 -1325
rect 2595 -1355 2645 -1325
rect 2675 -1355 2725 -1325
rect 2755 -1355 2805 -1325
rect 2835 -1355 2885 -1325
rect 2915 -1355 2965 -1325
rect 2995 -1355 3045 -1325
rect 3075 -1355 3205 -1325
rect 3235 -1355 3285 -1325
rect 3315 -1355 3365 -1325
rect 3395 -1355 3445 -1325
rect 3475 -1355 3525 -1325
rect 3555 -1355 3605 -1325
rect 3635 -1355 3685 -1325
rect 3715 -1355 3765 -1325
rect 2515 -1360 3765 -1355
rect 2515 -1430 2520 -1360
rect 2480 -1440 2520 -1430
rect 3760 -1430 3765 -1360
rect 3795 -1355 3845 -1325
rect 3875 -1355 3925 -1325
rect 3955 -1355 4005 -1325
rect 4035 -1355 4085 -1325
rect 4115 -1355 4165 -1325
rect 4195 -1355 4245 -1325
rect 4275 -1355 4325 -1325
rect 4355 -1355 4485 -1325
rect 4515 -1355 4565 -1325
rect 4595 -1355 4645 -1325
rect 4675 -1355 4725 -1325
rect 4755 -1355 4805 -1325
rect 4835 -1355 4885 -1325
rect 4915 -1355 4965 -1325
rect 4995 -1355 5045 -1325
rect 3795 -1360 5045 -1355
rect 3795 -1430 3800 -1360
rect 3760 -1440 3800 -1430
rect 5040 -1430 5045 -1360
rect 5075 -1430 5080 -1325
rect 5120 -1325 5240 -1320
rect 5120 -1355 5125 -1325
rect 5155 -1355 5205 -1325
rect 5235 -1355 5240 -1325
rect 5120 -1360 5240 -1355
rect 5040 -1440 5080 -1430
<< via2 >>
rect -75 130 -45 310
rect 1205 130 1235 310
rect 2485 130 2515 310
rect 3765 130 3795 310
rect 5045 130 5075 310
rect -235 -1035 -205 -1005
rect -155 -1035 -125 -1005
rect -75 -1035 -45 -1005
rect 5 -1035 35 -1005
rect 85 -1035 115 -1005
rect 165 -1035 195 -1005
rect 245 -1035 275 -1005
rect 325 -1035 355 -1005
rect 405 -1035 435 -1005
rect 485 -1035 515 -1005
rect 565 -1035 595 -1005
rect 645 -1035 675 -1005
rect 725 -1035 755 -1005
rect 805 -1035 835 -1005
rect 885 -1035 915 -1005
rect 965 -1035 995 -1005
rect 1045 -1035 1075 -1005
rect 1125 -1035 1155 -1005
rect 1205 -1035 1235 -1005
rect 1285 -1035 1315 -1005
rect 1365 -1035 1395 -1005
rect 1445 -1035 1475 -1005
rect 1525 -1035 1555 -1005
rect 1605 -1035 1635 -1005
rect 1685 -1035 1715 -1005
rect 1765 -1035 1795 -1005
rect 1845 -1035 1875 -1005
rect 1925 -1035 1955 -1005
rect 2005 -1035 2035 -1005
rect 2085 -1035 2115 -1005
rect 2165 -1035 2195 -1005
rect 2245 -1035 2275 -1005
rect 2325 -1035 2355 -1005
rect 2405 -1035 2435 -1005
rect 2485 -1035 2515 -1005
rect 2565 -1035 2595 -1005
rect 2645 -1035 2675 -1005
rect 2725 -1035 2755 -1005
rect 2805 -1035 2835 -1005
rect 2885 -1035 2915 -1005
rect 2965 -1035 2995 -1005
rect 3045 -1035 3075 -1005
rect 3125 -1035 3155 -1005
rect 3205 -1035 3235 -1005
rect 3285 -1035 3315 -1005
rect 3365 -1035 3395 -1005
rect 3445 -1035 3475 -1005
rect 3525 -1035 3555 -1005
rect 3605 -1035 3635 -1005
rect 3685 -1035 3715 -1005
rect 3765 -1035 3795 -1005
rect 3845 -1035 3875 -1005
rect 3925 -1035 3955 -1005
rect 4005 -1035 4035 -1005
rect 4085 -1035 4115 -1005
rect 4165 -1035 4195 -1005
rect 4245 -1035 4275 -1005
rect 4325 -1035 4355 -1005
rect 4405 -1035 4435 -1005
rect 4485 -1035 4515 -1005
rect 4565 -1035 4595 -1005
rect 4645 -1035 4675 -1005
rect 4725 -1035 4755 -1005
rect 4805 -1035 4835 -1005
rect 4885 -1035 4915 -1005
rect 4965 -1035 4995 -1005
rect 5045 -1035 5075 -1005
rect 5125 -1035 5155 -1005
rect 5205 -1035 5235 -1005
rect -235 -1195 -205 -1165
rect -155 -1195 -125 -1165
rect -75 -1195 -45 -1165
rect 5 -1195 35 -1165
rect 85 -1195 115 -1165
rect 165 -1195 195 -1165
rect 245 -1195 275 -1165
rect 325 -1195 355 -1165
rect 405 -1195 435 -1165
rect 485 -1195 515 -1165
rect 565 -1195 595 -1165
rect 645 -1195 675 -1165
rect 725 -1195 755 -1165
rect 805 -1195 835 -1165
rect 885 -1195 915 -1165
rect 965 -1195 995 -1165
rect 1045 -1195 1075 -1165
rect 1125 -1195 1155 -1165
rect 1205 -1195 1235 -1165
rect 1285 -1195 1315 -1165
rect 1365 -1195 1395 -1165
rect 1445 -1195 1475 -1165
rect 1525 -1195 1555 -1165
rect 1605 -1195 1635 -1165
rect 1685 -1195 1715 -1165
rect 1765 -1195 1795 -1165
rect 1845 -1195 1875 -1165
rect 1925 -1195 1955 -1165
rect 2005 -1195 2035 -1165
rect 2085 -1195 2115 -1165
rect 2165 -1195 2195 -1165
rect 2245 -1195 2275 -1165
rect 2325 -1195 2355 -1165
rect 2405 -1195 2435 -1165
rect 2485 -1195 2515 -1165
rect 2565 -1195 2595 -1165
rect 2645 -1195 2675 -1165
rect 2725 -1195 2755 -1165
rect 2805 -1195 2835 -1165
rect 2885 -1195 2915 -1165
rect 2965 -1195 2995 -1165
rect 3045 -1195 3075 -1165
rect 3125 -1195 3155 -1165
rect 3205 -1195 3235 -1165
rect 3285 -1195 3315 -1165
rect 3365 -1195 3395 -1165
rect 3445 -1195 3475 -1165
rect 3525 -1195 3555 -1165
rect 3605 -1195 3635 -1165
rect 3685 -1195 3715 -1165
rect 3765 -1195 3795 -1165
rect 3845 -1195 3875 -1165
rect 3925 -1195 3955 -1165
rect 4005 -1195 4035 -1165
rect 4085 -1195 4115 -1165
rect 4165 -1195 4195 -1165
rect 4245 -1195 4275 -1165
rect 4325 -1195 4355 -1165
rect 4405 -1195 4435 -1165
rect 4485 -1195 4515 -1165
rect 4565 -1195 4595 -1165
rect 4645 -1195 4675 -1165
rect 4725 -1195 4755 -1165
rect 4805 -1195 4835 -1165
rect 4885 -1195 4915 -1165
rect 4965 -1195 4995 -1165
rect 5045 -1195 5075 -1165
rect 5125 -1195 5155 -1165
rect 5205 -1195 5235 -1165
rect -235 -1355 -205 -1325
rect -155 -1355 -125 -1325
rect -75 -1350 -45 -1325
rect -75 -1430 -45 -1350
rect 5 -1355 35 -1325
rect 85 -1355 115 -1325
rect 165 -1355 195 -1325
rect 245 -1355 275 -1325
rect 325 -1355 355 -1325
rect 405 -1355 435 -1325
rect 485 -1355 515 -1325
rect 645 -1355 675 -1325
rect 725 -1355 755 -1325
rect 805 -1355 835 -1325
rect 885 -1355 915 -1325
rect 965 -1355 995 -1325
rect 1045 -1355 1075 -1325
rect 1125 -1355 1155 -1325
rect 1205 -1350 1235 -1325
rect 1205 -1430 1235 -1350
rect 1285 -1355 1315 -1325
rect 1365 -1355 1395 -1325
rect 1445 -1355 1475 -1325
rect 1525 -1355 1555 -1325
rect 1605 -1355 1635 -1325
rect 1685 -1355 1715 -1325
rect 1765 -1355 1795 -1325
rect 1925 -1355 1955 -1325
rect 2005 -1355 2035 -1325
rect 2085 -1355 2115 -1325
rect 2165 -1355 2195 -1325
rect 2245 -1355 2275 -1325
rect 2325 -1355 2355 -1325
rect 2405 -1355 2435 -1325
rect 2485 -1350 2515 -1325
rect 2485 -1430 2515 -1350
rect 2565 -1355 2595 -1325
rect 2645 -1355 2675 -1325
rect 2725 -1355 2755 -1325
rect 2805 -1355 2835 -1325
rect 2885 -1355 2915 -1325
rect 2965 -1355 2995 -1325
rect 3045 -1355 3075 -1325
rect 3205 -1355 3235 -1325
rect 3285 -1355 3315 -1325
rect 3365 -1355 3395 -1325
rect 3445 -1355 3475 -1325
rect 3525 -1355 3555 -1325
rect 3605 -1355 3635 -1325
rect 3685 -1355 3715 -1325
rect 3765 -1350 3795 -1325
rect 3765 -1430 3795 -1350
rect 3845 -1355 3875 -1325
rect 3925 -1355 3955 -1325
rect 4005 -1355 4035 -1325
rect 4085 -1355 4115 -1325
rect 4165 -1355 4195 -1325
rect 4245 -1355 4275 -1325
rect 4325 -1355 4355 -1325
rect 4485 -1355 4515 -1325
rect 4565 -1355 4595 -1325
rect 4645 -1355 4675 -1325
rect 4725 -1355 4755 -1325
rect 4805 -1355 4835 -1325
rect 4885 -1355 4915 -1325
rect 4965 -1355 4995 -1325
rect 5045 -1350 5075 -1325
rect 5045 -1430 5075 -1350
rect 5125 -1355 5155 -1325
rect 5205 -1355 5235 -1325
<< metal3 >>
rect -80 311 -40 320
rect -80 129 -76 311
rect -44 129 -40 311
rect -80 60 -40 129
rect 1200 311 1240 320
rect 1200 129 1204 311
rect 1236 129 1240 311
rect 1200 60 1240 129
rect 2480 311 2520 320
rect 2480 129 2484 311
rect 2516 129 2520 311
rect 2480 60 2520 129
rect 3760 311 3800 320
rect 3760 129 3764 311
rect 3796 129 3800 311
rect 3760 60 3800 129
rect 5040 311 5080 320
rect 5040 129 5044 311
rect 5076 129 5080 311
rect 5040 60 5080 129
rect -240 -1005 -200 -1000
rect -240 -1035 -235 -1005
rect -205 -1035 -200 -1005
rect -240 -1165 -200 -1035
rect -240 -1195 -235 -1165
rect -205 -1195 -200 -1165
rect -240 -1325 -200 -1195
rect -240 -1355 -235 -1325
rect -205 -1355 -200 -1325
rect -240 -1360 -200 -1355
rect -160 -1005 -120 -1000
rect -160 -1035 -155 -1005
rect -125 -1035 -120 -1005
rect -160 -1165 -120 -1035
rect -160 -1195 -155 -1165
rect -125 -1195 -120 -1165
rect -160 -1325 -120 -1195
rect -160 -1355 -155 -1325
rect -125 -1355 -120 -1325
rect -160 -1360 -120 -1355
rect -80 -1005 -40 -1000
rect -80 -1035 -75 -1005
rect -45 -1035 -40 -1005
rect -80 -1165 -40 -1035
rect -80 -1195 -75 -1165
rect -45 -1195 -40 -1165
rect -80 -1325 -40 -1195
rect -80 -1349 -75 -1325
rect -45 -1349 -40 -1325
rect -80 -1431 -76 -1349
rect -44 -1431 -40 -1349
rect 0 -1005 40 -1000
rect 0 -1035 5 -1005
rect 35 -1035 40 -1005
rect 0 -1165 40 -1035
rect 0 -1195 5 -1165
rect 35 -1195 40 -1165
rect 0 -1325 40 -1195
rect 0 -1355 5 -1325
rect 35 -1355 40 -1325
rect 0 -1360 40 -1355
rect 80 -1005 120 -1000
rect 80 -1035 85 -1005
rect 115 -1035 120 -1005
rect 80 -1165 120 -1035
rect 80 -1195 85 -1165
rect 115 -1195 120 -1165
rect 80 -1325 120 -1195
rect 80 -1355 85 -1325
rect 115 -1355 120 -1325
rect 80 -1360 120 -1355
rect 160 -1005 200 -1000
rect 160 -1035 165 -1005
rect 195 -1035 200 -1005
rect 160 -1165 200 -1035
rect 160 -1195 165 -1165
rect 195 -1195 200 -1165
rect 160 -1325 200 -1195
rect 160 -1355 165 -1325
rect 195 -1355 200 -1325
rect 160 -1360 200 -1355
rect 240 -1005 280 -1000
rect 240 -1035 245 -1005
rect 275 -1035 280 -1005
rect 240 -1165 280 -1035
rect 240 -1195 245 -1165
rect 275 -1195 280 -1165
rect 240 -1325 280 -1195
rect 240 -1355 245 -1325
rect 275 -1355 280 -1325
rect 240 -1360 280 -1355
rect 320 -1005 360 -1000
rect 320 -1035 325 -1005
rect 355 -1035 360 -1005
rect 320 -1165 360 -1035
rect 320 -1195 325 -1165
rect 355 -1195 360 -1165
rect 320 -1325 360 -1195
rect 320 -1355 325 -1325
rect 355 -1355 360 -1325
rect 320 -1360 360 -1355
rect 400 -1005 440 -1000
rect 400 -1035 405 -1005
rect 435 -1035 440 -1005
rect 400 -1165 440 -1035
rect 400 -1195 405 -1165
rect 435 -1195 440 -1165
rect 400 -1325 440 -1195
rect 400 -1355 405 -1325
rect 435 -1355 440 -1325
rect 400 -1360 440 -1355
rect 480 -1005 520 -1000
rect 480 -1035 485 -1005
rect 515 -1035 520 -1005
rect 480 -1165 520 -1035
rect 480 -1195 485 -1165
rect 515 -1195 520 -1165
rect 480 -1325 520 -1195
rect 560 -1005 600 -1000
rect 560 -1035 565 -1005
rect 595 -1035 600 -1005
rect 560 -1165 600 -1035
rect 560 -1195 565 -1165
rect 595 -1195 600 -1165
rect 560 -1200 600 -1195
rect 640 -1005 680 -1000
rect 640 -1035 645 -1005
rect 675 -1035 680 -1005
rect 640 -1165 680 -1035
rect 640 -1195 645 -1165
rect 675 -1195 680 -1165
rect 480 -1355 485 -1325
rect 515 -1355 520 -1325
rect 480 -1360 520 -1355
rect 640 -1325 680 -1195
rect 640 -1355 645 -1325
rect 675 -1355 680 -1325
rect 640 -1360 680 -1355
rect 720 -1005 760 -1000
rect 720 -1035 725 -1005
rect 755 -1035 760 -1005
rect 720 -1165 760 -1035
rect 720 -1195 725 -1165
rect 755 -1195 760 -1165
rect 720 -1325 760 -1195
rect 720 -1355 725 -1325
rect 755 -1355 760 -1325
rect 720 -1360 760 -1355
rect 800 -1005 840 -1000
rect 800 -1035 805 -1005
rect 835 -1035 840 -1005
rect 800 -1165 840 -1035
rect 800 -1195 805 -1165
rect 835 -1195 840 -1165
rect 800 -1325 840 -1195
rect 800 -1355 805 -1325
rect 835 -1355 840 -1325
rect 800 -1360 840 -1355
rect 880 -1005 920 -1000
rect 880 -1035 885 -1005
rect 915 -1035 920 -1005
rect 880 -1165 920 -1035
rect 880 -1195 885 -1165
rect 915 -1195 920 -1165
rect 880 -1325 920 -1195
rect 880 -1355 885 -1325
rect 915 -1355 920 -1325
rect 880 -1360 920 -1355
rect 960 -1005 1000 -1000
rect 960 -1035 965 -1005
rect 995 -1035 1000 -1005
rect 960 -1165 1000 -1035
rect 960 -1195 965 -1165
rect 995 -1195 1000 -1165
rect 960 -1325 1000 -1195
rect 960 -1355 965 -1325
rect 995 -1355 1000 -1325
rect 960 -1360 1000 -1355
rect 1040 -1005 1080 -1000
rect 1040 -1035 1045 -1005
rect 1075 -1035 1080 -1005
rect 1040 -1165 1080 -1035
rect 1040 -1195 1045 -1165
rect 1075 -1195 1080 -1165
rect 1040 -1325 1080 -1195
rect 1040 -1355 1045 -1325
rect 1075 -1355 1080 -1325
rect 1040 -1360 1080 -1355
rect 1120 -1005 1160 -1000
rect 1120 -1035 1125 -1005
rect 1155 -1035 1160 -1005
rect 1120 -1165 1160 -1035
rect 1120 -1195 1125 -1165
rect 1155 -1195 1160 -1165
rect 1120 -1325 1160 -1195
rect 1200 -1005 1240 -1000
rect 1200 -1035 1205 -1005
rect 1235 -1035 1240 -1005
rect 1200 -1165 1240 -1035
rect 1200 -1195 1205 -1165
rect 1235 -1195 1240 -1165
rect 1200 -1200 1240 -1195
rect 1280 -1005 1320 -1000
rect 1280 -1035 1285 -1005
rect 1315 -1035 1320 -1005
rect 1280 -1165 1320 -1035
rect 1280 -1195 1285 -1165
rect 1315 -1195 1320 -1165
rect 1120 -1355 1125 -1325
rect 1155 -1355 1160 -1325
rect 1120 -1360 1160 -1355
rect 1200 -1325 1240 -1320
rect 1200 -1349 1205 -1325
rect 1235 -1349 1240 -1325
rect -80 -1440 -40 -1431
rect 1200 -1431 1204 -1349
rect 1236 -1431 1240 -1349
rect 1280 -1325 1320 -1195
rect 1280 -1355 1285 -1325
rect 1315 -1355 1320 -1325
rect 1280 -1360 1320 -1355
rect 1360 -1005 1400 -1000
rect 1360 -1035 1365 -1005
rect 1395 -1035 1400 -1005
rect 1360 -1165 1400 -1035
rect 1360 -1195 1365 -1165
rect 1395 -1195 1400 -1165
rect 1360 -1325 1400 -1195
rect 1360 -1355 1365 -1325
rect 1395 -1355 1400 -1325
rect 1360 -1360 1400 -1355
rect 1440 -1005 1480 -1000
rect 1440 -1035 1445 -1005
rect 1475 -1035 1480 -1005
rect 1440 -1165 1480 -1035
rect 1440 -1195 1445 -1165
rect 1475 -1195 1480 -1165
rect 1440 -1325 1480 -1195
rect 1440 -1355 1445 -1325
rect 1475 -1355 1480 -1325
rect 1440 -1360 1480 -1355
rect 1520 -1005 1560 -1000
rect 1520 -1035 1525 -1005
rect 1555 -1035 1560 -1005
rect 1520 -1165 1560 -1035
rect 1520 -1195 1525 -1165
rect 1555 -1195 1560 -1165
rect 1520 -1325 1560 -1195
rect 1520 -1355 1525 -1325
rect 1555 -1355 1560 -1325
rect 1520 -1360 1560 -1355
rect 1600 -1005 1640 -1000
rect 1600 -1035 1605 -1005
rect 1635 -1035 1640 -1005
rect 1600 -1165 1640 -1035
rect 1600 -1195 1605 -1165
rect 1635 -1195 1640 -1165
rect 1600 -1325 1640 -1195
rect 1600 -1355 1605 -1325
rect 1635 -1355 1640 -1325
rect 1600 -1360 1640 -1355
rect 1680 -1005 1720 -1000
rect 1680 -1035 1685 -1005
rect 1715 -1035 1720 -1005
rect 1680 -1165 1720 -1035
rect 1680 -1195 1685 -1165
rect 1715 -1195 1720 -1165
rect 1680 -1325 1720 -1195
rect 1680 -1355 1685 -1325
rect 1715 -1355 1720 -1325
rect 1680 -1360 1720 -1355
rect 1760 -1005 1800 -1000
rect 1760 -1035 1765 -1005
rect 1795 -1035 1800 -1005
rect 1760 -1165 1800 -1035
rect 1760 -1195 1765 -1165
rect 1795 -1195 1800 -1165
rect 1760 -1325 1800 -1195
rect 1840 -1005 1880 -1000
rect 1840 -1035 1845 -1005
rect 1875 -1035 1880 -1005
rect 1840 -1165 1880 -1035
rect 1840 -1195 1845 -1165
rect 1875 -1195 1880 -1165
rect 1840 -1200 1880 -1195
rect 1920 -1005 1960 -1000
rect 1920 -1035 1925 -1005
rect 1955 -1035 1960 -1005
rect 1920 -1165 1960 -1035
rect 1920 -1195 1925 -1165
rect 1955 -1195 1960 -1165
rect 1760 -1355 1765 -1325
rect 1795 -1355 1800 -1325
rect 1760 -1360 1800 -1355
rect 1920 -1325 1960 -1195
rect 1920 -1355 1925 -1325
rect 1955 -1355 1960 -1325
rect 1920 -1360 1960 -1355
rect 2000 -1005 2040 -1000
rect 2000 -1035 2005 -1005
rect 2035 -1035 2040 -1005
rect 2000 -1165 2040 -1035
rect 2000 -1195 2005 -1165
rect 2035 -1195 2040 -1165
rect 2000 -1325 2040 -1195
rect 2000 -1355 2005 -1325
rect 2035 -1355 2040 -1325
rect 2000 -1360 2040 -1355
rect 2080 -1005 2120 -1000
rect 2080 -1035 2085 -1005
rect 2115 -1035 2120 -1005
rect 2080 -1165 2120 -1035
rect 2080 -1195 2085 -1165
rect 2115 -1195 2120 -1165
rect 2080 -1325 2120 -1195
rect 2080 -1355 2085 -1325
rect 2115 -1355 2120 -1325
rect 2080 -1360 2120 -1355
rect 2160 -1005 2200 -1000
rect 2160 -1035 2165 -1005
rect 2195 -1035 2200 -1005
rect 2160 -1165 2200 -1035
rect 2160 -1195 2165 -1165
rect 2195 -1195 2200 -1165
rect 2160 -1325 2200 -1195
rect 2160 -1355 2165 -1325
rect 2195 -1355 2200 -1325
rect 2160 -1360 2200 -1355
rect 2240 -1005 2280 -1000
rect 2240 -1035 2245 -1005
rect 2275 -1035 2280 -1005
rect 2240 -1165 2280 -1035
rect 2240 -1195 2245 -1165
rect 2275 -1195 2280 -1165
rect 2240 -1325 2280 -1195
rect 2240 -1355 2245 -1325
rect 2275 -1355 2280 -1325
rect 2240 -1360 2280 -1355
rect 2320 -1005 2360 -1000
rect 2320 -1035 2325 -1005
rect 2355 -1035 2360 -1005
rect 2320 -1165 2360 -1035
rect 2320 -1195 2325 -1165
rect 2355 -1195 2360 -1165
rect 2320 -1325 2360 -1195
rect 2320 -1355 2325 -1325
rect 2355 -1355 2360 -1325
rect 2320 -1360 2360 -1355
rect 2400 -1005 2440 -1000
rect 2400 -1035 2405 -1005
rect 2435 -1035 2440 -1005
rect 2400 -1165 2440 -1035
rect 2400 -1195 2405 -1165
rect 2435 -1195 2440 -1165
rect 2400 -1325 2440 -1195
rect 2480 -1005 2520 -1000
rect 2480 -1035 2485 -1005
rect 2515 -1035 2520 -1005
rect 2480 -1165 2520 -1035
rect 2480 -1195 2485 -1165
rect 2515 -1195 2520 -1165
rect 2480 -1200 2520 -1195
rect 2560 -1005 2600 -1000
rect 2560 -1035 2565 -1005
rect 2595 -1035 2600 -1005
rect 2560 -1165 2600 -1035
rect 2560 -1195 2565 -1165
rect 2595 -1195 2600 -1165
rect 2400 -1355 2405 -1325
rect 2435 -1355 2440 -1325
rect 2400 -1360 2440 -1355
rect 2480 -1325 2520 -1320
rect 2480 -1349 2485 -1325
rect 2515 -1349 2520 -1325
rect 1200 -1440 1240 -1431
rect 2480 -1431 2484 -1349
rect 2516 -1431 2520 -1349
rect 2560 -1325 2600 -1195
rect 2560 -1355 2565 -1325
rect 2595 -1355 2600 -1325
rect 2560 -1360 2600 -1355
rect 2640 -1005 2680 -1000
rect 2640 -1035 2645 -1005
rect 2675 -1035 2680 -1005
rect 2640 -1165 2680 -1035
rect 2640 -1195 2645 -1165
rect 2675 -1195 2680 -1165
rect 2640 -1325 2680 -1195
rect 2640 -1355 2645 -1325
rect 2675 -1355 2680 -1325
rect 2640 -1360 2680 -1355
rect 2720 -1005 2760 -1000
rect 2720 -1035 2725 -1005
rect 2755 -1035 2760 -1005
rect 2720 -1165 2760 -1035
rect 2720 -1195 2725 -1165
rect 2755 -1195 2760 -1165
rect 2720 -1325 2760 -1195
rect 2720 -1355 2725 -1325
rect 2755 -1355 2760 -1325
rect 2720 -1360 2760 -1355
rect 2800 -1005 2840 -1000
rect 2800 -1035 2805 -1005
rect 2835 -1035 2840 -1005
rect 2800 -1165 2840 -1035
rect 2800 -1195 2805 -1165
rect 2835 -1195 2840 -1165
rect 2800 -1325 2840 -1195
rect 2800 -1355 2805 -1325
rect 2835 -1355 2840 -1325
rect 2800 -1360 2840 -1355
rect 2880 -1005 2920 -1000
rect 2880 -1035 2885 -1005
rect 2915 -1035 2920 -1005
rect 2880 -1165 2920 -1035
rect 2880 -1195 2885 -1165
rect 2915 -1195 2920 -1165
rect 2880 -1325 2920 -1195
rect 2880 -1355 2885 -1325
rect 2915 -1355 2920 -1325
rect 2880 -1360 2920 -1355
rect 2960 -1005 3000 -1000
rect 2960 -1035 2965 -1005
rect 2995 -1035 3000 -1005
rect 2960 -1165 3000 -1035
rect 2960 -1195 2965 -1165
rect 2995 -1195 3000 -1165
rect 2960 -1325 3000 -1195
rect 2960 -1355 2965 -1325
rect 2995 -1355 3000 -1325
rect 2960 -1360 3000 -1355
rect 3040 -1005 3080 -1000
rect 3040 -1035 3045 -1005
rect 3075 -1035 3080 -1005
rect 3040 -1165 3080 -1035
rect 3040 -1195 3045 -1165
rect 3075 -1195 3080 -1165
rect 3040 -1325 3080 -1195
rect 3120 -1005 3160 -1000
rect 3120 -1035 3125 -1005
rect 3155 -1035 3160 -1005
rect 3120 -1165 3160 -1035
rect 3120 -1195 3125 -1165
rect 3155 -1195 3160 -1165
rect 3120 -1200 3160 -1195
rect 3200 -1005 3240 -1000
rect 3200 -1035 3205 -1005
rect 3235 -1035 3240 -1005
rect 3200 -1165 3240 -1035
rect 3200 -1195 3205 -1165
rect 3235 -1195 3240 -1165
rect 3040 -1355 3045 -1325
rect 3075 -1355 3080 -1325
rect 3040 -1360 3080 -1355
rect 3200 -1325 3240 -1195
rect 3200 -1355 3205 -1325
rect 3235 -1355 3240 -1325
rect 3200 -1360 3240 -1355
rect 3280 -1005 3320 -1000
rect 3280 -1035 3285 -1005
rect 3315 -1035 3320 -1005
rect 3280 -1165 3320 -1035
rect 3280 -1195 3285 -1165
rect 3315 -1195 3320 -1165
rect 3280 -1325 3320 -1195
rect 3280 -1355 3285 -1325
rect 3315 -1355 3320 -1325
rect 3280 -1360 3320 -1355
rect 3360 -1005 3400 -1000
rect 3360 -1035 3365 -1005
rect 3395 -1035 3400 -1005
rect 3360 -1165 3400 -1035
rect 3360 -1195 3365 -1165
rect 3395 -1195 3400 -1165
rect 3360 -1325 3400 -1195
rect 3360 -1355 3365 -1325
rect 3395 -1355 3400 -1325
rect 3360 -1360 3400 -1355
rect 3440 -1005 3480 -1000
rect 3440 -1035 3445 -1005
rect 3475 -1035 3480 -1005
rect 3440 -1165 3480 -1035
rect 3440 -1195 3445 -1165
rect 3475 -1195 3480 -1165
rect 3440 -1325 3480 -1195
rect 3440 -1355 3445 -1325
rect 3475 -1355 3480 -1325
rect 3440 -1360 3480 -1355
rect 3520 -1005 3560 -1000
rect 3520 -1035 3525 -1005
rect 3555 -1035 3560 -1005
rect 3520 -1165 3560 -1035
rect 3520 -1195 3525 -1165
rect 3555 -1195 3560 -1165
rect 3520 -1325 3560 -1195
rect 3520 -1355 3525 -1325
rect 3555 -1355 3560 -1325
rect 3520 -1360 3560 -1355
rect 3600 -1005 3640 -1000
rect 3600 -1035 3605 -1005
rect 3635 -1035 3640 -1005
rect 3600 -1165 3640 -1035
rect 3600 -1195 3605 -1165
rect 3635 -1195 3640 -1165
rect 3600 -1325 3640 -1195
rect 3600 -1355 3605 -1325
rect 3635 -1355 3640 -1325
rect 3600 -1360 3640 -1355
rect 3680 -1005 3720 -1000
rect 3680 -1035 3685 -1005
rect 3715 -1035 3720 -1005
rect 3680 -1165 3720 -1035
rect 3680 -1195 3685 -1165
rect 3715 -1195 3720 -1165
rect 3680 -1325 3720 -1195
rect 3760 -1005 3800 -1000
rect 3760 -1035 3765 -1005
rect 3795 -1035 3800 -1005
rect 3760 -1165 3800 -1035
rect 3760 -1195 3765 -1165
rect 3795 -1195 3800 -1165
rect 3760 -1200 3800 -1195
rect 3840 -1005 3880 -1000
rect 3840 -1035 3845 -1005
rect 3875 -1035 3880 -1005
rect 3840 -1165 3880 -1035
rect 3840 -1195 3845 -1165
rect 3875 -1195 3880 -1165
rect 3680 -1355 3685 -1325
rect 3715 -1355 3720 -1325
rect 3680 -1360 3720 -1355
rect 3760 -1325 3800 -1320
rect 3760 -1349 3765 -1325
rect 3795 -1349 3800 -1325
rect 2480 -1440 2520 -1431
rect 3760 -1431 3764 -1349
rect 3796 -1431 3800 -1349
rect 3840 -1325 3880 -1195
rect 3840 -1355 3845 -1325
rect 3875 -1355 3880 -1325
rect 3840 -1360 3880 -1355
rect 3920 -1005 3960 -1000
rect 3920 -1035 3925 -1005
rect 3955 -1035 3960 -1005
rect 3920 -1165 3960 -1035
rect 3920 -1195 3925 -1165
rect 3955 -1195 3960 -1165
rect 3920 -1325 3960 -1195
rect 3920 -1355 3925 -1325
rect 3955 -1355 3960 -1325
rect 3920 -1360 3960 -1355
rect 4000 -1005 4040 -1000
rect 4000 -1035 4005 -1005
rect 4035 -1035 4040 -1005
rect 4000 -1165 4040 -1035
rect 4000 -1195 4005 -1165
rect 4035 -1195 4040 -1165
rect 4000 -1325 4040 -1195
rect 4000 -1355 4005 -1325
rect 4035 -1355 4040 -1325
rect 4000 -1360 4040 -1355
rect 4080 -1005 4120 -1000
rect 4080 -1035 4085 -1005
rect 4115 -1035 4120 -1005
rect 4080 -1165 4120 -1035
rect 4080 -1195 4085 -1165
rect 4115 -1195 4120 -1165
rect 4080 -1325 4120 -1195
rect 4080 -1355 4085 -1325
rect 4115 -1355 4120 -1325
rect 4080 -1360 4120 -1355
rect 4160 -1005 4200 -1000
rect 4160 -1035 4165 -1005
rect 4195 -1035 4200 -1005
rect 4160 -1165 4200 -1035
rect 4160 -1195 4165 -1165
rect 4195 -1195 4200 -1165
rect 4160 -1325 4200 -1195
rect 4160 -1355 4165 -1325
rect 4195 -1355 4200 -1325
rect 4160 -1360 4200 -1355
rect 4240 -1005 4280 -1000
rect 4240 -1035 4245 -1005
rect 4275 -1035 4280 -1005
rect 4240 -1165 4280 -1035
rect 4240 -1195 4245 -1165
rect 4275 -1195 4280 -1165
rect 4240 -1325 4280 -1195
rect 4240 -1355 4245 -1325
rect 4275 -1355 4280 -1325
rect 4240 -1360 4280 -1355
rect 4320 -1005 4360 -1000
rect 4320 -1035 4325 -1005
rect 4355 -1035 4360 -1005
rect 4320 -1165 4360 -1035
rect 4320 -1195 4325 -1165
rect 4355 -1195 4360 -1165
rect 4320 -1325 4360 -1195
rect 4400 -1005 4440 -1000
rect 4400 -1035 4405 -1005
rect 4435 -1035 4440 -1005
rect 4400 -1165 4440 -1035
rect 4400 -1195 4405 -1165
rect 4435 -1195 4440 -1165
rect 4400 -1200 4440 -1195
rect 4480 -1005 4520 -1000
rect 4480 -1035 4485 -1005
rect 4515 -1035 4520 -1005
rect 4480 -1165 4520 -1035
rect 4480 -1195 4485 -1165
rect 4515 -1195 4520 -1165
rect 4320 -1355 4325 -1325
rect 4355 -1355 4360 -1325
rect 4320 -1360 4360 -1355
rect 4480 -1325 4520 -1195
rect 4480 -1355 4485 -1325
rect 4515 -1355 4520 -1325
rect 4480 -1360 4520 -1355
rect 4560 -1005 4600 -1000
rect 4560 -1035 4565 -1005
rect 4595 -1035 4600 -1005
rect 4560 -1165 4600 -1035
rect 4560 -1195 4565 -1165
rect 4595 -1195 4600 -1165
rect 4560 -1325 4600 -1195
rect 4560 -1355 4565 -1325
rect 4595 -1355 4600 -1325
rect 4560 -1360 4600 -1355
rect 4640 -1005 4680 -1000
rect 4640 -1035 4645 -1005
rect 4675 -1035 4680 -1005
rect 4640 -1165 4680 -1035
rect 4640 -1195 4645 -1165
rect 4675 -1195 4680 -1165
rect 4640 -1325 4680 -1195
rect 4640 -1355 4645 -1325
rect 4675 -1355 4680 -1325
rect 4640 -1360 4680 -1355
rect 4720 -1005 4760 -1000
rect 4720 -1035 4725 -1005
rect 4755 -1035 4760 -1005
rect 4720 -1165 4760 -1035
rect 4720 -1195 4725 -1165
rect 4755 -1195 4760 -1165
rect 4720 -1325 4760 -1195
rect 4720 -1355 4725 -1325
rect 4755 -1355 4760 -1325
rect 4720 -1360 4760 -1355
rect 4800 -1005 4840 -1000
rect 4800 -1035 4805 -1005
rect 4835 -1035 4840 -1005
rect 4800 -1165 4840 -1035
rect 4800 -1195 4805 -1165
rect 4835 -1195 4840 -1165
rect 4800 -1325 4840 -1195
rect 4800 -1355 4805 -1325
rect 4835 -1355 4840 -1325
rect 4800 -1360 4840 -1355
rect 4880 -1005 4920 -1000
rect 4880 -1035 4885 -1005
rect 4915 -1035 4920 -1005
rect 4880 -1165 4920 -1035
rect 4880 -1195 4885 -1165
rect 4915 -1195 4920 -1165
rect 4880 -1325 4920 -1195
rect 4880 -1355 4885 -1325
rect 4915 -1355 4920 -1325
rect 4880 -1360 4920 -1355
rect 4960 -1005 5000 -1000
rect 4960 -1035 4965 -1005
rect 4995 -1035 5000 -1005
rect 4960 -1165 5000 -1035
rect 4960 -1195 4965 -1165
rect 4995 -1195 5000 -1165
rect 4960 -1325 5000 -1195
rect 4960 -1355 4965 -1325
rect 4995 -1355 5000 -1325
rect 4960 -1360 5000 -1355
rect 5040 -1005 5080 -1000
rect 5040 -1035 5045 -1005
rect 5075 -1035 5080 -1005
rect 5040 -1165 5080 -1035
rect 5040 -1195 5045 -1165
rect 5075 -1195 5080 -1165
rect 5040 -1325 5080 -1195
rect 5040 -1349 5045 -1325
rect 5075 -1349 5080 -1325
rect 3760 -1440 3800 -1431
rect 5040 -1431 5044 -1349
rect 5076 -1431 5080 -1349
rect 5120 -1005 5160 -1000
rect 5120 -1035 5125 -1005
rect 5155 -1035 5160 -1005
rect 5120 -1165 5160 -1035
rect 5120 -1195 5125 -1165
rect 5155 -1195 5160 -1165
rect 5120 -1325 5160 -1195
rect 5120 -1355 5125 -1325
rect 5155 -1355 5160 -1325
rect 5120 -1360 5160 -1355
rect 5200 -1005 5240 -1000
rect 5200 -1035 5205 -1005
rect 5235 -1035 5240 -1005
rect 5200 -1165 5240 -1035
rect 5200 -1195 5205 -1165
rect 5235 -1195 5240 -1165
rect 5200 -1325 5240 -1195
rect 5200 -1355 5205 -1325
rect 5235 -1355 5240 -1325
rect 5200 -1360 5240 -1355
rect 5040 -1440 5080 -1431
<< via3 >>
rect -76 310 -44 311
rect -76 130 -75 310
rect -75 130 -45 310
rect -45 130 -44 310
rect -76 129 -44 130
rect 1204 310 1236 311
rect 1204 130 1205 310
rect 1205 130 1235 310
rect 1235 130 1236 310
rect 1204 129 1236 130
rect 2484 310 2516 311
rect 2484 130 2485 310
rect 2485 130 2515 310
rect 2515 130 2516 310
rect 2484 129 2516 130
rect 3764 310 3796 311
rect 3764 130 3765 310
rect 3765 130 3795 310
rect 3795 130 3796 310
rect 3764 129 3796 130
rect 5044 310 5076 311
rect 5044 130 5045 310
rect 5045 130 5075 310
rect 5075 130 5076 310
rect 5044 129 5076 130
rect -76 -1430 -75 -1349
rect -75 -1430 -45 -1349
rect -45 -1430 -44 -1349
rect -76 -1431 -44 -1430
rect 1204 -1430 1205 -1349
rect 1205 -1430 1235 -1349
rect 1235 -1430 1236 -1349
rect 1204 -1431 1236 -1430
rect 2484 -1430 2485 -1349
rect 2485 -1430 2515 -1349
rect 2515 -1430 2516 -1349
rect 2484 -1431 2516 -1430
rect 3764 -1430 3765 -1349
rect 3765 -1430 3795 -1349
rect 3795 -1430 3796 -1349
rect 3764 -1431 3796 -1430
rect 5044 -1430 5045 -1349
rect 5045 -1430 5075 -1349
rect 5075 -1430 5076 -1349
rect 5044 -1431 5076 -1430
<< metal4 >>
rect -240 311 5080 320
rect -240 280 -76 311
rect -44 280 1204 311
rect 1236 280 2484 311
rect 2516 280 3764 311
rect 3796 280 5044 311
rect 5076 280 5080 311
rect -240 160 -120 280
rect 0 160 1160 280
rect 1280 160 2440 280
rect 2560 160 3720 280
rect 3840 160 5000 280
rect -240 129 -76 160
rect -44 129 1204 160
rect 1236 129 2484 160
rect 2516 129 3764 160
rect 3796 129 5044 160
rect 5076 129 5080 160
rect -240 120 5080 129
rect 5120 120 5240 320
rect -240 -1349 5240 -1320
rect -240 -1431 -76 -1349
rect -44 -1360 1204 -1349
rect -44 -1431 520 -1360
rect -240 -1480 520 -1431
rect 640 -1431 1204 -1360
rect 1236 -1360 2484 -1349
rect 1236 -1431 1800 -1360
rect 640 -1480 1800 -1431
rect 1920 -1431 2484 -1360
rect 2516 -1360 3764 -1349
rect 2516 -1431 3080 -1360
rect 1920 -1480 3080 -1431
rect 3200 -1431 3764 -1360
rect 3796 -1360 5044 -1349
rect 3796 -1431 4360 -1360
rect 3200 -1480 4360 -1431
rect 4480 -1431 5044 -1360
rect 5076 -1431 5240 -1349
rect 4480 -1480 5240 -1431
rect -240 -1520 5240 -1480
<< via4 >>
rect -120 160 -76 280
rect -76 160 -44 280
rect -44 160 0 280
rect 1160 160 1204 280
rect 1204 160 1236 280
rect 1236 160 1280 280
rect 2440 160 2484 280
rect 2484 160 2516 280
rect 2516 160 2560 280
rect 3720 160 3764 280
rect 3764 160 3796 280
rect 3796 160 3840 280
rect 5000 160 5044 280
rect 5044 160 5076 280
rect 5076 160 5120 280
rect 520 -1480 640 -1360
rect 1800 -1480 1920 -1360
rect 3080 -1480 3200 -1360
rect 4360 -1480 4480 -1360
<< metal5 >>
rect -160 280 40 520
rect -160 160 -120 280
rect 0 160 40 280
rect -160 -1520 40 160
rect 480 -1360 680 520
rect 480 -1480 520 -1360
rect 640 -1480 680 -1360
rect 480 -1520 680 -1480
rect 1120 280 1320 520
rect 1120 160 1160 280
rect 1280 160 1320 280
rect 1120 -1520 1320 160
rect 1760 -1360 1960 520
rect 1760 -1480 1800 -1360
rect 1920 -1480 1960 -1360
rect 1760 -1520 1960 -1480
rect 2400 280 2600 520
rect 2400 160 2440 280
rect 2560 160 2600 280
rect 2400 -1520 2600 160
rect 3040 -1360 3240 520
rect 3040 -1480 3080 -1360
rect 3200 -1480 3240 -1360
rect 3040 -1520 3240 -1480
rect 3680 280 3880 520
rect 3680 160 3720 280
rect 3840 160 3880 280
rect 3680 -1520 3880 160
rect 4320 -1360 4520 520
rect 4320 -1480 4360 -1360
rect 4480 -1480 4520 -1360
rect 4320 -1520 4520 -1480
rect 4960 280 5160 520
rect 4960 160 5000 280
rect 5120 160 5160 280
rect 4960 -1520 5160 160
<< labels >>
rlabel locali 2480 0 2520 40 0 xp
rlabel metal2 5200 -400 5240 -360 0 gp
port 0 nsew
rlabel metal2 5200 -720 5240 -680 0 dp
port 1 nsew
rlabel metal2 5200 -800 5240 -760 0 out
port 2 nsew
rlabel metal2 5200 -880 5240 -840 0 dn
port 3 nsew
rlabel metal2 5200 -1120 5240 -1080 0 gn
port 4 nsew
rlabel metal2 5200 -1280 5240 -1240 0 xn
port 5 nsew
rlabel metal5 -160 480 40 520 0 vdda
port 6 nsew
rlabel metal5 480 480 680 520 0 vssa
port 7 nsew
rlabel metal1 240 -1440 280 -1340 0 n1
rlabel metal1 880 -1440 920 -1340 0 n2
rlabel metal1 1520 -1440 1560 -1340 0 n3
rlabel metal1 2160 -1440 2200 -1340 0 n4
rlabel metal1 2800 -1440 2840 -1340 0 n5
rlabel metal1 3440 -1440 3480 -1340 0 n6
rlabel metal1 4080 -1440 4120 -1340 0 n7
rlabel metal1 4720 -1440 4760 -1340 0 n8
rlabel metal1 240 60 280 360 0 p1
rlabel metal1 880 60 920 360 0 p2
rlabel metal1 1520 60 1560 360 0 p3
rlabel metal1 2160 60 2200 360 0 p4
rlabel metal1 2800 60 2840 360 0 p5
rlabel metal1 3440 60 3480 360 0 p6
rlabel metal1 4080 60 4120 360 0 p7
rlabel metal1 4720 60 4760 360 0 p8
<< end >>
