* operational amplifier buffer testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "../mag/opamp.spice"

* supply voltages
vdda vdda 0 1.8
vssa vssa 0 0.0
egnda gnda vssa vdda vssa 0.5

* input signals
vin in gnda dc 0 ac 1 SINE(0 0.9 100 0 0 0)
IB ib vss 10n


* DUT
Xdut out in out ib vdda gnda vssa opamp 
CL out gnda 1p
IL out gnda 0

.save v(in) v(out) v(ib) v(Xdut.x) i(vdda) i(egnda) i(vssa) v(Xdut.b) v(Xdut.c)
.option gmin=1e-15
.control

	op
	print ib i(vdda)
	
	dc il -300u 300u 10u
	plot v(out) v(Xdut.b) v(Xdut.c)
	plot i(vdda) i(gnda) i(vssa)
	
	wrdata ../data/opamp_tb_load_v.txt v(out) v(Xdut.b) v(Xdut.c)
	wrdata ../data/opamp_tb_load_i.txt i(vdda) i(egnda) i(vssa)
	

.endc

.end
