magic
tech sky130A
timestamp 1633696558
<< nwell >>
rect -370 -140 570 2690
<< pmoslvt >>
rect -300 2310 500 2610
rect -300 1980 500 2280
rect -300 1650 500 1950
rect -300 1320 500 1620
rect -300 990 500 1290
rect -300 660 500 960
rect -300 330 500 630
rect -300 0 500 300
<< pdiff >>
rect -350 2600 -300 2610
rect -350 2320 -340 2600
rect -310 2320 -300 2600
rect -350 2310 -300 2320
rect 500 2600 550 2610
rect 500 2320 510 2600
rect 540 2320 550 2600
rect 500 2310 550 2320
rect -350 2270 -300 2280
rect -350 1990 -340 2270
rect -310 1990 -300 2270
rect -350 1980 -300 1990
rect 500 2270 550 2280
rect 500 1990 510 2270
rect 540 1990 550 2270
rect 500 1980 550 1990
rect -350 1940 -300 1950
rect -350 1660 -340 1940
rect -310 1660 -300 1940
rect -350 1650 -300 1660
rect 500 1940 550 1950
rect 500 1660 510 1940
rect 540 1660 550 1940
rect 500 1650 550 1660
rect -350 1610 -300 1620
rect -350 1330 -340 1610
rect -310 1330 -300 1610
rect -350 1320 -300 1330
rect 500 1610 550 1620
rect 500 1330 510 1610
rect 540 1330 550 1610
rect 500 1320 550 1330
rect -350 1280 -300 1290
rect -350 1000 -340 1280
rect -310 1000 -300 1280
rect -350 990 -300 1000
rect 500 1280 550 1290
rect 500 1000 510 1280
rect 540 1000 550 1280
rect 500 990 550 1000
rect -350 950 -300 960
rect -350 670 -340 950
rect -310 670 -300 950
rect -350 660 -300 670
rect 500 950 550 960
rect 500 670 510 950
rect 540 670 550 950
rect 500 660 550 670
rect -350 620 -300 630
rect -350 340 -340 620
rect -310 340 -300 620
rect -350 330 -300 340
rect 500 620 550 630
rect 500 340 510 620
rect 540 340 550 620
rect 500 330 550 340
rect -350 290 -300 300
rect -350 10 -340 290
rect -310 10 -300 290
rect -350 0 -300 10
rect 500 290 550 300
rect 500 10 510 290
rect 540 10 550 290
rect 500 0 550 10
<< pdiffc >>
rect -340 2320 -310 2600
rect 510 2320 540 2600
rect -340 1990 -310 2270
rect 510 1990 540 2270
rect -340 1660 -310 1940
rect 510 1660 540 1940
rect -340 1330 -310 1610
rect 510 1330 540 1610
rect -340 1000 -310 1280
rect 510 1000 540 1280
rect -340 670 -310 950
rect 510 670 540 950
rect -340 340 -310 620
rect 510 340 540 620
rect -340 10 -310 290
rect 510 10 540 290
<< nsubdiff >>
rect -350 2640 -300 2670
rect 500 2640 540 2670
<< nsubdiffcont >>
rect -300 2640 500 2670
<< poly >>
rect -300 2610 500 2630
rect -300 2280 500 2310
rect -300 1950 500 1980
rect -300 1620 500 1650
rect -300 1290 500 1320
rect -300 960 500 990
rect -300 630 500 660
rect -300 300 500 330
rect -300 -30 500 0
rect -300 -60 -280 -30
rect 480 -60 500 -30
rect -300 -70 500 -60
<< polycont >>
rect -280 -60 480 -30
<< locali >>
rect -350 2640 -300 2670
rect 500 2640 540 2670
rect -340 2600 -310 2610
rect -340 2270 -310 2320
rect 510 2600 540 2610
rect 510 2310 540 2320
rect -340 1980 -310 1990
rect 510 2270 540 2280
rect -340 1940 -310 1950
rect -340 1610 -310 1660
rect 510 1940 540 1990
rect 510 1650 540 1660
rect -340 1320 -310 1330
rect 510 1610 540 1620
rect -340 1280 -310 1290
rect -340 950 -310 1000
rect 510 1280 540 1330
rect 510 990 540 1000
rect -340 660 -310 670
rect 510 950 540 960
rect -340 620 -310 630
rect -340 290 -310 340
rect 510 620 540 670
rect 510 330 540 340
rect -340 0 -310 10
rect 510 290 540 300
rect 510 0 540 10
rect -290 -60 -280 -30
rect 480 -60 490 -30
<< viali >>
rect 510 2320 540 2600
rect 510 10 540 290
rect -280 -60 -250 -30
<< metal1 >>
rect 510 2610 540 2690
rect 500 2600 550 2610
rect 500 2320 510 2600
rect 540 2320 550 2600
rect 500 2310 550 2320
rect 500 290 550 300
rect 500 10 510 290
rect 540 10 550 290
rect 500 0 550 10
rect -290 -30 -240 -20
rect -290 -60 -280 -30
rect -250 -60 -240 -30
rect -290 -70 -240 -60
rect -280 -140 -250 -70
rect 510 -140 540 0
<< labels >>
rlabel metal1 520 -110 530 -100 1 D
port 1 n
rlabel metal1 -270 -110 -260 -100 1 G
port 2 n
rlabel metal1 520 2650 530 2660 1 S
port 3 n
rlabel locali -330 2290 -320 2300 1 x1
rlabel locali 520 1960 530 1970 1 x2
rlabel locali -330 1630 -320 1640 1 x3
rlabel locali 520 1300 530 1310 1 x4
rlabel locali -330 970 -320 980 1 x5
rlabel locali 520 640 530 650 1 x6
rlabel locali -330 310 -320 320 1 x7
rlabel locali -330 2650 -320 2660 1 B
port 4 n
<< end >>
