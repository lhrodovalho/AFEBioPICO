**.subckt LNA_TB
X1 net1 MINUS1 OUT IBIAS VSS VDD LNA_OPAMP
XC4 OUT MINUS1 sky130_fd_pr__cap_mim_m3_1 W=22 L=22 MF=1 m=1
XC2 MINUS1 VM sky130_fd_pr__cap_mim_m3_1 W=22 L=22 MF=10 m=10
R2 OUT MINUS1 10E12 m=1
XC1 net1 GND sky130_fd_pr__cap_mim_m3_1 W=22 L=22 MF=1 m=1
XC3 net1 VP sky130_fd_pr__cap_mim_m3_1 W=22 L=22 MF=10 m=10
R1 net1 GND 10E12 m=1
V1 VDD GND 0.9
V4 IN GND AC 1
V3 VSS GND -0.9
I1 IBIAS GND 20n
C5 OUT GND 1p m=1
E1 VP GND IN GND 0.5
E2 VM GND IN GND -.5
**** begin user architecture code


.lib /usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.param mc_mm_switch=0





.option gmin=1E-14

.control

******************OP Simulation*************************************
op
print OUT
print MINUS1
********************************************************************


*******************DC Simulation************************************
*dc V2 0.85 0.95 10u
*plot OUT
*plot deriv(OUT)
********************************************************************


********************AC Simulation***********************************
ac dec 100 0.01 1MEG
plot db(OUT)
********************************************************************


********************Transient Simulation****************************
*tran 1m 2
*plot VP VM OUT
********************************************************************

********************Noise Simulation********************************
*set sqrnoise
noise v(out) V4 dec 100 50m 100
*setplot noise1
*plot log(inoise_spectrum)
*plot onoise_spectrum

print inoise_total
*print onoise_total
********************************************************************
.endc


**** end user architecture code
**.ends

* expanding   symbol:  LNA/LNA_OPAMP.sym # of pins=6
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/LNA/LNA_OPAMP.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/LNA/LNA_OPAMP.sch
.subckt LNA_OPAMP  PLUS MINUS OUT IBIAS VSS VDD
*.iopin VDD
*.iopin VSS
*.iopin PLUS
*.iopin MINUS
*.iopin OUT
*.iopin IBIAS
x9 OUT xp VSS VSS n1_32
x7 VDD net1 net1 VDD p1_32
x8 VDD net1 OUT VDD p1_32
x3 net2 PLUS xp VDD p1_32
x4 net2 MINUS xn VDD p1_32
x5 net1 xn VSS VSS n1_32
x6 xp xp VSS VSS n1_32
x10 xn xn VSS VSS n1_32
x1 IBIAS IBIAS VDD VDD p1_32
x2 net2 IBIAS VDD VDD p1_32
x11 net2 IBIAS VDD VDD p1_32
.ends


* expanding   symbol:  ARRAY/n1_32.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_32.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_32.sch
.subckt n1_32  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_16
xs X G S B n1_16
.ends


* expanding   symbol:  ARRAY/p1_32.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_32.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_32.sch
.subckt p1_32  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_16
xd D G X B p1_16
.ends


* expanding   symbol:  n1_16.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_16.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_16.sch
.subckt n1_16  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_8
xs X G S B n1_8
.ends


* expanding   symbol:  p1_16.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_16.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_16.sch
.subckt p1_16  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_8
xd D G X B p1_8
.ends


* expanding   symbol:  n1_8.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_8.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_8.sch
.subckt n1_8  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_4
xs X G S B n1_4
.ends


* expanding   symbol:  p1_8.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_8.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_8.sch
.subckt p1_8  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_4
xd D G X B p1_4
.ends


* expanding   symbol:  n1_4.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_4.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_4.sch
.subckt n1_4  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_2
xs X G S B n1_2
.ends


* expanding   symbol:  p1_4.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_4.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_4.sch
.subckt p1_4  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_2
xd D G X B p1_2
.ends


* expanding   symbol:  ARRAY/n1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_2.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_2.sch
.subckt n1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xd D G X B n1_1
xs X G S B n1_1
.ends


* expanding   symbol:  ARRAY/p1_2.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_2.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_2.sch
.subckt p1_2  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
xs X G S B p1_1
xd D G X B p1_1
.ends


* expanding   symbol:  n1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_1.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/n1_1.sch
.subckt n1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8_lvt L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
.ends


* expanding   symbol:  p1_1.sym # of pins=4
* sym_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_1.sym
* sch_path: /home/rodovalho/git/AFEBioPICO/xschem/ARRAY/p1_1.sch
.subckt p1_1  D  G  S  B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8_lvt L=8 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
.ends

.GLOBAL GND
** flattened .save nodes
.end
