magic
tech sky130A
timestamp 1633734961
<< metal3 >>
rect 9140 6520 11460 6540
rect 9140 6400 10240 6520
rect 10360 6400 11460 6520
rect 9140 6380 11460 6400
rect 9140 6200 11460 6220
rect 9140 5200 10240 6200
rect 10360 5200 11460 6200
rect 9140 5180 11460 5200
rect 9140 5000 11460 5020
rect 9140 4000 10240 5000
rect 10360 4000 11460 5000
rect 9140 3980 11460 4000
rect 9140 3800 11460 3820
rect 9140 2800 10240 3800
rect 10360 2800 11460 3800
rect 9140 2780 11460 2800
rect 9140 2600 11460 2620
rect 9140 1600 10240 2600
rect 10360 1600 11460 2600
rect 9140 1580 11460 1600
rect 9140 1400 11460 1420
rect 9140 400 10240 1400
rect 10360 400 11460 1400
rect 9140 380 11460 400
rect 9140 200 11460 220
rect 9140 -800 10240 200
rect 10360 -800 11460 200
rect 9140 -820 11460 -800
rect 9140 -1000 11460 -980
rect 9140 -2000 10240 -1000
rect 10360 -2000 11460 -1000
rect 9140 -2020 11460 -2000
rect 9140 -2200 11460 -2180
rect 9140 -3200 10240 -2200
rect 10360 -3200 11460 -2200
rect 9140 -3220 11460 -3200
rect 9140 -3400 11460 -3380
rect 9140 -4400 10240 -3400
rect 10360 -4400 11460 -3400
rect 9140 -4420 11460 -4400
rect 9140 -4600 11460 -4580
rect 9140 -4720 10240 -4600
rect 10360 -4720 11460 -4600
rect 9140 -4740 11460 -4720
<< via3 >>
rect 10240 6400 10360 6520
rect 10240 5200 10360 6200
rect 10240 4000 10360 5000
rect 10240 2800 10360 3800
rect 10240 1600 10360 2600
rect 10240 400 10360 1400
rect 10240 -800 10360 200
rect 10240 -2000 10360 -1000
rect 10240 -3200 10360 -2200
rect 10240 -4400 10360 -3400
rect 10240 -4720 10360 -4600
<< mimcap >>
rect 9160 6400 10160 6520
rect 10440 6400 11440 6520
rect 9160 5200 10160 6200
rect 10440 5200 11440 6200
rect 9160 4000 10160 5000
rect 10440 4000 11440 5000
rect 9160 2800 10160 3800
rect 10440 2800 11440 3800
rect 9160 1600 10160 2600
rect 10440 1600 11440 2600
rect 9160 400 10160 1400
rect 10440 400 11440 1400
rect 9160 -800 10160 200
rect 10440 -800 11440 200
rect 9160 -2000 10160 -1000
rect 10440 -2000 11440 -1000
rect 9160 -3200 10160 -2200
rect 10440 -3200 11440 -2200
rect 9160 -4400 10160 -3400
rect 10440 -4400 11440 -3400
rect 9160 -4720 10160 -4600
rect 10440 -4720 11440 -4600
<< metal4 >>
rect 7540 7480 13060 7500
rect 7540 7360 7560 7480
rect 7680 7360 8200 7480
rect 8320 7360 8840 7480
rect 8960 7360 11640 7480
rect 11760 7360 12280 7480
rect 12400 7360 12920 7480
rect 13040 7360 13060 7480
rect 7540 7340 13060 7360
rect 7540 7160 13060 7180
rect 7540 7040 10240 7160
rect 10360 7040 13060 7160
rect 7540 7020 13060 7040
rect 7540 6840 13060 6860
rect 7540 6720 7560 6840
rect 7680 6720 8200 6840
rect 8320 6720 8840 6840
rect 8960 6720 11640 6840
rect 11760 6720 12280 6840
rect 12400 6720 12920 6840
rect 13040 6720 13060 6840
rect 7540 6700 13060 6720
rect 9140 6520 11460 6540
rect 9140 6400 10240 6520
rect 10360 6400 11460 6520
rect 9140 6380 11460 6400
rect 8500 6200 10180 6220
rect 8500 5200 8520 6200
rect 8640 5200 10180 6200
rect 8500 5180 10180 5200
rect 10220 6200 10380 6220
rect 10220 5200 10240 6200
rect 10360 5200 10380 6200
rect 10220 5180 10380 5200
rect 10420 6200 12100 6220
rect 10420 5200 11960 6200
rect 12080 5200 12100 6200
rect 10420 5180 12100 5200
rect 8500 5000 10180 5020
rect 8500 4000 8520 5000
rect 8640 4000 10180 5000
rect 8500 3980 10180 4000
rect 10220 5000 10380 5020
rect 10220 4000 10240 5000
rect 10360 4000 10380 5000
rect 10220 3980 10380 4000
rect 10420 5000 12100 5020
rect 10420 4000 11960 5000
rect 12080 4000 12100 5000
rect 10420 3980 12100 4000
rect 8500 3800 10180 3820
rect 8500 2800 8520 3800
rect 8640 2800 10180 3800
rect 8500 2780 10180 2800
rect 10220 3800 10380 3820
rect 10220 2800 10240 3800
rect 10360 2800 10380 3800
rect 10220 2780 10380 2800
rect 10420 3800 12100 3820
rect 10420 2800 11960 3800
rect 12080 2800 12100 3800
rect 10420 2780 12100 2800
rect 8500 2600 10180 2620
rect 8500 1600 8520 2600
rect 8640 1600 10180 2600
rect 8500 1580 10180 1600
rect 10220 2600 10380 2620
rect 10220 1600 10240 2600
rect 10360 1600 10380 2600
rect 10220 1580 10380 1600
rect 10420 2600 12100 2620
rect 10420 1600 11960 2600
rect 12080 1600 12100 2600
rect 10420 1580 12100 1600
rect 7860 1400 10180 1420
rect 7860 400 7880 1400
rect 8000 400 10180 1400
rect 7860 380 10180 400
rect 10220 1400 10380 1420
rect 10220 400 10240 1400
rect 10360 400 10380 1400
rect 10220 380 10380 400
rect 10420 1400 12740 1420
rect 10420 400 12600 1400
rect 12720 400 12740 1400
rect 10420 380 12740 400
rect 8500 200 10180 220
rect 8500 -800 8520 200
rect 8640 -800 10180 200
rect 8500 -820 10180 -800
rect 10220 200 10380 220
rect 10220 -800 10240 200
rect 10360 -800 10380 200
rect 10220 -820 10380 -800
rect 10420 200 12100 220
rect 10420 -800 11960 200
rect 12080 -800 12100 200
rect 10420 -820 12100 -800
rect 8500 -1000 10180 -980
rect 8500 -2000 8520 -1000
rect 8640 -2000 10180 -1000
rect 8500 -2020 10180 -2000
rect 10220 -1000 10380 -980
rect 10220 -2000 10240 -1000
rect 10360 -2000 10380 -1000
rect 10220 -2020 10380 -2000
rect 10420 -1000 12100 -980
rect 10420 -2000 11960 -1000
rect 12080 -2000 12100 -1000
rect 10420 -2020 12100 -2000
rect 8500 -2200 10180 -2180
rect 8500 -3200 8520 -2200
rect 8640 -3200 10180 -2200
rect 8500 -3220 10180 -3200
rect 10220 -2200 10380 -2180
rect 10220 -3200 10240 -2200
rect 10360 -3200 10380 -2200
rect 10220 -3220 10380 -3200
rect 10420 -2200 12100 -2180
rect 10420 -3200 11960 -2200
rect 12080 -3200 12100 -2200
rect 10420 -3220 12100 -3200
rect 8500 -3400 10180 -3380
rect 8500 -4400 8520 -3400
rect 8640 -4400 10180 -3400
rect 8500 -4420 10180 -4400
rect 10220 -3400 10380 -3380
rect 10220 -4400 10240 -3400
rect 10360 -4400 10380 -3400
rect 10220 -4420 10380 -4400
rect 10420 -3400 12100 -3380
rect 10420 -4400 11960 -3400
rect 12080 -4400 12100 -3400
rect 10420 -4420 12100 -4400
rect 9140 -4600 11460 -4580
rect 9140 -4720 10240 -4600
rect 10360 -4720 11460 -4600
rect 9140 -4740 11460 -4720
rect 7540 -4920 13060 -4900
rect 7540 -5040 7560 -4920
rect 7680 -5040 8200 -4920
rect 8320 -5040 8840 -4920
rect 8960 -5040 11640 -4920
rect 11760 -5040 12280 -4920
rect 12400 -5040 12920 -4920
rect 13040 -5040 13060 -4920
rect 7540 -5060 13060 -5040
rect 7540 -5240 10220 -5220
rect 7540 -5360 8520 -5240
rect 8640 -5360 10220 -5240
rect 7540 -5380 10220 -5360
rect 10380 -5240 13060 -5220
rect 10380 -5360 11960 -5240
rect 12080 -5360 13060 -5240
rect 10380 -5380 13060 -5360
rect 7540 -5560 13060 -5540
rect 7540 -5680 7560 -5560
rect 7680 -5680 8200 -5560
rect 8320 -5680 8840 -5560
rect 8960 -5680 11640 -5560
rect 11760 -5680 12280 -5560
rect 12400 -5680 12920 -5560
rect 13040 -5680 13060 -5560
rect 7540 -5700 13060 -5680
rect 7540 -5880 10220 -5860
rect 7540 -6000 7880 -5880
rect 8000 -6000 10220 -5880
rect 7540 -6020 10220 -6000
rect 10380 -5880 13060 -5860
rect 10380 -6000 12600 -5880
rect 12720 -6000 13060 -5880
rect 10380 -6020 13060 -6000
rect 7540 -6200 13060 -6180
rect 7540 -6320 7560 -6200
rect 7680 -6320 8200 -6200
rect 8320 -6320 8840 -6200
rect 8960 -6320 11640 -6200
rect 11760 -6320 12280 -6200
rect 12400 -6320 12920 -6200
rect 13040 -6320 13060 -6200
rect 7540 -6340 13060 -6320
<< via4 >>
rect 7560 7360 7680 7480
rect 8200 7360 8320 7480
rect 8840 7360 8960 7480
rect 11640 7360 11760 7480
rect 12280 7360 12400 7480
rect 12920 7360 13040 7480
rect 10240 7040 10360 7160
rect 7560 6720 7680 6840
rect 8200 6720 8320 6840
rect 8840 6720 8960 6840
rect 11640 6720 11760 6840
rect 12280 6720 12400 6840
rect 12920 6720 13040 6840
rect 10240 6400 10360 6520
rect 8520 5200 8640 6200
rect 10240 5200 10360 6200
rect 11960 5200 12080 6200
rect 8520 4000 8640 5000
rect 10240 4000 10360 5000
rect 11960 4000 12080 5000
rect 8520 2800 8640 3800
rect 10240 2800 10360 3800
rect 11960 2800 12080 3800
rect 8520 1600 8640 2600
rect 10240 1600 10360 2600
rect 11960 1600 12080 2600
rect 7880 400 8000 1400
rect 10240 400 10360 1400
rect 12600 400 12720 1400
rect 8520 -800 8640 200
rect 10240 -800 10360 200
rect 11960 -800 12080 200
rect 8520 -2000 8640 -1000
rect 10240 -2000 10360 -1000
rect 11960 -2000 12080 -1000
rect 8520 -3200 8640 -2200
rect 10240 -3200 10360 -2200
rect 11960 -3200 12080 -2200
rect 8520 -4400 8640 -3400
rect 10240 -4400 10360 -3400
rect 11960 -4400 12080 -3400
rect 10240 -4720 10360 -4600
rect 7560 -5040 7680 -4920
rect 8200 -5040 8320 -4920
rect 8840 -5040 8960 -4920
rect 11640 -5040 11760 -4920
rect 12280 -5040 12400 -4920
rect 12920 -5040 13040 -4920
rect 8520 -5360 8640 -5240
rect 11960 -5360 12080 -5240
rect 7560 -5680 7680 -5560
rect 8200 -5680 8320 -5560
rect 8840 -5680 8960 -5560
rect 11640 -5680 11760 -5560
rect 12280 -5680 12400 -5560
rect 12920 -5680 13040 -5560
rect 7880 -6000 8000 -5880
rect 12600 -6000 12720 -5880
rect 7560 -6320 7680 -6200
rect 8200 -6320 8320 -6200
rect 8840 -6320 8960 -6200
rect 11640 -6320 11760 -6200
rect 12280 -6320 12400 -6200
rect 12920 -6320 13040 -6200
<< mimcap2 >>
rect 9160 6400 10160 6520
rect 10440 6400 11440 6520
rect 9160 6190 10160 6200
rect 9160 5210 9170 6190
rect 10150 5210 10160 6190
rect 9160 5200 10160 5210
rect 10440 6190 11440 6200
rect 10440 5210 10450 6190
rect 11430 5210 11440 6190
rect 10440 5200 11440 5210
rect 9160 4990 10160 5000
rect 9160 4010 9170 4990
rect 10150 4010 10160 4990
rect 9160 4000 10160 4010
rect 10440 4990 11440 5000
rect 10440 4010 10450 4990
rect 11430 4010 11440 4990
rect 10440 4000 11440 4010
rect 9160 3790 10160 3800
rect 9160 2810 9170 3790
rect 10150 2810 10160 3790
rect 9160 2800 10160 2810
rect 10440 3790 11440 3800
rect 10440 2810 10450 3790
rect 11430 2810 11440 3790
rect 10440 2800 11440 2810
rect 9160 2590 10160 2600
rect 9160 1610 9170 2590
rect 10150 1610 10160 2590
rect 9160 1600 10160 1610
rect 10440 2590 11440 2600
rect 10440 1610 10450 2590
rect 11430 1610 11440 2590
rect 10440 1600 11440 1610
rect 9160 1390 10160 1400
rect 9160 410 9170 1390
rect 10150 410 10160 1390
rect 9160 400 10160 410
rect 10440 1390 11440 1400
rect 10440 410 10450 1390
rect 11430 410 11440 1390
rect 10440 400 11440 410
rect 9160 190 10160 200
rect 9160 -790 9170 190
rect 10150 -790 10160 190
rect 9160 -800 10160 -790
rect 10440 190 11440 200
rect 10440 -790 10450 190
rect 11430 -790 11440 190
rect 10440 -800 11440 -790
rect 9160 -1010 10160 -1000
rect 9160 -1990 9170 -1010
rect 10150 -1990 10160 -1010
rect 9160 -2000 10160 -1990
rect 10440 -1010 11440 -1000
rect 10440 -1990 10450 -1010
rect 11430 -1990 11440 -1010
rect 10440 -2000 11440 -1990
rect 9160 -2210 10160 -2200
rect 9160 -3190 9170 -2210
rect 10150 -3190 10160 -2210
rect 9160 -3200 10160 -3190
rect 10440 -2210 11440 -2200
rect 10440 -3190 10450 -2210
rect 11430 -3190 11440 -2210
rect 10440 -3200 11440 -3190
rect 9160 -3410 10160 -3400
rect 9160 -4390 9170 -3410
rect 10150 -4390 10160 -3410
rect 9160 -4400 10160 -4390
rect 10440 -3410 11440 -3400
rect 10440 -4390 10450 -3410
rect 11430 -4390 11440 -3410
rect 10440 -4400 11440 -4390
rect 9160 -4720 10160 -4600
rect 10440 -4720 11440 -4600
<< mimcap2contact >>
rect 9170 5210 10150 6190
rect 10450 5210 11430 6190
rect 9170 4010 10150 4990
rect 10450 4010 11430 4990
rect 9170 2810 10150 3790
rect 10450 2810 11430 3790
rect 9170 1610 10150 2590
rect 10450 1610 11430 2590
rect 9170 410 10150 1390
rect 10450 410 11430 1390
rect 9170 -790 10150 190
rect 10450 -790 11430 190
rect 9170 -1990 10150 -1010
rect 10450 -1990 11430 -1010
rect 9170 -3190 10150 -2210
rect 10450 -3190 11430 -2210
rect 9170 -4390 10150 -3410
rect 10450 -4390 11430 -3410
<< metal5 >>
rect 7540 7480 7700 7500
rect 7540 7360 7560 7480
rect 7680 7360 7700 7480
rect 7540 6840 7700 7360
rect 7540 6720 7560 6840
rect 7680 6720 7700 6840
rect 7540 -4920 7700 6720
rect 8180 7480 8340 7500
rect 8180 7360 8200 7480
rect 8320 7360 8340 7480
rect 8180 6840 8340 7360
rect 8180 6720 8200 6840
rect 8320 6720 8340 6840
rect 7540 -5040 7560 -4920
rect 7680 -5040 7700 -4920
rect 7540 -5560 7700 -5040
rect 7540 -5680 7560 -5560
rect 7680 -5680 7700 -5560
rect 7540 -6200 7700 -5680
rect 7540 -6320 7560 -6200
rect 7680 -6320 7700 -6200
rect 7540 -6340 7700 -6320
rect 7860 1400 8020 6710
rect 7860 400 7880 1400
rect 8000 400 8020 1400
rect 7860 -5880 8020 400
rect 7860 -6000 7880 -5880
rect 8000 -6000 8020 -5880
rect 7860 -6340 8020 -6000
rect 8180 -4920 8340 6720
rect 8180 -5040 8200 -4920
rect 8320 -5040 8340 -4920
rect 8180 -5560 8340 -5040
rect 8180 -5680 8200 -5560
rect 8320 -5680 8340 -5560
rect 8180 -6200 8340 -5680
rect 8180 -6320 8200 -6200
rect 8320 -6320 8340 -6200
rect 8180 -6340 8340 -6320
rect 8500 6200 8660 7500
rect 8500 5200 8520 6200
rect 8640 5200 8660 6200
rect 8500 5000 8660 5200
rect 8500 4000 8520 5000
rect 8640 4000 8660 5000
rect 8500 3800 8660 4000
rect 8500 2800 8520 3800
rect 8640 2800 8660 3800
rect 8500 2600 8660 2800
rect 8500 1600 8520 2600
rect 8640 1600 8660 2600
rect 8500 200 8660 1600
rect 8500 -800 8520 200
rect 8640 -800 8660 200
rect 8500 -1000 8660 -800
rect 8500 -2000 8520 -1000
rect 8640 -2000 8660 -1000
rect 8500 -2200 8660 -2000
rect 8500 -3200 8520 -2200
rect 8640 -3200 8660 -2200
rect 8500 -3400 8660 -3200
rect 8500 -4400 8520 -3400
rect 8640 -4400 8660 -3400
rect 8500 -5240 8660 -4400
rect 8500 -5360 8520 -5240
rect 8640 -5360 8660 -5240
rect 8500 -6340 8660 -5360
rect 8820 7480 8980 7500
rect 8820 7360 8840 7480
rect 8960 7360 8980 7480
rect 8820 6840 8980 7360
rect 8820 6720 8840 6840
rect 8960 6720 8980 6840
rect 8820 -4920 8980 6720
rect 10220 7160 10380 7500
rect 10220 7040 10240 7160
rect 10360 7040 10380 7160
rect 10220 6540 10380 7040
rect 11620 7480 11780 7500
rect 11620 7360 11640 7480
rect 11760 7360 11780 7480
rect 11620 6840 11780 7360
rect 11620 6720 11640 6840
rect 11760 6720 11780 6840
rect 9140 6520 11460 6540
rect 9140 6400 10240 6520
rect 10360 6400 11460 6520
rect 9140 6380 11460 6400
rect 10220 6220 10380 6380
rect 9140 6200 11460 6220
rect 9140 6190 10240 6200
rect 9140 5210 9170 6190
rect 10150 5210 10240 6190
rect 9140 5200 10240 5210
rect 10360 6190 11460 6200
rect 10360 5210 10450 6190
rect 11430 5210 11460 6190
rect 10360 5200 11460 5210
rect 9140 5180 11460 5200
rect 10220 5020 10380 5180
rect 9140 5000 11460 5020
rect 9140 4990 10240 5000
rect 9140 4010 9170 4990
rect 10150 4010 10240 4990
rect 9140 4000 10240 4010
rect 10360 4990 11460 5000
rect 10360 4010 10450 4990
rect 11430 4010 11460 4990
rect 10360 4000 11460 4010
rect 9140 3980 11460 4000
rect 10220 3820 10380 3980
rect 9140 3800 11460 3820
rect 9140 3790 10240 3800
rect 9140 2810 9170 3790
rect 10150 2810 10240 3790
rect 9140 2800 10240 2810
rect 10360 3790 11460 3800
rect 10360 2810 10450 3790
rect 11430 2810 11460 3790
rect 10360 2800 11460 2810
rect 9140 2780 11460 2800
rect 10220 2620 10380 2780
rect 9140 2600 11460 2620
rect 9140 2590 10240 2600
rect 9140 1610 9170 2590
rect 10150 1610 10240 2590
rect 9140 1600 10240 1610
rect 10360 2590 11460 2600
rect 10360 1610 10450 2590
rect 11430 1610 11460 2590
rect 10360 1600 11460 1610
rect 9140 1580 11460 1600
rect 10220 1420 10380 1580
rect 9140 1400 11460 1420
rect 9140 1390 10240 1400
rect 9140 410 9170 1390
rect 10150 410 10240 1390
rect 9140 400 10240 410
rect 10360 1390 11460 1400
rect 10360 410 10450 1390
rect 11430 410 11460 1390
rect 10360 400 11460 410
rect 9140 380 11460 400
rect 10220 220 10380 380
rect 9140 200 11460 220
rect 9140 190 10240 200
rect 9140 -790 9170 190
rect 10150 -790 10240 190
rect 9140 -800 10240 -790
rect 10360 190 11460 200
rect 10360 -790 10450 190
rect 11430 -790 11460 190
rect 10360 -800 11460 -790
rect 9140 -820 11460 -800
rect 10220 -980 10380 -820
rect 9140 -1000 11460 -980
rect 9140 -1010 10240 -1000
rect 9140 -1990 9170 -1010
rect 10150 -1990 10240 -1010
rect 9140 -2000 10240 -1990
rect 10360 -1010 11460 -1000
rect 10360 -1990 10450 -1010
rect 11430 -1990 11460 -1010
rect 10360 -2000 11460 -1990
rect 9140 -2020 11460 -2000
rect 10220 -2180 10380 -2020
rect 9140 -2200 11460 -2180
rect 9140 -2210 10240 -2200
rect 9140 -3190 9170 -2210
rect 10150 -3190 10240 -2210
rect 9140 -3200 10240 -3190
rect 10360 -2210 11460 -2200
rect 10360 -3190 10450 -2210
rect 11430 -3190 11460 -2210
rect 10360 -3200 11460 -3190
rect 9140 -3220 11460 -3200
rect 10220 -3380 10380 -3220
rect 9140 -3400 11460 -3380
rect 9140 -3410 10240 -3400
rect 9140 -4390 9170 -3410
rect 10150 -4390 10240 -3410
rect 9140 -4400 10240 -4390
rect 10360 -3410 11460 -3400
rect 10360 -4390 10450 -3410
rect 11430 -4390 11460 -3410
rect 10360 -4400 11460 -4390
rect 9140 -4420 11460 -4400
rect 10220 -4580 10380 -4420
rect 9140 -4600 11460 -4580
rect 9140 -4720 10240 -4600
rect 10360 -4720 11460 -4600
rect 9140 -4740 11460 -4720
rect 8820 -5040 8840 -4920
rect 8960 -5040 8980 -4920
rect 8820 -5560 8980 -5040
rect 8820 -5680 8840 -5560
rect 8960 -5680 8980 -5560
rect 8820 -6200 8980 -5680
rect 8820 -6320 8840 -6200
rect 8960 -6320 8980 -6200
rect 8820 -6340 8980 -6320
rect 10220 -6340 10380 -4740
rect 11620 -4920 11780 6720
rect 12260 7480 12420 7500
rect 12260 7360 12280 7480
rect 12400 7360 12420 7480
rect 12260 6840 12420 7360
rect 12260 6720 12280 6840
rect 12400 6720 12420 6840
rect 11620 -5040 11640 -4920
rect 11760 -5040 11780 -4920
rect 11620 -5560 11780 -5040
rect 11620 -5680 11640 -5560
rect 11760 -5680 11780 -5560
rect 11620 -6200 11780 -5680
rect 11620 -6320 11640 -6200
rect 11760 -6320 11780 -6200
rect 11620 -6340 11780 -6320
rect 11940 6200 12100 6700
rect 11940 5200 11960 6200
rect 12080 5200 12100 6200
rect 11940 5000 12100 5200
rect 11940 4000 11960 5000
rect 12080 4000 12100 5000
rect 11940 3800 12100 4000
rect 11940 2800 11960 3800
rect 12080 2800 12100 3800
rect 11940 2600 12100 2800
rect 11940 1600 11960 2600
rect 12080 1600 12100 2600
rect 11940 200 12100 1600
rect 11940 -800 11960 200
rect 12080 -800 12100 200
rect 11940 -1000 12100 -800
rect 11940 -2000 11960 -1000
rect 12080 -2000 12100 -1000
rect 11940 -2200 12100 -2000
rect 11940 -3200 11960 -2200
rect 12080 -3200 12100 -2200
rect 11940 -3400 12100 -3200
rect 11940 -4400 11960 -3400
rect 12080 -4400 12100 -3400
rect 11940 -5240 12100 -4400
rect 11940 -5360 11960 -5240
rect 12080 -5360 12100 -5240
rect 11940 -6340 12100 -5360
rect 12260 -4920 12420 6720
rect 12900 7480 13060 7500
rect 12900 7360 12920 7480
rect 13040 7360 13060 7480
rect 12900 6840 13060 7360
rect 12900 6720 12920 6840
rect 13040 6720 13060 6840
rect 12260 -5040 12280 -4920
rect 12400 -5040 12420 -4920
rect 12260 -5560 12420 -5040
rect 12260 -5680 12280 -5560
rect 12400 -5680 12420 -5560
rect 12260 -6200 12420 -5680
rect 12260 -6320 12280 -6200
rect 12400 -6320 12420 -6200
rect 12260 -6340 12420 -6320
rect 12580 1400 12740 6700
rect 12580 400 12600 1400
rect 12720 400 12740 1400
rect 12580 -5880 12740 400
rect 12580 -6000 12600 -5880
rect 12720 -6000 12740 -5880
rect 12580 -6340 12740 -6000
rect 12900 -4920 13060 6720
rect 12900 -5040 12920 -4920
rect 13040 -5040 13060 -4920
rect 12900 -5560 13060 -5040
rect 12900 -5680 12920 -5560
rect 13040 -5680 13060 -5560
rect 12900 -6200 13060 -5680
rect 12900 -6320 12920 -6200
rect 13040 -6320 13060 -6200
rect 12900 -6340 13060 -6320
<< labels >>
rlabel metal5 10220 7340 10380 7500 1 A
port 1 n
rlabel metal5 11940 -6340 12100 -6180 1 B
port 2 n
rlabel metal5 12580 -6340 12740 -6180 1 C
port 3 n
rlabel metal5 12900 -6340 13060 -6180 1 gnd
port 4 n
<< end >>
