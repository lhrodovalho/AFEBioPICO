* lna-ota buffer testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "lna_ota.spice"
.include "pseudo.spice"
.include "pseudo_bias4x.spice"
.include "cap_1_10.spice"
.include "n8_1.spice"

.subckt cap2x_1_10 A B C gnd
	x1 A B C GND cap_1_10
	x2 A B C GND cap_1_10
.ends

.subckt cap4x_1_10 A B C gnd
	x1 A B C GND cap2x_1_10
	x2 A B C GND cap2x_1_10
.ends

.subckt cap8x_1_10 A B C gnd
	x1 A B C GND cap4x_1_10
	x2 A B C GND cap4x_1_10
.ends

.subckt inv0 in out vdda vssa
xp out in vdda vdda vssa p1_8
xn out in vssa vssa n1_8
.ends

.subckt inv in out vdda vssa
xps xp  in vdda vdda vssa p1_8
xpd out in xp   vdda vssa p8_1
xnd out in xn   vssa n8_1
xns xn  in vssa vssa n1_8
.ends


.subckt ota ip im op om vdda vssa
xap ip om vdda vssa inv
xam im op vdda vssa inv
xbp ip om  vdda vssa inv
xbm im op  vdda vssa inv
xcp om om vdda vssa inv
xcm op op vdda vssa inv
xdp op om  vdda vssa inv
xdm om op  vdda vssa inv
.ends

.subckt ota2 ip im op om vdda vssa
xap ip om vdda vssa inv
xam im op vdda vssa inv
xbp om x  vdda vssa inv
xbm op x  vdda vssa inv
xcp x  x  vdda vssa inv
xcm x  x  vdda vssa inv
xd  x  y  vdda vssa inv
xe  y  y  vdda vssa inv
xfp y  om vdda vssa inv
xfm y  op vdda vssa inv
.ends

.subckt load ip im vdda vssa
xap ip x  vdda vssa inv
xam im x  vdda vssa inv
xbp x  x  vdda vssa inv
xbm x  x  vdda vssa inv
xc  x  y  vdda vssa inv
xd  y  y  vdda vssa inv
xep y  ip vdda vssa inv
xem y  im vdda vssa inv
.ends

.subckt load2 ip im vdda vssa
xap ip ip vdda vssa inv
xam im im vdda vssa inv
xep ip im vdda vssa inv
xem im ip vdda vssa inv
.ends


* supply voltages
vdda	vdda 0 1.2
vgnda	gnda 0 0.6
vssa	vssa 0 0.0

* input signals
vin	in gnda dc 0 ac 1 SINE(0 10m 1 0 0 0)
einp	ip gnda in gnda  0.5
einm	im gnda in gnda -0.5

* DUT

.subckt lna ip im op om vdda vssa
xamp xp xm op om vdda vssa ota2
cip im xm 10p
cfp xm op 1p
*rfp xm gnda 1T

egnda gnda vssa vdda vssa 0.5

cim ip xp 10p
cfm xp om 1p
*rfm xp gnda 1T

xload xp xm vdda vssa load2

	.subckt p1_1 D G S B
		X1 D G S B sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=8e+06u
	.ends

.ends

x0 ip im op om vdda vssa lna

eout out gnda op om 1
CL out gnda 10p

.ic v(x0.xp)=0.6
.ic v(x0.xm)=0.6

.option gmin=1e-14
.option scale=1e-6
.control

	op
	
	tran 1m 2 1
	plot in out
    
.endc

.end
