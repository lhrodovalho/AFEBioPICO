magic
tech sky130A
timestamp 1633868591
<< nwell >>
rect 6310 4820 6370 4840
rect 6400 4820 6430 4840
rect 9110 4820 9140 4840
rect 10970 4820 11000 4840
rect 11900 4820 11930 4840
rect 14690 4820 14720 4840
rect 16550 4820 16580 4840
rect 16600 4820 16670 4840
rect 6310 4790 16670 4820
rect 6310 2060 6370 4790
rect 16600 4710 16670 4790
rect 16610 2060 16670 4710
rect 6310 2030 6380 2060
rect 6310 2010 6370 2030
rect 7390 2010 7420 2040
rect 8320 2010 8350 2040
rect 9250 2010 9280 2040
rect 10180 2010 10210 2040
rect 11110 2010 11140 2040
rect 12040 2010 12070 2040
rect 12970 2010 13000 2040
rect 13900 2010 13930 2040
rect 14830 2010 14860 2040
rect 15760 2010 15790 2040
rect 16510 2030 16670 2060
rect 16610 2010 16670 2030
rect 6310 0 6370 20
rect 6310 -30 6470 0
rect 7190 -10 7220 20
rect 8120 -10 8150 20
rect 9050 -10 9080 20
rect 9980 -10 10010 20
rect 10910 -10 10940 20
rect 11840 -10 11870 20
rect 12770 -10 12800 20
rect 13700 -10 13730 20
rect 14630 -10 14660 20
rect 15560 -10 15590 20
rect 16610 0 16670 20
rect 16600 -30 16670 0
rect 6310 -2680 6370 -30
rect 6310 -2760 6380 -2680
rect 16540 -2760 16590 -2750
rect 16610 -2760 16670 -30
rect 6310 -2790 16670 -2760
rect 6310 -2810 6380 -2790
rect 11050 -2810 11080 -2790
rect 11980 -2810 12010 -2790
rect 13840 -2810 13870 -2790
rect 16540 -2800 16590 -2790
rect 16550 -2810 16580 -2800
rect 16610 -2810 16670 -2790
<< psubdiff >>
rect 6260 4860 6310 4890
rect 16670 4860 16720 4890
rect 6260 4840 6290 4860
rect 16690 4840 16720 4860
rect 6260 -2830 6290 -2810
rect 16690 -2830 16720 -2810
rect 6260 -2860 6310 -2830
rect 16670 -2860 16720 -2830
<< nsubdiff >>
rect 6330 4790 16650 4820
rect 6330 4770 6360 4790
rect 6330 2060 6360 2080
rect 16620 4770 16650 4790
rect 16620 2060 16650 2080
rect 6330 2030 6380 2060
rect 16510 2030 16650 2060
rect 6330 -30 6470 0
rect 16600 -30 16650 0
rect 6330 -50 6360 -30
rect 6330 -2760 6360 -2740
rect 16620 -50 16650 -30
rect 16620 -2760 16650 -2740
rect 6330 -2790 16650 -2760
<< psubdiffcont >>
rect 6310 4860 16670 4890
rect 6260 -2810 6290 4840
rect 16690 -2810 16720 4840
rect 6310 -2860 16670 -2830
<< nsubdiffcont >>
rect 6330 2080 6360 4770
rect 16620 2080 16650 4770
rect 6380 2030 16510 2060
rect 6470 -30 16600 0
rect 6330 -2740 6360 -50
rect 16620 -2740 16650 -50
<< locali >>
rect 6260 4860 6310 4890
rect 16670 4860 16720 4890
rect 6260 4840 6290 4860
rect 16690 4840 16720 4860
rect 6330 4790 6400 4820
rect 6430 4790 16650 4820
rect 6330 4770 6360 4790
rect 6330 2060 6360 2080
rect 16620 4770 16650 4790
rect 16620 2060 16650 2080
rect 6330 2030 6380 2060
rect 16510 2030 16650 2060
rect 6330 -30 6470 0
rect 16600 -30 16650 0
rect 6330 -50 6360 -30
rect 6330 -2760 6360 -2740
rect 16620 -50 16650 -30
rect 16620 -2760 16650 -2740
rect 6330 -2790 6400 -2760
rect 6430 -2790 16550 -2760
rect 16580 -2790 16650 -2760
rect 6260 -2830 6290 -2810
rect 16690 -2830 16720 -2810
rect 6260 -2860 6310 -2830
rect 16670 -2860 16720 -2830
<< viali >>
rect 6400 4790 6430 4820
rect 6260 1310 6290 1390
rect 6260 640 6290 720
rect 6400 -2790 6430 -2760
rect 16550 -2790 16580 -2760
<< metal1 >>
rect 6400 4940 6430 4950
rect 6400 4830 6430 4860
rect 7250 4940 7280 4950
rect 6390 4820 6440 4830
rect 6390 4790 6400 4820
rect 6430 4790 6440 4820
rect 7250 4810 7280 4860
rect 9110 4940 9140 4950
rect 6390 4780 6440 4790
rect 6400 2060 6430 4780
rect 6400 1940 6430 2030
rect 6400 1820 6430 1910
rect 6400 1700 6430 1790
rect 6400 1580 6430 1670
rect 6400 1460 6430 1550
rect 6250 1390 6300 1400
rect 6250 1310 6260 1390
rect 6290 1310 6300 1390
rect 6250 1300 6300 1310
rect 6400 1270 6430 1430
rect 6400 1150 6430 1240
rect 6400 1030 6430 1120
rect 6400 910 6430 1000
rect 6400 790 6430 880
rect 6250 720 6300 730
rect 6250 640 6260 720
rect 6290 640 6300 720
rect 6250 630 6300 640
rect 6400 600 6430 760
rect 6400 540 6430 570
rect 6460 2000 6490 2040
rect 6400 480 6430 510
rect 6400 360 6430 450
rect 6400 240 6430 330
rect 6400 120 6430 210
rect 6400 0 6430 90
rect 6460 60 6490 1970
rect 7330 1390 7360 4760
rect 7330 1300 7360 1310
rect 7390 1880 7420 2040
rect 7330 720 7360 730
rect 6460 20 6490 30
rect 7190 60 7220 70
rect 7190 -10 7220 30
rect 6400 -2750 6430 -30
rect 6390 -2760 6440 -2750
rect 6390 -2790 6400 -2760
rect 6430 -2790 6440 -2760
rect 6390 -2800 6440 -2790
rect 6400 -2830 6430 -2800
rect 6400 -2920 6430 -2910
rect 7250 -2830 7280 20
rect 7330 -2790 7360 640
rect 7390 180 7420 1850
rect 8180 1760 8210 4840
rect 9110 4810 9140 4860
rect 10970 4940 11000 4950
rect 10970 4810 11000 4860
rect 11900 4940 11930 4950
rect 11900 4810 11930 4860
rect 12830 4940 12860 4950
rect 12830 4840 12860 4860
rect 14690 4940 14720 4950
rect 14690 4810 14720 4860
rect 15700 4940 15730 4950
rect 8320 2000 8350 2040
rect 8320 1960 8350 1970
rect 8180 1720 8210 1730
rect 9110 1760 9140 2040
rect 7390 140 7420 150
rect 8120 970 8150 980
rect 8120 -90 8150 940
rect 8180 850 8210 860
rect 8180 -10 8210 820
rect 8260 850 8290 860
rect 8260 20 8290 820
rect 9110 300 9140 1730
rect 9190 1390 9220 2040
rect 9190 1300 9220 1310
rect 9250 1640 9280 2040
rect 9110 260 9140 270
rect 9190 720 9220 730
rect 9050 60 9080 70
rect 9050 -40 9080 30
rect 9190 -2730 9220 640
rect 9250 420 9280 1610
rect 10040 1520 10070 2150
rect 10180 2000 10210 2040
rect 10180 1960 10210 1970
rect 10040 1480 10070 1490
rect 10970 1520 11000 2010
rect 11050 2000 11080 2010
rect 11050 1960 11080 1970
rect 11110 2000 11140 2040
rect 11110 1960 11140 1970
rect 12040 2000 12070 2040
rect 12040 1960 12070 1970
rect 9250 380 9280 390
rect 9980 1210 10010 1220
rect 9980 -10 10010 1180
rect 10040 1090 10070 1100
rect 10040 20 10070 1060
rect 10120 1090 10150 1100
rect 10120 -10 10150 1060
rect 10970 540 11000 1490
rect 12830 1090 12860 2040
rect 12830 1050 12860 1060
rect 12910 1090 12940 2010
rect 12970 1210 13000 2040
rect 13760 1390 13790 2150
rect 13900 2000 13930 2040
rect 13900 1960 13930 1970
rect 13760 1300 13790 1310
rect 12970 1170 13000 1180
rect 12910 1050 12940 1060
rect 14690 850 14720 2010
rect 14690 810 14720 820
rect 14770 850 14800 2040
rect 14830 970 14860 2120
rect 15620 1400 15650 4820
rect 15700 4750 15730 4860
rect 16550 4940 16580 4950
rect 15760 2000 15790 2040
rect 15760 1960 15790 1970
rect 15620 1290 15650 1300
rect 14830 930 14860 940
rect 14770 810 14800 820
rect 13760 720 13790 730
rect 10970 500 11000 510
rect 11980 540 12010 550
rect 10910 60 10940 70
rect 10910 -10 10940 30
rect 11840 60 11870 70
rect 11840 -10 11870 30
rect 11900 60 11930 70
rect 11900 20 11930 30
rect 11980 20 12010 510
rect 12910 540 12940 550
rect 12770 60 12800 70
rect 12770 -10 12800 30
rect 12910 -120 12940 510
rect 13700 420 13730 430
rect 13700 -10 13730 390
rect 13760 20 13790 640
rect 15620 720 15650 730
rect 13840 300 13870 310
rect 13840 20 13870 270
rect 14770 300 14800 310
rect 14630 60 14660 70
rect 14630 -10 14660 30
rect 7250 -2920 7280 -2910
rect 8260 -2830 8290 -2750
rect 8260 -2920 8290 -2910
rect 10120 -2830 10150 -2730
rect 10120 -2920 10150 -2910
rect 11050 -2830 11080 -2780
rect 11050 -2920 11080 -2910
rect 11980 -2830 12010 -2780
rect 11980 -2920 12010 -2910
rect 13840 -2830 13870 -2780
rect 14770 -2810 14800 270
rect 15560 180 15590 190
rect 15560 -10 15590 150
rect 15620 20 15650 640
rect 16490 60 16520 70
rect 16490 -10 16520 30
rect 16550 -2750 16580 4860
rect 16540 -2760 16590 -2750
rect 13840 -2920 13870 -2910
rect 15700 -2830 15730 -2780
rect 16540 -2790 16550 -2760
rect 16580 -2790 16590 -2760
rect 16540 -2800 16590 -2790
rect 15700 -2920 15730 -2910
rect 16550 -2830 16580 -2800
rect 16550 -2920 16580 -2910
<< via1 >>
rect 6400 4860 6430 4940
rect 7250 4860 7280 4940
rect 9110 4860 9140 4940
rect 6400 2030 6430 2060
rect 6400 1910 6430 1940
rect 6400 1790 6430 1820
rect 6400 1670 6430 1700
rect 6400 1550 6430 1580
rect 6400 1430 6430 1460
rect 6260 1310 6290 1390
rect 6400 1240 6430 1270
rect 6400 1120 6430 1150
rect 6400 1000 6430 1030
rect 6400 880 6430 910
rect 6400 760 6430 790
rect 6260 640 6290 720
rect 6400 570 6430 600
rect 6460 1970 6490 2000
rect 6400 450 6430 480
rect 6400 330 6430 360
rect 6400 210 6430 240
rect 6400 90 6430 120
rect 7330 1310 7360 1390
rect 7390 1850 7420 1880
rect 7330 640 7360 720
rect 6460 30 6490 60
rect 7190 30 7220 60
rect 6400 -30 6430 0
rect 6400 -2910 6430 -2830
rect 10970 4860 11000 4940
rect 11900 4860 11930 4940
rect 12830 4860 12860 4940
rect 14690 4860 14720 4940
rect 15700 4860 15730 4940
rect 8320 1970 8350 2000
rect 8180 1730 8210 1760
rect 9110 1730 9140 1760
rect 7390 150 7420 180
rect 8120 940 8150 970
rect 8180 820 8210 850
rect 8260 820 8290 850
rect 9190 1310 9220 1390
rect 9250 1610 9280 1640
rect 9110 270 9140 300
rect 9190 640 9220 720
rect 9050 30 9080 60
rect 10180 1970 10210 2000
rect 10040 1490 10070 1520
rect 11050 1970 11080 2000
rect 11110 1970 11140 2000
rect 12040 1970 12070 2000
rect 10970 1490 11000 1520
rect 9250 390 9280 420
rect 9980 1180 10010 1210
rect 10040 1060 10070 1090
rect 10120 1060 10150 1090
rect 12830 1060 12860 1090
rect 13900 1970 13930 2000
rect 13760 1310 13790 1390
rect 12970 1180 13000 1210
rect 12910 1060 12940 1090
rect 14690 820 14720 850
rect 16550 4860 16580 4940
rect 15760 1970 15790 2000
rect 15620 1300 15650 1400
rect 14830 940 14860 970
rect 14770 820 14800 850
rect 13760 640 13790 720
rect 10970 510 11000 540
rect 11980 510 12010 540
rect 10910 30 10940 60
rect 11840 30 11870 60
rect 11900 30 11930 60
rect 12910 510 12940 540
rect 12770 30 12800 60
rect 13700 390 13730 420
rect 15620 640 15650 720
rect 13840 270 13870 300
rect 14770 270 14800 300
rect 14630 30 14660 60
rect 7250 -2910 7280 -2830
rect 8260 -2910 8290 -2830
rect 10120 -2910 10150 -2830
rect 11050 -2910 11080 -2830
rect 11980 -2910 12010 -2830
rect 15560 150 15590 180
rect 16490 30 16520 60
rect 13840 -2910 13870 -2830
rect 15700 -2910 15730 -2830
rect 16550 -2910 16580 -2830
<< metal2 >>
rect 6250 4940 16730 4950
rect 6250 4860 6400 4940
rect 6430 4860 7250 4940
rect 7280 4860 9110 4940
rect 9140 4860 10970 4940
rect 11000 4860 11900 4940
rect 11930 4860 12830 4940
rect 12860 4860 14690 4940
rect 14720 4860 15700 4940
rect 15730 4860 16550 4940
rect 16580 4860 16730 4940
rect 6250 4850 16730 4860
rect 6250 2030 6400 2060
rect 6430 2030 16510 2060
rect 6250 1970 6460 2000
rect 6490 1970 8320 2000
rect 8350 1970 10180 2000
rect 10210 1970 11050 2000
rect 11080 1970 11110 2000
rect 11140 1970 12040 2000
rect 12070 1970 13900 2000
rect 13930 1970 15760 2000
rect 15790 1970 16720 2000
rect 6260 1910 6400 1940
rect 6430 1910 16720 1940
rect 6250 1850 7390 1880
rect 7420 1850 16720 1880
rect 6260 1790 6400 1820
rect 6430 1790 16720 1820
rect 6250 1730 8180 1760
rect 8210 1730 9110 1760
rect 9140 1730 16720 1760
rect 6260 1670 6400 1700
rect 6430 1670 16720 1700
rect 6250 1610 9250 1640
rect 9280 1610 16720 1640
rect 6260 1550 6400 1580
rect 6430 1550 16720 1580
rect 6250 1490 10040 1520
rect 10070 1490 10970 1520
rect 11000 1490 16720 1520
rect 6260 1430 6400 1460
rect 6430 1430 16730 1460
rect 6250 1390 15620 1400
rect 6250 1310 6260 1390
rect 6290 1310 7330 1390
rect 7360 1310 9190 1390
rect 9220 1310 13760 1390
rect 13790 1310 15620 1390
rect 6250 1300 15620 1310
rect 15650 1300 16730 1400
rect 6260 1240 6400 1270
rect 6430 1240 16730 1270
rect 6250 1180 9980 1210
rect 10010 1180 12970 1210
rect 13000 1180 16730 1210
rect 6260 1120 6400 1150
rect 6430 1120 16730 1150
rect 6250 1060 10040 1090
rect 10070 1060 10120 1090
rect 10150 1060 12830 1090
rect 12860 1060 12910 1090
rect 12940 1060 16730 1090
rect 6260 1000 6400 1030
rect 6430 1000 16730 1030
rect 6250 940 8120 970
rect 8150 940 14830 970
rect 14860 940 16730 970
rect 6260 880 6400 910
rect 6430 880 16730 910
rect 6250 820 8180 850
rect 8210 820 8260 850
rect 8290 820 14690 850
rect 14720 820 14770 850
rect 14800 820 16730 850
rect 6260 760 6400 790
rect 6430 760 16730 790
rect 6250 720 16730 730
rect 6250 640 6260 720
rect 6290 640 7330 720
rect 7360 640 9190 720
rect 9220 640 13760 720
rect 13790 640 15620 720
rect 15650 640 16730 720
rect 6250 630 16730 640
rect 6260 570 6400 600
rect 6430 570 16730 600
rect 6260 510 10970 540
rect 11000 510 11980 540
rect 12010 510 12910 540
rect 12940 510 16730 540
rect 6260 450 6400 480
rect 6430 450 16730 480
rect 6260 390 9250 420
rect 9280 390 13700 420
rect 13730 390 16730 420
rect 6260 330 6400 360
rect 6430 330 16730 360
rect 6260 270 9110 300
rect 9140 270 13840 300
rect 13870 270 14770 300
rect 14800 270 16730 300
rect 6260 210 6400 240
rect 6430 210 16730 240
rect 6260 150 7390 180
rect 7420 150 15560 180
rect 15590 150 16730 180
rect 6260 90 6400 120
rect 6430 90 16730 120
rect 6260 30 6460 60
rect 6490 30 7190 60
rect 7220 30 9050 60
rect 9080 30 10910 60
rect 10940 30 11840 60
rect 11870 30 11900 60
rect 11930 30 12770 60
rect 12800 30 14630 60
rect 14660 30 16490 60
rect 16520 30 16730 60
rect 6260 -30 6400 0
rect 6430 -30 16730 0
rect 6260 -2830 16730 -2820
rect 6260 -2910 6400 -2830
rect 6430 -2910 7250 -2830
rect 7280 -2910 8260 -2830
rect 8290 -2910 10120 -2830
rect 10150 -2910 11050 -2830
rect 11080 -2910 11980 -2830
rect 12010 -2910 13840 -2830
rect 13870 -2910 15700 -2830
rect 15730 -2910 16550 -2830
rect 16580 -2910 16730 -2830
rect 6260 -2920 16730 -2910
use p8_1  p8_1_7
timestamp 1633783901
transform -1 0 6940 0 -1 -120
box -370 -140 570 2690
use p1_8  p1_8_6
timestamp 1633696558
transform -1 0 12520 0 -1 -120
box -370 -140 570 2690
use p8_1  p8_1_10
timestamp 1633783901
transform -1 0 11590 0 -1 -120
box -370 -140 570 2690
use p1_8  p1_8_5
timestamp 1633696558
transform -1 0 10660 0 -1 -120
box -370 -140 570 2690
use p8_1  p8_1_9
timestamp 1633783901
transform -1 0 9730 0 -1 -120
box -370 -140 570 2690
use p8_1  p8_1_8
timestamp 1633783901
transform -1 0 7870 0 -1 -120
box -370 -140 570 2690
use p1_8  p1_8_4
timestamp 1633696558
transform -1 0 8800 0 -1 -120
box -370 -140 570 2690
use p8_1  p8_1_12
timestamp 1633783901
transform -1 0 15310 0 -1 -120
box -370 -140 570 2690
use p8_1  p8_1_13
timestamp 1633783901
transform -1 0 16240 0 -1 -120
box -370 -140 570 2690
use p1_8  p1_8_7
timestamp 1633696558
transform -1 0 14380 0 -1 -120
box -370 -140 570 2690
use p8_1  p8_1_11
timestamp 1633783901
transform -1 0 13450 0 -1 -120
box -370 -140 570 2690
use p8_1  p8_1_0
timestamp 1633783901
transform 1 0 6740 0 1 2150
box -370 -140 570 2690
use p8_1  p8_1_1
timestamp 1633783901
transform 1 0 7670 0 1 2150
box -370 -140 570 2690
use p8_1  p8_1_2
timestamp 1633783901
transform 1 0 9530 0 1 2150
box -370 -140 570 2690
use p1_8  p1_8_0
timestamp 1633696558
transform 1 0 8600 0 1 2150
box -370 -140 570 2690
use p8_1  p8_1_3
timestamp 1633783901
transform 1 0 11390 0 1 2150
box -370 -140 570 2690
use p1_8  p1_8_1
timestamp 1633696558
transform 1 0 10460 0 1 2150
box -370 -140 570 2690
use p1_8  p1_8_2
timestamp 1633696558
transform 1 0 12320 0 1 2150
box -370 -140 570 2690
use p8_1  p8_1_6
timestamp 1633783901
transform 1 0 16040 0 1 2150
box -370 -140 570 2690
use p8_1  p8_1_4
timestamp 1633783901
transform 1 0 13250 0 1 2150
box -370 -140 570 2690
use p8_1  p8_1_5
timestamp 1633783901
transform 1 0 15110 0 1 2150
box -370 -140 570 2690
use p1_8  p1_8_3
timestamp 1633696558
transform 1 0 14180 0 1 2150
box -370 -140 570 2690
<< labels >>
rlabel metal2 6250 1970 6260 2000 3 ib
port 1 e
rlabel metal2 6250 1850 6260 1880 3 ga
port 2 e
rlabel metal2 6250 1730 6260 1760 3 da
port 3 e
rlabel metal2 6250 1610 6260 1640 3 gb
port 4 e
rlabel metal2 6250 1490 6260 1520 3 db
port 5 e
rlabel metal2 6250 1180 6260 1210 3 gc
port 7 e
rlabel metal2 6250 1060 6260 1090 3 dc
port 8 e
rlabel metal2 6250 940 6260 970 3 gd
port 9 e
rlabel metal2 6250 820 6260 850 3 dd
port 10 e
rlabel metal2 6250 4850 6260 4950 3 vdda
port 11 e
rlabel metal2 6250 1300 6260 1400 3 gnd
port 12 e
<< end >>
