magic
tech sky130A
magscale 1 2
timestamp 1630377360
<< error_s >>
rect 5244 1644 5302 1650
rect 5244 1610 5256 1644
rect 5244 1604 5302 1610
rect 5244 1450 5302 1456
rect 5244 1416 5256 1450
rect 5244 1410 5302 1416
<< nmos >>
rect -200 1820 1600 2020
rect -200 1560 1600 1760
rect -200 1300 1600 1500
rect -200 1040 1600 1240
rect -200 780 1600 980
rect -200 520 1600 720
rect -200 260 1600 460
rect -200 0 1600 200
<< ndiff >>
rect -320 1980 -200 2020
rect -320 1860 -300 1980
rect -220 1860 -200 1980
rect -320 1820 -200 1860
rect 1600 1980 1720 2020
rect 1600 1860 1620 1980
rect 1700 1860 1720 1980
rect 1600 1820 1720 1860
rect -320 1720 -200 1760
rect -320 1600 -300 1720
rect -220 1600 -200 1720
rect -320 1560 -200 1600
rect 1600 1720 1720 1760
rect 1600 1600 1620 1720
rect 1700 1600 1720 1720
rect 1600 1560 1720 1600
rect -320 1460 -200 1500
rect -320 1340 -300 1460
rect -220 1340 -200 1460
rect -320 1300 -200 1340
rect 1600 1460 1720 1500
rect 1600 1340 1620 1460
rect 1700 1340 1720 1460
rect 1600 1300 1720 1340
rect -320 1200 -200 1240
rect -320 1080 -300 1200
rect -220 1080 -200 1200
rect -320 1040 -200 1080
rect 1600 1200 1720 1240
rect 1600 1080 1620 1200
rect 1700 1080 1720 1200
rect 1600 1040 1720 1080
rect -320 940 -200 980
rect -320 820 -300 940
rect -220 820 -200 940
rect -320 780 -200 820
rect 1600 940 1720 980
rect 1600 820 1620 940
rect 1700 820 1720 940
rect 1600 780 1720 820
rect -320 680 -200 720
rect -320 560 -300 680
rect -220 560 -200 680
rect -320 520 -200 560
rect 1600 680 1720 720
rect 1600 560 1620 680
rect 1700 560 1720 680
rect 1600 520 1720 560
rect -320 420 -200 460
rect -320 300 -300 420
rect -220 300 -200 420
rect -320 260 -200 300
rect 1600 420 1720 460
rect 1600 300 1620 420
rect 1700 300 1720 420
rect 1600 260 1720 300
rect -320 160 -200 200
rect -320 40 -300 160
rect -220 40 -200 160
rect -320 0 -200 40
rect 1600 160 1720 200
rect 1600 40 1620 160
rect 1700 40 1720 160
rect 1600 0 1720 40
<< ndiffc >>
rect -300 1860 -220 1980
rect 1620 1860 1700 1980
rect -300 1600 -220 1720
rect 1620 1600 1700 1720
rect -300 1340 -220 1460
rect 1620 1340 1700 1460
rect -300 1080 -220 1200
rect 1620 1080 1700 1200
rect -300 820 -220 940
rect 1620 820 1700 940
rect -300 560 -220 680
rect 1620 560 1700 680
rect -300 300 -220 420
rect 1620 300 1700 420
rect -300 40 -220 160
rect 1620 40 1700 160
<< psubdiff >>
rect -320 -140 -280 -60
rect 1680 -140 1720 -60
<< psubdiffcont >>
rect -280 -140 1680 -60
<< poly >>
rect -200 2140 1600 2160
rect -200 2080 -180 2140
rect 1580 2080 1600 2140
rect -200 2020 1600 2080
rect -200 1760 1600 1820
rect -200 1500 1600 1560
rect -200 1240 1600 1300
rect -200 980 1600 1040
rect -200 720 1600 780
rect -200 460 1600 520
rect -200 200 1600 260
rect -200 -40 1600 0
<< polycont >>
rect -180 2080 1580 2140
<< locali >>
rect -200 2080 -180 2140
rect 1580 2080 1600 2140
rect -300 1980 -220 2020
rect -300 1720 -220 1860
rect -300 1460 -220 1600
rect -300 1200 -220 1340
rect -300 940 -220 1080
rect -300 680 -220 820
rect -300 420 -220 560
rect -300 160 -220 300
rect -300 0 -220 40
rect 1620 1980 1700 2020
rect 1620 1720 1700 1860
rect 1620 1460 1700 1600
rect 1620 1200 1700 1340
rect 1620 940 1700 1080
rect 1620 680 1700 820
rect 1620 420 1700 560
rect 1620 160 1700 300
rect 1620 0 1700 40
rect -320 -140 -280 -60
rect 1680 -140 1720 -60
use sky130_fd_pr__nfet_01v8_E5V3SC  sky130_fd_pr__nfet_01v8_E5V3SC_0
timestamp 1630377360
transform 1 0 5273 0 1 1530
box -73 -130 73 130
use sky130_fd_pr__nfet_01v8_lvt_L8NDKD  sky130_fd_pr__nfet_01v8_lvt_L8NDKD_0
timestamp 1630377360
transform 1 0 6543 0 1 1457
box -996 -310 996 310
use sky130_fd_pr__rf_npn_05v5_W1p00L1p00  sky130_fd_pr__rf_npn_05v5_W1p00L1p00_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1621640962
transform 1 0 2200 0 1 600
box 0 0 1724 1724
<< labels >>
rlabel ndiffc 1660 1920 1660 1920 1 D
port 1 n
rlabel locali -180 2120 -180 2120 1 G
port 2 n
rlabel locali -260 220 -260 220 1 S
port 3 n
rlabel locali -300 -100 -300 -100 1 B
port 4 n
<< end >>
