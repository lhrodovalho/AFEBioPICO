* OpAmp open-loop dc testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "../mag/opamp_core.spice"

* supply voltages
vdda  vdda 0 dc 1.8 pulse(1.7 1.8 1m 100u 100u 10 1)
*vdda  vdda 0 dc 1.8
vssa  vssa 0 0.0


* DUT
x0 j in out ib q vdda bp vddx gnda vssa xn xp x y z opamp_core
ib vdda ib 1n
cl out gnda 100p
rf out j    9Meg
ri j   gnda 1Meg

* input signals
egnda gnda vssa ib vssa 1
vin in gnda dc 0 ac 1 pulse(-50m 50m 0 10u 10u 50m 100m)

*.option method="Gear"
.option gmin=1e-15
.control

	op	
	print i(vdda) v(q) v(ib)
	
	ac dec 100 1m 1Meg
	plot vdb(out)
	plot phase(out)*180/PI

	tran 100u 400m
	plot in out q ib
.endc

.end
